

module b22_C_gen_AntiSAT_k_128_6 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390;

  NAND2_X1 U7211 ( .A1(n14010), .A2(n14201), .ZN(n13998) );
  AND2_X1 U7212 ( .A1(n15002), .A2(n12246), .ZN(n12267) );
  AND2_X1 U7213 ( .A1(n7050), .A2(n6527), .ZN(n15001) );
  BUF_X2 U7214 ( .A(n10703), .Z(n6468) );
  AND3_X1 U7215 ( .A1(n6513), .A2(n6938), .A3(n6936), .ZN(n14225) );
  AND2_X1 U7216 ( .A1(n8968), .A2(n11332), .ZN(n6486) );
  OAI21_X1 U7218 ( .B1(n7683), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U7219 ( .A1(n14225), .A2(n14614), .ZN(n13490) );
  INV_X2 U7220 ( .A(n11477), .ZN(n11410) );
  OR2_X1 U7221 ( .A1(n13946), .A2(n13950), .ZN(n13947) );
  INV_X1 U7222 ( .A(n12233), .ZN(n15097) );
  OR2_X1 U7223 ( .A1(n15001), .A2(n12245), .ZN(n15002) );
  NAND2_X1 U7224 ( .A1(n11077), .A2(n11082), .ZN(n12451) );
  NOR2_X1 U7225 ( .A1(n6512), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U7226 ( .A1(n11991), .A2(n11990), .ZN(n12000) );
  INV_X1 U7227 ( .A(n11743), .ZN(n8948) );
  NAND2_X1 U7228 ( .A1(n11176), .A2(n11175), .ZN(n11466) );
  OAI211_X1 U7229 ( .C1(n11335), .C2(n9285), .A(n9284), .B(n9283), .ZN(n13498)
         );
  XNOR2_X1 U7230 ( .A(n11925), .B(n11924), .ZN(n14216) );
  NAND4_X1 U7231 ( .A1(n8954), .A2(n8953), .A3(n8952), .A4(n8951), .ZN(n12894)
         );
  INV_X1 U7232 ( .A(n13601), .ZN(n14188) );
  OR2_X1 U7233 ( .A1(n11641), .A2(n10139), .ZN(n14713) );
  AOI21_X2 U7234 ( .B1(n10295), .B2(n12015), .A(n6927), .ZN(n10450) );
  OAI21_X2 U7235 ( .B1(n10280), .B2(n12013), .A(n6541), .ZN(n10295) );
  AOI21_X2 U7236 ( .B1(n13824), .B2(n14699), .A(n13823), .ZN(n14059) );
  NAND2_X2 U7237 ( .A1(n8207), .A2(n8263), .ZN(n10965) );
  NAND4_X2 U7238 ( .A1(n8987), .A2(n8986), .A3(n8985), .A4(n8984), .ZN(n12895)
         );
  NAND3_X2 U7239 ( .A1(n6528), .A2(n7809), .A3(n7811), .ZN(n12233) );
  AOI21_X2 U7240 ( .B1(n15061), .B2(n7185), .A(n7184), .ZN(n7183) );
  NOR2_X2 U7241 ( .A1(n13947), .A2(n13601), .ZN(n7211) );
  AND2_X2 U7242 ( .A1(n14224), .A2(n11335), .ZN(n13601) );
  NAND2_X1 U7243 ( .A1(n9054), .A2(n9053), .ZN(n6463) );
  NAND2_X1 U7244 ( .A1(n9054), .A2(n9053), .ZN(n9589) );
  NOR2_X2 U7245 ( .A1(n6519), .A2(n14475), .ZN(n14482) );
  XNOR2_X2 U7246 ( .A(n8442), .B(n8441), .ZN(n9097) );
  OAI21_X2 U7247 ( .B1(n8447), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8442) );
  XNOR2_X2 U7248 ( .A(n6863), .B(n8900), .ZN(n8902) );
  NAND2_X2 U7249 ( .A1(n11928), .A2(n11927), .ZN(n13256) );
  INV_X2 U7250 ( .A(n14016), .ZN(n6464) );
  INV_X2 U7251 ( .A(n11782), .ZN(n11984) );
  INV_X4 U7252 ( .A(n11276), .ZN(n11436) );
  NAND4_X1 U7253 ( .A1(n9616), .A2(n9615), .A3(n9614), .A4(n9613), .ZN(n13728)
         );
  INV_X4 U7254 ( .A(n13520), .ZN(n6465) );
  INV_X4 U7255 ( .A(n11276), .ZN(n11459) );
  CLKBUF_X2 U7256 ( .A(P2_U3947), .Z(n6467) );
  CLKBUF_X2 U7257 ( .A(n8277), .Z(n12051) );
  INV_X1 U7259 ( .A(n13638), .ZN(n11483) );
  CLKBUF_X2 U7260 ( .A(n12402), .Z(n6480) );
  INV_X2 U7261 ( .A(n11632), .ZN(n13639) );
  NAND2_X2 U7262 ( .A1(n9055), .A2(n9050), .ZN(n13638) );
  XNOR2_X1 U7263 ( .A(n8069), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12402) );
  CLKBUF_X2 U7264 ( .A(n9051), .Z(n9050) );
  OR2_X1 U7265 ( .A1(n6534), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8209) );
  NOR2_X1 U7266 ( .A1(n8435), .A2(n8434), .ZN(n8436) );
  INV_X1 U7267 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8599) );
  OAI21_X1 U7268 ( .B1(n12419), .B2(n12579), .A(n12418), .ZN(n6913) );
  MUX2_X1 U7269 ( .A(n14166), .B(n14165), .S(n14713), .Z(n14167) );
  NOR2_X1 U7270 ( .A1(n12645), .A2(n6915), .ZN(n12717) );
  NOR2_X1 U7271 ( .A1(n12641), .A2(n6533), .ZN(n12714) );
  NAND2_X1 U7272 ( .A1(n12442), .A2(n6550), .ZN(n12645) );
  AND2_X1 U7273 ( .A1(n12646), .A2(n15148), .ZN(n6915) );
  NAND2_X1 U7274 ( .A1(n13478), .A2(n13479), .ZN(n13477) );
  NAND2_X1 U7275 ( .A1(n13415), .A2(n11418), .ZN(n13478) );
  OAI211_X1 U7276 ( .C1(n12424), .C2(n8189), .A(n15099), .B(n12423), .ZN(
        n12426) );
  NAND2_X1 U7277 ( .A1(n12839), .A2(n11670), .ZN(n12798) );
  NAND2_X1 U7278 ( .A1(n12165), .A2(n6697), .ZN(n7416) );
  NAND2_X1 U7279 ( .A1(n8174), .A2(n6830), .ZN(n12438) );
  NAND2_X1 U7280 ( .A1(n12488), .A2(n11071), .ZN(n12464) );
  AOI21_X1 U7281 ( .B1(n7128), .B2(n15007), .A(n7125), .ZN(n12403) );
  NOR2_X1 U7282 ( .A1(n12380), .A2(n12379), .ZN(n12384) );
  AND2_X1 U7283 ( .A1(n12380), .A2(n12379), .ZN(n7166) );
  NAND2_X1 U7284 ( .A1(n12518), .A2(n8104), .ZN(n12507) );
  NAND2_X1 U7285 ( .A1(n8091), .A2(n6828), .ZN(n12518) );
  AND2_X1 U7286 ( .A1(n7329), .A2(n7331), .ZN(n14379) );
  OR2_X1 U7287 ( .A1(n12293), .A2(n12698), .ZN(n7028) );
  AND2_X1 U7288 ( .A1(n13933), .A2(n7384), .ZN(n7383) );
  NAND2_X1 U7289 ( .A1(n6917), .A2(n6644), .ZN(n12582) );
  XNOR2_X1 U7290 ( .A(n12330), .B(n12331), .ZN(n12293) );
  NAND2_X1 U7291 ( .A1(n7162), .A2(n7161), .ZN(n12292) );
  NAND2_X1 U7292 ( .A1(n6658), .A2(n6525), .ZN(n7277) );
  NOR2_X1 U7293 ( .A1(n6952), .A2(n14473), .ZN(n14476) );
  OR2_X1 U7294 ( .A1(n12296), .A2(n12297), .ZN(n6658) );
  NAND2_X1 U7295 ( .A1(n10925), .A2(n13549), .ZN(n11614) );
  OAI21_X1 U7296 ( .B1(n14353), .B2(n7990), .A(n7989), .ZN(n12618) );
  OAI21_X1 U7297 ( .B1(n12105), .B2(n8310), .A(n8309), .ZN(n12159) );
  NAND2_X1 U7298 ( .A1(n6825), .A2(n7975), .ZN(n14353) );
  OR2_X1 U7299 ( .A1(n12274), .A2(n12275), .ZN(n7280) );
  OAI21_X1 U7300 ( .B1(n9788), .B2(n7286), .A(n7284), .ZN(n9910) );
  OAI21_X1 U7301 ( .B1(n7174), .B2(n6647), .A(n6645), .ZN(n10754) );
  NAND2_X1 U7302 ( .A1(n7959), .A2(n7958), .ZN(n10750) );
  NAND2_X1 U7303 ( .A1(n10106), .A2(n10105), .ZN(n10255) );
  AND2_X1 U7304 ( .A1(n6753), .A2(n6593), .ZN(n10321) );
  NAND2_X1 U7305 ( .A1(n8225), .A2(n11002), .ZN(n15035) );
  AOI21_X1 U7306 ( .B1(n7580), .B2(n7578), .A(n7577), .ZN(n10666) );
  AND2_X1 U7307 ( .A1(n14984), .A2(n14985), .ZN(n14987) );
  OR2_X1 U7308 ( .A1(n14390), .A2(n7206), .ZN(n7205) );
  AND2_X1 U7309 ( .A1(n14979), .A2(n10575), .ZN(n12241) );
  NAND2_X1 U7310 ( .A1(n10271), .A2(n6696), .ZN(n12068) );
  OAI21_X1 U7311 ( .B1(n14579), .B2(n6573), .A(n7409), .ZN(n14560) );
  NAND2_X1 U7312 ( .A1(n10466), .A2(n10465), .ZN(n11866) );
  NAND2_X1 U7313 ( .A1(n10461), .A2(n10460), .ZN(n11860) );
  NAND2_X1 U7314 ( .A1(n7118), .A2(n10308), .ZN(n11851) );
  OAI21_X1 U7315 ( .B1(n9469), .B2(n6859), .A(n6858), .ZN(n9626) );
  NAND2_X1 U7316 ( .A1(n7158), .A2(n7157), .ZN(n10236) );
  NAND2_X1 U7317 ( .A1(n6518), .A2(n7045), .ZN(n7158) );
  INV_X2 U7318 ( .A(n9837), .ZN(n14016) );
  AOI21_X1 U7319 ( .B1(n7422), .B2(n9895), .A(n6700), .ZN(n7421) );
  OAI21_X1 U7320 ( .B1(n8687), .B2(n6840), .A(n6838), .ZN(n9002) );
  NAND2_X1 U7321 ( .A1(n8923), .A2(n8899), .ZN(n12877) );
  OR2_X1 U7322 ( .A1(n14962), .A2(n9866), .ZN(n7069) );
  OR2_X1 U7323 ( .A1(n9035), .A2(n9034), .ZN(n9260) );
  INV_X2 U7324 ( .A(n13155), .ZN(n6466) );
  AND2_X1 U7325 ( .A1(n9185), .A2(n9073), .ZN(n9094) );
  NAND2_X1 U7326 ( .A1(n9645), .A2(n9644), .ZN(n11826) );
  NAND2_X1 U7327 ( .A1(n14937), .A2(n14938), .ZN(n14936) );
  OAI21_X1 U7328 ( .B1(n6979), .B2(n12051), .A(n15089), .ZN(n6978) );
  NOR2_X1 U7329 ( .A1(n14960), .A2(n14961), .ZN(n14962) );
  INV_X1 U7330 ( .A(n12824), .ZN(n14836) );
  INV_X1 U7331 ( .A(n6469), .ZN(n6472) );
  INV_X4 U7332 ( .A(n9289), .ZN(n11367) );
  NAND4_X1 U7333 ( .A1(n7918), .A2(n7917), .A3(n7916), .A4(n7915), .ZN(n15024)
         );
  NAND2_X1 U7334 ( .A1(n9576), .A2(n9575), .ZN(n14602) );
  CLKBUF_X2 U7335 ( .A(n11051), .Z(n6476) );
  INV_X1 U7336 ( .A(n9327), .ZN(n11579) );
  CLKBUF_X3 U7337 ( .A(n9327), .Z(n11736) );
  NAND2_X1 U7338 ( .A1(n8519), .A2(n8518), .ZN(n8537) );
  NAND4_X2 U7339 ( .A1(n9133), .A2(n9132), .A3(n9131), .A4(n9130), .ZN(n14636)
         );
  NAND2_X2 U7340 ( .A1(n13490), .A2(n9838), .ZN(n11477) );
  INV_X4 U7341 ( .A(n11234), .ZN(n11276) );
  NAND4_X2 U7342 ( .A1(n9060), .A2(n9059), .A3(n9058), .A4(n9057), .ZN(n13732)
         );
  AND3_X1 U7343 ( .A1(n7832), .A2(n7831), .A3(n7830), .ZN(n9898) );
  AND2_X1 U7344 ( .A1(n6688), .A2(n6606), .ZN(n12760) );
  AND2_X1 U7345 ( .A1(n7723), .A2(n12768), .ZN(n7807) );
  NOR2_X1 U7346 ( .A1(n9280), .A2(n9079), .ZN(n9081) );
  XNOR2_X1 U7347 ( .A(n8205), .B(n8204), .ZN(n10853) );
  NAND2_X1 U7348 ( .A1(n6977), .A2(n6975), .ZN(n14614) );
  XNOR2_X1 U7349 ( .A(n8445), .B(n8444), .ZN(n9095) );
  NOR2_X2 U7350 ( .A1(n9463), .A2(n12003), .ZN(n13332) );
  NAND2_X2 U7351 ( .A1(n9140), .A2(n8945), .ZN(n8096) );
  AND2_X2 U7352 ( .A1(n9054), .A2(n9050), .ZN(n11632) );
  NAND2_X1 U7353 ( .A1(n6997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6996) );
  NAND2_X2 U7354 ( .A1(n13365), .A2(n8622), .ZN(n8968) );
  NAND2_X2 U7355 ( .A1(n8213), .A2(n8212), .ZN(n9140) );
  NAND3_X1 U7356 ( .A1(n7369), .A2(n7368), .A3(n7370), .ZN(n9054) );
  NAND2_X1 U7357 ( .A1(n8203), .A2(n8202), .ZN(n8263) );
  NAND2_X1 U7358 ( .A1(n8210), .A2(n8209), .ZN(n9452) );
  NAND2_X1 U7359 ( .A1(n9046), .A2(n7373), .ZN(n7368) );
  OR2_X1 U7360 ( .A1(n9046), .A2(n7374), .ZN(n7369) );
  NAND2_X1 U7361 ( .A1(n8244), .A2(n8243), .ZN(n10372) );
  INV_X1 U7362 ( .A(n8209), .ZN(n8203) );
  NAND2_X1 U7363 ( .A1(n7016), .A2(n7014), .ZN(n13365) );
  INV_X1 U7364 ( .A(n9047), .ZN(n9046) );
  NAND2_X2 U7365 ( .A1(n8902), .A2(n7022), .ZN(n11743) );
  XNOR2_X1 U7366 ( .A(n6794), .B(n8901), .ZN(n7022) );
  NAND2_X1 U7367 ( .A1(n7531), .A2(n8755), .ZN(n9045) );
  NAND2_X1 U7368 ( .A1(n7962), .A2(n7582), .ZN(n7978) );
  INV_X4 U7369 ( .A(n8945), .ZN(n11332) );
  INV_X2 U7370 ( .A(n8494), .ZN(n8945) );
  AND2_X2 U7371 ( .A1(n6948), .A2(n6947), .ZN(n8494) );
  AND2_X1 U7372 ( .A1(n7582), .A2(n7581), .ZN(n6496) );
  OAI21_X1 U7373 ( .B1(n7372), .B2(n14210), .A(n7371), .ZN(n7370) );
  NAND2_X1 U7374 ( .A1(n7027), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7814) );
  AND3_X1 U7375 ( .A1(n8400), .A2(n8399), .A3(n8398), .ZN(n8781) );
  AND3_X1 U7376 ( .A1(n8569), .A2(n8555), .A3(n8551), .ZN(n8780) );
  AND3_X1 U7377 ( .A1(n7614), .A2(n7613), .A3(n7612), .ZN(n8401) );
  AND2_X1 U7378 ( .A1(n7706), .A2(n7707), .ZN(n7582) );
  AND3_X1 U7379 ( .A1(n7214), .A2(n7213), .A3(n7212), .ZN(n7390) );
  NAND4_X1 U7380 ( .A1(n10809), .A2(n7095), .A3(n7094), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6948) );
  NAND4_X1 U7381 ( .A1(n15184), .A2(n7093), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6947) );
  INV_X4 U7382 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7383 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8822) );
  XNOR2_X1 U7384 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14285) );
  INV_X1 U7385 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6973) );
  INV_X1 U7386 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7993) );
  NOR2_X1 U7387 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7614) );
  NOR2_X1 U7388 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8400) );
  NOR2_X1 U7389 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7613) );
  INV_X1 U7390 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8202) );
  NOR2_X1 U7391 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7705) );
  NOR2_X1 U7392 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7704) );
  NOR2_X1 U7393 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n7212) );
  NOR2_X1 U7394 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n7213) );
  NOR2_X1 U7395 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n7214) );
  INV_X1 U7396 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8204) );
  INV_X1 U7397 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8441) );
  INV_X1 U7398 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8569) );
  INV_X1 U7399 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8264) );
  INV_X1 U7400 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8551) );
  NOR2_X1 U7401 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7710) );
  NOR2_X1 U7402 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8398) );
  NOR2_X1 U7403 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n7709) );
  INV_X4 U7404 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7405 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8602) );
  NOR2_X1 U7406 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7556) );
  NOR2_X1 U7407 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8399) );
  NAND2_X1 U7408 ( .A1(n13407), .A2(n13406), .ZN(n13456) );
  AOI21_X2 U7409 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n9498), .A(n9497), .ZN(
        n9499) );
  AOI22_X2 U7410 ( .A1(n12133), .A2(n12132), .B1(n12570), .B2(n8320), .ZN(
        n12185) );
  INV_X1 U7411 ( .A(n11938), .ZN(n6469) );
  INV_X1 U7412 ( .A(n6469), .ZN(n6470) );
  INV_X2 U7413 ( .A(n6469), .ZN(n6471) );
  CLKBUF_X1 U7414 ( .A(n8341), .Z(n6473) );
  BUF_X4 U7415 ( .A(n8341), .Z(n6474) );
  INV_X1 U7416 ( .A(n8277), .ZN(n8341) );
  AOI211_X2 U7417 ( .C1(n12457), .C2(n15099), .A(n12456), .B(n12455), .ZN(
        n12651) );
  BUF_X2 U7418 ( .A(n11051), .Z(n6475) );
  NAND2_X1 U7419 ( .A1(n10960), .A2(n11160), .ZN(n11051) );
  NOR2_X2 U7420 ( .A1(n13998), .A2(n13981), .ZN(n13979) );
  XNOR2_X2 U7421 ( .A(n10255), .B(SI_22_), .ZN(n11333) );
  XNOR2_X2 U7422 ( .A(n7786), .B(n7716), .ZN(n8212) );
  OR3_X4 U7423 ( .A1(n9097), .A2(n10747), .A3(n9095), .ZN(n9122) );
  CLKBUF_X1 U7424 ( .A(n7807), .Z(n6478) );
  BUF_X4 U7425 ( .A(n7807), .Z(n6479) );
  AND2_X4 U7426 ( .A1(n12048), .A2(n12768), .ZN(n7806) );
  BUF_X4 U7427 ( .A(n7805), .Z(n6481) );
  BUF_X4 U7428 ( .A(n7805), .Z(n6482) );
  NAND2_X1 U7429 ( .A1(n11906), .A2(n7655), .ZN(n7654) );
  INV_X1 U7430 ( .A(n10988), .ZN(n7185) );
  NAND2_X1 U7431 ( .A1(n10973), .A2(n10972), .ZN(n6958) );
  NOR2_X1 U7432 ( .A1(n12433), .A2(n6831), .ZN(n6830) );
  INV_X1 U7433 ( .A(n8173), .ZN(n6831) );
  OAI21_X1 U7434 ( .B1(n7824), .B2(n7338), .A(n7840), .ZN(n6777) );
  AOI21_X1 U7435 ( .B1(n8671), .B2(n6850), .A(n6571), .ZN(n6847) );
  INV_X1 U7436 ( .A(n9885), .ZN(n7157) );
  NAND2_X1 U7437 ( .A1(n7069), .A2(n7068), .ZN(n10223) );
  INV_X1 U7438 ( .A(n9868), .ZN(n7068) );
  NAND2_X1 U7439 ( .A1(n15010), .A2(n15009), .ZN(n15008) );
  AND2_X1 U7440 ( .A1(n11091), .A2(n8232), .ZN(n12421) );
  OR2_X1 U7441 ( .A1(n12681), .A2(n8322), .ZN(n11040) );
  NOR2_X1 U7442 ( .A1(n13987), .A2(n7393), .ZN(n7392) );
  AOI21_X1 U7443 ( .B1(n7248), .B2(n7250), .A(n7246), .ZN(n7245) );
  AOI22_X1 U7444 ( .A1(n12894), .A2(n11782), .B1(n11801), .B2(n11902), .ZN(
        n11802) );
  NAND2_X1 U7445 ( .A1(n7641), .A2(n7647), .ZN(n7646) );
  INV_X1 U7446 ( .A(n11802), .ZN(n7641) );
  INV_X1 U7447 ( .A(n11803), .ZN(n7647) );
  NAND2_X1 U7448 ( .A1(n6999), .A2(n6998), .ZN(n6990) );
  INV_X1 U7449 ( .A(n11813), .ZN(n6998) );
  MUX2_X1 U7450 ( .A(n14437), .B(n14390), .S(n6465), .Z(n13576) );
  AND2_X1 U7451 ( .A1(n11861), .A2(n11862), .ZN(n7635) );
  NOR2_X1 U7452 ( .A1(n6885), .A2(n11854), .ZN(n6884) );
  NAND2_X1 U7453 ( .A1(n7634), .A2(n7633), .ZN(n7632) );
  INV_X1 U7454 ( .A(n11862), .ZN(n7634) );
  INV_X1 U7455 ( .A(n11861), .ZN(n7633) );
  INV_X1 U7456 ( .A(n11904), .ZN(n7653) );
  AOI21_X1 U7457 ( .B1(n11070), .B2(n6491), .A(n6565), .ZN(n11072) );
  OAI21_X1 U7458 ( .B1(n11068), .B2(n11067), .A(n11066), .ZN(n7348) );
  INV_X1 U7459 ( .A(n7618), .ZN(n7617) );
  OAI21_X1 U7460 ( .B1(n7623), .B2(n11916), .A(n7619), .ZN(n7618) );
  NAND2_X1 U7461 ( .A1(n7622), .A2(n7620), .ZN(n7619) );
  INV_X1 U7462 ( .A(n7624), .ZN(n7623) );
  AND2_X1 U7463 ( .A1(n9941), .A2(n11812), .ZN(n7482) );
  AND2_X1 U7464 ( .A1(n13645), .A2(n13656), .ZN(n13487) );
  NAND2_X1 U7465 ( .A1(n7062), .A2(n7060), .ZN(n14234) );
  NAND2_X1 U7466 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7061), .ZN(n7060) );
  NAND2_X1 U7467 ( .A1(n14284), .A2(n14283), .ZN(n7062) );
  INV_X1 U7468 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7061) );
  XNOR2_X1 U7469 ( .A(n6474), .B(n10083), .ZN(n8286) );
  OR2_X1 U7470 ( .A1(n12061), .A2(n12440), .ZN(n11091) );
  OR2_X1 U7471 ( .A1(n12648), .A2(n12472), .ZN(n11077) );
  OR2_X1 U7472 ( .A1(n12665), .A2(n12523), .ZN(n11069) );
  OR2_X1 U7473 ( .A1(n12536), .A2(n12522), .ZN(n11056) );
  OR2_X1 U7474 ( .A1(n12752), .A2(n8315), .ZN(n11034) );
  INV_X1 U7475 ( .A(n7179), .ZN(n7178) );
  INV_X1 U7476 ( .A(n7177), .ZN(n7176) );
  OAI21_X1 U7477 ( .B1(n7180), .B2(n7178), .A(n11011), .ZN(n7177) );
  NAND2_X1 U7478 ( .A1(n6484), .A2(n7962), .ZN(n8249) );
  INV_X1 U7479 ( .A(n7575), .ZN(n7573) );
  NAND2_X1 U7480 ( .A1(n8068), .A2(n7769), .ZN(n7770) );
  AND2_X1 U7481 ( .A1(n9330), .A2(n9328), .ZN(n7471) );
  NOR2_X1 U7482 ( .A1(n7503), .A2(n10596), .ZN(n7502) );
  NAND2_X1 U7483 ( .A1(n8904), .A2(n8902), .ZN(n8955) );
  INV_X1 U7484 ( .A(n7022), .ZN(n8904) );
  OR2_X1 U7485 ( .A1(n13267), .A2(n12776), .ZN(n13017) );
  NAND2_X1 U7486 ( .A1(n13157), .A2(n13034), .ZN(n7451) );
  NAND2_X1 U7487 ( .A1(n13208), .A2(n7477), .ZN(n6903) );
  NOR2_X1 U7488 ( .A1(n6789), .A2(n6785), .ZN(n6784) );
  INV_X1 U7489 ( .A(n7673), .ZN(n6785) );
  INV_X1 U7490 ( .A(n7455), .ZN(n6789) );
  INV_X1 U7491 ( .A(n12896), .ZN(n9224) );
  AND2_X1 U7492 ( .A1(n11957), .A2(n9685), .ZN(n11762) );
  NAND2_X1 U7493 ( .A1(n7666), .A2(n8415), .ZN(n7138) );
  AND2_X1 U7494 ( .A1(n7140), .A2(n7139), .ZN(n8613) );
  NOR2_X1 U7495 ( .A1(n13850), .A2(n13830), .ZN(n7199) );
  NAND2_X1 U7496 ( .A1(n7386), .A2(n7385), .ZN(n7384) );
  INV_X1 U7497 ( .A(n7388), .ZN(n7385) );
  NOR2_X1 U7498 ( .A1(n13944), .A2(n7242), .ZN(n7241) );
  INV_X1 U7499 ( .A(n11603), .ZN(n7242) );
  OR2_X1 U7500 ( .A1(n14145), .A2(n14445), .ZN(n7207) );
  INV_X1 U7501 ( .A(n9051), .ZN(n9053) );
  OR2_X1 U7502 ( .A1(n13731), .A2(n10110), .ZN(n13494) );
  INV_X1 U7503 ( .A(n13487), .ZN(n9838) );
  INV_X1 U7504 ( .A(n8757), .ZN(n7531) );
  OAI21_X1 U7505 ( .B1(n10745), .B2(n10744), .A(n10746), .ZN(n11169) );
  XNOR2_X1 U7506 ( .A(n9717), .B(SI_20_), .ZN(n9716) );
  INV_X1 U7507 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9072) );
  INV_X1 U7508 ( .A(n6839), .ZN(n6838) );
  OAI21_X1 U7509 ( .B1(n6840), .B2(n7595), .A(n8996), .ZN(n6839) );
  NAND2_X1 U7510 ( .A1(n8687), .A2(n7598), .ZN(n8776) );
  AOI21_X1 U7511 ( .B1(n8580), .B2(n7593), .A(n6566), .ZN(n7592) );
  AND2_X1 U7512 ( .A1(n8335), .A2(n6698), .ZN(n6697) );
  INV_X1 U7513 ( .A(n8336), .ZN(n6698) );
  NAND2_X1 U7514 ( .A1(n12165), .A2(n8335), .ZN(n8337) );
  XNOR2_X1 U7515 ( .A(n12231), .B(n8286), .ZN(n10011) );
  NAND2_X1 U7516 ( .A1(n6701), .A2(n12232), .ZN(n7423) );
  INV_X1 U7517 ( .A(n8285), .ZN(n6701) );
  OAI21_X1 U7518 ( .B1(n9365), .B2(n14909), .A(n9146), .ZN(n9359) );
  OAI22_X1 U7519 ( .A1(n9307), .A2(n9306), .B1(n9178), .B2(n9319), .ZN(n14923)
         );
  NAND2_X1 U7520 ( .A1(n14923), .A2(n14922), .ZN(n14921) );
  AND2_X1 U7521 ( .A1(n9882), .A2(n9881), .ZN(n9883) );
  NAND2_X1 U7522 ( .A1(n10225), .A2(n7132), .ZN(n6811) );
  NAND2_X1 U7523 ( .A1(n10227), .A2(n10226), .ZN(n7132) );
  AND2_X1 U7524 ( .A1(n7054), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7052) );
  AND2_X1 U7525 ( .A1(n7122), .A2(n7121), .ZN(n15010) );
  NAND2_X1 U7526 ( .A1(n7133), .A2(n6631), .ZN(n12303) );
  AND2_X1 U7527 ( .A1(n12292), .A2(n12300), .ZN(n12330) );
  NAND2_X1 U7528 ( .A1(n7277), .A2(n12316), .ZN(n12349) );
  XNOR2_X1 U7529 ( .A(n7084), .B(n12371), .ZN(n12351) );
  NOR2_X1 U7530 ( .A1(n12351), .A2(n12350), .ZN(n12364) );
  AND2_X1 U7531 ( .A1(n12438), .A2(n8188), .ZN(n12424) );
  NAND2_X1 U7532 ( .A1(n12437), .A2(n12433), .ZN(n6984) );
  NAND2_X1 U7533 ( .A1(n8174), .A2(n8173), .ZN(n12437) );
  NAND2_X1 U7534 ( .A1(n12485), .A2(n11068), .ZN(n12488) );
  NOR2_X1 U7535 ( .A1(n12524), .A2(n6829), .ZN(n6828) );
  INV_X1 U7536 ( .A(n8090), .ZN(n6829) );
  NAND2_X1 U7537 ( .A1(n12563), .A2(n6553), .ZN(n12550) );
  NOR2_X1 U7538 ( .A1(n7942), .A2(n7579), .ZN(n7578) );
  NOR2_X1 U7539 ( .A1(n7944), .A2(n15019), .ZN(n7577) );
  INV_X1 U7540 ( .A(n7894), .ZN(n7579) );
  OAI211_X1 U7541 ( .C1(n10208), .C2(n6650), .A(n6649), .B(n11128), .ZN(n10397) );
  INV_X1 U7542 ( .A(n7819), .ZN(n7558) );
  INV_X1 U7543 ( .A(n12397), .ZN(n8213) );
  NAND2_X1 U7544 ( .A1(n12438), .A2(n6542), .ZN(n12423) );
  INV_X1 U7545 ( .A(n8096), .ZN(n11108) );
  INV_X1 U7546 ( .A(n7010), .ZN(n8070) );
  INV_X1 U7547 ( .A(n9140), .ZN(n8136) );
  OAI22_X1 U7548 ( .A1(n11099), .A2(n11098), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n12049), .ZN(n11106) );
  XNOR2_X1 U7549 ( .A(n7722), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U7550 ( .A1(n7721), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7722) );
  NOR2_X1 U7551 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(n7575), .ZN(n7574) );
  OAI21_X1 U7552 ( .B1(n8161), .B2(n7779), .A(n7780), .ZN(n8176) );
  NAND2_X1 U7553 ( .A1(n7351), .A2(n11302), .ZN(n7350) );
  INV_X1 U7554 ( .A(n8051), .ZN(n7340) );
  OAI21_X1 U7555 ( .B1(n7757), .B2(n6765), .A(n6763), .ZN(n8018) );
  INV_X1 U7556 ( .A(n6764), .ZN(n6763) );
  OAI21_X1 U7557 ( .B1(n7756), .B2(n6765), .A(n7354), .ZN(n6764) );
  AOI21_X1 U7558 ( .B1(n7356), .B2(n7758), .A(n7355), .ZN(n7354) );
  AND2_X1 U7559 ( .A1(n7736), .A2(n7735), .ZN(n7840) );
  NAND2_X1 U7560 ( .A1(n7825), .A2(n7824), .ZN(n7827) );
  CLKBUF_X2 U7561 ( .A(n8955), .Z(n11962) );
  BUF_X1 U7562 ( .A(n11726), .Z(n6950) );
  NAND2_X1 U7563 ( .A1(n6888), .A2(n7022), .ZN(n11726) );
  INV_X1 U7564 ( .A(n8902), .ZN(n6888) );
  OR2_X1 U7565 ( .A1(n7022), .A2(n8902), .ZN(n8956) );
  NOR2_X1 U7566 ( .A1(n8554), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U7567 ( .A1(n13069), .A2(n13068), .ZN(n13016) );
  OR2_X1 U7568 ( .A1(n6796), .A2(n13267), .ZN(n13061) );
  INV_X1 U7569 ( .A(n13077), .ZN(n13068) );
  AOI21_X1 U7570 ( .B1(n13146), .B2(n13150), .A(n7678), .ZN(n13134) );
  NAND2_X1 U7571 ( .A1(n6924), .A2(n6923), .ZN(n7450) );
  NAND2_X1 U7572 ( .A1(n13187), .A2(n13030), .ZN(n6923) );
  NAND2_X1 U7573 ( .A1(n13177), .A2(n13031), .ZN(n6924) );
  AND2_X1 U7574 ( .A1(n6905), .A2(n6904), .ZN(n13208) );
  NAND2_X1 U7575 ( .A1(n13323), .A2(n13025), .ZN(n6904) );
  OR2_X1 U7576 ( .A1(n7150), .A2(n13025), .ZN(n7674) );
  AND2_X1 U7577 ( .A1(n13331), .A2(n11187), .ZN(n7499) );
  AOI21_X1 U7578 ( .B1(n10876), .B2(n10875), .A(n6922), .ZN(n10879) );
  NOR2_X1 U7579 ( .A1(n13331), .A2(n12883), .ZN(n6922) );
  OR2_X1 U7580 ( .A1(n11851), .A2(n12886), .ZN(n10521) );
  NAND2_X1 U7581 ( .A1(n6582), .A2(n6489), .ZN(n7520) );
  AND2_X1 U7582 ( .A1(n11851), .A2(n11853), .ZN(n7525) );
  INV_X1 U7583 ( .A(n7526), .ZN(n7523) );
  NAND2_X1 U7584 ( .A1(n14878), .A2(n7527), .ZN(n7526) );
  AND2_X1 U7585 ( .A1(n14878), .A2(n12887), .ZN(n7439) );
  CLKBUF_X2 U7586 ( .A(n6486), .Z(n11951) );
  NAND2_X1 U7587 ( .A1(n9918), .A2(n14836), .ZN(n7461) );
  NAND2_X1 U7588 ( .A1(n9919), .A2(n7462), .ZN(n7460) );
  OR2_X1 U7589 ( .A1(n14836), .A2(n9918), .ZN(n7462) );
  NAND2_X1 U7590 ( .A1(n11258), .A2(n6486), .ZN(n10878) );
  NOR2_X1 U7591 ( .A1(n6886), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n7140) );
  AND2_X1 U7592 ( .A1(n8785), .A2(n8817), .ZN(n12948) );
  NAND2_X1 U7593 ( .A1(n7612), .A2(n8456), .ZN(n8546) );
  INV_X1 U7594 ( .A(n13723), .ZN(n10649) );
  NAND2_X1 U7595 ( .A1(n9573), .A2(n7287), .ZN(n13389) );
  NOR2_X1 U7596 ( .A1(n13387), .A2(n7288), .ZN(n7287) );
  INV_X1 U7597 ( .A(n9572), .ZN(n7288) );
  NAND2_X1 U7598 ( .A1(n10384), .A2(n7290), .ZN(n10507) );
  NOR2_X1 U7599 ( .A1(n10387), .A2(n7291), .ZN(n7290) );
  INV_X1 U7600 ( .A(n10383), .ZN(n7291) );
  NAND2_X1 U7601 ( .A1(n7325), .A2(n7328), .ZN(n7324) );
  INV_X1 U7602 ( .A(n14386), .ZN(n7325) );
  NAND2_X1 U7603 ( .A1(n7199), .A2(n7198), .ZN(n13811) );
  NOR2_X1 U7604 ( .A1(n13842), .A2(n6520), .ZN(n13825) );
  NAND2_X1 U7605 ( .A1(n13825), .A2(n13818), .ZN(n13829) );
  NOR2_X1 U7606 ( .A1(n13844), .A2(n13843), .ZN(n13842) );
  NAND2_X1 U7607 ( .A1(n13967), .A2(n11603), .ZN(n7240) );
  INV_X1 U7608 ( .A(n13669), .ZN(n7252) );
  NAND2_X1 U7609 ( .A1(n11225), .A2(n11224), .ZN(n13981) );
  AOI21_X1 U7610 ( .B1(n7402), .B2(n13688), .A(n6551), .ZN(n7401) );
  NAND2_X1 U7611 ( .A1(n14024), .A2(n11599), .ZN(n14007) );
  OR2_X1 U7612 ( .A1(n14145), .A2(n14374), .ZN(n13562) );
  OAI21_X1 U7613 ( .B1(n10718), .B2(n10717), .A(n10716), .ZN(n10760) );
  NAND2_X1 U7614 ( .A1(n7413), .A2(n14578), .ZN(n7412) );
  NAND2_X2 U7615 ( .A1(n11594), .A2(n14496), .ZN(n11335) );
  OAI21_X1 U7616 ( .B1(n11466), .B2(n7603), .A(n7601), .ZN(n11922) );
  AOI21_X1 U7617 ( .B1(n7604), .B2(n7602), .A(n6634), .ZN(n7601) );
  INV_X1 U7618 ( .A(n7604), .ZN(n7603) );
  XNOR2_X1 U7619 ( .A(n7119), .B(n7682), .ZN(n10607) );
  NAND2_X1 U7620 ( .A1(n8776), .A2(n8775), .ZN(n7119) );
  AND2_X1 U7621 ( .A1(n6721), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14286) );
  INV_X1 U7622 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6721) );
  AND2_X1 U7623 ( .A1(n6728), .A2(n6583), .ZN(n14303) );
  NAND2_X1 U7624 ( .A1(n6726), .A2(n6724), .ZN(n6723) );
  INV_X1 U7625 ( .A(n7278), .ZN(n10562) );
  NAND2_X1 U7626 ( .A1(n6934), .A2(n6465), .ZN(n6933) );
  NAND2_X1 U7627 ( .A1(n13488), .A2(n13672), .ZN(n6934) );
  NAND2_X1 U7628 ( .A1(n13672), .A2(n13520), .ZN(n6932) );
  INV_X1 U7629 ( .A(n11783), .ZN(n6992) );
  OAI21_X1 U7630 ( .B1(n6709), .B2(n13510), .A(n13509), .ZN(n6708) );
  NAND2_X1 U7631 ( .A1(n6882), .A2(n6881), .ZN(n11815) );
  NAND2_X1 U7632 ( .A1(n13525), .A2(n7543), .ZN(n7542) );
  NAND2_X1 U7633 ( .A1(n6685), .A2(n13527), .ZN(n6684) );
  INV_X1 U7634 ( .A(n13527), .ZN(n6686) );
  NAND2_X1 U7635 ( .A1(n7540), .A2(n7538), .ZN(n7537) );
  AND2_X1 U7636 ( .A1(n7541), .A2(n13540), .ZN(n7540) );
  INV_X1 U7637 ( .A(n11834), .ZN(n6994) );
  AND2_X1 U7638 ( .A1(n6873), .A2(n6585), .ZN(n6872) );
  INV_X1 U7639 ( .A(n7534), .ZN(n7533) );
  AOI21_X1 U7640 ( .B1(n13593), .B2(n13594), .A(n7535), .ZN(n7534) );
  INV_X1 U7641 ( .A(n13591), .ZN(n7535) );
  OR2_X1 U7642 ( .A1(n11871), .A2(n11872), .ZN(n11873) );
  AND2_X1 U7643 ( .A1(n11887), .A2(n7662), .ZN(n7658) );
  NAND2_X1 U7644 ( .A1(n11880), .A2(n11881), .ZN(n7662) );
  NAND2_X1 U7645 ( .A1(n7661), .A2(n7660), .ZN(n7659) );
  INV_X1 U7646 ( .A(n11884), .ZN(n7661) );
  NAND2_X1 U7647 ( .A1(n6942), .A2(n6941), .ZN(n13599) );
  NAND2_X1 U7648 ( .A1(n7553), .A2(n13602), .ZN(n7552) );
  INV_X1 U7649 ( .A(n13603), .ZN(n7553) );
  INV_X1 U7650 ( .A(n13605), .ZN(n6943) );
  INV_X1 U7651 ( .A(n13609), .ZN(n6969) );
  NAND2_X1 U7652 ( .A1(n13613), .A2(n6949), .ZN(n7549) );
  INV_X1 U7653 ( .A(n13612), .ZN(n6949) );
  AOI21_X1 U7654 ( .B1(n6869), .B2(n6868), .A(n6504), .ZN(n6867) );
  INV_X1 U7655 ( .A(n11897), .ZN(n6868) );
  NAND2_X1 U7656 ( .A1(n11899), .A2(n11898), .ZN(n6869) );
  NAND2_X1 U7657 ( .A1(n11901), .A2(n11900), .ZN(n6870) );
  NAND2_X1 U7658 ( .A1(n6675), .A2(n6674), .ZN(n13623) );
  AOI21_X1 U7659 ( .B1(n6676), .B2(n6679), .A(n6485), .ZN(n6674) );
  NAND2_X1 U7660 ( .A1(n13616), .A2(n6676), .ZN(n6675) );
  AND2_X1 U7661 ( .A1(n13617), .A2(n6680), .ZN(n6679) );
  INV_X1 U7662 ( .A(n11944), .ZN(n7628) );
  INV_X1 U7663 ( .A(n11943), .ZN(n7627) );
  AND2_X1 U7664 ( .A1(n7617), .A2(n6879), .ZN(n6878) );
  NAND2_X1 U7665 ( .A1(n11913), .A2(n6880), .ZN(n6879) );
  NAND2_X1 U7666 ( .A1(n7617), .A2(n7621), .ZN(n7615) );
  NOR2_X1 U7667 ( .A1(n7622), .A2(n6549), .ZN(n7621) );
  OR2_X1 U7668 ( .A1(n14614), .A2(n14225), .ZN(n6972) );
  INV_X1 U7669 ( .A(n6853), .ZN(n9717) );
  AOI21_X1 U7670 ( .B1(n9469), .B2(n6856), .A(n6854), .ZN(n6853) );
  NOR2_X1 U7671 ( .A1(n9625), .A2(n6857), .ZN(n6856) );
  OAI21_X1 U7672 ( .B1(n9625), .B2(n6855), .A(n9632), .ZN(n6854) );
  NOR2_X1 U7673 ( .A1(n8692), .A2(n7599), .ZN(n7598) );
  INV_X1 U7674 ( .A(n8686), .ZN(n7599) );
  NAND2_X1 U7675 ( .A1(n7271), .A2(n14235), .ZN(n14236) );
  NAND2_X1 U7676 ( .A1(n14291), .A2(n14292), .ZN(n7271) );
  INV_X1 U7677 ( .A(n10658), .ZN(n7429) );
  NAND2_X1 U7678 ( .A1(n9308), .A2(n9158), .ZN(n9160) );
  NAND2_X1 U7679 ( .A1(n12303), .A2(n12302), .ZN(n12304) );
  NOR2_X1 U7680 ( .A1(n12304), .A2(n12305), .ZN(n12323) );
  AOI21_X1 U7681 ( .B1(n7280), .B2(n7279), .A(n7067), .ZN(n12317) );
  INV_X1 U7682 ( .A(n12301), .ZN(n7067) );
  INV_X1 U7683 ( .A(n12294), .ZN(n7279) );
  INV_X1 U7684 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15255) );
  AOI21_X1 U7685 ( .B1(n12372), .B2(n12371), .A(n12370), .ZN(n12396) );
  OAI21_X1 U7686 ( .B1(n11074), .B2(n11076), .A(n11077), .ZN(n7171) );
  OR2_X1 U7687 ( .A1(n12653), .A2(n12480), .ZN(n11080) );
  NAND2_X1 U7688 ( .A1(n8226), .A2(n11027), .ZN(n7191) );
  NAND2_X1 U7689 ( .A1(n10077), .A2(n10075), .ZN(n7572) );
  NAND2_X1 U7690 ( .A1(n12230), .A2(n15132), .ZN(n10987) );
  OR2_X1 U7691 ( .A1(n12417), .A2(n12427), .ZN(n11125) );
  NAND2_X1 U7692 ( .A1(n15058), .A2(n7879), .ZN(n10398) );
  OR2_X1 U7693 ( .A1(n11100), .A2(SI_2_), .ZN(n7817) );
  NAND2_X1 U7694 ( .A1(n8249), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7134) );
  OR2_X1 U7695 ( .A1(n7774), .A2(n11664), .ZN(n7776) );
  INV_X1 U7696 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7714) );
  INV_X1 U7697 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7708) );
  INV_X1 U7698 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7707) );
  INV_X1 U7699 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7706) );
  INV_X1 U7700 ( .A(n7734), .ZN(n7338) );
  NOR2_X1 U7701 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n9145) );
  INV_X1 U7702 ( .A(n12774), .ZN(n7114) );
  NAND2_X1 U7703 ( .A1(n6752), .A2(n7108), .ZN(n11190) );
  NAND2_X1 U7704 ( .A1(n7500), .A2(n6548), .ZN(n7108) );
  NAND2_X1 U7705 ( .A1(n7104), .A2(n6558), .ZN(n6752) );
  INV_X1 U7706 ( .A(n13017), .ZN(n7513) );
  INV_X1 U7707 ( .A(n13007), .ZN(n6902) );
  INV_X1 U7708 ( .A(n13224), .ZN(n7454) );
  NOR2_X1 U7709 ( .A1(n9946), .A2(n11820), .ZN(n7152) );
  INV_X1 U7710 ( .A(n12006), .ZN(n7468) );
  NOR2_X1 U7711 ( .A1(n7482), .A2(n6897), .ZN(n6896) );
  OR2_X1 U7712 ( .A1(n12007), .A2(n7482), .ZN(n6898) );
  NAND2_X1 U7713 ( .A1(n9923), .A2(n9924), .ZN(n6895) );
  NAND2_X1 U7714 ( .A1(n8612), .A2(n7669), .ZN(n7668) );
  INV_X1 U7715 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8612) );
  NAND3_X1 U7716 ( .A1(n7013), .A2(n8413), .A3(n8412), .ZN(n6886) );
  AND3_X1 U7717 ( .A1(n8409), .A2(n8408), .A3(n8407), .ZN(n8412) );
  AND2_X1 U7718 ( .A1(n7136), .A2(n7135), .ZN(n8413) );
  NAND2_X1 U7719 ( .A1(n8404), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8421) );
  OR2_X1 U7720 ( .A1(n8617), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n8404) );
  OR2_X1 U7721 ( .A1(n8568), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U7722 ( .A1(n13454), .A2(n11351), .ZN(n7313) );
  NAND2_X1 U7723 ( .A1(n11267), .A2(n11266), .ZN(n7328) );
  NOR2_X1 U7724 ( .A1(n7220), .A2(n14561), .ZN(n7216) );
  NAND2_X1 U7725 ( .A1(n13683), .A2(n7219), .ZN(n7218) );
  INV_X1 U7726 ( .A(n10334), .ZN(n7219) );
  NOR2_X1 U7727 ( .A1(n14684), .A2(n14570), .ZN(n7204) );
  AND2_X1 U7728 ( .A1(n13676), .A2(n10093), .ZN(n7223) );
  INV_X1 U7729 ( .A(n9832), .ZN(n7225) );
  AND2_X1 U7730 ( .A1(n13674), .A2(n13673), .ZN(n7377) );
  INV_X1 U7731 ( .A(n9845), .ZN(n7378) );
  INV_X1 U7732 ( .A(n7227), .ZN(n7234) );
  AOI21_X1 U7733 ( .B1(n9045), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_28__SCAN_IN), .ZN(n7227) );
  INV_X1 U7734 ( .A(n14614), .ZN(n13489) );
  OAI21_X1 U7735 ( .B1(n11169), .B2(n11168), .A(n11172), .ZN(n11445) );
  OAI21_X1 U7736 ( .B1(n10532), .B2(n7600), .A(n10535), .ZN(n10745) );
  INV_X1 U7737 ( .A(n10533), .ZN(n7600) );
  INV_X1 U7738 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8438) );
  INV_X1 U7739 ( .A(n8752), .ZN(n8439) );
  AND2_X1 U7740 ( .A1(n7588), .A2(n9009), .ZN(n7587) );
  NAND2_X1 U7741 ( .A1(n9005), .A2(n7589), .ZN(n7588) );
  NAND2_X1 U7742 ( .A1(n6841), .A2(n8819), .ZN(n6840) );
  INV_X1 U7743 ( .A(n7596), .ZN(n7595) );
  OAI21_X1 U7744 ( .B1(n7598), .B2(n7597), .A(n7682), .ZN(n7596) );
  OR2_X1 U7745 ( .A1(n8787), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8788) );
  XNOR2_X1 U7746 ( .A(n8517), .B(SI_5_), .ZN(n8524) );
  XNOR2_X1 U7747 ( .A(n14236), .B(n7270), .ZN(n14281) );
  INV_X1 U7748 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7270) );
  OAI21_X1 U7749 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14249), .A(n14248), .ZN(
        n14312) );
  NAND2_X1 U7750 ( .A1(n12068), .A2(n12067), .ZN(n12066) );
  OR2_X1 U7751 ( .A1(n8058), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U7752 ( .A1(n12151), .A2(n12150), .ZN(n7419) );
  NAND2_X1 U7753 ( .A1(n8316), .A2(n7434), .ZN(n7433) );
  NAND2_X1 U7754 ( .A1(n12209), .A2(n8315), .ZN(n8316) );
  NAND2_X1 U7755 ( .A1(n11217), .A2(n8314), .ZN(n7434) );
  OR2_X1 U7756 ( .A1(n9894), .A2(n9895), .ZN(n7424) );
  OAI21_X1 U7757 ( .B1(n12151), .B2(n7418), .A(n6681), .ZN(n8334) );
  AOI21_X1 U7758 ( .B1(n7417), .B2(n6683), .A(n6682), .ZN(n6681) );
  INV_X1 U7759 ( .A(n8332), .ZN(n6682) );
  INV_X1 U7760 ( .A(n12150), .ZN(n6683) );
  INV_X1 U7761 ( .A(n12167), .ZN(n6699) );
  AND4_X1 U7762 ( .A1(n8063), .A2(n8062), .A3(n8061), .A4(n8060), .ZN(n8322)
         );
  NAND2_X1 U7763 ( .A1(n6814), .A2(n6813), .ZN(n14914) );
  OR2_X1 U7764 ( .A1(n6812), .A2(n6815), .ZN(n6814) );
  NAND2_X1 U7765 ( .A1(n6812), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6813) );
  INV_X1 U7766 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U7767 ( .A1(n9309), .A2(n9310), .ZN(n9308) );
  NAND2_X1 U7768 ( .A1(n9361), .A2(n9146), .ZN(n9314) );
  OAI21_X1 U7769 ( .B1(n9177), .B2(P3_REG2_REG_2__SCAN_IN), .A(n7085), .ZN(
        n9315) );
  NAND2_X1 U7770 ( .A1(n9314), .A2(n9315), .ZN(n9313) );
  NAND2_X1 U7771 ( .A1(n7031), .A2(n14924), .ZN(n7030) );
  INV_X1 U7772 ( .A(n9160), .ZN(n7031) );
  INV_X1 U7773 ( .A(n9148), .ZN(n9149) );
  NAND2_X1 U7774 ( .A1(n14921), .A2(n9179), .ZN(n9180) );
  NAND2_X1 U7775 ( .A1(n9180), .A2(n9181), .ZN(n9489) );
  AND2_X1 U7776 ( .A1(n7033), .A2(n7032), .ZN(n9497) );
  INV_X1 U7777 ( .A(n9162), .ZN(n7032) );
  OR2_X1 U7778 ( .A1(n9503), .A2(n9502), .ZN(n9882) );
  NAND2_X1 U7779 ( .A1(n14936), .A2(n9491), .ZN(n9492) );
  NAND2_X1 U7780 ( .A1(n9492), .A2(n9493), .ZN(n9874) );
  NAND2_X1 U7781 ( .A1(n14952), .A2(n9876), .ZN(n9877) );
  NAND2_X1 U7782 ( .A1(n9877), .A2(n9878), .ZN(n10225) );
  NAND2_X1 U7783 ( .A1(n7057), .A2(n6515), .ZN(n7156) );
  AND2_X1 U7784 ( .A1(n10236), .A2(n10235), .ZN(n10570) );
  NAND2_X1 U7785 ( .A1(n7156), .A2(n7155), .ZN(n14979) );
  INV_X1 U7786 ( .A(n14975), .ZN(n7155) );
  OR2_X1 U7787 ( .A1(n14970), .A2(n14969), .ZN(n14967) );
  NOR2_X1 U7788 ( .A1(n12257), .A2(n6817), .ZN(n6816) );
  INV_X1 U7789 ( .A(n12255), .ZN(n6817) );
  OR2_X1 U7790 ( .A1(n12268), .A2(n12269), .ZN(n7162) );
  NAND2_X1 U7791 ( .A1(n12306), .A2(n6809), .ZN(n6808) );
  INV_X1 U7792 ( .A(n12308), .ZN(n6809) );
  XNOR2_X1 U7793 ( .A(n12317), .B(n12331), .ZN(n12296) );
  NAND2_X1 U7794 ( .A1(n7028), .A2(n6526), .ZN(n7154) );
  NAND2_X1 U7795 ( .A1(n7154), .A2(n7153), .ZN(n12344) );
  INV_X1 U7796 ( .A(n12335), .ZN(n7153) );
  NAND2_X1 U7797 ( .A1(n6808), .A2(n6807), .ZN(n6806) );
  INV_X1 U7798 ( .A(n12323), .ZN(n6807) );
  NAND2_X1 U7799 ( .A1(n6805), .A2(n12355), .ZN(n12358) );
  NAND2_X1 U7800 ( .A1(n6806), .A2(n6640), .ZN(n6805) );
  AND2_X1 U7801 ( .A1(n12344), .A2(n12343), .ZN(n12376) );
  NAND2_X1 U7802 ( .A1(n6656), .A2(n11075), .ZN(n12452) );
  NAND2_X1 U7803 ( .A1(n12464), .A2(n11074), .ZN(n6656) );
  NAND2_X1 U7804 ( .A1(n7698), .A2(n15209), .ZN(n8164) );
  OR2_X1 U7805 ( .A1(n8122), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U7806 ( .A1(n6651), .A2(n11069), .ZN(n12500) );
  AND3_X1 U7807 ( .A1(n8089), .A2(n8088), .A3(n8087), .ZN(n12522) );
  NAND2_X1 U7808 ( .A1(n12677), .A2(n12571), .ZN(n7009) );
  AND2_X1 U7809 ( .A1(n8227), .A2(n6643), .ZN(n6642) );
  NAND2_X1 U7810 ( .A1(n12587), .A2(n11031), .ZN(n6643) );
  AND2_X1 U7811 ( .A1(n11034), .A2(n11024), .ZN(n12611) );
  AND4_X1 U7812 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8013), .ZN(n12620)
         );
  NAND2_X1 U7813 ( .A1(n7565), .A2(n7564), .ZN(n12622) );
  NAND2_X1 U7814 ( .A1(n10750), .A2(n11140), .ZN(n6825) );
  AND4_X1 U7815 ( .A1(n7988), .A2(n7987), .A3(n7986), .A4(n7985), .ZN(n12619)
         );
  INV_X1 U7816 ( .A(n6646), .ZN(n6645) );
  OAI21_X1 U7817 ( .B1(n7172), .B2(n6647), .A(n10955), .ZN(n6646) );
  INV_X1 U7818 ( .A(n11137), .ZN(n6647) );
  AOI21_X1 U7819 ( .B1(n7176), .B2(n7178), .A(n7173), .ZN(n7172) );
  INV_X1 U7820 ( .A(n11012), .ZN(n7173) );
  AND2_X1 U7821 ( .A1(n10955), .A2(n11014), .ZN(n11137) );
  NAND2_X1 U7822 ( .A1(n8297), .A2(n15152), .ZN(n7179) );
  NAND2_X1 U7823 ( .A1(n15024), .A2(n15048), .ZN(n7180) );
  INV_X1 U7824 ( .A(n8224), .ZN(n11128) );
  INV_X1 U7825 ( .A(n10995), .ZN(n7184) );
  NAND2_X1 U7826 ( .A1(n10214), .A2(n6834), .ZN(n15058) );
  AND2_X1 U7827 ( .A1(n11134), .A2(n7867), .ZN(n6834) );
  AND2_X1 U7828 ( .A1(n10988), .A2(n10987), .ZN(n11130) );
  NAND2_X1 U7829 ( .A1(n10208), .A2(n11130), .ZN(n10210) );
  INV_X1 U7830 ( .A(n15093), .ZN(n15072) );
  NAND2_X1 U7831 ( .A1(n9140), .A2(n7167), .ZN(n7795) );
  OR2_X1 U7832 ( .A1(n11100), .A2(n8460), .ZN(n7796) );
  NOR2_X1 U7833 ( .A1(n11332), .A2(n8459), .ZN(n7167) );
  NAND2_X1 U7834 ( .A1(n8363), .A2(n11093), .ZN(n15096) );
  NOR2_X2 U7835 ( .A1(n15094), .A2(n12707), .ZN(n15088) );
  AND2_X1 U7836 ( .A1(n11125), .A2(n11123), .ZN(n11147) );
  OAI21_X1 U7837 ( .B1(n8191), .B2(n8190), .A(n8192), .ZN(n11099) );
  INV_X1 U7838 ( .A(n8249), .ZN(n6695) );
  NOR2_X1 U7839 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6694) );
  NAND2_X1 U7840 ( .A1(n6770), .A2(n11374), .ZN(n8134) );
  INV_X1 U7841 ( .A(n8132), .ZN(n6770) );
  OAI21_X1 U7842 ( .B1(n7350), .B2(n6768), .A(n6766), .ZN(n8106) );
  INV_X1 U7843 ( .A(n6767), .ZN(n6766) );
  OAI21_X1 U7844 ( .B1(n7353), .B2(n6768), .A(n7772), .ZN(n6767) );
  INV_X1 U7845 ( .A(n8092), .ZN(n6768) );
  NAND2_X1 U7846 ( .A1(n7352), .A2(n11519), .ZN(n7351) );
  NAND2_X1 U7847 ( .A1(n7770), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7353) );
  INV_X1 U7848 ( .A(n7350), .ZN(n7349) );
  AND2_X1 U7849 ( .A1(n7767), .A2(n7766), .ZN(n8051) );
  AOI21_X1 U7850 ( .B1(n8035), .B2(n7344), .A(n7343), .ZN(n7342) );
  INV_X1 U7851 ( .A(n7765), .ZN(n7343) );
  INV_X1 U7852 ( .A(n7763), .ZN(n7344) );
  INV_X1 U7853 ( .A(n8035), .ZN(n7345) );
  AND2_X1 U7854 ( .A1(n7763), .A2(n7762), .ZN(n8017) );
  NAND2_X1 U7855 ( .A1(n7360), .A2(n7359), .ZN(n7358) );
  INV_X1 U7856 ( .A(n7992), .ZN(n7360) );
  INV_X1 U7857 ( .A(n7759), .ZN(n7357) );
  OAI21_X1 U7858 ( .B1(n7935), .B2(n6757), .A(n6755), .ZN(n7961) );
  INV_X1 U7859 ( .A(n7751), .ZN(n6757) );
  AOI21_X1 U7860 ( .B1(n6756), .B2(n7751), .A(n6621), .ZN(n6755) );
  AND2_X1 U7861 ( .A1(n7750), .A2(n7749), .ZN(n7932) );
  OAI21_X1 U7862 ( .B1(n7887), .B2(n7743), .A(n7744), .ZN(n7907) );
  AND2_X1 U7863 ( .A1(n7734), .A2(n7733), .ZN(n7824) );
  NAND2_X1 U7864 ( .A1(n6776), .A2(n7732), .ZN(n7825) );
  AOI21_X1 U7865 ( .B1(n7484), .B2(n7117), .A(n7116), .ZN(n7115) );
  INV_X1 U7866 ( .A(n11706), .ZN(n7116) );
  INV_X1 U7867 ( .A(n12797), .ZN(n7117) );
  AND2_X1 U7868 ( .A1(n7485), .A2(n7114), .ZN(n7113) );
  INV_X1 U7869 ( .A(n12838), .ZN(n7483) );
  NAND2_X1 U7870 ( .A1(n11660), .A2(n11580), .ZN(n7090) );
  NAND2_X1 U7871 ( .A1(n11574), .A2(n11573), .ZN(n7092) );
  AND2_X1 U7872 ( .A1(n7471), .A2(n9329), .ZN(n9560) );
  NAND4_X1 U7873 ( .A1(n6751), .A2(n6750), .A3(n6568), .A4(n9707), .ZN(n9708)
         );
  NAND2_X1 U7874 ( .A1(n7120), .A2(n7506), .ZN(n7503) );
  NAND2_X1 U7875 ( .A1(n10319), .A2(n10309), .ZN(n7120) );
  NAND2_X1 U7876 ( .A1(n10321), .A2(n10319), .ZN(n7504) );
  AND2_X1 U7877 ( .A1(n7504), .A2(n7502), .ZN(n10594) );
  OR2_X1 U7878 ( .A1(n11500), .A2(n11499), .ZN(n11501) );
  XNOR2_X1 U7879 ( .A(n11190), .B(n11189), .ZN(n11650) );
  AND4_X1 U7880 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n12799) );
  NOR2_X1 U7882 ( .A1(n11743), .A2(n8957), .ZN(n6929) );
  NAND3_X1 U7883 ( .A1(n8926), .A2(n8927), .A3(n8925), .ZN(n11768) );
  OR2_X1 U7884 ( .A1(n8956), .A2(n8924), .ZN(n8925) );
  NOR2_X1 U7885 ( .A1(n6935), .A2(n7020), .ZN(n8927) );
  AND2_X1 U7886 ( .A1(n6827), .A2(n6826), .ZN(n9251) );
  NAND2_X1 U7887 ( .A1(n10172), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U7888 ( .A1(n14738), .A2(n12936), .ZN(n12937) );
  NAND2_X1 U7889 ( .A1(n14792), .A2(n12945), .ZN(n12967) );
  AND2_X1 U7890 ( .A1(n7507), .A2(n13251), .ZN(n6981) );
  INV_X1 U7891 ( .A(n7508), .ZN(n7507) );
  OAI21_X1 U7892 ( .B1(n7514), .B2(n7512), .A(n7509), .ZN(n7508) );
  NAND2_X1 U7893 ( .A1(n13044), .A2(n7513), .ZN(n7509) );
  AND2_X1 U7894 ( .A1(n7514), .A2(n13044), .ZN(n7511) );
  OR2_X1 U7895 ( .A1(n13044), .A2(n7513), .ZN(n7512) );
  NOR2_X1 U7896 ( .A1(n13271), .A2(n13276), .ZN(n6795) );
  NAND2_X1 U7897 ( .A1(n6790), .A2(n6926), .ZN(n13055) );
  NAND2_X1 U7898 ( .A1(n13271), .A2(n12880), .ZN(n6926) );
  XNOR2_X1 U7899 ( .A(n13271), .B(n13042), .ZN(n13077) );
  OR2_X1 U7900 ( .A1(n13037), .A2(n13036), .ZN(n7677) );
  AND2_X1 U7901 ( .A1(n13008), .A2(n7677), .ZN(n7465) );
  OR2_X1 U7902 ( .A1(n13114), .A2(n13115), .ZN(n13116) );
  NAND2_X1 U7903 ( .A1(n13134), .A2(n13133), .ZN(n13132) );
  OR2_X1 U7904 ( .A1(n7447), .A2(n7444), .ZN(n7443) );
  INV_X1 U7905 ( .A(n7451), .ZN(n7444) );
  NAND2_X1 U7906 ( .A1(n7450), .A2(n7445), .ZN(n7440) );
  OAI21_X1 U7907 ( .B1(n7450), .B2(n7442), .A(n7441), .ZN(n13128) );
  INV_X1 U7908 ( .A(n7443), .ZN(n7442) );
  AOI21_X1 U7909 ( .B1(n7443), .B2(n7446), .A(n13133), .ZN(n7441) );
  AOI21_X1 U7910 ( .B1(n13164), .B2(n13033), .A(n13005), .ZN(n13146) );
  NAND2_X1 U7911 ( .A1(n13173), .A2(n12848), .ZN(n7452) );
  NOR2_X1 U7912 ( .A1(n13150), .A2(n7448), .ZN(n7447) );
  INV_X1 U7913 ( .A(n7452), .ZN(n7448) );
  AOI21_X1 U7914 ( .B1(n7479), .B2(n7478), .A(n6502), .ZN(n7477) );
  INV_X1 U7915 ( .A(n13001), .ZN(n7478) );
  NAND2_X1 U7916 ( .A1(n6786), .A2(n13028), .ZN(n13177) );
  INV_X1 U7917 ( .A(n7674), .ZN(n7456) );
  NAND2_X1 U7918 ( .A1(n7498), .A2(n12882), .ZN(n7497) );
  OR2_X1 U7919 ( .A1(n13223), .A2(n13224), .ZN(n6905) );
  NAND2_X1 U7920 ( .A1(n13024), .A2(n7673), .ZN(n13221) );
  NAND2_X1 U7921 ( .A1(n13221), .A2(n13224), .ZN(n13220) );
  NAND2_X1 U7922 ( .A1(n10837), .A2(n7680), .ZN(n10839) );
  NAND2_X1 U7923 ( .A1(n10481), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10887) );
  NAND2_X1 U7924 ( .A1(n6783), .A2(n6782), .ZN(n10876) );
  OR2_X1 U7925 ( .A1(n11866), .A2(n12884), .ZN(n6782) );
  NAND2_X1 U7926 ( .A1(n6779), .A2(n6539), .ZN(n6783) );
  OR2_X1 U7927 ( .A1(n10194), .A2(n10193), .ZN(n10469) );
  OR2_X1 U7928 ( .A1(n10523), .A2(n11853), .ZN(n7681) );
  NAND2_X1 U7929 ( .A1(n7522), .A2(n6489), .ZN(n7521) );
  INV_X1 U7930 ( .A(n12014), .ZN(n7522) );
  AND2_X1 U7931 ( .A1(n11837), .A2(n11839), .ZN(n6927) );
  AOI21_X1 U7932 ( .B1(n10049), .B2(n10048), .A(n6524), .ZN(n10280) );
  NAND2_X1 U7933 ( .A1(n7460), .A2(n6545), .ZN(n9937) );
  NAND2_X1 U7934 ( .A1(n9805), .A2(n9804), .ZN(n9919) );
  NAND2_X1 U7935 ( .A1(n9924), .A2(n9806), .ZN(n12005) );
  XNOR2_X1 U7936 ( .A(n14829), .B(n12894), .ZN(n12006) );
  AND2_X1 U7937 ( .A1(n9423), .A2(n9414), .ZN(n10032) );
  MUX2_X1 U7938 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13369), .S(n8968), .Z(n13244)
         );
  INV_X1 U7939 ( .A(n13332), .ZN(n13243) );
  AOI21_X1 U7940 ( .B1(n6892), .B2(n6891), .A(n13058), .ZN(n13268) );
  NAND2_X1 U7941 ( .A1(n13057), .A2(n13056), .ZN(n6891) );
  NAND2_X1 U7942 ( .A1(n11495), .A2(n6486), .ZN(n11497) );
  NAND2_X1 U7943 ( .A1(n10696), .A2(n11951), .ZN(n10461) );
  NAND2_X1 U7944 ( .A1(n10547), .A2(n11951), .ZN(n10180) );
  INV_X1 U7945 ( .A(n11837), .ZN(n14868) );
  NAND2_X1 U7946 ( .A1(n9574), .A2(n6486), .ZN(n8946) );
  AOI21_X1 U7947 ( .B1(n11507), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n6532), .ZN(
        n7146) );
  NOR2_X1 U7948 ( .A1(n7668), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7667) );
  INV_X1 U7949 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8900) );
  NOR2_X1 U7950 ( .A1(n7669), .A2(n7012), .ZN(n7011) );
  INV_X1 U7951 ( .A(n7141), .ZN(n8616) );
  XNOR2_X1 U7952 ( .A(n8416), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8887) );
  INV_X1 U7953 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U7954 ( .A1(n7139), .A2(n6483), .ZN(n8894) );
  NAND2_X1 U7955 ( .A1(n8414), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9021) );
  NOR2_X1 U7956 ( .A1(n8587), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8675) );
  INV_X1 U7957 ( .A(n8782), .ZN(n8554) );
  AND2_X1 U7958 ( .A1(n9083), .A2(n9082), .ZN(n9087) );
  XNOR2_X1 U7959 ( .A(n7289), .B(n11410), .ZN(n9088) );
  NAND2_X1 U7960 ( .A1(n9084), .A2(n6667), .ZN(n7289) );
  NAND2_X1 U7961 ( .A1(n6668), .A2(n9068), .ZN(n6667) );
  AOI21_X1 U7962 ( .B1(n13438), .B2(n13437), .A(n6665), .ZN(n13407) );
  AND2_X1 U7963 ( .A1(n11314), .A2(n11315), .ZN(n6665) );
  NAND2_X1 U7964 ( .A1(n14379), .A2(n7672), .ZN(n11255) );
  NOR2_X1 U7965 ( .A1(n10934), .A2(n10933), .ZN(n11272) );
  NAND2_X1 U7966 ( .A1(n7315), .A2(n7304), .ZN(n7303) );
  INV_X1 U7967 ( .A(n7310), .ZN(n7304) );
  AOI21_X1 U7968 ( .B1(n6487), .B2(n7312), .A(n7311), .ZN(n7310) );
  INV_X1 U7969 ( .A(n7314), .ZN(n7312) );
  NAND2_X1 U7970 ( .A1(n13389), .A2(n9584), .ZN(n9786) );
  NAND2_X1 U7971 ( .A1(n10507), .A2(n10506), .ZN(n10641) );
  AND2_X1 U7972 ( .A1(n9067), .A2(n9066), .ZN(n9187) );
  INV_X1 U7973 ( .A(n7335), .ZN(n7334) );
  AOI21_X1 U7974 ( .B1(n10920), .B2(n7334), .A(n13449), .ZN(n7333) );
  NAND2_X1 U7975 ( .A1(n7318), .A2(n7322), .ZN(n13467) );
  AND2_X1 U7976 ( .A1(n13469), .A2(n7323), .ZN(n7322) );
  OR2_X1 U7977 ( .A1(n6490), .A2(n7327), .ZN(n7323) );
  NAND2_X1 U7978 ( .A1(n9783), .A2(n9782), .ZN(n9788) );
  XNOR2_X1 U7979 ( .A(n11255), .B(n11256), .ZN(n14422) );
  AND2_X1 U7980 ( .A1(n13706), .A2(n13666), .ZN(n6967) );
  OAI21_X1 U7981 ( .B1(n13649), .B2(n6704), .A(n6703), .ZN(n6951) );
  NAND2_X1 U7982 ( .A1(n13652), .A2(n13651), .ZN(n6703) );
  NOR2_X1 U7983 ( .A1(n13652), .A2(n13651), .ZN(n6704) );
  AOI22_X1 U7984 ( .A1(n13634), .A2(n13633), .B1(n6931), .B2(n13632), .ZN(
        n13649) );
  INV_X1 U7985 ( .A(n7199), .ZN(n13831) );
  INV_X1 U7986 ( .A(n13695), .ZN(n13843) );
  AND3_X1 U7987 ( .A1(n11606), .A2(n11607), .A3(n6516), .ZN(n7262) );
  NAND2_X1 U7988 ( .A1(n11606), .A2(n11607), .ZN(n13877) );
  OR2_X1 U7989 ( .A1(n13893), .A2(n13897), .ZN(n7263) );
  AND2_X1 U7990 ( .A1(n13913), .A2(n11623), .ZN(n13898) );
  INV_X1 U7991 ( .A(n7237), .ZN(n7236) );
  OAI21_X1 U7992 ( .B1(n7239), .B2(n7241), .A(n13930), .ZN(n7237) );
  NAND2_X1 U7993 ( .A1(n13966), .A2(n7241), .ZN(n7235) );
  AND2_X1 U7994 ( .A1(n7389), .A2(n11620), .ZN(n7388) );
  INV_X1 U7995 ( .A(n13953), .ZN(n13944) );
  NAND2_X1 U7996 ( .A1(n7243), .A2(n11619), .ZN(n13964) );
  INV_X1 U7997 ( .A(n13966), .ZN(n7243) );
  AOI21_X1 U7998 ( .B1(n7251), .B2(n11600), .A(n7249), .ZN(n7248) );
  INV_X1 U7999 ( .A(n13586), .ZN(n7249) );
  AOI21_X1 U8000 ( .B1(n7401), .B2(n7398), .A(n7397), .ZN(n7396) );
  OR2_X1 U8001 ( .A1(n11614), .A2(n7399), .ZN(n7394) );
  NOR2_X1 U8002 ( .A1(n7206), .A2(n14123), .ZN(n7397) );
  AND2_X1 U8003 ( .A1(n13562), .A2(n13686), .ZN(n7402) );
  OR2_X1 U8004 ( .A1(n11614), .A2(n13688), .ZN(n7403) );
  AOI21_X1 U8005 ( .B1(n7257), .B2(n13685), .A(n6537), .ZN(n7255) );
  INV_X1 U8006 ( .A(n7257), .ZN(n7256) );
  NAND2_X1 U8007 ( .A1(n10701), .A2(n13685), .ZN(n10773) );
  NAND2_X1 U8008 ( .A1(n10760), .A2(n10759), .ZN(n10762) );
  OR2_X1 U8009 ( .A1(n10622), .A2(n10621), .ZN(n10624) );
  NOR2_X1 U8010 ( .A1(n10605), .A2(n7407), .ZN(n7406) );
  INV_X1 U8011 ( .A(n10550), .ZN(n7407) );
  NAND2_X1 U8012 ( .A1(n7405), .A2(n7404), .ZN(n10771) );
  NOR2_X1 U8013 ( .A1(n13684), .A2(n7686), .ZN(n7404) );
  NAND2_X1 U8014 ( .A1(n10338), .A2(n10337), .ZN(n14702) );
  AND2_X1 U8015 ( .A1(n14559), .A2(n10350), .ZN(n10351) );
  NAND2_X1 U8016 ( .A1(n10351), .A2(n7220), .ZN(n10551) );
  NAND2_X1 U8017 ( .A1(n10328), .A2(n10327), .ZN(n14562) );
  AND2_X1 U8018 ( .A1(n6529), .A2(n13679), .ZN(n7411) );
  OR2_X1 U8019 ( .A1(n9997), .A2(n9996), .ZN(n9999) );
  NAND2_X1 U8020 ( .A1(n9831), .A2(n9830), .ZN(n10087) );
  INV_X1 U8021 ( .A(n13674), .ZN(n10093) );
  AND2_X1 U8022 ( .A1(n14633), .A2(n13656), .ZN(n14604) );
  NAND2_X1 U8023 ( .A1(n11376), .A2(n11375), .ZN(n13903) );
  NAND2_X1 U8024 ( .A1(n11318), .A2(n11317), .ZN(n13950) );
  AND2_X1 U8025 ( .A1(n11233), .A2(n11232), .ZN(n14124) );
  NAND2_X1 U8026 ( .A1(n10929), .A2(n10928), .ZN(n14145) );
  AND2_X1 U8027 ( .A1(n9127), .A2(n11594), .ZN(n14635) );
  NOR2_X1 U8028 ( .A1(n14225), .A2(n13645), .ZN(n14633) );
  NAND2_X1 U8029 ( .A1(n9099), .A2(n9098), .ZN(n10946) );
  XNOR2_X1 U8030 ( .A(n11922), .B(n11181), .ZN(n13635) );
  NAND2_X1 U8031 ( .A1(n9045), .A2(n7233), .ZN(n7232) );
  NOR2_X1 U8032 ( .A1(n8756), .A2(n6937), .ZN(n7233) );
  INV_X1 U8033 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8755) );
  INV_X1 U8034 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8430) );
  INV_X1 U8035 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U8036 ( .A1(n8432), .A2(n6973), .ZN(n8435) );
  INV_X1 U8037 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U8038 ( .A1(n8439), .A2(n7336), .ZN(n8447) );
  AND2_X1 U8039 ( .A1(n7337), .A2(n8438), .ZN(n7336) );
  AND2_X1 U8040 ( .A1(n8440), .A2(n6939), .ZN(n7337) );
  INV_X1 U8041 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8440) );
  INV_X1 U8042 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9042) );
  NOR2_X1 U8043 ( .A1(n8433), .A2(n6937), .ZN(n6702) );
  XNOR2_X1 U8044 ( .A(n9524), .B(n9523), .ZN(n11505) );
  NOR2_X1 U8045 ( .A1(n9197), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U8046 ( .A1(n9470), .A2(n9072), .ZN(n9473) );
  NAND2_X1 U8047 ( .A1(n6849), .A2(n8598), .ZN(n8672) );
  NAND2_X1 U8048 ( .A1(n8596), .A2(n8595), .ZN(n6849) );
  NAND2_X1 U8049 ( .A1(n7594), .A2(n8538), .ZN(n8581) );
  NAND2_X1 U8050 ( .A1(n8537), .A2(n8536), .ZN(n7594) );
  AOI21_X1 U8051 ( .B1(n14336), .B2(n14290), .A(n14333), .ZN(n14294) );
  NAND2_X1 U8052 ( .A1(n14241), .A2(n14240), .ZN(n14304) );
  AOI21_X1 U8053 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14253), .A(n14252), .ZN(
        n14276) );
  OAI21_X1 U8054 ( .B1(n14469), .B2(n7066), .A(n6735), .ZN(n14318) );
  OR2_X1 U8055 ( .A1(n14470), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6735) );
  AND2_X1 U8056 ( .A1(n14470), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7066) );
  OAI22_X1 U8057 ( .A1(n14321), .A2(n14259), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n14258), .ZN(n14273) );
  AND2_X1 U8058 ( .A1(n7266), .A2(n14485), .ZN(n14328) );
  AND2_X1 U8059 ( .A1(n14489), .A2(n14491), .ZN(n14330) );
  AND3_X1 U8060 ( .A1(n7893), .A2(n7892), .A3(n7891), .ZN(n12069) );
  NAND2_X1 U8061 ( .A1(n8121), .A2(n8120), .ZN(n12501) );
  OR2_X1 U8062 ( .A1(n11100), .A2(SI_3_), .ZN(n7832) );
  NAND2_X1 U8063 ( .A1(n7788), .A2(n7787), .ZN(n12061) );
  NAND2_X1 U8064 ( .A1(n8281), .A2(n8279), .ZN(n9403) );
  NAND2_X1 U8065 ( .A1(n12051), .A2(n7017), .ZN(n8279) );
  NOR2_X1 U8066 ( .A1(n7018), .A2(n7430), .ZN(n7017) );
  NAND2_X1 U8067 ( .A1(n8098), .A2(n8097), .ZN(n12526) );
  OR2_X1 U8068 ( .A1(n7010), .A2(n15361), .ZN(n8097) );
  OR2_X1 U8069 ( .A1(n9633), .A2(n8096), .ZN(n8098) );
  INV_X1 U8070 ( .A(n12223), .ZN(n12472) );
  AND3_X1 U8071 ( .A1(n7848), .A2(n7847), .A3(n7846), .ZN(n10083) );
  NAND2_X1 U8072 ( .A1(n8084), .A2(n8083), .ZN(n12536) );
  NAND2_X1 U8073 ( .A1(n8359), .A2(n8358), .ZN(n12203) );
  INV_X1 U8074 ( .A(n12522), .ZN(n12548) );
  AND2_X1 U8075 ( .A1(n14983), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7160) );
  NOR2_X1 U8076 ( .A1(n9144), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14909) );
  XNOR2_X1 U8077 ( .A(n9175), .B(n9365), .ZN(n9353) );
  NOR2_X1 U8078 ( .A1(n14914), .A2(n14915), .ZN(n14912) );
  INV_X1 U8079 ( .A(n7158), .ZN(n9886) );
  AND2_X1 U8080 ( .A1(n7077), .A2(n7080), .ZN(n12236) );
  NAND2_X1 U8081 ( .A1(n6505), .A2(n7079), .ZN(n7078) );
  OAI211_X1 U8082 ( .C1(n14999), .C2(n7073), .A(n7072), .B(n7070), .ZN(n12240)
         );
  NAND2_X1 U8083 ( .A1(n7074), .A2(n12280), .ZN(n7073) );
  AOI21_X1 U8084 ( .B1(n6627), .B2(n14998), .A(n7071), .ZN(n7070) );
  NAND2_X1 U8085 ( .A1(n14999), .A2(n6627), .ZN(n7072) );
  NOR2_X1 U8086 ( .A1(n12240), .A2(n14360), .ZN(n12274) );
  OR2_X1 U8087 ( .A1(n12345), .A2(n12346), .ZN(n7034) );
  XNOR2_X1 U8088 ( .A(n12376), .B(n7035), .ZN(n12345) );
  INV_X1 U8089 ( .A(n7084), .ZN(n12363) );
  NAND2_X1 U8090 ( .A1(n7165), .A2(n6821), .ZN(n6820) );
  AOI21_X1 U8091 ( .B1(n14983), .B2(n12395), .A(n12375), .ZN(n6821) );
  OAI21_X1 U8092 ( .B1(n12384), .B2(n7166), .A(n15005), .ZN(n7165) );
  AOI21_X1 U8093 ( .B1(n6987), .B2(n6986), .A(n14911), .ZN(n6819) );
  NAND2_X1 U8094 ( .A1(n12373), .A2(n12374), .ZN(n6986) );
  INV_X1 U8095 ( .A(n12394), .ZN(n6987) );
  NAND2_X1 U8096 ( .A1(n12426), .A2(n7024), .ZN(n12641) );
  NOR2_X1 U8097 ( .A1(n7025), .A2(n6615), .ZN(n7024) );
  NAND2_X1 U8098 ( .A1(n8057), .A2(n8056), .ZN(n12681) );
  NAND2_X1 U8099 ( .A1(n8042), .A2(n8041), .ZN(n12689) );
  NAND2_X1 U8100 ( .A1(n9699), .A2(n15053), .ZN(n15107) );
  NAND2_X1 U8101 ( .A1(n11110), .A2(n11109), .ZN(n12633) );
  NAND2_X1 U8102 ( .A1(n12765), .A2(n11108), .ZN(n11110) );
  OR2_X1 U8103 ( .A1(n7010), .A2(n15347), .ZN(n8177) );
  OR2_X1 U8104 ( .A1(n10375), .A2(n8136), .ZN(n12725) );
  NAND2_X1 U8105 ( .A1(n8010), .A2(n8009), .ZN(n12752) );
  INV_X1 U8106 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n6689) );
  NOR2_X1 U8107 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), .ZN(
        n6832) );
  NAND2_X1 U8108 ( .A1(n7905), .A2(n7904), .ZN(n10234) );
  NAND2_X1 U8109 ( .A1(n11590), .A2(n11580), .ZN(n11662) );
  XNOR2_X1 U8110 ( .A(n7092), .B(n11660), .ZN(n11590) );
  AND4_X1 U8111 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n13006) );
  NAND2_X1 U8112 ( .A1(n10171), .A2(n10170), .ZN(n10266) );
  NAND2_X1 U8113 ( .A1(n11724), .A2(n11723), .ZN(n13267) );
  NAND2_X1 U8114 ( .A1(n9222), .A2(n8970), .ZN(n9373) );
  AND2_X1 U8115 ( .A1(n9223), .A2(n8969), .ZN(n8970) );
  XNOR2_X1 U8116 ( .A(n10458), .B(n10456), .ZN(n10319) );
  NAND2_X1 U8117 ( .A1(n10607), .A2(n11951), .ZN(n7118) );
  NAND2_X1 U8118 ( .A1(n7086), .A2(n11209), .ZN(n11502) );
  NAND2_X1 U8119 ( .A1(n11268), .A2(n6486), .ZN(n11196) );
  NAND2_X1 U8120 ( .A1(n11521), .A2(n11520), .ZN(n13309) );
  AND2_X1 U8121 ( .A1(n8960), .A2(n8959), .ZN(n13020) );
  OAI21_X1 U8122 ( .B1(n11995), .B2(n12000), .A(n11999), .ZN(n12037) );
  NAND4_X1 U8123 ( .A1(n9552), .A2(n9551), .A3(n9550), .A4(n9549), .ZN(n12892)
         );
  NAND2_X1 U8124 ( .A1(n6498), .A2(n8910), .ZN(n12898) );
  OR2_X1 U8125 ( .A1(n8956), .A2(n8903), .ZN(n8909) );
  NAND2_X1 U8126 ( .A1(n14765), .A2(n12941), .ZN(n14776) );
  NAND2_X1 U8127 ( .A1(n14776), .A2(n14775), .ZN(n14774) );
  XNOR2_X1 U8128 ( .A(n13055), .B(n13056), .ZN(n13269) );
  INV_X1 U8129 ( .A(n13246), .ZN(n13239) );
  NAND2_X1 U8130 ( .A1(n6798), .A2(n8968), .ZN(n6797) );
  OAI21_X1 U8131 ( .B1(n9079), .B2(n8945), .A(n6576), .ZN(n6798) );
  OAI211_X1 U8132 ( .C1(n13269), .C2(n13337), .A(n13268), .B(n6803), .ZN(
        n13341) );
  NOR2_X1 U8133 ( .A1(n13266), .A2(n6804), .ZN(n6803) );
  AND2_X1 U8134 ( .A1(n13267), .A2(n14879), .ZN(n6804) );
  NAND2_X1 U8135 ( .A1(n13467), .A2(n6666), .ZN(n13398) );
  AND2_X1 U8136 ( .A1(n13399), .A2(n13397), .ZN(n6666) );
  NAND2_X1 U8137 ( .A1(n11468), .A2(n11467), .ZN(n13830) );
  NAND2_X1 U8138 ( .A1(n11260), .A2(n11259), .ZN(n14390) );
  NAND2_X1 U8139 ( .A1(n11258), .A2(n6468), .ZN(n11260) );
  NAND2_X1 U8140 ( .A1(n14422), .A2(n14421), .ZN(n14420) );
  XNOR2_X1 U8141 ( .A(n9786), .B(n9784), .ZN(n9783) );
  INV_X1 U8142 ( .A(n14196), .ZN(n13973) );
  NAND2_X1 U8143 ( .A1(n10700), .A2(n10699), .ZN(n13550) );
  INV_X1 U8144 ( .A(n13724), .ZN(n14404) );
  INV_X1 U8145 ( .A(n14410), .ZN(n14431) );
  INV_X1 U8146 ( .A(n13592), .ZN(n13719) );
  NAND2_X1 U8147 ( .A1(n13655), .A2(n13654), .ZN(n14040) );
  AND2_X1 U8148 ( .A1(n13829), .A2(n13828), .ZN(n14061) );
  INV_X1 U8149 ( .A(n14201), .ZN(n14001) );
  NOR2_X1 U8150 ( .A1(n6538), .A2(n9081), .ZN(n6669) );
  NAND2_X1 U8151 ( .A1(n10947), .A2(n9116), .ZN(n14599) );
  INV_X1 U8152 ( .A(n10143), .ZN(n9116) );
  INV_X1 U8153 ( .A(n13830), .ZN(n14168) );
  INV_X1 U8154 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14287) );
  XNOR2_X1 U8155 ( .A(n14288), .B(n6738), .ZN(n15389) );
  INV_X1 U8156 ( .A(n14297), .ZN(n6730) );
  NAND2_X1 U8157 ( .A1(n6722), .A2(n14311), .ZN(n6726) );
  NAND2_X1 U8158 ( .A1(n14309), .A2(n14310), .ZN(n6722) );
  NAND2_X1 U8159 ( .A1(n14309), .A2(n6543), .ZN(n6725) );
  XNOR2_X1 U8160 ( .A(n6523), .B(n7265), .ZN(n14341) );
  INV_X1 U8161 ( .A(n14314), .ZN(n7265) );
  NAND2_X1 U8162 ( .A1(n14343), .A2(n14344), .ZN(n14342) );
  NAND2_X1 U8163 ( .A1(n6736), .A2(n14342), .ZN(n14469) );
  OAI21_X1 U8164 ( .B1(n14343), .B2(n14344), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n6736) );
  NOR2_X1 U8165 ( .A1(n14318), .A2(n14319), .ZN(n14472) );
  OR2_X1 U8166 ( .A1(n14330), .A2(n14329), .ZN(n14348) );
  NOR2_X1 U8167 ( .A1(n15182), .A2(n15183), .ZN(n7065) );
  INV_X1 U8168 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15184) );
  INV_X1 U8169 ( .A(n7065), .ZN(n7274) );
  NAND2_X1 U8170 ( .A1(n7276), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U8171 ( .A1(n15182), .A2(n15183), .ZN(n7276) );
  NAND2_X1 U8172 ( .A1(n6933), .A2(n6932), .ZN(n13492) );
  AND2_X1 U8173 ( .A1(n7644), .A2(n11809), .ZN(n7643) );
  INV_X1 U8174 ( .A(n11809), .ZN(n6989) );
  NAND2_X1 U8175 ( .A1(n13516), .A2(n13519), .ZN(n6705) );
  NOR2_X1 U8176 ( .A1(n13519), .A2(n13516), .ZN(n6706) );
  OAI22_X1 U8177 ( .A1(n13514), .A2(n6552), .B1(n13513), .B2(n7545), .ZN(
        n13517) );
  INV_X1 U8178 ( .A(n13526), .ZN(n7543) );
  INV_X1 U8179 ( .A(n11823), .ZN(n7640) );
  OR2_X1 U8180 ( .A1(n7547), .A2(n13530), .ZN(n7546) );
  OAI21_X1 U8181 ( .B1(n6687), .B2(n6575), .A(n6500), .ZN(n7023) );
  INV_X1 U8182 ( .A(n13529), .ZN(n7547) );
  INV_X1 U8183 ( .A(n13539), .ZN(n7541) );
  INV_X1 U8184 ( .A(n13540), .ZN(n7539) );
  OR3_X1 U8185 ( .A1(n13547), .A2(n13546), .A3(n13575), .ZN(n13581) );
  INV_X1 U8186 ( .A(n11840), .ZN(n7637) );
  INV_X1 U8187 ( .A(n11857), .ZN(n6885) );
  NAND2_X1 U8188 ( .A1(n6530), .A2(n7533), .ZN(n7532) );
  NAND2_X1 U8189 ( .A1(n11872), .A2(n7631), .ZN(n7630) );
  NAND2_X1 U8190 ( .A1(n7635), .A2(n7632), .ZN(n7631) );
  INV_X1 U8191 ( .A(n11881), .ZN(n7664) );
  INV_X1 U8192 ( .A(n11885), .ZN(n7660) );
  INV_X1 U8193 ( .A(n13597), .ZN(n6941) );
  INV_X1 U8194 ( .A(n13602), .ZN(n7554) );
  AOI21_X1 U8195 ( .B1(n6622), .B2(n11887), .A(n6503), .ZN(n7656) );
  INV_X1 U8196 ( .A(n13604), .ZN(n6716) );
  NOR2_X1 U8197 ( .A1(n6943), .A2(n13604), .ZN(n6717) );
  NAND2_X1 U8198 ( .A1(n7551), .A2(n7552), .ZN(n13606) );
  NAND2_X1 U8199 ( .A1(n7654), .A2(n11903), .ZN(n7651) );
  OR2_X1 U8200 ( .A1(n11914), .A2(n11915), .ZN(n7625) );
  AND2_X1 U8201 ( .A1(n7650), .A2(n11903), .ZN(n7649) );
  INV_X1 U8202 ( .A(n7625), .ZN(n7620) );
  INV_X1 U8203 ( .A(n13615), .ZN(n6680) );
  NAND2_X1 U8204 ( .A1(n13614), .A2(n13612), .ZN(n7550) );
  AND2_X1 U8205 ( .A1(n6540), .A2(n6677), .ZN(n6676) );
  NAND2_X1 U8206 ( .A1(n6678), .A2(n13615), .ZN(n6677) );
  NAND2_X1 U8207 ( .A1(n6866), .A2(n6865), .ZN(n11909) );
  NOR2_X1 U8208 ( .A1(n7649), .A2(n7648), .ZN(n6865) );
  NAND2_X1 U8209 ( .A1(n6870), .A2(n6867), .ZN(n6866) );
  NOR2_X1 U8210 ( .A1(n7655), .A2(n11906), .ZN(n7648) );
  NOR2_X1 U8211 ( .A1(n6495), .A2(n11917), .ZN(n7622) );
  NAND2_X1 U8212 ( .A1(n7348), .A2(n6476), .ZN(n7347) );
  INV_X1 U8213 ( .A(n8118), .ZN(n7365) );
  INV_X1 U8214 ( .A(n7773), .ZN(n7362) );
  AND2_X1 U8215 ( .A1(n11942), .A2(n12029), .ZN(n11975) );
  AOI21_X1 U8216 ( .B1(n9631), .B2(n9630), .A(n9629), .ZN(n9632) );
  NAND2_X1 U8217 ( .A1(n6859), .A2(n6858), .ZN(n6855) );
  INV_X1 U8218 ( .A(n6858), .ZN(n6857) );
  NAND2_X1 U8219 ( .A1(n12232), .A2(n15120), .ZN(n10980) );
  INV_X1 U8220 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7581) );
  OAI21_X1 U8221 ( .B1(n8106), .B2(n7363), .A(n7361), .ZN(n7774) );
  INV_X1 U8222 ( .A(n7364), .ZN(n7363) );
  AOI21_X1 U8223 ( .B1(n7364), .B2(n7362), .A(n6636), .ZN(n7361) );
  AOI21_X1 U8224 ( .B1(n8105), .B2(n7773), .A(n7365), .ZN(n7364) );
  INV_X1 U8225 ( .A(n12790), .ZN(n7099) );
  NAND2_X1 U8226 ( .A1(n6514), .A2(n7501), .ZN(n7105) );
  NAND2_X1 U8227 ( .A1(n6514), .A2(n10321), .ZN(n7104) );
  NAND2_X1 U8228 ( .A1(n6877), .A2(n6878), .ZN(n7616) );
  NAND2_X1 U8229 ( .A1(n7628), .A2(n7627), .ZN(n7626) );
  NAND2_X1 U8230 ( .A1(n11975), .A2(n7607), .ZN(n7606) );
  NOR2_X1 U8231 ( .A1(n11977), .A2(n11976), .ZN(n7607) );
  INV_X1 U8232 ( .A(n7668), .ZN(n7666) );
  NOR2_X1 U8233 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7135) );
  NOR2_X1 U8234 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7136) );
  NOR2_X1 U8235 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8411) );
  NOR2_X1 U8236 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8410) );
  NAND2_X1 U8237 ( .A1(n13628), .A2(n13627), .ZN(n13630) );
  AND2_X1 U8238 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9609) );
  NAND2_X1 U8239 ( .A1(n10439), .A2(n10254), .ZN(n6844) );
  AOI21_X1 U8240 ( .B1(n6843), .B2(n10439), .A(n6619), .ZN(n6842) );
  AND2_X1 U8241 ( .A1(n6860), .A2(n15257), .ZN(n6859) );
  OR2_X1 U8242 ( .A1(n6860), .A2(n15257), .ZN(n6858) );
  NAND2_X1 U8243 ( .A1(n9002), .A2(n7587), .ZN(n7586) );
  AOI21_X1 U8244 ( .B1(n7587), .B2(n9004), .A(n7585), .ZN(n7584) );
  INV_X1 U8245 ( .A(n9190), .ZN(n7585) );
  INV_X1 U8246 ( .A(n9001), .ZN(n7589) );
  INV_X1 U8247 ( .A(n8775), .ZN(n7597) );
  INV_X1 U8248 ( .A(n6846), .ZN(n6845) );
  OAI21_X1 U8249 ( .B1(n8595), .B2(n6850), .A(n8671), .ZN(n6846) );
  INV_X1 U8250 ( .A(n8598), .ZN(n6850) );
  INV_X1 U8251 ( .A(n8538), .ZN(n7593) );
  OAI21_X1 U8252 ( .B1(n11332), .B2(n7002), .A(n7001), .ZN(n8582) );
  NAND2_X1 U8253 ( .A1(n11332), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7001) );
  OAI21_X1 U8254 ( .B1(n11332), .B2(n8523), .A(n6862), .ZN(n6861) );
  NAND2_X1 U8255 ( .A1(n11332), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6862) );
  INV_X1 U8256 ( .A(n8507), .ZN(n8501) );
  AND2_X1 U8257 ( .A1(n12140), .A2(n8347), .ZN(n8387) );
  NAND2_X1 U8258 ( .A1(n7415), .A2(n12139), .ZN(n8389) );
  NAND2_X1 U8259 ( .A1(n7416), .A2(n12479), .ZN(n7415) );
  OR2_X1 U8260 ( .A1(n10585), .A2(n10586), .ZN(n7122) );
  XNOR2_X1 U8261 ( .A(n12725), .B(n7366), .ZN(n11065) );
  INV_X1 U8262 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15199) );
  INV_X1 U8263 ( .A(n8003), .ZN(n7561) );
  OR2_X1 U8264 ( .A1(n7945), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U8265 ( .A1(n10980), .A2(n10979), .ZN(n7833) );
  NAND2_X1 U8266 ( .A1(n15071), .A2(n9898), .ZN(n10979) );
  NAND2_X1 U8267 ( .A1(n7572), .A2(n7850), .ZN(n10212) );
  NAND2_X1 U8268 ( .A1(n12759), .A2(n8449), .ZN(n9693) );
  NAND2_X1 U8269 ( .A1(n7714), .A2(n7576), .ZN(n7575) );
  INV_X1 U8270 ( .A(n7761), .ZN(n7355) );
  INV_X1 U8271 ( .A(n7356), .ZN(n6765) );
  NAND2_X1 U8272 ( .A1(n7754), .A2(n7753), .ZN(n7755) );
  NAND2_X1 U8273 ( .A1(n7961), .A2(n7752), .ZN(n7754) );
  INV_X1 U8274 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7702) );
  NOR2_X1 U8275 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7703) );
  INV_X1 U8276 ( .A(n7750), .ZN(n6756) );
  AND2_X1 U8277 ( .A1(n7496), .A2(n12829), .ZN(n6748) );
  INV_X1 U8278 ( .A(n7100), .ZN(n7098) );
  NAND2_X1 U8279 ( .A1(n7103), .A2(n7099), .ZN(n7097) );
  NAND2_X1 U8280 ( .A1(n14871), .A2(n8965), .ZN(n9327) );
  INV_X1 U8281 ( .A(n11762), .ZN(n8965) );
  NAND2_X1 U8282 ( .A1(n7684), .A2(n6747), .ZN(n6749) );
  OR2_X1 U8283 ( .A1(n11983), .A2(n11982), .ZN(n7670) );
  NOR2_X1 U8284 ( .A1(n11726), .A2(n14889), .ZN(n6935) );
  NOR2_X1 U8285 ( .A1(n13263), .A2(n13267), .ZN(n7144) );
  AND2_X1 U8286 ( .A1(n11710), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n11727) );
  OR2_X1 U8287 ( .A1(n13276), .A2(n12799), .ZN(n13012) );
  OR2_X1 U8288 ( .A1(n13323), .A2(n13328), .ZN(n7149) );
  OR2_X1 U8289 ( .A1(n7498), .A2(n13023), .ZN(n7673) );
  INV_X1 U8290 ( .A(n7458), .ZN(n6778) );
  INV_X1 U8291 ( .A(n10674), .ZN(n7519) );
  AND2_X1 U8292 ( .A1(n9532), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9540) );
  AND2_X1 U8293 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9334) );
  AND2_X1 U8294 ( .A1(n9334), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9532) );
  NOR2_X1 U8295 ( .A1(n13056), .A2(n7515), .ZN(n7514) );
  INV_X1 U8296 ( .A(n13015), .ZN(n7515) );
  NAND2_X1 U8297 ( .A1(n6801), .A2(n6800), .ZN(n13195) );
  AND2_X1 U8298 ( .A1(n6921), .A2(n6802), .ZN(n6801) );
  INV_X1 U8299 ( .A(n7149), .ZN(n6802) );
  NOR2_X1 U8300 ( .A1(n13318), .A2(n7148), .ZN(n6921) );
  OR2_X1 U8301 ( .A1(n14847), .A2(n11822), .ZN(n9953) );
  NOR2_X1 U8302 ( .A1(n9737), .A2(n11801), .ZN(n9809) );
  NAND2_X1 U8303 ( .A1(n7147), .A2(n11790), .ZN(n9737) );
  INV_X1 U8304 ( .A(n10040), .ZN(n7147) );
  INV_X1 U8305 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8892) );
  NOR2_X1 U8306 ( .A1(n13378), .A2(n11331), .ZN(n7314) );
  INV_X1 U8307 ( .A(n13427), .ZN(n7311) );
  INV_X1 U8308 ( .A(n9068), .ZN(n11476) );
  NOR2_X1 U8309 ( .A1(n7327), .A2(n7320), .ZN(n7319) );
  INV_X1 U8310 ( .A(n7328), .ZN(n7320) );
  NOR2_X1 U8311 ( .A1(n11305), .A2(n13439), .ZN(n11319) );
  INV_X1 U8312 ( .A(n11616), .ZN(n7393) );
  INV_X1 U8313 ( .A(n7248), .ZN(n7247) );
  NAND2_X1 U8314 ( .A1(n11289), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U8315 ( .A1(n7401), .A2(n7400), .ZN(n7399) );
  INV_X1 U8316 ( .A(n11615), .ZN(n7400) );
  NOR2_X1 U8317 ( .A1(n7402), .A2(n11615), .ZN(n7398) );
  NOR2_X1 U8318 ( .A1(n13559), .A2(n7258), .ZN(n7257) );
  INV_X1 U8319 ( .A(n10719), .ZN(n7258) );
  NOR2_X1 U8320 ( .A1(n7203), .A2(n14702), .ZN(n7202) );
  INV_X1 U8321 ( .A(n7204), .ZN(n7203) );
  AND2_X1 U8322 ( .A1(n9609), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9790) );
  AOI21_X1 U8323 ( .B1(n11465), .B2(n11179), .A(n7605), .ZN(n7604) );
  INV_X1 U8324 ( .A(n11610), .ZN(n7605) );
  INV_X1 U8325 ( .A(n11179), .ZN(n7602) );
  INV_X1 U8326 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7093) );
  INV_X1 U8327 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7095) );
  AND2_X1 U8328 ( .A1(n8755), .A2(n8756), .ZN(n7530) );
  INV_X1 U8329 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U8330 ( .A1(n8602), .A2(n8423), .ZN(n8712) );
  INV_X1 U8331 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8423) );
  XNOR2_X1 U8332 ( .A(n10534), .B(SI_24_), .ZN(n10532) );
  NAND2_X1 U8333 ( .A1(n9719), .A2(n9718), .ZN(n10103) );
  NAND2_X1 U8334 ( .A1(n9716), .A2(n9715), .ZN(n9719) );
  NAND2_X1 U8335 ( .A1(n9002), .A2(n9001), .ZN(n9204) );
  OR2_X1 U8336 ( .A1(n8542), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U8337 ( .A1(n6861), .A2(SI_6_), .ZN(n8538) );
  XNOR2_X1 U8338 ( .A(n6861), .B(SI_6_), .ZN(n8535) );
  INV_X1 U8339 ( .A(n8524), .ZN(n8516) );
  AND2_X1 U8340 ( .A1(n9216), .A2(n8521), .ZN(n8540) );
  NOR2_X1 U8341 ( .A1(n8531), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9216) );
  OAI21_X1 U8342 ( .B1(n8494), .B2(n8499), .A(n6954), .ZN(n8507) );
  NAND2_X1 U8343 ( .A1(n8494), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U8344 ( .A1(n8486), .A2(n8485), .ZN(n8504) );
  INV_X1 U8345 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8427) );
  NOR2_X2 U8346 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8454) );
  OAI21_X1 U8347 ( .B1(n8494), .B2(n7611), .A(n7610), .ZN(n8484) );
  NAND2_X1 U8348 ( .A1(n8494), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7610) );
  XNOR2_X1 U8349 ( .A(n14234), .B(n7059), .ZN(n14291) );
  INV_X1 U8350 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7059) );
  NAND2_X1 U8351 ( .A1(n7064), .A2(n14238), .ZN(n14239) );
  NAND2_X1 U8352 ( .A1(n14281), .A2(n14237), .ZN(n7064) );
  XNOR2_X1 U8353 ( .A(n14239), .B(n7063), .ZN(n14299) );
  INV_X1 U8354 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7063) );
  AOI22_X1 U8355 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14243), .B1(n14304), .B2(
        n14242), .ZN(n14245) );
  OR2_X1 U8356 ( .A1(n14243), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14242) );
  INV_X1 U8357 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14243) );
  OAI21_X1 U8358 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14255), .A(n14254), .ZN(
        n14316) );
  NAND2_X1 U8359 ( .A1(n8289), .A2(n12229), .ZN(n6696) );
  OAI21_X1 U8360 ( .B1(n12090), .B2(n7428), .A(n7425), .ZN(n10780) );
  AOI21_X1 U8361 ( .B1(n7427), .B2(n7426), .A(n6567), .ZN(n7425) );
  INV_X1 U8362 ( .A(n12089), .ZN(n7426) );
  INV_X1 U8363 ( .A(n8043), .ZN(n7692) );
  NAND2_X1 U8364 ( .A1(n12090), .A2(n12089), .ZN(n12088) );
  OR2_X1 U8365 ( .A1(n8349), .A2(n12196), .ZN(n12198) );
  NAND2_X1 U8366 ( .A1(n11215), .A2(n8314), .ZN(n12119) );
  OR2_X1 U8367 ( .A1(n7997), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U8368 ( .A1(n7691), .A2(n15320), .ZN(n8028) );
  INV_X1 U8369 ( .A(n8011), .ZN(n7691) );
  NAND2_X1 U8370 ( .A1(n6762), .A2(n6761), .ZN(n6760) );
  NOR2_X1 U8371 ( .A1(n11150), .A2(n11124), .ZN(n6761) );
  NAND2_X1 U8372 ( .A1(n11126), .A2(n11125), .ZN(n6762) );
  NAND2_X1 U8373 ( .A1(n12633), .A2(n11149), .ZN(n7195) );
  AOI21_X1 U8374 ( .B1(n11120), .B2(n6956), .A(n11151), .ZN(n11156) );
  OR2_X1 U8375 ( .A1(n9359), .A2(n15109), .ZN(n9361) );
  NAND2_X1 U8376 ( .A1(n6812), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7124) );
  NAND2_X1 U8377 ( .A1(n12369), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7123) );
  NAND2_X1 U8378 ( .A1(n9313), .A2(n9147), .ZN(n6659) );
  NAND2_X1 U8379 ( .A1(n6659), .A2(n9173), .ZN(n9148) );
  NAND2_X1 U8380 ( .A1(n9482), .A2(n9481), .ZN(n6663) );
  OR2_X1 U8381 ( .A1(n14941), .A2(n14942), .ZN(n7282) );
  NAND2_X1 U8382 ( .A1(n6577), .A2(n7038), .ZN(n7045) );
  NOR2_X1 U8383 ( .A1(n7044), .A2(n15175), .ZN(n7037) );
  NAND2_X1 U8384 ( .A1(n9882), .A2(n7040), .ZN(n7036) );
  NOR2_X1 U8385 ( .A1(n7042), .A2(n7041), .ZN(n7040) );
  INV_X1 U8386 ( .A(n9881), .ZN(n7042) );
  NAND2_X1 U8387 ( .A1(n7039), .A2(n7041), .ZN(n7038) );
  INV_X1 U8388 ( .A(n9882), .ZN(n7039) );
  NAND2_X1 U8389 ( .A1(n9874), .A2(n9875), .ZN(n14953) );
  AND2_X1 U8390 ( .A1(n9864), .A2(n9863), .ZN(n9865) );
  NAND2_X1 U8391 ( .A1(n10236), .A2(n6614), .ZN(n7051) );
  NAND2_X1 U8392 ( .A1(n7056), .A2(n7055), .ZN(n7054) );
  INV_X1 U8393 ( .A(n10235), .ZN(n7056) );
  NAND2_X1 U8394 ( .A1(n6810), .A2(n10582), .ZN(n14984) );
  NAND2_X1 U8395 ( .A1(n6811), .A2(n10581), .ZN(n6810) );
  NAND2_X1 U8396 ( .A1(n10223), .A2(n10222), .ZN(n7278) );
  INV_X1 U8397 ( .A(n7122), .ZN(n12250) );
  NAND2_X1 U8398 ( .A1(n14979), .A2(n7048), .ZN(n7046) );
  NAND2_X1 U8399 ( .A1(n7082), .A2(n14969), .ZN(n7079) );
  INV_X1 U8400 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12110) );
  NOR2_X1 U8401 ( .A1(n7163), .A2(n7075), .ZN(n7071) );
  INV_X1 U8402 ( .A(n14998), .ZN(n7074) );
  NAND2_X1 U8403 ( .A1(n12349), .A2(n12348), .ZN(n7084) );
  NOR2_X1 U8404 ( .A1(n12427), .A2(n15096), .ZN(n7025) );
  AOI21_X1 U8405 ( .B1(n7170), .B2(n11076), .A(n11083), .ZN(n7169) );
  INV_X1 U8406 ( .A(n7171), .ZN(n7170) );
  NAND2_X1 U8407 ( .A1(n7697), .A2(n7696), .ZN(n8150) );
  INV_X1 U8408 ( .A(n11065), .ZN(n12486) );
  NAND2_X1 U8409 ( .A1(n7695), .A2(n7694), .ZN(n8109) );
  OR2_X1 U8410 ( .A1(n8109), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U8411 ( .A1(n6652), .A2(n11061), .ZN(n12512) );
  AND2_X1 U8412 ( .A1(n11069), .A2(n11064), .ZN(n12511) );
  NAND2_X1 U8413 ( .A1(n7693), .A2(n15199), .ZN(n8085) );
  INV_X1 U8414 ( .A(n8073), .ZN(n7693) );
  OR2_X1 U8415 ( .A1(n8085), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8099) );
  OR2_X1 U8416 ( .A1(n12689), .A2(n12570), .ZN(n12560) );
  NAND2_X1 U8417 ( .A1(n12582), .A2(n8050), .ZN(n12566) );
  NAND2_X1 U8418 ( .A1(n12599), .A2(n11035), .ZN(n12588) );
  NAND2_X1 U8419 ( .A1(n12588), .A2(n12587), .ZN(n12590) );
  OAI21_X1 U8420 ( .B1(n12618), .B2(n7562), .A(n7560), .ZN(n12596) );
  INV_X1 U8421 ( .A(n7563), .ZN(n7562) );
  AOI21_X1 U8422 ( .B1(n7563), .B2(n7561), .A(n6564), .ZN(n7560) );
  AOI21_X1 U8423 ( .B1(n12629), .B2(n8003), .A(n6557), .ZN(n7563) );
  AOI21_X1 U8424 ( .B1(n7189), .B2(n7188), .A(n7187), .ZN(n7186) );
  INV_X1 U8425 ( .A(n11027), .ZN(n7188) );
  INV_X1 U8426 ( .A(n11034), .ZN(n7187) );
  AND2_X1 U8427 ( .A1(n11036), .A2(n11035), .ZN(n12600) );
  NAND2_X1 U8428 ( .A1(n7688), .A2(n12110), .ZN(n7983) );
  INV_X1 U8429 ( .A(n7968), .ZN(n7688) );
  NAND2_X1 U8430 ( .A1(n7690), .A2(n7689), .ZN(n7997) );
  INV_X1 U8431 ( .A(n7983), .ZN(n7690) );
  OR2_X1 U8432 ( .A1(n10957), .A2(n11028), .ZN(n14352) );
  NAND2_X1 U8433 ( .A1(n10754), .A2(n10753), .ZN(n10752) );
  INV_X1 U8434 ( .A(n12227), .ZN(n14356) );
  AND2_X1 U8435 ( .A1(n15018), .A2(n15022), .ZN(n15019) );
  AND2_X1 U8436 ( .A1(n7895), .A2(n15348), .ZN(n7913) );
  NAND2_X1 U8437 ( .A1(n7913), .A2(n7912), .ZN(n7926) );
  AND2_X1 U8438 ( .A1(n11002), .A2(n11003), .ZN(n11129) );
  NAND2_X1 U8439 ( .A1(n7580), .A2(n7894), .ZN(n15037) );
  NOR2_X1 U8440 ( .A1(n7880), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7895) );
  AND2_X1 U8441 ( .A1(n7866), .A2(n7850), .ZN(n7571) );
  OR2_X1 U8442 ( .A1(n7868), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7880) );
  INV_X1 U8443 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7852) );
  INV_X1 U8444 ( .A(n7833), .ZN(n11133) );
  NAND2_X1 U8445 ( .A1(n7818), .A2(n6958), .ZN(n15077) );
  NAND2_X1 U8446 ( .A1(n15090), .A2(n15089), .ZN(n15092) );
  AND2_X1 U8447 ( .A1(n9690), .A2(n6477), .ZN(n10861) );
  AOI21_X1 U8448 ( .B1(n12428), .B2(n8045), .A(n7728), .ZN(n12440) );
  NAND2_X1 U8449 ( .A1(n8268), .A2(n11154), .ZN(n15099) );
  INV_X1 U8450 ( .A(n15160), .ZN(n15156) );
  NAND2_X1 U8451 ( .A1(n7783), .A2(n7782), .ZN(n8191) );
  OR2_X1 U8452 ( .A1(n8176), .A2(n7781), .ZN(n7783) );
  NAND2_X1 U8453 ( .A1(n6769), .A2(n7778), .ZN(n8161) );
  NAND2_X1 U8454 ( .A1(n8147), .A2(n7777), .ZN(n6769) );
  NAND2_X1 U8455 ( .A1(n8134), .A2(n7776), .ZN(n8147) );
  XNOR2_X1 U8456 ( .A(n8265), .B(n8264), .ZN(n9141) );
  OAI21_X1 U8457 ( .B1(n8263), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8265) );
  AND2_X1 U8458 ( .A1(n7769), .A2(n7768), .ZN(n8065) );
  NAND2_X1 U8459 ( .A1(n8024), .A2(n8023), .ZN(n7438) );
  AND2_X1 U8460 ( .A1(n8023), .A2(n7437), .ZN(n7436) );
  INV_X1 U8461 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U8462 ( .A1(n7757), .A2(n7756), .ZN(n7992) );
  XNOR2_X1 U8463 ( .A(n7755), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n7976) );
  AND2_X1 U8464 ( .A1(n7748), .A2(n7747), .ZN(n7920) );
  AND2_X1 U8465 ( .A1(n7746), .A2(n7745), .ZN(n7906) );
  NOR2_X1 U8466 ( .A1(n7902), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7937) );
  OR2_X1 U8467 ( .A1(n7901), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7902) );
  AND2_X1 U8468 ( .A1(n7744), .A2(n7742), .ZN(n7886) );
  AND2_X1 U8469 ( .A1(n6775), .A2(n6774), .ZN(n7859) );
  NAND2_X1 U8470 ( .A1(n6777), .A2(n7736), .ZN(n6775) );
  NOR2_X1 U8471 ( .A1(n7338), .A2(n6773), .ZN(n6772) );
  AND2_X1 U8472 ( .A1(n7738), .A2(n7737), .ZN(n7858) );
  INV_X1 U8473 ( .A(n9145), .ZN(n7027) );
  XNOR2_X1 U8474 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7794) );
  NAND2_X1 U8475 ( .A1(n8911), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7803) );
  NOR2_X1 U8476 ( .A1(n7501), .A2(n10319), .ZN(n7500) );
  INV_X1 U8477 ( .A(n7502), .ZN(n7501) );
  INV_X1 U8478 ( .A(n7487), .ZN(n7103) );
  AOI21_X1 U8479 ( .B1(n7487), .B2(n7102), .A(n7101), .ZN(n7100) );
  INV_X1 U8480 ( .A(n11528), .ZN(n7101) );
  INV_X1 U8481 ( .A(n12782), .ZN(n7102) );
  NOR2_X1 U8482 ( .A1(n12847), .A2(n7488), .ZN(n7487) );
  INV_X1 U8483 ( .A(n12781), .ZN(n7488) );
  NAND2_X1 U8484 ( .A1(n12783), .A2(n12782), .ZN(n7489) );
  NAND2_X1 U8485 ( .A1(n6744), .A2(n6743), .ZN(n11570) );
  INV_X1 U8486 ( .A(n7096), .ZN(n6743) );
  NAND2_X1 U8487 ( .A1(n12783), .A2(n6535), .ZN(n6744) );
  OAI21_X1 U8488 ( .B1(n7098), .B2(n7097), .A(n11541), .ZN(n7096) );
  INV_X1 U8489 ( .A(n11547), .ZN(n11548) );
  OR2_X1 U8490 ( .A1(n10266), .A2(n10267), .ZN(n6753) );
  XNOR2_X1 U8491 ( .A(n9327), .B(n14814), .ZN(n9372) );
  INV_X1 U8492 ( .A(n9565), .ZN(n7492) );
  NAND2_X1 U8493 ( .A1(n12798), .A2(n12797), .ZN(n7486) );
  NOR2_X1 U8494 ( .A1(n8919), .A2(n14803), .ZN(n8923) );
  AND2_X1 U8495 ( .A1(n12042), .A2(n11957), .ZN(n8960) );
  NAND2_X1 U8496 ( .A1(n6742), .A2(n6556), .ZN(n8617) );
  INV_X1 U8497 ( .A(n8894), .ZN(n6742) );
  INV_X1 U8498 ( .A(n6950), .ZN(n11958) );
  OR2_X1 U8499 ( .A1(n11741), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8985) );
  AOI21_X1 U8500 ( .B1(n12901), .B2(n12900), .A(n12899), .ZN(n12903) );
  AOI21_X1 U8501 ( .B1(n8728), .B2(n8727), .A(n8726), .ZN(n8725) );
  NOR2_X1 U8502 ( .A1(n9027), .A2(n6822), .ZN(n12919) );
  AND2_X1 U8503 ( .A1(n9643), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6822) );
  OR2_X1 U8504 ( .A1(n9031), .A2(n9030), .ZN(n6827) );
  NAND2_X1 U8505 ( .A1(n14755), .A2(n12938), .ZN(n12939) );
  INV_X1 U8506 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8893) );
  XNOR2_X1 U8507 ( .A(n12970), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n12978) );
  NOR2_X1 U8508 ( .A1(n12969), .A2(n12968), .ZN(n12970) );
  OAI21_X1 U8509 ( .B1(n13092), .B2(n13041), .A(n13040), .ZN(n13078) );
  NAND2_X1 U8510 ( .A1(n13102), .A2(n13090), .ZN(n13086) );
  AND2_X1 U8511 ( .A1(n13012), .A2(n13013), .ZN(n13091) );
  NAND2_X1 U8512 ( .A1(n6799), .A2(n13037), .ZN(n13122) );
  AOI21_X1 U8513 ( .B1(n13115), .B2(n6902), .A(n6521), .ZN(n6899) );
  NAND2_X1 U8514 ( .A1(n13115), .A2(n13133), .ZN(n6901) );
  NAND2_X1 U8515 ( .A1(n6903), .A2(n7476), .ZN(n13004) );
  AOI21_X1 U8516 ( .B1(n7477), .B2(n7480), .A(n13178), .ZN(n7476) );
  NAND2_X1 U8517 ( .A1(n6788), .A2(n7453), .ZN(n6787) );
  NAND2_X1 U8518 ( .A1(n13024), .A2(n6784), .ZN(n6788) );
  NOR2_X1 U8519 ( .A1(n13000), .A2(n13318), .ZN(n7457) );
  NOR2_X1 U8520 ( .A1(n11197), .A2(n12960), .ZN(n11510) );
  INV_X1 U8521 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n12960) );
  NOR3_X1 U8522 ( .A1(n7149), .A2(n10896), .A3(n13318), .ZN(n13211) );
  NOR2_X1 U8523 ( .A1(n10896), .A2(n7149), .ZN(n13229) );
  NOR2_X1 U8524 ( .A1(n10469), .A2(n10467), .ZN(n10481) );
  NAND2_X1 U8525 ( .A1(n7517), .A2(n6887), .ZN(n10837) );
  AOI21_X1 U8526 ( .B1(n7521), .B2(n7518), .A(n10673), .ZN(n7517) );
  NAND2_X1 U8527 ( .A1(n10450), .A2(n7518), .ZN(n6887) );
  AND2_X1 U8528 ( .A1(n7520), .A2(n7519), .ZN(n7518) );
  NAND2_X1 U8529 ( .A1(n11860), .A2(n12885), .ZN(n7458) );
  NAND2_X1 U8530 ( .A1(n6907), .A2(n6780), .ZN(n6779) );
  NOR2_X1 U8531 ( .A1(n6781), .A2(n7459), .ZN(n6780) );
  NOR2_X1 U8532 ( .A1(n11860), .A2(n12885), .ZN(n7459) );
  INV_X1 U8533 ( .A(n10521), .ZN(n6781) );
  AND2_X1 U8534 ( .A1(n10525), .A2(n10685), .ZN(n10680) );
  NOR2_X1 U8535 ( .A1(n10445), .A2(n11851), .ZN(n10525) );
  OR2_X1 U8536 ( .A1(n10184), .A2(n10183), .ZN(n10194) );
  OR2_X1 U8537 ( .A1(n14868), .A2(n11839), .ZN(n7675) );
  OR2_X1 U8538 ( .A1(n10299), .A2(n14878), .ZN(n10445) );
  NAND2_X1 U8539 ( .A1(n10288), .A2(n14868), .ZN(n10299) );
  NAND2_X1 U8540 ( .A1(n7152), .A2(n14853), .ZN(n10055) );
  INV_X1 U8541 ( .A(n7152), .ZN(n10054) );
  AND2_X1 U8542 ( .A1(n9809), .A2(n14836), .ZN(n9930) );
  NAND2_X1 U8543 ( .A1(n9731), .A2(n12006), .ZN(n9805) );
  XNOR2_X1 U8544 ( .A(n12895), .B(n11786), .ZN(n12008) );
  NAND2_X1 U8545 ( .A1(n13242), .A2(n14822), .ZN(n10040) );
  NAND2_X1 U8546 ( .A1(n11507), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U8547 ( .A1(n13249), .A2(n6953), .ZN(n9422) );
  NOR2_X1 U8548 ( .A1(n14814), .A2(n13244), .ZN(n13242) );
  NAND2_X1 U8549 ( .A1(n6940), .A2(n13241), .ZN(n13240) );
  NAND2_X1 U8550 ( .A1(n6906), .A2(n13244), .ZN(n9454) );
  OR2_X1 U8551 ( .A1(n11957), .A2(n12042), .ZN(n9463) );
  NAND2_X1 U8552 ( .A1(n6898), .A2(n6894), .ZN(n9957) );
  AND2_X1 U8553 ( .A1(n6895), .A2(n12007), .ZN(n9940) );
  INV_X1 U8554 ( .A(n14867), .ZN(n14879) );
  AND2_X1 U8555 ( .A1(n8887), .A2(n8879), .ZN(n14799) );
  NAND2_X1 U8556 ( .A1(n7141), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8615) );
  OAI21_X1 U8557 ( .B1(n8419), .B2(n8421), .A(n8420), .ZN(n10258) );
  XNOR2_X1 U8558 ( .A(n7473), .B(P2_IR_REG_21__SCAN_IN), .ZN(n11957) );
  OAI21_X1 U8559 ( .B1(n8894), .B2(P2_IR_REG_20__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7473) );
  INV_X1 U8560 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8911) );
  AOI21_X1 U8561 ( .B1(n13370), .B2(n11441), .A(n11464), .ZN(n7298) );
  INV_X1 U8562 ( .A(n7298), .ZN(n7295) );
  INV_X1 U8563 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U8564 ( .A1(n7309), .A2(n6487), .ZN(n13428) );
  NAND2_X1 U8565 ( .A1(n13456), .A2(n7314), .ZN(n7309) );
  NOR2_X1 U8566 ( .A1(n9982), .A2(n9981), .ZN(n9990) );
  AND2_X1 U8567 ( .A1(n10541), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U8568 ( .A1(n10612), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10709) );
  INV_X1 U8569 ( .A(n11336), .ZN(n11337) );
  NOR2_X1 U8570 ( .A1(n10356), .A2(n10355), .ZN(n10541) );
  OR2_X1 U8571 ( .A1(n10341), .A2(n10340), .ZN(n10356) );
  NAND2_X1 U8572 ( .A1(n7299), .A2(n7300), .ZN(n13415) );
  AOI21_X1 U8573 ( .B1(n7302), .B2(n7308), .A(n7301), .ZN(n7300) );
  INV_X1 U8574 ( .A(n13416), .ZN(n7301) );
  OR2_X1 U8575 ( .A1(n10722), .A2(n10721), .ZN(n10934) );
  OR2_X1 U8576 ( .A1(n10709), .A2(n10708), .ZN(n10722) );
  AND3_X1 U8577 ( .A1(n13642), .A2(n13641), .A3(n13640), .ZN(n13806) );
  INV_X1 U8578 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14292) );
  INV_X1 U8579 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14300) );
  NAND2_X1 U8580 ( .A1(n6974), .A2(n6973), .ZN(n9197) );
  INV_X1 U8581 ( .A(n9010), .ZN(n6974) );
  AOI21_X1 U8582 ( .B1(n7262), .B2(n13897), .A(n7261), .ZN(n7260) );
  INV_X1 U8583 ( .A(n11607), .ZN(n7261) );
  NAND2_X1 U8584 ( .A1(n7209), .A2(n7208), .ZN(n13881) );
  NAND2_X1 U8585 ( .A1(n7211), .A2(n7210), .ZN(n13902) );
  AOI21_X1 U8586 ( .B1(n7383), .B2(n7387), .A(n6570), .ZN(n7381) );
  INV_X1 U8587 ( .A(n7211), .ZN(n13935) );
  NOR3_X1 U8588 ( .A1(n10764), .A2(n7207), .A3(n14390), .ZN(n14027) );
  OAI21_X1 U8589 ( .B1(n11598), .B2(n11597), .A(n11596), .ZN(n14022) );
  NOR2_X1 U8590 ( .A1(n10764), .A2(n7207), .ZN(n14025) );
  AND2_X1 U8591 ( .A1(n14586), .A2(n7200), .ZN(n10625) );
  NOR2_X1 U8592 ( .A1(n14416), .A2(n7201), .ZN(n7200) );
  INV_X1 U8593 ( .A(n7202), .ZN(n7201) );
  NAND2_X1 U8594 ( .A1(n7215), .A2(n7217), .ZN(n10622) );
  AND2_X1 U8595 ( .A1(n7218), .A2(n10554), .ZN(n7217) );
  NAND2_X1 U8596 ( .A1(n14562), .A2(n7216), .ZN(n7215) );
  OR2_X1 U8597 ( .A1(n7411), .A2(n7410), .ZN(n7409) );
  INV_X1 U8598 ( .A(n10348), .ZN(n7410) );
  NAND2_X1 U8599 ( .A1(n14586), .A2(n7204), .ZN(n14571) );
  NAND2_X1 U8600 ( .A1(n14586), .A2(n10003), .ZN(n14569) );
  AND2_X1 U8601 ( .A1(n14588), .A2(n14676), .ZN(n14586) );
  NAND2_X1 U8602 ( .A1(n7222), .A2(n7224), .ZN(n14577) );
  AOI21_X1 U8603 ( .B1(n13676), .B2(n7225), .A(n6559), .ZN(n7224) );
  NAND2_X1 U8604 ( .A1(n10087), .A2(n7223), .ZN(n7222) );
  AND2_X1 U8605 ( .A1(n9790), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U8606 ( .A1(n7376), .A2(n7375), .ZN(n9997) );
  AOI21_X1 U8607 ( .B1(n7378), .B2(n13674), .A(n6563), .ZN(n7375) );
  NAND2_X1 U8608 ( .A1(n10018), .A2(n7377), .ZN(n7376) );
  NOR2_X1 U8609 ( .A1(n10089), .A2(n13515), .ZN(n14588) );
  NAND2_X1 U8610 ( .A1(n7379), .A2(n9845), .ZN(n10094) );
  NAND2_X1 U8611 ( .A1(n7197), .A2(n14671), .ZN(n10089) );
  OR2_X1 U8612 ( .A1(n10124), .A2(n13498), .ZN(n14603) );
  NOR2_X1 U8613 ( .A1(n14603), .A2(n14602), .ZN(n14606) );
  XNOR2_X1 U8614 ( .A(n14636), .B(n13498), .ZN(n13496) );
  AND2_X1 U8615 ( .A1(n13832), .A2(n13831), .ZN(n14057) );
  INV_X1 U8616 ( .A(n14701), .ZN(n14691) );
  OR2_X1 U8617 ( .A1(n9839), .A2(n13489), .ZN(n14647) );
  OR3_X1 U8618 ( .A1(n9836), .A2(n9835), .A3(n9834), .ZN(n11641) );
  NAND2_X1 U8619 ( .A1(n9113), .A2(n9112), .ZN(n11638) );
  INV_X1 U8620 ( .A(n14708), .ZN(n14639) );
  INV_X1 U8621 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U8622 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n7374) );
  AND2_X1 U8623 ( .A1(n14210), .A2(n9048), .ZN(n7373) );
  NOR2_X1 U8624 ( .A1(n9048), .A2(n6937), .ZN(n7372) );
  NAND2_X1 U8625 ( .A1(n14210), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7371) );
  XNOR2_X1 U8626 ( .A(n11611), .B(n11610), .ZN(n11931) );
  OAI21_X1 U8627 ( .B1(n11466), .B2(n11465), .A(n11179), .ZN(n11611) );
  XNOR2_X1 U8628 ( .A(n11466), .B(n11465), .ZN(n11721) );
  XNOR2_X1 U8629 ( .A(n11445), .B(n11444), .ZN(n13364) );
  INV_X1 U8630 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8754) );
  XNOR2_X1 U8631 ( .A(n8753), .B(P1_IR_REG_21__SCAN_IN), .ZN(n13645) );
  OR2_X1 U8632 ( .A1(n9002), .A2(n9004), .ZN(n7583) );
  INV_X1 U8633 ( .A(n6837), .ZN(n8997) );
  AOI21_X1 U8634 ( .B1(n8687), .B2(n7595), .A(n6840), .ZN(n6837) );
  NAND2_X1 U8635 ( .A1(n8687), .A2(n8686), .ZN(n8693) );
  NAND2_X1 U8636 ( .A1(n8454), .A2(n8427), .ZN(n8520) );
  XNOR2_X1 U8637 ( .A(n8484), .B(n8460), .ZN(n8483) );
  OAI21_X1 U8638 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n14232), .A(n14231), .ZN(
        n14284) );
  XNOR2_X1 U8639 ( .A(n14281), .B(n14237), .ZN(n14282) );
  NAND2_X1 U8640 ( .A1(n7268), .A2(n14306), .ZN(n14308) );
  AOI21_X1 U8641 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14251), .A(n14250), .ZN(
        n14277) );
  NOR2_X1 U8642 ( .A1(n14313), .A2(n14312), .ZN(n14250) );
  AOI21_X1 U8643 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14516), .A(n14256), .ZN(
        n14321) );
  NOR2_X1 U8644 ( .A1(n14317), .A2(n14316), .ZN(n14256) );
  AND2_X1 U8645 ( .A1(n12139), .A2(n12479), .ZN(n7414) );
  NAND2_X1 U8646 ( .A1(n7416), .A2(n12139), .ZN(n12075) );
  AND3_X1 U8647 ( .A1(n7941), .A2(n7940), .A3(n7939), .ZN(n10785) );
  NOR2_X1 U8648 ( .A1(n9403), .A2(n6978), .ZN(n9401) );
  INV_X1 U8649 ( .A(n8280), .ZN(n6979) );
  NAND2_X1 U8650 ( .A1(n7419), .A2(n8329), .ZN(n12098) );
  NOR2_X1 U8651 ( .A1(n8287), .A2(n12231), .ZN(n6700) );
  INV_X1 U8652 ( .A(n7432), .ZN(n7431) );
  OAI21_X1 U8653 ( .B1(n7433), .B2(n8314), .A(n8317), .ZN(n7432) );
  NAND2_X1 U8654 ( .A1(n7424), .A2(n7422), .ZN(n10009) );
  AND2_X1 U8655 ( .A1(n7424), .A2(n7423), .ZN(n10010) );
  NAND2_X1 U8656 ( .A1(n12088), .A2(n8295), .ZN(n10657) );
  NAND2_X1 U8657 ( .A1(n8324), .A2(n12571), .ZN(n8325) );
  INV_X1 U8658 ( .A(n8323), .ZN(n8324) );
  NAND2_X1 U8659 ( .A1(n8108), .A2(n8107), .ZN(n12665) );
  AND4_X1 U8660 ( .A1(n7931), .A2(n7930), .A3(n7929), .A4(n7928), .ZN(n12179)
         );
  AND4_X1 U8661 ( .A1(n7950), .A2(n7949), .A3(n7948), .A4(n7947), .ZN(n12173)
         );
  AND2_X1 U8662 ( .A1(n8157), .A2(n8156), .ZN(n12480) );
  OR2_X1 U8663 ( .A1(n8364), .A2(n8363), .ZN(n12213) );
  AND2_X1 U8664 ( .A1(n8362), .A2(n8363), .ZN(n12211) );
  INV_X1 U8665 ( .A(n12203), .ZN(n12219) );
  NAND2_X1 U8666 ( .A1(n8377), .A2(n8376), .ZN(n12217) );
  NAND2_X1 U8667 ( .A1(n6758), .A2(n7194), .ZN(n6911) );
  INV_X1 U8668 ( .A(n11154), .ZN(n7194) );
  XNOR2_X1 U8669 ( .A(n6759), .B(n6480), .ZN(n6758) );
  NAND2_X1 U8670 ( .A1(n6581), .A2(n6760), .ZN(n6759) );
  NAND2_X1 U8671 ( .A1(n11156), .A2(n11155), .ZN(n7192) );
  OR2_X1 U8672 ( .A1(n11152), .A2(n11153), .ZN(n7193) );
  NOR2_X1 U8673 ( .A1(n11148), .A2(n11149), .ZN(n6957) );
  INV_X1 U8674 ( .A(n11119), .ZN(n12407) );
  NAND2_X1 U8675 ( .A1(n8187), .A2(n8186), .ZN(n12425) );
  NAND2_X1 U8676 ( .A1(n8171), .A2(n8170), .ZN(n12223) );
  INV_X1 U8677 ( .A(n12480), .ZN(n12224) );
  INV_X1 U8678 ( .A(n8322), .ZN(n12584) );
  INV_X1 U8679 ( .A(n12619), .ZN(n12226) );
  INV_X1 U8680 ( .A(n12173), .ZN(n15025) );
  NAND2_X1 U8681 ( .A1(n7805), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7791) );
  NAND2_X1 U8682 ( .A1(n7030), .A2(n9159), .ZN(n14926) );
  OAI21_X1 U8683 ( .B1(n9173), .B2(n6659), .A(n9148), .ZN(n14928) );
  NOR2_X1 U8684 ( .A1(n14928), .A2(n14929), .ZN(n14930) );
  OR2_X1 U8685 ( .A1(n9151), .A2(n9150), .ZN(n9482) );
  XNOR2_X1 U8686 ( .A(n6663), .B(n6662), .ZN(n14941) );
  NAND2_X1 U8687 ( .A1(n6661), .A2(n6660), .ZN(n9864) );
  AOI21_X1 U8688 ( .B1(n7281), .B2(n14942), .A(n9484), .ZN(n6660) );
  NAND2_X1 U8689 ( .A1(n14941), .A2(n7281), .ZN(n6661) );
  XNOR2_X1 U8690 ( .A(n7278), .B(n7055), .ZN(n10224) );
  INV_X1 U8691 ( .A(n6811), .ZN(n10583) );
  INV_X1 U8692 ( .A(n7156), .ZN(n14976) );
  NAND2_X1 U8693 ( .A1(n14967), .A2(n7082), .ZN(n7081) );
  NOR2_X1 U8694 ( .A1(n12236), .A2(n6664), .ZN(n14999) );
  NOR2_X1 U8695 ( .A1(n14999), .A2(n14998), .ZN(n15000) );
  NAND2_X1 U8696 ( .A1(n15008), .A2(n12255), .ZN(n12256) );
  INV_X1 U8697 ( .A(n7162), .ZN(n12271) );
  INV_X1 U8698 ( .A(n7280), .ZN(n12295) );
  INV_X1 U8699 ( .A(n12282), .ZN(n7161) );
  INV_X1 U8700 ( .A(n6808), .ZN(n12322) );
  INV_X1 U8701 ( .A(n12306), .ZN(n12307) );
  INV_X1 U8702 ( .A(n7028), .ZN(n12332) );
  INV_X1 U8703 ( .A(n6658), .ZN(n12318) );
  INV_X1 U8704 ( .A(n7154), .ZN(n12336) );
  INV_X1 U8705 ( .A(n6806), .ZN(n12356) );
  INV_X1 U8706 ( .A(n7277), .ZN(n12320) );
  XNOR2_X1 U8707 ( .A(n7130), .B(n7129), .ZN(n7128) );
  INV_X1 U8708 ( .A(n12400), .ZN(n7129) );
  NOR2_X1 U8709 ( .A1(n12394), .A2(n7131), .ZN(n7130) );
  NAND2_X1 U8710 ( .A1(n7127), .A2(n7126), .ZN(n7125) );
  INV_X1 U8711 ( .A(n12401), .ZN(n7126) );
  NAND2_X1 U8712 ( .A1(n14983), .A2(n6480), .ZN(n7127) );
  NAND2_X1 U8713 ( .A1(n8091), .A2(n8090), .ZN(n12520) );
  NAND2_X1 U8714 ( .A1(n12563), .A2(n11040), .ZN(n12553) );
  NAND2_X1 U8715 ( .A1(n12622), .A2(n8003), .ZN(n12608) );
  AND2_X1 U8716 ( .A1(n7967), .A2(n7966), .ZN(n14366) );
  NAND2_X1 U8717 ( .A1(n7174), .A2(n7172), .ZN(n10668) );
  NAND2_X1 U8718 ( .A1(n8240), .A2(n9690), .ZN(n15080) );
  NAND2_X1 U8719 ( .A1(n7175), .A2(n7179), .ZN(n15016) );
  NAND2_X1 U8720 ( .A1(n15035), .A2(n7180), .ZN(n7175) );
  NAND2_X1 U8721 ( .A1(n6648), .A2(n7183), .ZN(n10395) );
  NAND2_X1 U8722 ( .A1(n10208), .A2(n7181), .ZN(n6648) );
  NAND2_X1 U8723 ( .A1(n10210), .A2(n10988), .ZN(n15062) );
  AND3_X1 U8724 ( .A1(n7865), .A2(n7864), .A3(n7863), .ZN(n10249) );
  INV_X1 U8725 ( .A(n9898), .ZN(n15120) );
  NOR2_X1 U8726 ( .A1(n10082), .A2(n15131), .ZN(n12627) );
  AOI21_X1 U8727 ( .B1(n12417), .B2(n7570), .A(n7569), .ZN(n7568) );
  NOR2_X1 U8728 ( .A1(n15181), .A2(n11756), .ZN(n7569) );
  INV_X1 U8729 ( .A(n12633), .ZN(n12710) );
  INV_X1 U8730 ( .A(n12637), .ZN(n12713) );
  AND2_X1 U8731 ( .A1(n12658), .A2(n12657), .ZN(n12723) );
  XNOR2_X1 U8732 ( .A(n6771), .B(n11107), .ZN(n12765) );
  OAI22_X1 U8733 ( .A1(n11106), .A2(n11105), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n14219), .ZN(n6771) );
  NAND2_X1 U8734 ( .A1(n7721), .A2(n7720), .ZN(n12768) );
  NAND2_X1 U8735 ( .A1(n8248), .A2(n6692), .ZN(n6691) );
  NOR2_X1 U8736 ( .A1(n6695), .A2(n6694), .ZN(n6693) );
  NOR2_X1 U8737 ( .A1(n8021), .A2(n7576), .ZN(n6692) );
  OAI21_X1 U8738 ( .B1(n7978), .B2(n7713), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8242) );
  NAND2_X1 U8739 ( .A1(n7712), .A2(n7671), .ZN(n7713) );
  NAND2_X1 U8740 ( .A1(n7367), .A2(n6509), .ZN(n10375) );
  NAND2_X1 U8741 ( .A1(n8135), .A2(n8945), .ZN(n7367) );
  OAI21_X1 U8742 ( .B1(n8106), .B2(n8105), .A(n7773), .ZN(n8119) );
  NAND2_X1 U8743 ( .A1(n8093), .A2(n8092), .ZN(n8095) );
  NAND2_X1 U8744 ( .A1(n7350), .A2(n7353), .ZN(n8093) );
  INV_X1 U8745 ( .A(SI_20_), .ZN(n15325) );
  NAND2_X1 U8746 ( .A1(n7349), .A2(n7353), .ZN(n8082) );
  NAND2_X1 U8747 ( .A1(n7351), .A2(n7353), .ZN(n8080) );
  INV_X1 U8748 ( .A(SI_19_), .ZN(n15267) );
  INV_X1 U8749 ( .A(SI_18_), .ZN(n15344) );
  OAI21_X1 U8750 ( .B1(n8020), .B2(n7345), .A(n7342), .ZN(n8052) );
  NAND2_X1 U8751 ( .A1(n8036), .A2(n8035), .ZN(n8038) );
  NAND2_X1 U8752 ( .A1(n8020), .A2(n7763), .ZN(n8036) );
  INV_X1 U8753 ( .A(SI_16_), .ZN(n15336) );
  NAND2_X1 U8754 ( .A1(n7358), .A2(n7356), .ZN(n8007) );
  NAND2_X1 U8755 ( .A1(n7358), .A2(n7759), .ZN(n8005) );
  INV_X1 U8756 ( .A(SI_15_), .ZN(n9208) );
  INV_X1 U8757 ( .A(SI_14_), .ZN(n15322) );
  NAND2_X1 U8758 ( .A1(n7978), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7994) );
  INV_X1 U8759 ( .A(n7978), .ZN(n7979) );
  INV_X1 U8760 ( .A(SI_13_), .ZN(n8999) );
  INV_X1 U8761 ( .A(SI_11_), .ZN(n8688) );
  NAND2_X1 U8762 ( .A1(n7935), .A2(n7750), .ZN(n7952) );
  XNOR2_X1 U8763 ( .A(n7890), .B(P3_IR_REG_7__SCAN_IN), .ZN(n14956) );
  NAND2_X1 U8764 ( .A1(n7827), .A2(n7734), .ZN(n7841) );
  NAND2_X1 U8765 ( .A1(n7556), .A2(n7555), .ZN(n7842) );
  INV_X1 U8766 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7159) );
  NAND2_X1 U8767 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7283) );
  OR2_X1 U8768 ( .A1(n10442), .A2(n8418), .ZN(n8920) );
  AND2_X1 U8769 ( .A1(n10258), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8891) );
  NAND2_X1 U8770 ( .A1(n9970), .A2(n11951), .ZN(n9637) );
  AND2_X1 U8771 ( .A1(n7109), .A2(n7106), .ZN(n11186) );
  INV_X1 U8772 ( .A(n7500), .ZN(n7109) );
  INV_X1 U8773 ( .A(n7107), .ZN(n7106) );
  OAI21_X1 U8774 ( .B1(n10321), .B2(n7501), .A(n6514), .ZN(n7107) );
  NAND2_X1 U8775 ( .A1(n12856), .A2(n6745), .ZN(n12783) );
  NAND2_X1 U8776 ( .A1(n11503), .A2(n6746), .ZN(n6745) );
  INV_X1 U8777 ( .A(n11504), .ZN(n6746) );
  AOI21_X1 U8778 ( .B1(n7113), .B2(n7115), .A(n7112), .ZN(n7111) );
  NOR2_X1 U8779 ( .A1(n11720), .A2(n11719), .ZN(n7112) );
  OAI21_X1 U8780 ( .B1(n12783), .B2(n7103), .A(n7100), .ZN(n12791) );
  NAND2_X1 U8781 ( .A1(n11674), .A2(n11673), .ZN(n13282) );
  NAND2_X1 U8782 ( .A1(n9769), .A2(n6486), .ZN(n9557) );
  NAND2_X1 U8783 ( .A1(n7494), .A2(n12829), .ZN(n12818) );
  OR2_X1 U8784 ( .A1(n9560), .A2(n9559), .ZN(n7494) );
  OAI211_X1 U8785 ( .C1(n11574), .C2(n6488), .A(n7088), .B(n7087), .ZN(n12839)
         );
  INV_X1 U8786 ( .A(n7089), .ZN(n7088) );
  OAI21_X1 U8787 ( .B1(n11573), .B2(n6488), .A(n7483), .ZN(n7089) );
  NAND2_X1 U8788 ( .A1(n11662), .A2(n11661), .ZN(n12837) );
  NAND2_X1 U8789 ( .A1(n7092), .A2(n7091), .ZN(n11661) );
  XNOR2_X1 U8790 ( .A(n12825), .B(n9554), .ZN(n9330) );
  NAND2_X1 U8791 ( .A1(n7472), .A2(n8992), .ZN(n9329) );
  INV_X1 U8792 ( .A(n9560), .ZN(n12832) );
  NAND2_X1 U8793 ( .A1(n7470), .A2(n9677), .ZN(n10171) );
  NAND2_X1 U8794 ( .A1(n9763), .A2(n9658), .ZN(n7470) );
  NAND2_X1 U8795 ( .A1(n9660), .A2(n9659), .ZN(n14860) );
  NAND2_X1 U8796 ( .A1(n10329), .A2(n11951), .ZN(n9660) );
  INV_X1 U8797 ( .A(n13241), .ZN(n8915) );
  NAND2_X1 U8798 ( .A1(n12898), .A2(n13244), .ZN(n13241) );
  AND2_X1 U8799 ( .A1(n8923), .A2(n12038), .ZN(n12871) );
  NAND2_X1 U8800 ( .A1(n7489), .A2(n12781), .ZN(n12846) );
  INV_X1 U8801 ( .A(n7503), .ZN(n7505) );
  XNOR2_X1 U8802 ( .A(n11570), .B(n11571), .ZN(n11566) );
  OR2_X1 U8803 ( .A1(n12877), .A2(n11702), .ZN(n12828) );
  INV_X1 U8804 ( .A(n6753), .ZN(n10265) );
  NAND2_X1 U8805 ( .A1(n11502), .A2(n7490), .ZN(n12856) );
  NOR2_X1 U8806 ( .A1(n12854), .A2(n7491), .ZN(n7490) );
  INV_X1 U8807 ( .A(n11501), .ZN(n7491) );
  NAND2_X1 U8808 ( .A1(n11502), .A2(n11501), .ZN(n12855) );
  NAND2_X1 U8809 ( .A1(n7493), .A2(n7495), .ZN(n9564) );
  AND2_X1 U8810 ( .A1(n7486), .A2(n7484), .ZN(n12867) );
  NAND2_X1 U8811 ( .A1(n7486), .A2(n11687), .ZN(n12866) );
  NOR2_X1 U8812 ( .A1(n11650), .A2(n11188), .ZN(n11659) );
  NAND2_X1 U8813 ( .A1(n8947), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12873) );
  NAND4_X1 U8814 ( .A1(n9342), .A2(n9341), .A3(n9340), .A4(n9339), .ZN(n12893)
         );
  NAND2_X1 U8815 ( .A1(n8982), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8958) );
  OAI22_X1 U8816 ( .A1(n11726), .A2(n14891), .B1(n8956), .B2(n10041), .ZN(
        n6930) );
  CLKBUF_X1 U8817 ( .A(n11768), .Z(n12897) );
  OAI22_X1 U8818 ( .A1(n8782), .A2(n6833), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        P2_IR_REG_3__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U8819 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6833) );
  NOR2_X1 U8820 ( .A1(n8736), .A2(n8735), .ZN(n8734) );
  AND2_X1 U8821 ( .A1(n6824), .A2(n6823), .ZN(n9027) );
  NAND2_X1 U8822 ( .A1(n8765), .A2(n8764), .ZN(n6824) );
  INV_X1 U8823 ( .A(n8763), .ZN(n6823) );
  OAI21_X1 U8824 ( .B1(n8725), .B2(n8701), .A(n8700), .ZN(n8765) );
  INV_X1 U8825 ( .A(n6827), .ZN(n9248) );
  AOI21_X1 U8826 ( .B1(n9387), .B2(n9386), .A(n9385), .ZN(n12931) );
  NAND2_X1 U8827 ( .A1(n9251), .A2(n9250), .ZN(n9387) );
  AOI21_X1 U8828 ( .B1(n12933), .B2(n12932), .A(n12931), .ZN(n14740) );
  XNOR2_X1 U8829 ( .A(n12937), .B(n14752), .ZN(n14756) );
  NAND2_X1 U8830 ( .A1(n14756), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14755) );
  NAND2_X1 U8831 ( .A1(n14774), .A2(n6639), .ZN(n14794) );
  XNOR2_X1 U8832 ( .A(n12967), .B(n12972), .ZN(n12946) );
  NOR2_X1 U8833 ( .A1(n12946), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n12969) );
  OAI21_X1 U8834 ( .B1(n12978), .B2(n14733), .A(n6836), .ZN(n6835) );
  NAND2_X1 U8835 ( .A1(n12979), .A2(n14785), .ZN(n6836) );
  XNOR2_X1 U8836 ( .A(n13046), .B(n13045), .ZN(n13261) );
  AND2_X1 U8837 ( .A1(n13267), .A2(n13043), .ZN(n6925) );
  NAND2_X1 U8838 ( .A1(n7510), .A2(n6981), .ZN(n6980) );
  INV_X1 U8839 ( .A(n13061), .ZN(n13062) );
  AOI21_X1 U8840 ( .B1(n13071), .B2(n13251), .A(n13070), .ZN(n13273) );
  NAND2_X1 U8841 ( .A1(n13116), .A2(n7677), .ZN(n13099) );
  NAND2_X1 U8842 ( .A1(n13132), .A2(n13007), .ZN(n13110) );
  NAND2_X1 U8843 ( .A1(n7440), .A2(n7443), .ZN(n13130) );
  NAND2_X1 U8844 ( .A1(n11545), .A2(n11544), .ZN(n13157) );
  NAND2_X1 U8845 ( .A1(n7449), .A2(n7452), .ZN(n13149) );
  NAND2_X1 U8846 ( .A1(n7450), .A2(n13163), .ZN(n7449) );
  INV_X1 U8847 ( .A(n7450), .ZN(n13162) );
  NAND2_X1 U8848 ( .A1(n7475), .A2(n7477), .ZN(n13179) );
  OR2_X1 U8849 ( .A1(n13208), .A2(n7480), .ZN(n7475) );
  NAND2_X1 U8850 ( .A1(n11505), .A2(n6486), .ZN(n11509) );
  AND2_X1 U8851 ( .A1(n7481), .A2(n6492), .ZN(n13191) );
  NAND2_X1 U8852 ( .A1(n13208), .A2(n13001), .ZN(n7481) );
  AND2_X1 U8853 ( .A1(n13220), .A2(n7455), .ZN(n13205) );
  NAND2_X1 U8854 ( .A1(n13220), .A2(n7674), .ZN(n13206) );
  INV_X1 U8855 ( .A(n6905), .ZN(n13222) );
  CLKBUF_X1 U8856 ( .A(n10880), .Z(n10840) );
  NAND2_X1 U8857 ( .A1(n10926), .A2(n6486), .ZN(n10834) );
  NAND2_X1 U8858 ( .A1(n10704), .A2(n6486), .ZN(n10466) );
  NAND2_X1 U8859 ( .A1(n6907), .A2(n10521), .ZN(n10683) );
  NAND2_X1 U8860 ( .A1(n7516), .A2(n7520), .ZN(n10675) );
  OR2_X1 U8861 ( .A1(n10450), .A2(n7521), .ZN(n7516) );
  NAND2_X1 U8862 ( .A1(n7524), .A2(n7526), .ZN(n10522) );
  OR2_X1 U8863 ( .A1(n10450), .A2(n12014), .ZN(n7524) );
  NAND2_X1 U8864 ( .A1(n10174), .A2(n10173), .ZN(n11837) );
  NAND2_X1 U8865 ( .A1(n10335), .A2(n6486), .ZN(n10174) );
  NAND2_X1 U8866 ( .A1(n9976), .A2(n11951), .ZN(n9645) );
  NAND2_X1 U8867 ( .A1(n7460), .A2(n7461), .ZN(n9921) );
  NAND2_X1 U8868 ( .A1(n13155), .A2(n9736), .ZN(n13231) );
  INV_X1 U8869 ( .A(n13245), .ZN(n13159) );
  CLKBUF_X1 U8870 ( .A(n9413), .Z(n11781) );
  INV_X1 U8871 ( .A(n13231), .ZN(n13248) );
  AND2_X1 U8872 ( .A1(n13155), .A2(n8963), .ZN(n13245) );
  AND2_X1 U8873 ( .A1(n13155), .A2(n9807), .ZN(n13246) );
  AND2_X2 U8874 ( .A1(n9432), .A2(n9431), .ZN(n14908) );
  NAND2_X1 U8875 ( .A1(n6793), .A2(n6791), .ZN(n13340) );
  NOR2_X1 U8876 ( .A1(n13022), .A2(n6792), .ZN(n6791) );
  NAND2_X1 U8877 ( .A1(n13261), .A2(n14850), .ZN(n6793) );
  INV_X1 U8878 ( .A(n13264), .ZN(n6792) );
  AND2_X2 U8879 ( .A1(n9432), .A2(n14802), .ZN(n14887) );
  AND2_X1 U8880 ( .A1(n8920), .A2(n8891), .ZN(n14805) );
  INV_X1 U8881 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U8882 ( .A1(n13355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6794) );
  NAND2_X1 U8883 ( .A1(n6864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6863) );
  NOR2_X1 U8884 ( .A1(n8616), .A2(n7015), .ZN(n7014) );
  NAND2_X1 U8885 ( .A1(n7466), .A2(n7011), .ZN(n7016) );
  NOR2_X1 U8886 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7015) );
  XNOR2_X1 U8887 ( .A(n8407), .B(n8405), .ZN(n10442) );
  NAND2_X1 U8888 ( .A1(n8420), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8405) );
  XNOR2_X1 U8889 ( .A(n8896), .B(n8895), .ZN(n9685) );
  INV_X1 U8890 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9214) );
  INV_X1 U8891 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9022) );
  INV_X1 U8892 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8697) );
  INV_X1 U8893 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8677) );
  INV_X1 U8894 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8610) );
  INV_X1 U8895 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8590) );
  INV_X1 U8896 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8567) );
  INV_X1 U8897 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n8562) );
  INV_X1 U8898 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8574) );
  INV_X1 U8899 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9326) );
  INV_X1 U8900 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U8901 ( .A1(n8458), .A2(n8546), .ZN(n8967) );
  NAND2_X1 U8902 ( .A1(n10160), .A2(n10159), .ZN(n10384) );
  XNOR2_X1 U8903 ( .A(n6673), .B(n13370), .ZN(n13371) );
  NAND2_X1 U8904 ( .A1(n13477), .A2(n11442), .ZN(n6673) );
  NAND2_X1 U8905 ( .A1(n6522), .A2(n7332), .ZN(n7331) );
  INV_X1 U8906 ( .A(n7333), .ZN(n7332) );
  NAND2_X1 U8907 ( .A1(n6670), .A2(n10645), .ZN(n14408) );
  NAND2_X1 U8908 ( .A1(n10641), .A2(n10640), .ZN(n6670) );
  NAND2_X1 U8909 ( .A1(n9573), .A2(n9572), .ZN(n13388) );
  NAND2_X1 U8910 ( .A1(n10384), .A2(n10383), .ZN(n10386) );
  INV_X1 U8911 ( .A(n10110), .ZN(n6668) );
  NOR2_X1 U8912 ( .A1(n10919), .A2(n10920), .ZN(n11239) );
  NAND2_X1 U8913 ( .A1(n9788), .A2(n9787), .ZN(n9902) );
  NAND2_X1 U8914 ( .A1(n7326), .A2(n7324), .ZN(n14396) );
  NAND2_X1 U8915 ( .A1(n7305), .A2(n7303), .ZN(n13430) );
  NAND2_X1 U8916 ( .A1(n7307), .A2(n7306), .ZN(n7305) );
  INV_X1 U8917 ( .A(n13456), .ZN(n7307) );
  OR2_X1 U8918 ( .A1(n9125), .A2(n9124), .ZN(n13462) );
  NAND2_X1 U8919 ( .A1(n13398), .A2(n6617), .ZN(n13438) );
  NAND2_X1 U8920 ( .A1(n10919), .A2(n7334), .ZN(n7330) );
  NOR2_X1 U8921 ( .A1(n11239), .A2(n7335), .ZN(n13450) );
  AOI21_X1 U8922 ( .B1(n13456), .B2(n13455), .A(n13454), .ZN(n13458) );
  OR3_X1 U8923 ( .A1(n9125), .A2(n9127), .A3(n14701), .ZN(n14410) );
  NAND2_X1 U8924 ( .A1(n7321), .A2(n14394), .ZN(n13468) );
  NAND2_X1 U8925 ( .A1(n7326), .A2(n6490), .ZN(n7321) );
  INV_X1 U8926 ( .A(n7285), .ZN(n7284) );
  INV_X1 U8927 ( .A(n9901), .ZN(n7286) );
  AND4_X1 U8928 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n14428) );
  NOR2_X1 U8929 ( .A1(n13710), .A2(n13709), .ZN(n6964) );
  INV_X1 U8930 ( .A(n13714), .ZN(n6945) );
  OR2_X1 U8931 ( .A1(n9122), .A2(n10949), .ZN(n13721) );
  OR2_X1 U8932 ( .A1(n13638), .A2(n10119), .ZN(n9075) );
  INV_X1 U8933 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n10809) );
  XNOR2_X1 U8934 ( .A(n13810), .B(n14040), .ZN(n13804) );
  NAND2_X1 U8935 ( .A1(n13637), .A2(n13636), .ZN(n13815) );
  NOR2_X1 U8936 ( .A1(n13830), .A2(n13372), .ZN(n7003) );
  INV_X1 U8937 ( .A(n13819), .ZN(n7004) );
  XNOR2_X1 U8938 ( .A(n6852), .B(n6851), .ZN(n14056) );
  INV_X1 U8939 ( .A(n13696), .ZN(n6851) );
  NAND2_X1 U8940 ( .A1(n13829), .A2(n6536), .ZN(n6852) );
  INV_X1 U8941 ( .A(n13822), .ZN(n13823) );
  INV_X1 U8942 ( .A(n13618), .ZN(n14066) );
  INV_X1 U8943 ( .A(n13842), .ZN(n13846) );
  INV_X1 U8944 ( .A(n13877), .ZN(n13887) );
  NAND2_X1 U8945 ( .A1(n7263), .A2(n7262), .ZN(n13886) );
  AND2_X1 U8946 ( .A1(n7263), .A2(n6516), .ZN(n13888) );
  NAND2_X1 U8947 ( .A1(n7235), .A2(n7238), .ZN(n13931) );
  NAND2_X1 U8948 ( .A1(n7382), .A2(n7386), .ZN(n13934) );
  NAND2_X1 U8949 ( .A1(n13960), .A2(n7388), .ZN(n7382) );
  NAND2_X1 U8950 ( .A1(n13960), .A2(n11620), .ZN(n13954) );
  NAND2_X1 U8951 ( .A1(n13964), .A2(n11603), .ZN(n13945) );
  NAND2_X1 U8952 ( .A1(n7244), .A2(n7248), .ZN(n13988) );
  NAND2_X1 U8953 ( .A1(n14007), .A2(n7251), .ZN(n7244) );
  NAND2_X1 U8954 ( .A1(n11617), .A2(n11616), .ZN(n13978) );
  NAND2_X1 U8955 ( .A1(n7253), .A2(n13669), .ZN(n13991) );
  NAND2_X1 U8956 ( .A1(n7254), .A2(n13670), .ZN(n7253) );
  INV_X1 U8957 ( .A(n14007), .ZN(n7254) );
  NAND2_X1 U8958 ( .A1(n7395), .A2(n7401), .ZN(n14005) );
  NAND2_X1 U8959 ( .A1(n11614), .A2(n7402), .ZN(n7395) );
  NAND2_X1 U8960 ( .A1(n7403), .A2(n7402), .ZN(n14020) );
  NAND2_X1 U8961 ( .A1(n7403), .A2(n13562), .ZN(n14018) );
  NAND2_X1 U8962 ( .A1(n10773), .A2(n10702), .ZN(n10924) );
  NAND2_X1 U8963 ( .A1(n10707), .A2(n10706), .ZN(n14445) );
  NAND2_X1 U8964 ( .A1(n10762), .A2(n10719), .ZN(n10930) );
  AND2_X1 U8965 ( .A1(n7405), .A2(n7408), .ZN(n10611) );
  NAND2_X1 U8966 ( .A1(n10610), .A2(n10609), .ZN(n13538) );
  NAND2_X1 U8967 ( .A1(n10551), .A2(n10550), .ZN(n10606) );
  NAND2_X1 U8968 ( .A1(n7221), .A2(n10334), .ZN(n10553) );
  NAND2_X1 U8969 ( .A1(n14562), .A2(n10333), .ZN(n7221) );
  NAND2_X1 U8970 ( .A1(n10332), .A2(n10331), .ZN(n14570) );
  NAND2_X1 U8971 ( .A1(n7412), .A2(n7411), .ZN(n10349) );
  NAND2_X1 U8972 ( .A1(n7226), .A2(n9832), .ZN(n9969) );
  NAND2_X1 U8973 ( .A1(n10087), .A2(n10093), .ZN(n7226) );
  INV_X1 U8974 ( .A(n14609), .ZN(n14035) );
  NAND2_X1 U8975 ( .A1(n6464), .A2(n14613), .ZN(n13982) );
  AND2_X1 U8976 ( .A1(n14042), .A2(n14041), .ZN(n14156) );
  INV_X1 U8977 ( .A(n13815), .ZN(n14163) );
  NAND2_X1 U8978 ( .A1(n11421), .A2(n11420), .ZN(n14174) );
  AND2_X1 U8979 ( .A1(n11304), .A2(n11303), .ZN(n14196) );
  AND2_X1 U8980 ( .A1(n11286), .A2(n11285), .ZN(n14201) );
  INV_X1 U8981 ( .A(n13538), .ZN(n10819) );
  INV_X1 U8982 ( .A(n13515), .ZN(n10147) );
  INV_X2 U8983 ( .A(n14713), .ZN(n14714) );
  NAND2_X1 U8984 ( .A1(n9046), .A2(n9048), .ZN(n14213) );
  OAI21_X1 U8985 ( .B1(n11922), .B2(n11921), .A(n11920), .ZN(n11925) );
  NOR2_X1 U8986 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7228) );
  NOR2_X1 U8987 ( .A1(n9045), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n6672) );
  INV_X1 U8988 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U8989 ( .A1(n8447), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8445) );
  OAI21_X1 U8990 ( .B1(n11333), .B2(n7609), .A(n10256), .ZN(n10440) );
  XNOR2_X1 U8991 ( .A(n11334), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14224) );
  OR2_X1 U8992 ( .A1(n11333), .A2(n11332), .ZN(n11334) );
  NAND2_X1 U8993 ( .A1(n6937), .A2(n6939), .ZN(n6936) );
  OR2_X1 U8994 ( .A1(n8751), .A2(n6939), .ZN(n6938) );
  XNOR2_X1 U8995 ( .A(n9043), .B(n9042), .ZN(n13656) );
  NOR2_X1 U8996 ( .A1(n8437), .A2(n6976), .ZN(n6975) );
  NAND2_X1 U8997 ( .A1(n9473), .A2(n6702), .ZN(n6977) );
  NOR2_X1 U8998 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6976) );
  INV_X1 U8999 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9199) );
  INV_X1 U9000 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9013) );
  INV_X1 U9001 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9026) );
  INV_X1 U9002 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10697) );
  INV_X1 U9003 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8790) );
  INV_X1 U9004 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8717) );
  INV_X1 U9005 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8681) );
  INV_X1 U9006 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8605) );
  INV_X1 U9007 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8593) );
  INV_X1 U9008 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U9009 ( .A1(n6737), .A2(n14289), .ZN(n14335) );
  NAND2_X1 U9010 ( .A1(n15389), .A2(n15390), .ZN(n6737) );
  NOR2_X1 U9011 ( .A1(n14335), .A2(n14334), .ZN(n14333) );
  XNOR2_X1 U9012 ( .A(n14303), .B(n7269), .ZN(n14339) );
  INV_X1 U9013 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7269) );
  XNOR2_X1 U9014 ( .A(n14308), .B(n7267), .ZN(n15386) );
  INV_X1 U9015 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7267) );
  NAND2_X1 U9016 ( .A1(n7264), .A2(n14315), .ZN(n14343) );
  NOR2_X1 U9017 ( .A1(n14472), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U9018 ( .A1(n7058), .A2(n6741), .ZN(n14486) );
  NAND2_X1 U9019 ( .A1(n14482), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7058) );
  OR2_X1 U9020 ( .A1(n14327), .A2(n14328), .ZN(n14492) );
  NAND2_X1 U9021 ( .A1(n14492), .A2(n14493), .ZN(n14489) );
  NAND2_X1 U9022 ( .A1(n14346), .A2(n14348), .ZN(n15182) );
  OAI21_X1 U9023 ( .B1(n12719), .B2(n12214), .A(n8380), .ZN(n8381) );
  AOI21_X1 U9024 ( .B1(n14913), .B2(n14912), .A(n7160), .ZN(n14917) );
  INV_X1 U9025 ( .A(n7069), .ZN(n9869) );
  INV_X1 U9026 ( .A(n7034), .ZN(n12377) );
  NAND2_X1 U9027 ( .A1(n7164), .A2(n6818), .ZN(P3_U3200) );
  OR2_X1 U9028 ( .A1(n12381), .A2(n14990), .ZN(n7164) );
  NOR2_X1 U9029 ( .A1(n6820), .A2(n6819), .ZN(n6818) );
  INV_X1 U9030 ( .A(n6913), .ZN(n6912) );
  INV_X1 U9031 ( .A(n6960), .ZN(n6959) );
  OAI22_X1 U9032 ( .A1(n12716), .A2(n12705), .B1(n15181), .B2(n12643), .ZN(
        n6960) );
  OAI21_X1 U9033 ( .B1(n12717), .B2(n6961), .A(n6620), .ZN(P3_U3486) );
  OR2_X1 U9034 ( .A1(n15181), .A2(n12647), .ZN(n6985) );
  NAND2_X1 U9035 ( .A1(n12444), .A2(n7570), .ZN(n7008) );
  INV_X1 U9036 ( .A(n6963), .ZN(n6962) );
  OAI22_X1 U9037 ( .A1(n12716), .A2(n12757), .B1(n15164), .B2(n12715), .ZN(
        n6963) );
  AOI21_X1 U9038 ( .B1(n12444), .B2(n8273), .A(n7006), .ZN(n7005) );
  NOR2_X1 U9039 ( .A1(n15164), .A2(n12718), .ZN(n7006) );
  NAND2_X1 U9040 ( .A1(n6920), .A2(n6918), .ZN(P2_U3233) );
  AOI21_X1 U9041 ( .B1(n6835), .B2(n8963), .A(n6919), .ZN(n6918) );
  OR2_X1 U9042 ( .A1(n12980), .A2(n8963), .ZN(n6920) );
  OAI21_X1 U9043 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n12982), .A(n12981), .ZN(
        n6919) );
  NAND2_X1 U9044 ( .A1(n13341), .A2(n14887), .ZN(n6890) );
  NAND2_X1 U9045 ( .A1(n14420), .A2(n6511), .ZN(n14385) );
  INV_X1 U9046 ( .A(n6909), .ZN(n6908) );
  OAI22_X1 U9047 ( .A1(n14168), .A2(n14155), .B1(n14062), .B2(n14730), .ZN(
        n6909) );
  NAND2_X1 U9048 ( .A1(n6729), .A2(n6731), .ZN(n15383) );
  NAND2_X1 U9049 ( .A1(n6726), .A2(n6725), .ZN(n14340) );
  NOR2_X1 U9050 ( .A1(n14469), .A2(n14470), .ZN(n14468) );
  NOR2_X1 U9051 ( .A1(n14482), .A2(n14481), .ZN(n14480) );
  INV_X1 U9052 ( .A(n14348), .ZN(n14347) );
  XNOR2_X1 U9053 ( .A(n6739), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  OR2_X1 U9054 ( .A1(n6740), .A2(n7065), .ZN(n6739) );
  AND2_X1 U9055 ( .A1(n15182), .A2(n15183), .ZN(n6740) );
  XNOR2_X1 U9056 ( .A(n6531), .B(n15186), .ZN(n7272) );
  NAND2_X1 U9057 ( .A1(n7275), .A2(n7274), .ZN(n7273) );
  INV_X1 U9058 ( .A(n6510), .ZN(n11938) );
  NAND2_X1 U9059 ( .A1(n6574), .A2(n14420), .ZN(n7326) );
  AND4_X1 U9060 ( .A1(n8403), .A2(n8402), .A3(n8892), .A4(n8406), .ZN(n6483)
         );
  AND4_X1 U9061 ( .A1(n7712), .A2(n6496), .A3(n7671), .A4(n7573), .ZN(n6484)
         );
  AND2_X1 U9062 ( .A1(n13619), .A2(n7536), .ZN(n6485) );
  AND2_X1 U9063 ( .A1(n13377), .A2(n7313), .ZN(n6487) );
  INV_X1 U9064 ( .A(n6479), .ZN(n8142) );
  INV_X1 U9065 ( .A(n13987), .ZN(n7246) );
  INV_X1 U9066 ( .A(n13683), .ZN(n7220) );
  AND2_X1 U9067 ( .A1(n11660), .A2(n7090), .ZN(n6488) );
  AND2_X1 U9068 ( .A1(n7724), .A2(n7723), .ZN(n7797) );
  OR2_X1 U9069 ( .A1(n11851), .A2(n11853), .ZN(n6489) );
  INV_X1 U9070 ( .A(n15071), .ZN(n12232) );
  AND2_X1 U9071 ( .A1(n7962), .A2(n7706), .ZN(n7964) );
  INV_X1 U9072 ( .A(n13173), .ZN(n13304) );
  AND2_X1 U9073 ( .A1(n11532), .A2(n11531), .ZN(n13173) );
  XNOR2_X1 U9074 ( .A(n7134), .B(P3_IR_REG_27__SCAN_IN), .ZN(n12397) );
  INV_X1 U9075 ( .A(n12234), .ZN(n7018) );
  INV_X1 U9076 ( .A(n14390), .ZN(n14205) );
  AND2_X1 U9077 ( .A1(n7324), .A2(n6629), .ZN(n6490) );
  INV_X1 U9078 ( .A(n7480), .ZN(n7479) );
  NAND2_X1 U9079 ( .A1(n6578), .A2(n6492), .ZN(n7480) );
  AND2_X1 U9080 ( .A1(n12499), .A2(n11069), .ZN(n6491) );
  NAND2_X1 U9081 ( .A1(n13213), .A2(n13000), .ZN(n6492) );
  OR4_X1 U9082 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(n6493) );
  AND2_X1 U9083 ( .A1(n13260), .A2(n7144), .ZN(n6494) );
  INV_X1 U9084 ( .A(n10632), .ZN(n8267) );
  NAND2_X1 U9085 ( .A1(n6693), .A2(n6691), .ZN(n10632) );
  AND2_X1 U9086 ( .A1(n11914), .A2(n11915), .ZN(n6495) );
  NAND2_X1 U9087 ( .A1(n10834), .A2(n10833), .ZN(n13331) );
  INV_X1 U9088 ( .A(n11860), .ZN(n10685) );
  INV_X1 U9089 ( .A(n7387), .ZN(n7386) );
  NOR2_X1 U9090 ( .A1(n13944), .A2(n11622), .ZN(n7387) );
  AND2_X1 U9091 ( .A1(n11578), .A2(n11577), .ZN(n12983) );
  INV_X1 U9092 ( .A(n12983), .ZN(n13292) );
  NAND2_X1 U9093 ( .A1(n10180), .A2(n10179), .ZN(n14878) );
  OR2_X1 U9094 ( .A1(n13523), .A2(n13524), .ZN(n6497) );
  AND3_X1 U9095 ( .A1(n8907), .A2(n8908), .A3(n8909), .ZN(n6498) );
  INV_X1 U9096 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7716) );
  AND2_X1 U9097 ( .A1(n7568), .A2(n6961), .ZN(n6499) );
  AND2_X1 U9098 ( .A1(n11509), .A2(n11508), .ZN(n13202) );
  INV_X1 U9099 ( .A(n13202), .ZN(n7148) );
  AND2_X1 U9100 ( .A1(n6579), .A2(n6684), .ZN(n6500) );
  OR2_X1 U9101 ( .A1(n11815), .A2(n11814), .ZN(n6501) );
  AND2_X1 U9102 ( .A1(n7148), .A2(n13002), .ZN(n6502) );
  NOR2_X1 U9103 ( .A1(n12710), .A2(n12407), .ZN(n11151) );
  INV_X1 U9104 ( .A(n11151), .ZN(n7196) );
  INV_X1 U9105 ( .A(n11660), .ZN(n7091) );
  NAND2_X1 U9106 ( .A1(n10878), .A2(n10877), .ZN(n13328) );
  INV_X1 U9107 ( .A(n13328), .ZN(n7498) );
  NOR2_X1 U9108 ( .A1(n11889), .A2(n11888), .ZN(n6503) );
  AND2_X1 U9109 ( .A1(n7652), .A2(n7651), .ZN(n6504) );
  INV_X1 U9110 ( .A(n12444), .ZN(n12719) );
  NAND2_X1 U9111 ( .A1(n8178), .A2(n8177), .ZN(n12444) );
  AND2_X1 U9112 ( .A1(n7083), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6505) );
  AND2_X1 U9113 ( .A1(n8274), .A2(n6630), .ZN(n6506) );
  AND2_X1 U9114 ( .A1(n7049), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U9115 ( .A1(n8916), .A2(n9685), .ZN(n9459) );
  AND2_X1 U9116 ( .A1(n7493), .A2(n6637), .ZN(n6508) );
  NAND2_X1 U9117 ( .A1(n8267), .A2(n6690), .ZN(n8639) );
  OR2_X1 U9118 ( .A1(n8945), .A2(SI_24_), .ZN(n6509) );
  NOR2_X1 U9119 ( .A1(n12253), .A2(n12237), .ZN(n7076) );
  INV_X1 U9120 ( .A(n7076), .ZN(n7075) );
  OR2_X1 U9121 ( .A1(n11757), .A2(n12042), .ZN(n6510) );
  NAND2_X1 U9122 ( .A1(n8149), .A2(n8148), .ZN(n12653) );
  OR2_X1 U9123 ( .A1(n11257), .A2(n11256), .ZN(n6511) );
  NAND2_X1 U9124 ( .A1(n8018), .A2(n8017), .ZN(n8020) );
  AND4_X1 U9125 ( .A1(n7857), .A2(n7856), .A3(n7855), .A4(n7854), .ZN(n15055)
         );
  INV_X1 U9126 ( .A(n14578), .ZN(n14576) );
  OR2_X1 U9127 ( .A1(n7978), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n6512) );
  INV_X1 U9128 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U9129 ( .A1(n8163), .A2(n8162), .ZN(n12648) );
  NAND2_X1 U9130 ( .A1(n11933), .A2(n11932), .ZN(n13263) );
  OR2_X1 U9131 ( .A1(n8750), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6513) );
  NOR2_X1 U9132 ( .A1(n10479), .A2(n10478), .ZN(n6514) );
  XNOR2_X1 U9133 ( .A(n7862), .B(P3_IR_REG_5__SCAN_IN), .ZN(n14940) );
  INV_X1 U9134 ( .A(n14940), .ZN(n6662) );
  NAND2_X1 U9135 ( .A1(n11447), .A2(n11446), .ZN(n13618) );
  OR2_X1 U9136 ( .A1(n10571), .A2(n10570), .ZN(n6515) );
  OR2_X1 U9137 ( .A1(n13903), .A2(n13924), .ZN(n6516) );
  INV_X1 U9138 ( .A(n6958), .ZN(n15074) );
  AND2_X1 U9139 ( .A1(n7416), .A2(n7414), .ZN(n6517) );
  XNOR2_X1 U9140 ( .A(n8618), .B(P2_IR_REG_22__SCAN_IN), .ZN(n12042) );
  OR2_X1 U9141 ( .A1(n14956), .A2(n9883), .ZN(n6518) );
  AOI21_X1 U9142 ( .B1(n7455), .B2(n7454), .A(n7457), .ZN(n7453) );
  AND2_X1 U9143 ( .A1(n14322), .A2(n14478), .ZN(n6519) );
  NOR2_X1 U9144 ( .A1(n13618), .A2(n13820), .ZN(n6520) );
  INV_X1 U9145 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8555) );
  AND2_X1 U9146 ( .A1(n13287), .A2(n13036), .ZN(n6521) );
  NOR2_X1 U9147 ( .A1(n14376), .A2(n14377), .ZN(n6522) );
  AND2_X1 U9148 ( .A1(n6723), .A2(n6725), .ZN(n6523) );
  AND2_X1 U9149 ( .A1(n11826), .A2(n9958), .ZN(n6524) );
  OR2_X1 U9150 ( .A1(n12331), .A2(n12317), .ZN(n6525) );
  OR2_X1 U9151 ( .A1(n12331), .A2(n12330), .ZN(n6526) );
  OR2_X1 U9152 ( .A1(n12251), .A2(n12241), .ZN(n6527) );
  INV_X1 U9153 ( .A(n10032), .ZN(n7021) );
  AND2_X1 U9154 ( .A1(n7810), .A2(n7808), .ZN(n6528) );
  NAND2_X1 U9155 ( .A1(n14585), .A2(n10390), .ZN(n6529) );
  OAI211_X1 U9156 ( .C1(n9140), .C2(n9365), .A(n7796), .B(n7795), .ZN(n15101)
         );
  INV_X1 U9157 ( .A(n15101), .ZN(n7430) );
  NAND2_X1 U9158 ( .A1(n11196), .A2(n11195), .ZN(n13323) );
  INV_X1 U9159 ( .A(n13323), .ZN(n7150) );
  INV_X1 U9160 ( .A(n7239), .ZN(n7238) );
  OAI22_X1 U9161 ( .A1(n13944), .A2(n7240), .B1(n13950), .B2(n13718), .ZN(
        n7239) );
  OR2_X1 U9162 ( .A1(n13593), .A2(n13594), .ZN(n6530) );
  INV_X1 U9163 ( .A(n15082), .ZN(n6657) );
  NAND2_X1 U9164 ( .A1(n8145), .A2(n8144), .ZN(n12469) );
  INV_X1 U9165 ( .A(n12469), .ZN(n7366) );
  XNOR2_X1 U9166 ( .A(n15380), .B(n15379), .ZN(n6531) );
  AND2_X1 U9167 ( .A1(n11506), .A2(n12905), .ZN(n6532) );
  NAND2_X1 U9168 ( .A1(n8946), .A2(n7146), .ZN(n11786) );
  AND2_X1 U9169 ( .A1(n12642), .A2(n15160), .ZN(n6533) );
  NAND2_X1 U9170 ( .A1(n11666), .A2(n11665), .ZN(n13287) );
  INV_X1 U9171 ( .A(n11812), .ZN(n14841) );
  INV_X1 U9172 ( .A(n15044), .ZN(n10659) );
  INV_X1 U9173 ( .A(n13912), .ZN(n13914) );
  INV_X1 U9174 ( .A(n13684), .ZN(n10717) );
  OR2_X1 U9175 ( .A1(n7978), .A2(n8201), .ZN(n6534) );
  AND2_X1 U9176 ( .A1(n7100), .A2(n7099), .ZN(n6535) );
  XNOR2_X1 U9177 ( .A(n13903), .B(n13924), .ZN(n13897) );
  INV_X1 U9178 ( .A(n8221), .ZN(n7567) );
  OR2_X1 U9179 ( .A1(n14168), .A2(n13372), .ZN(n6536) );
  NAND2_X1 U9180 ( .A1(n13102), .A2(n6795), .ZN(n6796) );
  NAND2_X1 U9181 ( .A1(n10549), .A2(n10548), .ZN(n14416) );
  OR2_X1 U9182 ( .A1(n7844), .A2(n6655), .ZN(n6654) );
  INV_X1 U9183 ( .A(n6654), .ZN(n7962) );
  AND2_X1 U9184 ( .A1(n14445), .A2(n14147), .ZN(n6537) );
  AND2_X1 U9185 ( .A1(n12560), .A2(n11041), .ZN(n12587) );
  INV_X1 U9186 ( .A(n12587), .ZN(n6644) );
  NAND2_X1 U9187 ( .A1(n11613), .A2(n11612), .ZN(n13629) );
  INV_X1 U9188 ( .A(n13629), .ZN(n7198) );
  MUX2_X2 U9189 ( .A(n13664), .B(n13665), .S(n13643), .Z(n13520) );
  NOR2_X1 U9190 ( .A1(n11335), .A2(n13736), .ZN(n6538) );
  INV_X1 U9191 ( .A(n14311), .ZN(n6727) );
  INV_X1 U9192 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8021) );
  NAND3_X1 U9193 ( .A1(n9215), .A2(n8436), .A3(n8431), .ZN(n9041) );
  NOR2_X1 U9194 ( .A1(n10832), .A2(n6778), .ZN(n6539) );
  OR2_X1 U9195 ( .A1(n7536), .A2(n13619), .ZN(n6540) );
  OR2_X1 U9196 ( .A1(n10284), .A2(n12889), .ZN(n6541) );
  INV_X1 U9197 ( .A(n13318), .ZN(n13213) );
  NAND2_X1 U9198 ( .A1(n11497), .A2(n11496), .ZN(n13318) );
  AND2_X1 U9199 ( .A1(n8189), .A2(n8188), .ZN(n6542) );
  INV_X1 U9200 ( .A(n7209), .ZN(n13901) );
  NOR2_X1 U9201 ( .A1(n13902), .A2(n13903), .ZN(n7209) );
  AND2_X1 U9202 ( .A1(n14310), .A2(n6727), .ZN(n6543) );
  INV_X1 U9203 ( .A(n7485), .ZN(n7484) );
  NAND2_X1 U9204 ( .A1(n11705), .A2(n11687), .ZN(n7485) );
  INV_X1 U9205 ( .A(n13022), .ZN(n13265) );
  AND2_X1 U9206 ( .A1(n7091), .A2(n11580), .ZN(n6544) );
  AND2_X1 U9207 ( .A1(n9920), .A2(n7461), .ZN(n6545) );
  AND2_X1 U9208 ( .A1(n11691), .A2(n11690), .ZN(n13090) );
  INV_X1 U9209 ( .A(n13090), .ZN(n13276) );
  OR2_X1 U9210 ( .A1(n8334), .A2(n8333), .ZN(n6546) );
  INV_X1 U9211 ( .A(n13528), .ZN(n6685) );
  AND2_X1 U9212 ( .A1(n13552), .A2(n7537), .ZN(n6547) );
  INV_X1 U9213 ( .A(n7446), .ZN(n7445) );
  NAND2_X1 U9214 ( .A1(n13163), .A2(n7451), .ZN(n7446) );
  INV_X1 U9215 ( .A(n7308), .ZN(n7306) );
  NAND2_X1 U9216 ( .A1(n7315), .A2(n6487), .ZN(n7308) );
  NAND2_X1 U9217 ( .A1(n11185), .A2(n11184), .ZN(n6548) );
  NOR2_X1 U9218 ( .A1(n6495), .A2(n11916), .ZN(n6549) );
  OR2_X1 U9219 ( .A1(n12644), .A2(n12453), .ZN(n6550) );
  AND2_X1 U9220 ( .A1(n14390), .A2(n14425), .ZN(n6551) );
  AND2_X1 U9221 ( .A1(n7545), .A2(n13513), .ZN(n6552) );
  INV_X1 U9222 ( .A(n7182), .ZN(n7181) );
  AND2_X1 U9223 ( .A1(n8228), .A2(n11040), .ZN(n6553) );
  NAND2_X1 U9224 ( .A1(n9160), .A2(n9173), .ZN(n9159) );
  OR2_X1 U9225 ( .A1(n11156), .A2(n15103), .ZN(n6554) );
  AND2_X1 U9226 ( .A1(n7608), .A2(n7606), .ZN(n6555) );
  AND2_X1 U9227 ( .A1(n8895), .A2(n8408), .ZN(n6556) );
  AND2_X1 U9228 ( .A1(n12752), .A2(n12620), .ZN(n6557) );
  INV_X1 U9229 ( .A(n7044), .ZN(n7043) );
  NOR2_X1 U9230 ( .A1(n9881), .A2(n14956), .ZN(n7044) );
  INV_X1 U9231 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8415) );
  AND2_X1 U9232 ( .A1(n7105), .A2(n6548), .ZN(n6558) );
  AND2_X1 U9233 ( .A1(n11061), .A2(n11060), .ZN(n12524) );
  NOR2_X1 U9234 ( .A1(n13727), .A2(n13515), .ZN(n6559) );
  AND2_X1 U9235 ( .A1(n13116), .A2(n7465), .ZN(n6560) );
  AND2_X1 U9236 ( .A1(n7449), .A2(n7447), .ZN(n6561) );
  AND2_X1 U9237 ( .A1(n7419), .A2(n7417), .ZN(n6562) );
  INV_X1 U9238 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7669) );
  NOR2_X1 U9239 ( .A1(n13728), .A2(n14671), .ZN(n6563) );
  NOR2_X1 U9240 ( .A1(n12752), .A2(n12620), .ZN(n6564) );
  AND2_X1 U9241 ( .A1(n12501), .A2(n12479), .ZN(n6565) );
  AND2_X1 U9242 ( .A1(n8582), .A2(SI_7_), .ZN(n6566) );
  INV_X1 U9243 ( .A(n13256), .ZN(n7145) );
  AND2_X1 U9244 ( .A1(n8298), .A2(n8297), .ZN(n6567) );
  INV_X1 U9245 ( .A(n10247), .ZN(n12231) );
  AND4_X1 U9246 ( .A1(n7839), .A2(n7838), .A3(n7837), .A4(n7836), .ZN(n10247)
         );
  INV_X1 U9247 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7576) );
  INV_X1 U9248 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6937) );
  OR2_X1 U9249 ( .A1(n7492), .A2(n9642), .ZN(n6568) );
  NAND4_X1 U9250 ( .A1(n8431), .A2(n8436), .A3(n7390), .A4(n9215), .ZN(n6569)
         );
  AND2_X1 U9251 ( .A1(n13601), .A2(n13921), .ZN(n6570) );
  AND2_X1 U9252 ( .A1(n8673), .A2(SI_9_), .ZN(n6571) );
  AND2_X1 U9253 ( .A1(n13522), .A2(n13521), .ZN(n6572) );
  NAND2_X1 U9254 ( .A1(n14578), .A2(n10348), .ZN(n6573) );
  INV_X1 U9255 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8523) );
  INV_X1 U9256 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8614) );
  AND2_X1 U9257 ( .A1(n6511), .A2(n7328), .ZN(n6574) );
  INV_X1 U9258 ( .A(n7190), .ZN(n7189) );
  INV_X1 U9259 ( .A(n7418), .ZN(n7417) );
  NAND2_X1 U9260 ( .A1(n8331), .A2(n8329), .ZN(n7418) );
  INV_X1 U9261 ( .A(n7428), .ZN(n7427) );
  NAND2_X1 U9262 ( .A1(n7429), .A2(n8295), .ZN(n7428) );
  AND2_X1 U9263 ( .A1(n13528), .A2(n6686), .ZN(n6575) );
  AND2_X1 U9264 ( .A1(n9080), .A2(n6669), .ZN(n10110) );
  AND2_X1 U9265 ( .A1(n11708), .A2(n11707), .ZN(n13076) );
  INV_X1 U9266 ( .A(n13076), .ZN(n13271) );
  AND2_X1 U9267 ( .A1(n11040), .A2(n11044), .ZN(n12565) );
  INV_X1 U9268 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U9269 ( .A1(n8945), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6576) );
  AND2_X1 U9270 ( .A1(n7036), .A2(n7037), .ZN(n6577) );
  OR2_X1 U9271 ( .A1(n7148), .A2(n13002), .ZN(n6578) );
  OR2_X1 U9272 ( .A1(n13529), .A2(n13531), .ZN(n6579) );
  NAND2_X1 U9273 ( .A1(n11955), .A2(n11954), .ZN(n12996) );
  MUX2_X1 U9274 ( .A(n13895), .B(n14078), .S(n13520), .Z(n13613) );
  OR2_X1 U9275 ( .A1(n11820), .A2(n11822), .ZN(n6580) );
  AND2_X1 U9276 ( .A1(n7196), .A2(n7195), .ZN(n6581) );
  INV_X1 U9277 ( .A(n7652), .ZN(n7650) );
  NAND2_X1 U9278 ( .A1(n7654), .A2(n7653), .ZN(n7652) );
  AND2_X1 U9279 ( .A1(n11271), .A2(n11270), .ZN(n14440) );
  INV_X1 U9280 ( .A(n14440), .ZN(n7206) );
  INV_X1 U9281 ( .A(n13426), .ZN(n7315) );
  OR2_X1 U9282 ( .A1(n7525), .A2(n7523), .ZN(n6582) );
  OR2_X1 U9283 ( .A1(n14302), .A2(n14301), .ZN(n6583) );
  OR2_X1 U9284 ( .A1(n14847), .A2(n12891), .ZN(n6584) );
  INV_X1 U9285 ( .A(n13686), .ZN(n14021) );
  OR2_X1 U9286 ( .A1(n11840), .A2(n7638), .ZN(n6585) );
  INV_X1 U9287 ( .A(n13008), .ZN(n13100) );
  AND2_X1 U9288 ( .A1(n7115), .A2(n7114), .ZN(n6586) );
  OR2_X1 U9289 ( .A1(n7035), .A2(n12376), .ZN(n6587) );
  OR2_X1 U9290 ( .A1(n12716), .A2(n12440), .ZN(n6588) );
  AND3_X1 U9291 ( .A1(n8430), .A2(n8429), .A3(n8428), .ZN(n6589) );
  AND2_X1 U9292 ( .A1(n11573), .A2(n6544), .ZN(n6590) );
  NOR2_X1 U9293 ( .A1(n13282), .A2(n13038), .ZN(n6591) );
  NOR2_X1 U9294 ( .A1(n11074), .A2(n12465), .ZN(n6592) );
  NOR2_X1 U9295 ( .A1(n10191), .A2(n10192), .ZN(n6593) );
  NOR2_X1 U9296 ( .A1(n8241), .A2(n7566), .ZN(n6594) );
  NOR2_X1 U9297 ( .A1(n13668), .A2(n13702), .ZN(n6595) );
  AND2_X1 U9298 ( .A1(n7667), .A2(n8900), .ZN(n6596) );
  AND2_X1 U9299 ( .A1(n11128), .A2(n10996), .ZN(n6597) );
  AND2_X1 U9300 ( .A1(n7646), .A2(n6989), .ZN(n6598) );
  INV_X1 U9301 ( .A(n13617), .ZN(n6678) );
  AND2_X1 U9302 ( .A1(n13548), .A2(n10702), .ZN(n6599) );
  AND2_X1 U9303 ( .A1(n12561), .A2(n8050), .ZN(n6600) );
  AND2_X1 U9304 ( .A1(n11058), .A2(n12524), .ZN(n6601) );
  INV_X1 U9305 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8406) );
  OR2_X1 U9306 ( .A1(n7640), .A2(n11819), .ZN(n6602) );
  AND2_X1 U9307 ( .A1(n6494), .A2(n13256), .ZN(n6603) );
  AND2_X1 U9308 ( .A1(n6522), .A2(n7334), .ZN(n6604) );
  AND2_X1 U9309 ( .A1(n7615), .A2(n7626), .ZN(n6605) );
  NAND2_X1 U9310 ( .A1(n10632), .A2(n10372), .ZN(n6606) );
  NAND2_X1 U9311 ( .A1(n7544), .A2(n13526), .ZN(n6607) );
  NAND2_X1 U9312 ( .A1(n7554), .A2(n13603), .ZN(n6608) );
  INV_X1 U9313 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6939) );
  AND2_X1 U9314 ( .A1(n7390), .A2(n8754), .ZN(n6609) );
  AND2_X1 U9315 ( .A1(n7303), .A2(n11394), .ZN(n7302) );
  NOR2_X1 U9316 ( .A1(n8241), .A2(n7567), .ZN(n6610) );
  INV_X1 U9317 ( .A(n9642), .ZN(n7496) );
  INV_X1 U9318 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7002) );
  OR2_X1 U9319 ( .A1(n11823), .A2(n11818), .ZN(n6611) );
  NOR2_X1 U9320 ( .A1(n13207), .A2(n7456), .ZN(n7455) );
  CLKBUF_X3 U9321 ( .A(n7797), .Z(n8045) );
  NAND2_X1 U9322 ( .A1(n9068), .A2(n9044), .ZN(n9289) );
  INV_X1 U9323 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7012) );
  INV_X1 U9324 ( .A(n12887), .ZN(n7527) );
  NAND2_X1 U9325 ( .A1(n11354), .A2(n11353), .ZN(n13918) );
  INV_X1 U9326 ( .A(n13918), .ZN(n7210) );
  INV_X1 U9327 ( .A(n14956), .ZN(n7041) );
  INV_X1 U9328 ( .A(n11905), .ZN(n7655) );
  NAND2_X1 U9329 ( .A1(n11397), .A2(n11396), .ZN(n14078) );
  INV_X1 U9330 ( .A(n14078), .ZN(n7208) );
  AND2_X1 U9331 ( .A1(n7330), .A2(n7333), .ZN(n6612) );
  INV_X1 U9332 ( .A(n11912), .ZN(n6880) );
  NOR2_X1 U9333 ( .A1(n8004), .A2(n7357), .ZN(n7356) );
  NOR2_X1 U9334 ( .A1(n12665), .A2(n12496), .ZN(n6613) );
  NAND2_X1 U9335 ( .A1(n8129), .A2(n8128), .ZN(n12509) );
  INV_X1 U9336 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7611) );
  AND2_X1 U9337 ( .A1(n10235), .A2(n10571), .ZN(n6614) );
  INV_X1 U9338 ( .A(n14394), .ZN(n7327) );
  AND2_X1 U9339 ( .A1(n12425), .A2(n15093), .ZN(n6615) );
  INV_X1 U9340 ( .A(n12890), .ZN(n9958) );
  NAND2_X1 U9341 ( .A1(n8116), .A2(n8115), .ZN(n12496) );
  INV_X1 U9342 ( .A(n12496), .ZN(n12523) );
  OR2_X1 U9343 ( .A1(n10764), .A2(n14445), .ZN(n6616) );
  OR2_X1 U9344 ( .A1(n11300), .A2(n11301), .ZN(n6617) );
  NOR3_X1 U9345 ( .A1(n13167), .A2(n13157), .A3(n13292), .ZN(n6799) );
  AND4_X1 U9346 ( .A1(n7873), .A2(n7872), .A3(n7871), .A4(n7870), .ZN(n10401)
         );
  INV_X1 U9347 ( .A(n6800), .ZN(n10896) );
  NOR2_X1 U9348 ( .A1(n10847), .A2(n13331), .ZN(n6800) );
  INV_X1 U9349 ( .A(n7251), .ZN(n7250) );
  NOR2_X1 U9350 ( .A1(n13587), .A2(n7252), .ZN(n7251) );
  INV_X1 U9351 ( .A(n7133), .ZN(n12283) );
  NAND2_X1 U9352 ( .A1(n15008), .A2(n6816), .ZN(n7133) );
  AND2_X1 U9353 ( .A1(n7489), .A2(n7487), .ZN(n6618) );
  AND2_X1 U9354 ( .A1(n10509), .A2(n10508), .ZN(n10639) );
  NOR2_X1 U9355 ( .A1(n10896), .A2(n13328), .ZN(n7151) );
  INV_X1 U9356 ( .A(n7758), .ZN(n7359) );
  AND2_X1 U9357 ( .A1(n9026), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7758) );
  AND4_X1 U9358 ( .A1(n7885), .A2(n7884), .A3(n7883), .A4(n7882), .ZN(n15056)
         );
  INV_X1 U9359 ( .A(n15056), .ZN(n12228) );
  NAND2_X1 U9360 ( .A1(n7539), .A2(n13539), .ZN(n7538) );
  INV_X1 U9361 ( .A(n7435), .ZN(n11215) );
  NOR2_X1 U9362 ( .A1(n11216), .A2(n11217), .ZN(n7435) );
  INV_X1 U9363 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U9364 ( .A1(n8194), .A2(n8193), .ZN(n12417) );
  NOR2_X1 U9365 ( .A1(n9200), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n9476) );
  AND2_X1 U9366 ( .A1(n10441), .A2(SI_23_), .ZN(n6619) );
  AND2_X1 U9367 ( .A1(n7008), .A2(n6985), .ZN(n6620) );
  NAND2_X1 U9368 ( .A1(n8072), .A2(n8071), .ZN(n12677) );
  AND2_X1 U9369 ( .A1(n8717), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U9370 ( .A1(n7663), .A2(n7659), .ZN(n6622) );
  OR2_X1 U9371 ( .A1(n11913), .A2(n6880), .ZN(n6623) );
  AND2_X1 U9372 ( .A1(n6779), .A2(n7458), .ZN(n6624) );
  OR2_X1 U9373 ( .A1(n7637), .A2(n11841), .ZN(n6625) );
  OR2_X1 U9374 ( .A1(n14969), .A2(n12251), .ZN(n6626) );
  NAND2_X2 U9375 ( .A1(n13332), .A2(n8963), .ZN(n9668) );
  INV_X1 U9376 ( .A(n6749), .ZN(n7495) );
  INV_X1 U9377 ( .A(n12705), .ZN(n7570) );
  OR2_X1 U9378 ( .A1(n7980), .A2(n7979), .ZN(n12280) );
  AND2_X1 U9379 ( .A1(n7163), .A2(n7075), .ZN(n6627) );
  INV_X2 U9380 ( .A(n15162), .ZN(n15164) );
  AND2_X1 U9381 ( .A1(n14586), .A2(n7202), .ZN(n6628) );
  AND2_X1 U9382 ( .A1(n11027), .A2(n11023), .ZN(n12629) );
  OR2_X1 U9383 ( .A1(n11281), .A2(n11280), .ZN(n6629) );
  OR2_X1 U9384 ( .A1(n15164), .A2(n8272), .ZN(n6630) );
  INV_X1 U9385 ( .A(n8613), .ZN(n8611) );
  NOR2_X1 U9386 ( .A1(n12285), .A2(n12284), .ZN(n6631) );
  INV_X1 U9387 ( .A(n10254), .ZN(n7609) );
  NAND2_X1 U9388 ( .A1(n10214), .A2(n7867), .ZN(n6632) );
  AND2_X1 U9389 ( .A1(n12088), .A2(n7427), .ZN(n6633) );
  AND2_X1 U9390 ( .A1(n11180), .A2(n15364), .ZN(n6634) );
  INV_X1 U9391 ( .A(n12280), .ZN(n7163) );
  AND3_X2 U9392 ( .A1(n10866), .A2(n10865), .A3(n10864), .ZN(n15181) );
  INV_X1 U9393 ( .A(n15181), .ZN(n6961) );
  OR2_X1 U9394 ( .A1(n8414), .A2(n6886), .ZN(n6635) );
  AND2_X1 U9395 ( .A1(n11576), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6636) );
  AND2_X1 U9396 ( .A1(n7495), .A2(n7492), .ZN(n6637) );
  AND2_X1 U9397 ( .A1(n7412), .A2(n6529), .ZN(n6638) );
  INV_X1 U9398 ( .A(n7686), .ZN(n7408) );
  INV_X2 U9399 ( .A(n14727), .ZN(n14730) );
  INV_X1 U9400 ( .A(n12371), .ZN(n7035) );
  XNOR2_X1 U9401 ( .A(n8972), .B(n9372), .ZN(n9222) );
  NAND2_X1 U9402 ( .A1(n6663), .A2(n6662), .ZN(n7281) );
  INV_X1 U9403 ( .A(n6953), .ZN(n6940) );
  INV_X1 U9404 ( .A(n9924), .ZN(n6897) );
  INV_X1 U9405 ( .A(n12898), .ZN(n6906) );
  NAND2_X1 U9406 ( .A1(n9380), .A2(n8981), .ZN(n8990) );
  NAND2_X1 U9407 ( .A1(n14606), .A2(n10021), .ZN(n10088) );
  INV_X1 U9408 ( .A(n10088), .ZN(n7197) );
  OR2_X1 U9409 ( .A1(n12953), .A2(n12942), .ZN(n6639) );
  NAND2_X1 U9410 ( .A1(n12326), .A2(n12347), .ZN(n6640) );
  INV_X1 U9411 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8419) );
  AND2_X1 U9412 ( .A1(n9419), .A2(n11997), .ZN(n13226) );
  INV_X1 U9413 ( .A(n13226), .ZN(n13251) );
  AND2_X1 U9414 ( .A1(n7282), .A2(n7281), .ZN(n6641) );
  INV_X1 U9415 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6738) );
  INV_X1 U9416 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6724) );
  AND2_X1 U9417 ( .A1(n9122), .A2(n8747), .ZN(n10947) );
  OR2_X1 U9418 ( .A1(n10236), .A2(n10571), .ZN(n7053) );
  INV_X1 U9419 ( .A(n10571), .ZN(n7055) );
  NAND2_X1 U9420 ( .A1(n12252), .A2(n12251), .ZN(n7121) );
  AOI21_X1 U9421 ( .B1(n14967), .B2(n10567), .A(n12251), .ZN(n6664) );
  OR2_X1 U9422 ( .A1(n14979), .A2(n12251), .ZN(n7047) );
  AND2_X1 U9423 ( .A1(n10575), .A2(n12251), .ZN(n7048) );
  OR2_X1 U9424 ( .A1(n10575), .A2(n12251), .ZN(n7049) );
  AND2_X1 U9425 ( .A1(n10567), .A2(n12251), .ZN(n7082) );
  OR2_X1 U9426 ( .A1(n10567), .A2(n12251), .ZN(n7083) );
  OAI21_X2 U9427 ( .B1(n12599), .B2(n6644), .A(n6642), .ZN(n12563) );
  NAND2_X1 U9428 ( .A1(n7182), .A2(n7183), .ZN(n6649) );
  INV_X1 U9429 ( .A(n7183), .ZN(n6650) );
  NAND2_X1 U9430 ( .A1(n8223), .A2(n10983), .ZN(n10208) );
  NAND2_X1 U9431 ( .A1(n12512), .A2(n11064), .ZN(n6651) );
  NAND2_X1 U9432 ( .A1(n12525), .A2(n11060), .ZN(n6652) );
  NOR2_X2 U9433 ( .A1(n6653), .A2(n6654), .ZN(n7715) );
  NAND3_X1 U9434 ( .A1(n7712), .A2(n6496), .A3(n7671), .ZN(n6653) );
  NAND3_X1 U9435 ( .A1(n7555), .A2(n7701), .A3(n7556), .ZN(n7844) );
  NAND4_X1 U9436 ( .A1(n7703), .A2(n7705), .A3(n7704), .A4(n7702), .ZN(n6655)
         );
  NAND3_X1 U9437 ( .A1(n7817), .A2(n7815), .A3(n7816), .ZN(n15082) );
  NAND2_X1 U9438 ( .A1(n6657), .A2(n15097), .ZN(n10972) );
  XNOR2_X1 U9439 ( .A(n6473), .B(n6657), .ZN(n8283) );
  AOI22_X1 U9440 ( .A1(n12193), .A2(n6657), .B1(n12211), .B2(n12232), .ZN(
        n9512) );
  NAND2_X2 U9441 ( .A1(n9140), .A2(n11332), .ZN(n11100) );
  XNOR2_X2 U9442 ( .A(n7283), .B(n7793), .ZN(n9365) );
  NOR2_X1 U9443 ( .A1(n10224), .A2(n10228), .ZN(n10563) );
  NAND2_X2 U9444 ( .A1(n7232), .A2(n6671), .ZN(n11594) );
  NOR2_X1 U9445 ( .A1(n6672), .A2(n7228), .ZN(n6671) );
  OAI21_X1 U9446 ( .B1(n6971), .B2(n6572), .A(n7542), .ZN(n6687) );
  NAND3_X1 U9447 ( .A1(n8267), .A2(n6689), .A3(n6690), .ZN(n6688) );
  NAND2_X1 U9448 ( .A1(n8247), .A2(n10495), .ZN(n6690) );
  OR2_X1 U9449 ( .A1(n8639), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8251) );
  NAND2_X2 U9450 ( .A1(n12066), .A2(n8292), .ZN(n12090) );
  NAND2_X2 U9451 ( .A1(n6699), .A2(n12523), .ZN(n12165) );
  AND2_X2 U9452 ( .A1(n7423), .A2(n10011), .ZN(n7422) );
  INV_X1 U9453 ( .A(n6951), .ZN(n13667) );
  OAI21_X1 U9454 ( .B1(n13517), .B2(n6706), .A(n6705), .ZN(n13523) );
  NAND2_X1 U9455 ( .A1(n6708), .A2(n6707), .ZN(n13514) );
  NAND2_X1 U9456 ( .A1(n6709), .A2(n13510), .ZN(n6707) );
  NAND2_X1 U9457 ( .A1(n13507), .A2(n6710), .ZN(n6709) );
  NAND3_X1 U9458 ( .A1(n6711), .A2(n13502), .A3(n13503), .ZN(n6710) );
  NAND3_X1 U9459 ( .A1(n13497), .A2(n13495), .A3(n13496), .ZN(n6711) );
  NAND2_X1 U9460 ( .A1(n6712), .A2(n6547), .ZN(n13584) );
  NAND2_X1 U9461 ( .A1(n6713), .A2(n7538), .ZN(n6712) );
  NAND2_X1 U9462 ( .A1(n6715), .A2(n6714), .ZN(n6713) );
  NAND2_X1 U9463 ( .A1(n13537), .A2(n13536), .ZN(n6714) );
  NAND2_X1 U9464 ( .A1(n13533), .A2(n13532), .ZN(n6715) );
  NAND2_X1 U9465 ( .A1(n13610), .A2(n13609), .ZN(n13608) );
  OAI22_X1 U9466 ( .A1(n13606), .A2(n6717), .B1(n6716), .B2(n13605), .ZN(
        n13610) );
  INV_X1 U9467 ( .A(n13598), .ZN(n6942) );
  NAND2_X1 U9468 ( .A1(n6718), .A2(n7532), .ZN(n13598) );
  NAND4_X1 U9469 ( .A1(n6720), .A2(n6530), .A3(n6719), .A4(n7246), .ZN(n6718)
         );
  NAND2_X1 U9470 ( .A1(n13588), .A2(n13587), .ZN(n6719) );
  OAI21_X1 U9471 ( .B1(n13588), .B2(n13586), .A(n13585), .ZN(n6720) );
  NAND3_X1 U9472 ( .A1(n6729), .A2(n6734), .A3(n6731), .ZN(n6728) );
  NAND2_X1 U9473 ( .A1(n14297), .A2(n14298), .ZN(n14302) );
  OAI21_X1 U9474 ( .B1(n6730), .B2(n6733), .A(n14301), .ZN(n6729) );
  NAND2_X1 U9475 ( .A1(n6732), .A2(n14297), .ZN(n6731) );
  NOR2_X1 U9476 ( .A1(n14301), .A2(n6733), .ZN(n6732) );
  INV_X1 U9477 ( .A(n14298), .ZN(n6733) );
  INV_X1 U9478 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6734) );
  OAI21_X1 U9479 ( .B1(n14486), .B2(n14487), .A(P2_ADDR_REG_15__SCAN_IN), .ZN(
        n7266) );
  OAI21_X1 U9480 ( .B1(n14482), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n14481), .ZN(
        n6741) );
  NAND2_X1 U9481 ( .A1(n7496), .A2(n6749), .ZN(n6751) );
  NAND2_X1 U9482 ( .A1(n9559), .A2(n12829), .ZN(n6747) );
  NAND3_X1 U9483 ( .A1(n7471), .A2(n6748), .A3(n9329), .ZN(n6750) );
  INV_X1 U9484 ( .A(n7803), .ZN(n6754) );
  NAND2_X1 U9485 ( .A1(n6754), .A2(n7794), .ZN(n7730) );
  NAND2_X1 U9486 ( .A1(n6776), .A2(n6772), .ZN(n6774) );
  NAND2_X1 U9487 ( .A1(n7732), .A2(n7736), .ZN(n6773) );
  NAND2_X1 U9488 ( .A1(n7813), .A2(n7812), .ZN(n6776) );
  NAND2_X1 U9489 ( .A1(n9730), .A2(n9729), .ZN(n9731) );
  INV_X1 U9490 ( .A(n6787), .ZN(n13190) );
  NAND2_X1 U9491 ( .A1(n6787), .A2(n13027), .ZN(n6786) );
  NAND2_X1 U9492 ( .A1(n13078), .A2(n13077), .ZN(n6790) );
  NAND2_X1 U9493 ( .A1(n7464), .A2(n7463), .ZN(n13092) );
  NAND3_X1 U9494 ( .A1(n7140), .A2(n7139), .A3(n6596), .ZN(n13355) );
  XNOR2_X1 U9495 ( .A(n11768), .B(n14814), .ZN(n6953) );
  INV_X1 U9496 ( .A(n6796), .ZN(n13072) );
  OAI21_X2 U9497 ( .B1(n8968), .B2(n8967), .A(n6797), .ZN(n14814) );
  NAND2_X2 U9498 ( .A1(n8968), .A2(n8945), .ZN(n11953) );
  NOR2_X1 U9499 ( .A1(n13167), .A2(n13157), .ZN(n13152) );
  INV_X1 U9500 ( .A(n6799), .ZN(n13138) );
  INV_X1 U9501 ( .A(n7715), .ZN(n8243) );
  CLKBUF_X1 U9502 ( .A(n12397), .Z(n6812) );
  INV_X2 U9503 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7612) );
  NAND2_X1 U9504 ( .A1(n14766), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n14765) );
  NAND2_X1 U9505 ( .A1(n12582), .A2(n6600), .ZN(n12568) );
  NAND2_X1 U9506 ( .A1(n7717), .A2(n7716), .ZN(n7718) );
  NAND2_X1 U9507 ( .A1(n7717), .A2(n6832), .ZN(n7721) );
  NAND2_X1 U9508 ( .A1(n7572), .A2(n7571), .ZN(n10214) );
  NAND2_X1 U9509 ( .A1(n7595), .A2(n7597), .ZN(n6841) );
  OAI21_X1 U9510 ( .B1(n11333), .B2(n6844), .A(n6842), .ZN(n10534) );
  INV_X1 U9511 ( .A(n10256), .ZN(n6843) );
  NAND2_X1 U9512 ( .A1(n8596), .A2(n6845), .ZN(n6848) );
  NAND2_X1 U9513 ( .A1(n6848), .A2(n6847), .ZN(n8684) );
  INV_X1 U9514 ( .A(n9468), .ZN(n6860) );
  NAND3_X1 U9515 ( .A1(n7140), .A2(n7139), .A3(n7667), .ZN(n6864) );
  NAND2_X1 U9516 ( .A1(n6871), .A2(n6625), .ZN(n11847) );
  NAND2_X1 U9517 ( .A1(n7636), .A2(n6872), .ZN(n6871) );
  NAND3_X1 U9518 ( .A1(n6876), .A2(n6875), .A3(n6874), .ZN(n6873) );
  INV_X1 U9519 ( .A(n11835), .ZN(n6874) );
  INV_X1 U9520 ( .A(n11830), .ZN(n6875) );
  INV_X1 U9521 ( .A(n11831), .ZN(n6876) );
  OR2_X1 U9522 ( .A1(n11831), .A2(n11830), .ZN(n11836) );
  NAND3_X1 U9523 ( .A1(n11911), .A2(n11910), .A3(n6623), .ZN(n6877) );
  NAND2_X1 U9524 ( .A1(n11815), .A2(n11814), .ZN(n6999) );
  OAI21_X1 U9525 ( .B1(n7642), .B2(n11804), .A(n6598), .ZN(n6881) );
  NAND2_X1 U9526 ( .A1(n6883), .A2(n11808), .ZN(n6882) );
  NAND2_X1 U9527 ( .A1(n7645), .A2(n7643), .ZN(n6883) );
  OAI22_X2 U9528 ( .A1(n11856), .A2(n6884), .B1(n11857), .B2(n11855), .ZN(
        n11863) );
  AOI21_X1 U9529 ( .B1(n11863), .B2(n7632), .A(n7630), .ZN(n7629) );
  NOR2_X1 U9530 ( .A1(n6886), .A2(n7138), .ZN(n7137) );
  NAND2_X1 U9531 ( .A1(n6890), .A2(n6889), .ZN(P2_U3495) );
  OR2_X1 U9532 ( .A1(n14887), .A2(n11731), .ZN(n6889) );
  AOI21_X1 U9533 ( .B1(n13016), .B2(n7514), .A(n13226), .ZN(n6892) );
  NAND2_X1 U9534 ( .A1(n6893), .A2(n6584), .ZN(n10049) );
  NAND3_X1 U9535 ( .A1(n6894), .A2(n6898), .A3(n6580), .ZN(n6893) );
  NAND2_X1 U9536 ( .A1(n9923), .A2(n6896), .ZN(n6894) );
  INV_X1 U9537 ( .A(n13134), .ZN(n6900) );
  OAI21_X1 U9538 ( .B1(n6900), .B2(n6901), .A(n6899), .ZN(n13096) );
  NOR2_X1 U9539 ( .A1(n10882), .A2(n7499), .ZN(n10884) );
  NAND2_X1 U9540 ( .A1(n9424), .A2(n12008), .ZN(n9725) );
  NAND2_X1 U9541 ( .A1(n8482), .A2(n8483), .ZN(n8486) );
  NAND2_X1 U9542 ( .A1(n11979), .A2(n11978), .ZN(n7608) );
  NAND2_X1 U9543 ( .A1(n8515), .A2(n8514), .ZN(n8525) );
  NAND2_X1 U9544 ( .A1(n9822), .A2(n11951), .ZN(n9530) );
  NAND2_X1 U9545 ( .A1(n8511), .A2(n8510), .ZN(n8530) );
  NOR2_X1 U9546 ( .A1(n6930), .A2(n6929), .ZN(n6928) );
  CLKBUF_X3 U9547 ( .A(n8956), .Z(n11741) );
  NAND2_X1 U9548 ( .A1(n10032), .A2(n10031), .ZN(n10030) );
  NAND2_X1 U9549 ( .A1(n9939), .A2(n9938), .ZN(n9954) );
  AOI21_X1 U9550 ( .B1(n10444), .B2(n10443), .A(n7439), .ZN(n10520) );
  AOI21_X1 U9551 ( .B1(n13055), .B2(n13056), .A(n6925), .ZN(n13046) );
  NAND2_X1 U9552 ( .A1(n10294), .A2(n7675), .ZN(n10444) );
  NAND2_X1 U9553 ( .A1(n10520), .A2(n7681), .ZN(n6907) );
  NAND2_X1 U9554 ( .A1(n10968), .A2(n10969), .ZN(n15090) );
  AOI21_X1 U9555 ( .B1(n12478), .B2(n8158), .A(n6592), .ZN(n12466) );
  OAI22_X1 U9556 ( .A1(n12596), .A2(n8034), .B1(n12127), .B2(n12583), .ZN(
        n12580) );
  NAND2_X1 U9557 ( .A1(n6928), .A2(n8958), .ZN(n12896) );
  NAND2_X1 U9558 ( .A1(n13014), .A2(n13013), .ZN(n13069) );
  NAND2_X1 U9559 ( .A1(n7137), .A2(n7474), .ZN(n7141) );
  NAND2_X1 U9560 ( .A1(n13011), .A2(n13010), .ZN(n13082) );
  NAND2_X1 U9561 ( .A1(n7018), .A2(n15101), .ZN(n10968) );
  AOI21_X2 U9562 ( .B1(n12507), .B2(n8117), .A(n6613), .ZN(n12495) );
  OAI21_X2 U9563 ( .B1(n12547), .B2(n8079), .A(n7009), .ZN(n12532) );
  INV_X1 U9564 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7094) );
  NAND2_X1 U9565 ( .A1(n12494), .A2(n8131), .ZN(n12478) );
  NAND2_X1 U9566 ( .A1(n7583), .A2(n7587), .ZN(n9191) );
  NAND2_X1 U9567 ( .A1(n13667), .A2(n6967), .ZN(n6966) );
  NAND2_X1 U9568 ( .A1(n13839), .A2(n11628), .ZN(n13819) );
  NAND2_X1 U9569 ( .A1(n13898), .A2(n13897), .ZN(n13896) );
  NAND2_X1 U9570 ( .A1(n6910), .A2(n6908), .ZN(P1_U3556) );
  OR2_X1 U9571 ( .A1(n14166), .A2(n14727), .ZN(n6910) );
  NAND2_X1 U9572 ( .A1(n8066), .A2(n8065), .ZN(n8068) );
  AND4_X2 U9573 ( .A1(n6911), .A2(n6554), .A3(n7192), .A4(n7193), .ZN(n11163)
         );
  AND2_X1 U9574 ( .A1(n8425), .A2(n8424), .ZN(n7317) );
  NAND2_X1 U9575 ( .A1(n9910), .A2(n9909), .ZN(n10155) );
  NAND2_X1 U9576 ( .A1(n8054), .A2(n7767), .ZN(n8066) );
  NOR2_X1 U9577 ( .A1(n11088), .A2(n12439), .ZN(n11094) );
  NAND2_X1 U9578 ( .A1(n12413), .A2(n15107), .ZN(n6914) );
  OAI21_X1 U9579 ( .B1(n11755), .B2(n15162), .A(n6506), .ZN(P3_U3456) );
  NAND3_X1 U9580 ( .A1(n6493), .A2(n7000), .A3(n6555), .ZN(n7026) );
  NAND2_X1 U9581 ( .A1(n6914), .A2(n6912), .ZN(P3_U3204) );
  NAND2_X1 U9582 ( .A1(n10067), .A2(n7834), .ZN(n10077) );
  NAND2_X1 U9583 ( .A1(n10398), .A2(n8224), .ZN(n7580) );
  NAND2_X1 U9584 ( .A1(n15092), .A2(n15073), .ZN(n7818) );
  NAND2_X1 U9585 ( .A1(n7559), .A2(n15077), .ZN(n10067) );
  OAI21_X1 U9586 ( .B1(n10979), .B2(n7558), .A(n7557), .ZN(n7559) );
  NAND2_X1 U9587 ( .A1(n12423), .A2(n6588), .ZN(n8200) );
  NAND2_X1 U9588 ( .A1(n12466), .A2(n8159), .ZN(n12450) );
  AND2_X1 U9589 ( .A1(n7792), .A2(n7789), .ZN(n6916) );
  NAND3_X2 U9590 ( .A1(n6916), .A2(n7790), .A3(n7791), .ZN(n12234) );
  INV_X1 U9591 ( .A(n12580), .ZN(n6917) );
  INV_X2 U9592 ( .A(n8955), .ZN(n8982) );
  INV_X1 U9593 ( .A(n13630), .ZN(n6931) );
  NAND2_X1 U9594 ( .A1(n7531), .A2(n7530), .ZN(n9047) );
  NAND2_X1 U9595 ( .A1(n7023), .A2(n7546), .ZN(n13534) );
  NAND2_X1 U9596 ( .A1(n6970), .A2(n6969), .ZN(n6968) );
  NAND2_X1 U9597 ( .A1(n10287), .A2(n10286), .ZN(n10294) );
  NAND2_X1 U9598 ( .A1(n10036), .A2(n9415), .ZN(n9417) );
  NAND2_X1 U9599 ( .A1(n13534), .A2(n13535), .ZN(n13533) );
  NAND2_X1 U9600 ( .A1(n13623), .A2(n13624), .ZN(n13622) );
  MUX2_X1 U9601 ( .A(n13500), .B(n13499), .S(n13498), .Z(n13501) );
  INV_X1 U9602 ( .A(n9041), .ZN(n8437) );
  NAND2_X1 U9603 ( .A1(n6944), .A2(n13713), .ZN(P1_U3242) );
  NAND2_X1 U9604 ( .A1(n6946), .A2(n6945), .ZN(n6944) );
  NAND3_X1 U9605 ( .A1(n6965), .A2(n6966), .A3(n6964), .ZN(n6946) );
  NAND2_X1 U9606 ( .A1(n10285), .A2(n7676), .ZN(n10287) );
  NAND2_X1 U9607 ( .A1(n10052), .A2(n9955), .ZN(n9956) );
  INV_X1 U9608 ( .A(n13610), .ZN(n6970) );
  XNOR2_X1 U9609 ( .A(n8496), .B(n8495), .ZN(n9574) );
  NAND2_X1 U9610 ( .A1(n12434), .A2(n12433), .ZN(n12436) );
  NAND2_X1 U9611 ( .A1(n9195), .A2(n9194), .ZN(n9469) );
  NAND2_X1 U9612 ( .A1(n8684), .A2(n8683), .ZN(n8687) );
  NAND2_X1 U9613 ( .A1(n7260), .A2(n7259), .ZN(n13859) );
  INV_X1 U9614 ( .A(n9454), .ZN(n13249) );
  NAND2_X1 U9615 ( .A1(n6951), .A2(n6595), .ZN(n6965) );
  OAI21_X2 U9616 ( .B1(n14351), .B2(n10957), .A(n10951), .ZN(n12630) );
  OAI21_X2 U9617 ( .B1(n12630), .B2(n7190), .A(n7186), .ZN(n12601) );
  NAND2_X1 U9618 ( .A1(n14341), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U9619 ( .A1(n14339), .A2(n14338), .ZN(n7268) );
  NAND2_X1 U9620 ( .A1(n14486), .A2(n14487), .ZN(n14485) );
  XNOR2_X1 U9621 ( .A(n7273), .B(n7272), .ZN(SUB_1596_U4) );
  NAND2_X1 U9622 ( .A1(n7341), .A2(n7339), .ZN(n8054) );
  NAND2_X1 U9623 ( .A1(n7741), .A2(n7740), .ZN(n7887) );
  NAND2_X1 U9624 ( .A1(n7907), .A2(n7906), .ZN(n7909) );
  XNOR2_X1 U9625 ( .A(n6955), .B(n9247), .ZN(n11152) );
  NAND3_X1 U9626 ( .A1(n7196), .A2(n6957), .A3(n6956), .ZN(n6955) );
  INV_X1 U9627 ( .A(n11150), .ZN(n6956) );
  XNOR2_X2 U9628 ( .A(n14188), .B(n13717), .ZN(n13930) );
  INV_X1 U9629 ( .A(n11130), .ZN(n7866) );
  OAI21_X1 U9630 ( .B1(n12714), .B2(n6961), .A(n6959), .ZN(P3_U3487) );
  OAI21_X1 U9631 ( .B1(n12714), .B2(n15162), .A(n6962), .ZN(P3_U3455) );
  NAND3_X1 U9632 ( .A1(n13611), .A2(n7549), .A3(n6968), .ZN(n7548) );
  NAND2_X1 U9633 ( .A1(n6497), .A2(n6607), .ZN(n6971) );
  NAND3_X1 U9634 ( .A1(n13600), .A2(n13599), .A3(n6608), .ZN(n7551) );
  NAND2_X1 U9635 ( .A1(n6972), .A2(n13490), .ZN(n13643) );
  AOI21_X1 U9636 ( .B1(n7465), .B2(n13115), .A(n6591), .ZN(n7463) );
  OAI22_X1 U9637 ( .A1(n9510), .A2(n9511), .B1(n12233), .B2(n8284), .ZN(n9894)
         );
  OAI22_X2 U9638 ( .A1(n12159), .A2(n8311), .B1(n12619), .B2(n8312), .ZN(
        n11216) );
  AOI22_X1 U9639 ( .A1(n10246), .A2(n10245), .B1(n15055), .B2(n8288), .ZN(
        n10273) );
  NAND2_X1 U9640 ( .A1(n15070), .A2(n15074), .ZN(n15069) );
  NAND2_X1 U9641 ( .A1(n15069), .A2(n10972), .ZN(n10062) );
  NAND2_X1 U9642 ( .A1(n12233), .A2(n15082), .ZN(n10973) );
  OAI21_X1 U9643 ( .B1(n6980), .B2(n6982), .A(n13021), .ZN(n13022) );
  NAND2_X1 U9644 ( .A1(n8948), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8926) );
  NOR2_X1 U9645 ( .A1(n13016), .A2(n7512), .ZN(n6982) );
  AOI21_X1 U9646 ( .B1(n6983), .B2(n15099), .A(n12441), .ZN(n12442) );
  NAND2_X1 U9647 ( .A1(n12438), .A2(n6984), .ZN(n6983) );
  NAND2_X1 U9648 ( .A1(n11059), .A2(n6601), .ZN(n11063) );
  NAND2_X1 U9649 ( .A1(n10997), .A2(n6597), .ZN(n11001) );
  MUX2_X2 U9650 ( .A(n11018), .B(n11017), .S(n11093), .Z(n11020) );
  AOI21_X1 U9651 ( .B1(n11073), .B2(n11093), .A(n12467), .ZN(n7346) );
  NAND2_X1 U9652 ( .A1(n14953), .A2(n14954), .ZN(n14952) );
  NOR2_X1 U9653 ( .A1(n14987), .A2(n10584), .ZN(n10585) );
  AOI22_X1 U9654 ( .A1(n9353), .A2(n14912), .B1(n9176), .B2(n9175), .ZN(n9307)
         );
  NAND2_X1 U9655 ( .A1(n9224), .A2(n9413), .ZN(n9423) );
  NAND2_X1 U9656 ( .A1(n6988), .A2(n11771), .ZN(n11778) );
  NAND2_X1 U9657 ( .A1(n11767), .A2(n11772), .ZN(n6988) );
  OR2_X1 U9658 ( .A1(n11847), .A2(n11846), .ZN(n7687) );
  NAND3_X1 U9659 ( .A1(n6501), .A2(n6990), .A3(n6611), .ZN(n7639) );
  AOI21_X1 U9660 ( .B1(n11829), .B2(n11828), .A(n11827), .ZN(n11831) );
  OAI21_X1 U9661 ( .B1(n11785), .B2(n11784), .A(n6991), .ZN(n11793) );
  NAND2_X1 U9662 ( .A1(n6993), .A2(n6992), .ZN(n6991) );
  NAND2_X1 U9663 ( .A1(n11785), .A2(n11784), .ZN(n6993) );
  NAND2_X2 U9664 ( .A1(n7019), .A2(n11956), .ZN(n14881) );
  NAND2_X1 U9665 ( .A1(n6995), .A2(n6994), .ZN(n7636) );
  NAND2_X1 U9666 ( .A1(n11836), .A2(n11835), .ZN(n6995) );
  NAND3_X2 U9667 ( .A1(n8781), .A2(n8401), .A3(n8780), .ZN(n8414) );
  XNOR2_X2 U9668 ( .A(n6996), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U9669 ( .A1(n9476), .A2(n8406), .ZN(n6997) );
  NAND2_X1 U9670 ( .A1(n11947), .A2(n11946), .ZN(n7000) );
  INV_X1 U9671 ( .A(n7644), .ZN(n7642) );
  AOI21_X1 U9672 ( .B1(n11847), .B2(n11846), .A(n11844), .ZN(n11845) );
  NAND2_X1 U9673 ( .A1(n10103), .A2(n10102), .ZN(n10106) );
  NAND2_X1 U9674 ( .A1(n11445), .A2(n11443), .ZN(n11176) );
  OAI22_X2 U9675 ( .A1(n7004), .A2(n7003), .B1(n14168), .B2(n14050), .ZN(
        n11629) );
  AOI21_X1 U9676 ( .B1(n7342), .B2(n7345), .A(n7340), .ZN(n7339) );
  NAND2_X1 U9677 ( .A1(n7007), .A2(n7005), .ZN(P3_U3454) );
  OR2_X1 U9678 ( .A1(n12717), .A2(n15162), .ZN(n7007) );
  NAND2_X1 U9679 ( .A1(n12532), .A2(n12538), .ZN(n8091) );
  NAND2_X1 U9680 ( .A1(n12495), .A2(n8130), .ZN(n12494) );
  NAND2_X1 U9681 ( .A1(n13016), .A2(n13015), .ZN(n13057) );
  NOR2_X1 U9682 ( .A1(n8955), .A2(n8629), .ZN(n7020) );
  AND2_X1 U9683 ( .A1(n8410), .A2(n8411), .ZN(n7013) );
  NAND2_X1 U9684 ( .A1(n12999), .A2(n7497), .ZN(n13223) );
  NAND2_X1 U9685 ( .A1(n8613), .A2(n8612), .ZN(n7466) );
  AND2_X2 U9686 ( .A1(n14915), .A2(n7793), .ZN(n7555) );
  XNOR2_X1 U9687 ( .A(n8277), .B(n7430), .ZN(n8278) );
  OAI21_X1 U9688 ( .B1(n12144), .B2(n12143), .A(n12203), .ZN(n12149) );
  INV_X1 U9689 ( .A(n9459), .ZN(n7019) );
  INV_X1 U9690 ( .A(n8414), .ZN(n7474) );
  NAND2_X1 U9691 ( .A1(n7616), .A2(n6605), .ZN(n11947) );
  NAND2_X1 U9692 ( .A1(n9422), .A2(n9421), .ZN(n10031) );
  AOI21_X1 U9693 ( .B1(n10881), .B2(n12883), .A(n10880), .ZN(n10882) );
  INV_X1 U9694 ( .A(n9413), .ZN(n14822) );
  INV_X1 U9695 ( .A(n13512), .ZN(n7545) );
  NAND2_X1 U9696 ( .A1(n10884), .A2(n10883), .ZN(n12999) );
  AOI22_X2 U9697 ( .A1(n8276), .A2(n9452), .B1(n8275), .B2(n12760), .ZN(n8277)
         );
  NAND2_X1 U9698 ( .A1(n6546), .A2(n8335), .ZN(n12167) );
  NAND2_X1 U9699 ( .A1(n7467), .A2(n9813), .ZN(n9923) );
  NAND2_X1 U9700 ( .A1(n7469), .A2(n7468), .ZN(n9812) );
  NAND2_X1 U9701 ( .A1(n7026), .A2(n7670), .ZN(n11991) );
  NAND2_X1 U9702 ( .A1(n7591), .A2(n7592), .ZN(n8596) );
  NOR2_X1 U9703 ( .A1(n8535), .A2(n8579), .ZN(n7590) );
  NAND2_X1 U9704 ( .A1(n7586), .A2(n7584), .ZN(n9195) );
  INV_X1 U9705 ( .A(n8201), .ZN(n7712) );
  NAND2_X1 U9706 ( .A1(n7029), .A2(n9159), .ZN(n7033) );
  NAND3_X1 U9707 ( .A1(n7030), .A2(P3_REG1_REG_3__SCAN_IN), .A3(n9159), .ZN(
        n7029) );
  INV_X1 U9708 ( .A(n7033), .ZN(n9163) );
  AND2_X2 U9709 ( .A1(n7034), .A2(n6587), .ZN(n12380) );
  NAND3_X1 U9710 ( .A1(n7038), .A2(n7043), .A3(n7036), .ZN(n14958) );
  INV_X1 U9711 ( .A(n7045), .ZN(n14957) );
  NAND3_X1 U9712 ( .A1(n7047), .A2(n7049), .A3(n7046), .ZN(n10576) );
  NAND3_X1 U9713 ( .A1(n7047), .A2(n6507), .A3(n7046), .ZN(n7050) );
  INV_X1 U9714 ( .A(n7050), .ZN(n12242) );
  NAND3_X1 U9715 ( .A1(n7053), .A2(n7054), .A3(n7051), .ZN(n10237) );
  NAND3_X1 U9716 ( .A1(n7053), .A2(n7052), .A3(n7051), .ZN(n7057) );
  INV_X1 U9717 ( .A(n7057), .ZN(n10572) );
  NOR2_X1 U9718 ( .A1(n15000), .A2(n7076), .ZN(n12273) );
  OR2_X1 U9719 ( .A1(n14970), .A2(n6626), .ZN(n7080) );
  AOI21_X1 U9720 ( .B1(n14970), .B2(n7082), .A(n7078), .ZN(n7077) );
  NAND3_X1 U9721 ( .A1(n7081), .A2(n7083), .A3(n7080), .ZN(n10568) );
  NAND2_X1 U9722 ( .A1(n9177), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7085) );
  XNOR2_X2 U9723 ( .A(n7814), .B(P3_IR_REG_2__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U9724 ( .A1(n11207), .A2(n11194), .ZN(n7086) );
  NAND2_X1 U9725 ( .A1(n12807), .A2(n12806), .ZN(n11207) );
  NAND2_X1 U9726 ( .A1(n11574), .A2(n6590), .ZN(n7087) );
  NAND2_X1 U9727 ( .A1(n12798), .A2(n6586), .ZN(n7110) );
  OAI21_X1 U9728 ( .B1(n12798), .B2(n7485), .A(n7115), .ZN(n12773) );
  NAND2_X1 U9729 ( .A1(n7110), .A2(n7111), .ZN(n11740) );
  MUX2_X1 U9730 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8945), .Z(n8517) );
  AND2_X1 U9731 ( .A1(n7124), .A2(n7123), .ZN(n9175) );
  AND2_X1 U9732 ( .A1(n12396), .A2(n12395), .ZN(n7131) );
  INV_X2 U9733 ( .A(n8414), .ZN(n7139) );
  AND2_X1 U9734 ( .A1(n13072), .A2(n7144), .ZN(n13047) );
  OR2_X1 U9735 ( .A1(n13072), .A2(n13256), .ZN(n7143) );
  NAND2_X1 U9736 ( .A1(n13072), .A2(n6494), .ZN(n12992) );
  OAI211_X1 U9737 ( .C1(n6494), .C2(n13256), .A(n7143), .B(n7142), .ZN(n12984)
         );
  NAND2_X1 U9738 ( .A1(n13072), .A2(n6603), .ZN(n7142) );
  INV_X1 U9739 ( .A(n7151), .ZN(n13230) );
  NOR2_X2 U9740 ( .A1(n13122), .A2(n13282), .ZN(n13102) );
  NOR2_X2 U9741 ( .A1(n10055), .A2(n14860), .ZN(n10288) );
  NAND3_X1 U9742 ( .A1(n14915), .A2(n7793), .A3(n7159), .ZN(n7828) );
  INV_X2 U9743 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n14915) );
  MUX2_X1 U9744 ( .A(n12772), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  MUX2_X1 U9745 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12772), .S(n9140), .Z(n9700)
         );
  NOR2_X2 U9746 ( .A1(n12247), .A2(n14365), .ZN(n12268) );
  XNOR2_X2 U9747 ( .A(n12267), .B(n7163), .ZN(n12247) );
  NAND2_X1 U9748 ( .A1(n7168), .A2(n7169), .ZN(n12434) );
  NAND2_X1 U9749 ( .A1(n12464), .A2(n7170), .ZN(n7168) );
  NAND2_X1 U9750 ( .A1(n15035), .A2(n7176), .ZN(n7174) );
  OAI21_X1 U9751 ( .B1(n11130), .B2(n7185), .A(n15061), .ZN(n7182) );
  OAI21_X1 U9752 ( .B1(n12630), .B2(n8226), .A(n11027), .ZN(n12612) );
  NAND2_X1 U9753 ( .A1(n12611), .A2(n7191), .ZN(n7190) );
  NOR2_X2 U9754 ( .A1(n13811), .A2(n13815), .ZN(n13810) );
  NOR3_X4 U9755 ( .A1(n10764), .A2(n7205), .A3(n7207), .ZN(n14010) );
  OAI211_X1 U9756 ( .C1(n7231), .C2(n7234), .A(n8945), .B(n7229), .ZN(n9280)
         );
  NAND2_X1 U9757 ( .A1(n7230), .A2(n14496), .ZN(n7229) );
  INV_X1 U9758 ( .A(n7232), .ZN(n7230) );
  INV_X1 U9759 ( .A(n14496), .ZN(n7231) );
  OAI21_X1 U9760 ( .B1(n13966), .B2(n7239), .A(n7236), .ZN(n13929) );
  OAI21_X1 U9761 ( .B1(n14007), .B2(n7247), .A(n7245), .ZN(n11602) );
  OAI21_X1 U9762 ( .B1(n10760), .B2(n7256), .A(n7255), .ZN(n11598) );
  NAND2_X1 U9763 ( .A1(n13893), .A2(n7262), .ZN(n7259) );
  INV_X1 U9764 ( .A(n7263), .ZN(n13892) );
  INV_X1 U9765 ( .A(n7282), .ZN(n14943) );
  OAI21_X1 U9766 ( .B1(n9787), .B2(n7286), .A(n9903), .ZN(n7285) );
  OAI211_X1 U9767 ( .C1(n13477), .C2(n7297), .A(n7294), .B(n7292), .ZN(n11494)
         );
  NAND2_X1 U9768 ( .A1(n13477), .A2(n7293), .ZN(n7292) );
  NOR2_X1 U9769 ( .A1(n7295), .A2(n11481), .ZN(n7293) );
  OAI22_X1 U9770 ( .A1(n7296), .A2(n7295), .B1(n11481), .B2(n7298), .ZN(n7294)
         );
  NOR2_X1 U9771 ( .A1(n11481), .A2(n13370), .ZN(n7296) );
  NAND2_X1 U9772 ( .A1(n13370), .A2(n11481), .ZN(n7297) );
  NAND2_X1 U9773 ( .A1(n13456), .A2(n7302), .ZN(n7299) );
  AND3_X4 U9774 ( .A1(n7316), .A2(n7317), .A3(n8426), .ZN(n9215) );
  AND4_X2 U9775 ( .A1(n8822), .A2(n8599), .A3(n8715), .A4(n8825), .ZN(n7316)
         );
  AND3_X2 U9776 ( .A1(n6589), .A2(n8454), .A3(n8427), .ZN(n8431) );
  NAND3_X1 U9777 ( .A1(n14420), .A2(n6511), .A3(n7319), .ZN(n7318) );
  NAND2_X1 U9778 ( .A1(n10919), .A2(n6604), .ZN(n7329) );
  AND2_X1 U9779 ( .A1(n11240), .A2(n11241), .ZN(n7335) );
  NAND2_X1 U9780 ( .A1(n8439), .A2(n8438), .ZN(n8750) );
  NAND2_X1 U9781 ( .A1(n8020), .A2(n7342), .ZN(n7341) );
  NAND2_X1 U9782 ( .A1(n7347), .A2(n7346), .ZN(n11085) );
  INV_X1 U9783 ( .A(n7770), .ZN(n7352) );
  NAND2_X1 U9784 ( .A1(n10018), .A2(n13673), .ZN(n7379) );
  NAND2_X1 U9785 ( .A1(n13960), .A2(n7383), .ZN(n7380) );
  NAND2_X1 U9786 ( .A1(n7380), .A2(n7381), .ZN(n13915) );
  INV_X1 U9787 ( .A(n11622), .ZN(n7389) );
  NAND4_X1 U9788 ( .A1(n9215), .A2(n6609), .A3(n8436), .A4(n8431), .ZN(n8757)
         );
  NAND2_X1 U9789 ( .A1(n10773), .A2(n6599), .ZN(n10925) );
  NAND2_X1 U9790 ( .A1(n11617), .A2(n7392), .ZN(n7391) );
  NAND2_X1 U9791 ( .A1(n7391), .A2(n11618), .ZN(n13959) );
  NAND2_X1 U9792 ( .A1(n7394), .A2(n7396), .ZN(n13992) );
  NAND2_X1 U9793 ( .A1(n10551), .A2(n7406), .ZN(n7405) );
  INV_X1 U9794 ( .A(n14579), .ZN(n7413) );
  NAND2_X2 U9795 ( .A1(n8337), .A2(n8336), .ZN(n12139) );
  NAND2_X1 U9796 ( .A1(n9894), .A2(n7422), .ZN(n7420) );
  NAND2_X1 U9797 ( .A1(n7420), .A2(n7421), .ZN(n10246) );
  INV_X1 U9798 ( .A(n7424), .ZN(n9893) );
  OAI21_X1 U9799 ( .B1(n11216), .B2(n7433), .A(n7431), .ZN(n8319) );
  NAND2_X1 U9800 ( .A1(n8024), .A2(n7436), .ZN(n7683) );
  NAND2_X1 U9801 ( .A1(n7438), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8039) );
  AND2_X1 U9802 ( .A1(n8025), .A2(n7438), .ZN(n12333) );
  NAND2_X1 U9803 ( .A1(n6486), .A2(n9594), .ZN(n9325) );
  NAND2_X1 U9804 ( .A1(n13114), .A2(n7465), .ZN(n7464) );
  NAND2_X1 U9805 ( .A1(n9812), .A2(n9814), .ZN(n7467) );
  NAND2_X1 U9806 ( .A1(n9725), .A2(n9724), .ZN(n7469) );
  INV_X1 U9807 ( .A(n8990), .ZN(n7472) );
  XNOR2_X1 U9808 ( .A(n11736), .B(n11801), .ZN(n12825) );
  NAND2_X1 U9809 ( .A1(n9560), .A2(n12829), .ZN(n7493) );
  NAND2_X1 U9810 ( .A1(n7504), .A2(n7505), .ZN(n10595) );
  OAI21_X1 U9811 ( .B1(n10321), .B2(n10309), .A(n10319), .ZN(n10457) );
  OR2_X1 U9812 ( .A1(n10458), .A2(n10459), .ZN(n7506) );
  NAND2_X1 U9813 ( .A1(n13016), .A2(n7511), .ZN(n7510) );
  NAND3_X1 U9814 ( .A1(n7529), .A2(n8975), .A3(n7528), .ZN(n9413) );
  NAND2_X1 U9815 ( .A1(n11506), .A2(n8974), .ZN(n7529) );
  NAND2_X1 U9816 ( .A1(n8431), .A2(n9215), .ZN(n9010) );
  INV_X1 U9817 ( .A(n13620), .ZN(n7536) );
  INV_X1 U9818 ( .A(n13525), .ZN(n7544) );
  NAND2_X1 U9819 ( .A1(n7548), .A2(n7550), .ZN(n13616) );
  NAND3_X1 U9820 ( .A1(n12232), .A2(n15120), .A3(n7819), .ZN(n7557) );
  NAND2_X1 U9821 ( .A1(n15077), .A2(n7819), .ZN(n10065) );
  INV_X1 U9822 ( .A(n12629), .ZN(n7564) );
  INV_X1 U9823 ( .A(n12618), .ZN(n7565) );
  AND2_X1 U9824 ( .A1(n8222), .A2(n6610), .ZN(n11755) );
  AOI21_X1 U9825 ( .B1(n8222), .B2(n6594), .A(n6499), .ZN(P3_U3488) );
  NAND2_X1 U9826 ( .A1(n7568), .A2(n8221), .ZN(n7566) );
  NAND2_X1 U9827 ( .A1(n8222), .A2(n8221), .ZN(n12413) );
  NAND2_X1 U9828 ( .A1(n7715), .A2(n7574), .ZN(n7785) );
  NAND2_X1 U9829 ( .A1(n7715), .A2(n7714), .ZN(n8248) );
  INV_X1 U9830 ( .A(n7785), .ZN(n7717) );
  NAND2_X1 U9831 ( .A1(n8537), .A2(n7590), .ZN(n7591) );
  OAI21_X1 U9832 ( .B1(n7625), .B2(n6495), .A(n11917), .ZN(n7624) );
  OAI21_X1 U9833 ( .B1(n11863), .B2(n7635), .A(n7632), .ZN(n11871) );
  INV_X1 U9834 ( .A(n7629), .ZN(n11870) );
  INV_X1 U9835 ( .A(n11841), .ZN(n7638) );
  NAND2_X1 U9836 ( .A1(n7639), .A2(n6602), .ZN(n11829) );
  NAND2_X1 U9837 ( .A1(n11802), .A2(n11803), .ZN(n7644) );
  NAND2_X1 U9838 ( .A1(n11804), .A2(n7646), .ZN(n7645) );
  NAND3_X1 U9839 ( .A1(n11874), .A2(n7658), .A3(n11873), .ZN(n7657) );
  AND2_X1 U9840 ( .A1(n7657), .A2(n7656), .ZN(n11894) );
  NAND2_X1 U9841 ( .A1(n7665), .A2(n7664), .ZN(n7663) );
  INV_X1 U9842 ( .A(n11880), .ZN(n7665) );
  NAND2_X1 U9843 ( .A1(n8437), .A2(n9042), .ZN(n8752) );
  INV_X1 U9844 ( .A(n11255), .ZN(n11257) );
  AND2_X4 U9845 ( .A1(n9122), .A2(n13487), .ZN(n11234) );
  INV_X1 U9846 ( .A(n12768), .ZN(n7724) );
  OR2_X1 U9847 ( .A1(n9095), .A2(P1_B_REG_SCAN_IN), .ZN(n9096) );
  AND2_X1 U9848 ( .A1(n12436), .A2(n12435), .ZN(n12644) );
  OAI22_X1 U9849 ( .A1(n13675), .A2(n10108), .B1(n13731), .B2(n6668), .ZN(
        n10122) );
  NAND2_X1 U9850 ( .A1(n8948), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8910) );
  OR2_X1 U9851 ( .A1(n8955), .A2(n8905), .ZN(n8908) );
  NAND2_X1 U9852 ( .A1(n10053), .A2(n12012), .ZN(n10052) );
  XNOR2_X1 U9853 ( .A(n10532), .B(n10533), .ZN(n11663) );
  NAND2_X1 U9854 ( .A1(n13240), .A2(n9412), .ZN(n10037) );
  NAND2_X1 U9855 ( .A1(n7139), .A2(n8892), .ZN(n9212) );
  AND2_X1 U9856 ( .A1(n6480), .A2(n9452), .ZN(n11121) );
  INV_X1 U9857 ( .A(n7723), .ZN(n12048) );
  NAND4_X2 U9858 ( .A1(n7801), .A2(n7800), .A3(n7799), .A4(n7798), .ZN(n15094)
         );
  INV_X2 U9859 ( .A(n15107), .ZN(n15068) );
  AND4_X1 U9860 ( .A1(n8204), .A2(n8202), .A3(n7711), .A4(n8264), .ZN(n7671)
         );
  NAND2_X1 U9861 ( .A1(n11251), .A2(n11250), .ZN(n7672) );
  OR2_X1 U9862 ( .A1(n10284), .A2(n10283), .ZN(n7676) );
  AND2_X1 U9863 ( .A1(n13298), .A2(n13034), .ZN(n7678) );
  OR2_X1 U9864 ( .A1(n13187), .A2(n13029), .ZN(n7679) );
  INV_X1 U9865 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7689) );
  OR2_X1 U9866 ( .A1(n10836), .A2(n12884), .ZN(n7680) );
  INV_X1 U9867 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7912) );
  AND2_X1 U9868 ( .A1(n11332), .A2(P2_U3088), .ZN(n10257) );
  AND2_X1 U9869 ( .A1(n8819), .A2(n8779), .ZN(n7682) );
  OR2_X1 U9870 ( .A1(n9563), .A2(n9562), .ZN(n7684) );
  AND2_X1 U9871 ( .A1(n13929), .A2(n11604), .ZN(n7685) );
  INV_X1 U9872 ( .A(n12007), .ZN(n9920) );
  AND2_X1 U9873 ( .A1(n14416), .A2(n10649), .ZN(n7686) );
  NAND2_X1 U9874 ( .A1(n8918), .A2(n13232), .ZN(n12875) );
  NAND2_X1 U9875 ( .A1(n12898), .A2(n11760), .ZN(n11764) );
  NAND2_X1 U9876 ( .A1(n12897), .A2(n11782), .ZN(n11774) );
  NAND2_X1 U9877 ( .A1(n11798), .A2(n11797), .ZN(n11804) );
  INV_X1 U9878 ( .A(n11854), .ZN(n11855) );
  INV_X1 U9879 ( .A(n11891), .ZN(n11892) );
  OAI21_X1 U9880 ( .B1(n11894), .B2(n11893), .A(n11892), .ZN(n11895) );
  AND2_X1 U9881 ( .A1(n11975), .A2(n11945), .ZN(n11946) );
  INV_X1 U9882 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7711) );
  OR2_X1 U9883 ( .A1(n11866), .A2(n11868), .ZN(n10838) );
  INV_X1 U9884 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8433) );
  INV_X1 U9885 ( .A(n12620), .ZN(n8315) );
  INV_X1 U9886 ( .A(n8099), .ZN(n7695) );
  INV_X1 U9887 ( .A(n14633), .ZN(n9044) );
  OR4_X1 U9888 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U9889 ( .A1(n9072), .A2(n8433), .ZN(n8434) );
  INV_X1 U9890 ( .A(n15024), .ZN(n8297) );
  INV_X1 U9891 ( .A(n12179), .ZN(n8302) );
  INV_X1 U9892 ( .A(n8137), .ZN(n7697) );
  INV_X1 U9893 ( .A(n12421), .ZN(n8189) );
  INV_X1 U9894 ( .A(n12499), .ZN(n8130) );
  INV_X1 U9895 ( .A(n12552), .ZN(n8228) );
  INV_X1 U9896 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7701) );
  INV_X1 U9897 ( .A(n11989), .ZN(n11990) );
  INV_X1 U9898 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9646) );
  INV_X1 U9899 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8408) );
  INV_X1 U9900 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9981) );
  INV_X1 U9901 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14233) );
  NAND2_X1 U9902 ( .A1(n12234), .A2(n7430), .ZN(n10969) );
  NAND2_X1 U9903 ( .A1(n12120), .A2(n12620), .ZN(n8317) );
  NAND2_X1 U9904 ( .A1(n8303), .A2(n8302), .ZN(n8304) );
  INV_X1 U9905 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15320) );
  OR2_X1 U9906 ( .A1(n8181), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8195) );
  OR2_X1 U9907 ( .A1(n8164), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8179) );
  INV_X1 U9908 ( .A(n12760), .ZN(n9691) );
  NOR2_X1 U9909 ( .A1(n8639), .A2(n8262), .ZN(n9694) );
  INV_X1 U9910 ( .A(n11727), .ZN(n11729) );
  INV_X1 U9911 ( .A(n8991), .ZN(n8992) );
  INV_X1 U9912 ( .A(n12868), .ZN(n11705) );
  NAND2_X1 U9913 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n11548), .ZN(n11558) );
  NOR2_X1 U9914 ( .A1(n9647), .A2(n9646), .ZN(n9662) );
  NAND2_X1 U9915 ( .A1(n13004), .A2(n7679), .ZN(n13164) );
  OR2_X1 U9916 ( .A1(n10887), .A2(n10886), .ZN(n11197) );
  INV_X1 U9917 ( .A(n12988), .ZN(n12858) );
  NAND2_X1 U9918 ( .A1(n10638), .A2(n10639), .ZN(n10644) );
  INV_X1 U9919 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U9920 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n11337), .ZN(n11357) );
  NAND2_X1 U9921 ( .A1(n9842), .A2(n9841), .ZN(n14594) );
  OR2_X1 U9922 ( .A1(n10946), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9101) );
  INV_X1 U9923 ( .A(n9280), .ZN(n10703) );
  INV_X1 U9924 ( .A(n13656), .ZN(n13664) );
  AND2_X1 U9925 ( .A1(n9840), .A2(n13493), .ZN(n10128) );
  OR2_X1 U9926 ( .A1(n9717), .A2(n15325), .ZN(n9718) );
  INV_X1 U9927 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n14232) );
  INV_X1 U9928 ( .A(n10779), .ZN(n8299) );
  INV_X1 U9929 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15348) );
  OR2_X1 U9930 ( .A1(n8028), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U9931 ( .A1(n7692), .A2(n15255), .ZN(n8058) );
  OR2_X1 U9932 ( .A1(n7010), .A2(n15358), .ZN(n8162) );
  INV_X1 U9933 ( .A(n8195), .ZN(n12408) );
  INV_X1 U9934 ( .A(n12571), .ZN(n12534) );
  INV_X1 U9935 ( .A(n12565), .ZN(n12561) );
  OR2_X1 U9936 ( .A1(n7926), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7945) );
  INV_X1 U9937 ( .A(n10965), .ZN(n10960) );
  AND2_X1 U9938 ( .A1(n10854), .A2(n11093), .ZN(n10857) );
  INV_X1 U9939 ( .A(n12225), .ZN(n14355) );
  INV_X1 U9940 ( .A(n15099), .ZN(n15075) );
  INV_X1 U9941 ( .A(n9693), .ZN(n8355) );
  AND2_X1 U9942 ( .A1(n7765), .A2(n7764), .ZN(n8035) );
  AND2_X1 U9943 ( .A1(n7732), .A2(n7731), .ZN(n7812) );
  NOR2_X1 U9944 ( .A1(n11659), .A2(n11191), .ZN(n12807) );
  OR2_X1 U9945 ( .A1(n11208), .A2(n11193), .ZN(n11194) );
  XNOR2_X1 U9946 ( .A(n11786), .B(n11579), .ZN(n9332) );
  OR2_X1 U9947 ( .A1(n9678), .A2(n9657), .ZN(n9658) );
  AND2_X1 U9948 ( .A1(n11522), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n11533) );
  AND2_X1 U9949 ( .A1(n11510), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n11522) );
  INV_X1 U9950 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10193) );
  INV_X1 U9951 ( .A(n13133), .ZN(n13129) );
  NOR2_X1 U9952 ( .A1(n10836), .A2(n11868), .ZN(n10832) );
  NAND2_X1 U9953 ( .A1(n12892), .A2(n11812), .ZN(n9936) );
  NAND2_X1 U9954 ( .A1(n14805), .A2(n8917), .ZN(n13232) );
  NAND2_X1 U9955 ( .A1(n8963), .A2(n9685), .ZN(n11993) );
  INV_X1 U9956 ( .A(n11866), .ZN(n10836) );
  NAND2_X1 U9957 ( .A1(n8419), .A2(n8421), .ZN(n8420) );
  OR2_X1 U9958 ( .A1(n8784), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8817) );
  INV_X1 U9959 ( .A(n14050), .ZN(n13372) );
  INV_X1 U9960 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10708) );
  AND2_X1 U9961 ( .A1(n11418), .A2(n11417), .ZN(n13416) );
  INV_X1 U9962 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10355) );
  OR2_X1 U9963 ( .A1(n13462), .A2(n14704), .ZN(n14427) );
  AND2_X1 U9964 ( .A1(n11287), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11289) );
  INV_X1 U9965 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14249) );
  INV_X1 U9966 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14255) );
  INV_X1 U9967 ( .A(n13688), .ZN(n11597) );
  NOR2_X1 U9968 ( .A1(n9604), .A2(P1_U3086), .ZN(n13711) );
  NAND2_X1 U9969 ( .A1(n14059), .A2(n14058), .ZN(n14060) );
  INV_X1 U9970 ( .A(n11335), .ZN(n11283) );
  INV_X1 U9971 ( .A(n13559), .ZN(n13689) );
  INV_X1 U9972 ( .A(n13722), .ZN(n14405) );
  INV_X1 U9973 ( .A(n14604), .ZN(n13980) );
  INV_X1 U9974 ( .A(n13502), .ZN(n14593) );
  NAND2_X1 U9975 ( .A1(n14604), .A2(n13489), .ZN(n10143) );
  OR2_X1 U9976 ( .A1(n9167), .A2(n9166), .ZN(n14974) );
  INV_X1 U9977 ( .A(n12213), .ZN(n12189) );
  AND2_X1 U9978 ( .A1(n11115), .A2(n11114), .ZN(n11119) );
  AND3_X1 U9979 ( .A1(n8103), .A2(n8102), .A3(n8101), .ZN(n12535) );
  INV_X1 U9980 ( .A(n14911), .ZN(n15007) );
  AND2_X1 U9981 ( .A1(n9164), .A2(n9143), .ZN(n14997) );
  AND2_X1 U9982 ( .A1(n8214), .A2(n11093), .ZN(n15093) );
  OR2_X1 U9983 ( .A1(n15080), .A2(n15083), .ZN(n15034) );
  INV_X1 U9984 ( .A(n12579), .ZN(n15065) );
  NAND2_X1 U9985 ( .A1(n10064), .A2(n10979), .ZN(n10076) );
  INV_X1 U9986 ( .A(n15131), .ZN(n15151) );
  AND2_X1 U9987 ( .A1(n9696), .A2(n9695), .ZN(n10864) );
  OR2_X1 U9988 ( .A1(n15080), .A2(n15148), .ZN(n15160) );
  AND2_X1 U9989 ( .A1(n11121), .A2(n10853), .ZN(n15148) );
  NAND2_X1 U9990 ( .A1(n10853), .A2(n10965), .ZN(n15131) );
  INV_X1 U9991 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7888) );
  AND2_X1 U9992 ( .A1(n14867), .A2(n8898), .ZN(n8899) );
  AOI21_X1 U9993 ( .B1(n12034), .B2(n7019), .A(n12033), .ZN(n12036) );
  AND4_X1 U9994 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(
        n13042) );
  AND3_X1 U9995 ( .A1(n11538), .A2(n11537), .A3(n11536), .ZN(n12848) );
  OR2_X1 U9996 ( .A1(n8632), .A2(n12039), .ZN(n14742) );
  INV_X1 U9997 ( .A(n14742), .ZN(n14785) );
  NAND2_X1 U9998 ( .A1(n13017), .A2(n12001), .ZN(n13056) );
  INV_X1 U9999 ( .A(n6466), .ZN(n13228) );
  OAI21_X2 U10000 ( .B1(n9458), .B2(n9457), .A(n13232), .ZN(n13155) );
  NAND2_X1 U10001 ( .A1(n11993), .A2(n8897), .ZN(n14867) );
  INV_X1 U10002 ( .A(n12996), .ZN(n13260) );
  INV_X1 U10003 ( .A(n14850), .ZN(n13337) );
  NAND2_X1 U10004 ( .A1(n14881), .A2(n14871), .ZN(n14850) );
  INV_X1 U10005 ( .A(n14881), .ZN(n14875) );
  AND2_X1 U10006 ( .A1(n11272), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11287) );
  INV_X1 U10007 ( .A(n13659), .ZN(n9127) );
  INV_X1 U10008 ( .A(n13462), .ZN(n14387) );
  NAND2_X1 U10009 ( .A1(n9117), .A2(n14599), .ZN(n14415) );
  AND2_X1 U10010 ( .A1(n11312), .A2(n11311), .ZN(n13592) );
  INV_X1 U10011 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14237) );
  INV_X1 U10012 ( .A(n14538), .ZN(n14545) );
  INV_X1 U10013 ( .A(n14536), .ZN(n14548) );
  NAND2_X1 U10014 ( .A1(n7685), .A2(n13912), .ZN(n13911) );
  OAI21_X1 U10015 ( .B1(n11641), .B2(n11638), .A(n14599), .ZN(n9837) );
  AND2_X1 U10016 ( .A1(n6464), .A2(n14614), .ZN(n14609) );
  INV_X1 U10017 ( .A(n13982), .ZN(n14601) );
  AND2_X1 U10018 ( .A1(n6464), .A2(n14699), .ZN(n14623) );
  OR2_X1 U10019 ( .A1(n9833), .A2(n9834), .ZN(n10145) );
  NAND2_X1 U10020 ( .A1(n14647), .A2(n14646), .ZN(n14708) );
  NAND2_X1 U10021 ( .A1(n9846), .A2(n13647), .ZN(n14699) );
  INV_X1 U10022 ( .A(n14646), .ZN(n14697) );
  AND2_X1 U10023 ( .A1(n8678), .A2(n8603), .ZN(n10330) );
  AND2_X1 U10024 ( .A1(n14318), .A2(n14319), .ZN(n14473) );
  INV_X1 U10025 ( .A(n14974), .ZN(n14996) );
  NAND2_X1 U10026 ( .A1(n8353), .A2(n8354), .ZN(n12064) );
  INV_X1 U10027 ( .A(n12217), .ZN(n12191) );
  AND2_X1 U10028 ( .A1(n11115), .A2(n8199), .ZN(n12427) );
  INV_X1 U10029 ( .A(P3_U3897), .ZN(n12235) );
  INV_X1 U10030 ( .A(n14983), .ZN(n14993) );
  INV_X1 U10031 ( .A(n14997), .ZN(n14990) );
  INV_X1 U10032 ( .A(n12627), .ZN(n15049) );
  NAND2_X1 U10033 ( .A1(n9686), .A2(n11121), .ZN(n15053) );
  NAND2_X1 U10034 ( .A1(n15181), .A2(n15151), .ZN(n12705) );
  INV_X1 U10035 ( .A(n12061), .ZN(n12716) );
  OR2_X1 U10036 ( .A1(n12691), .A2(n12690), .ZN(n12744) );
  OR2_X1 U10037 ( .A1(n15162), .A2(n15131), .ZN(n12757) );
  AND2_X1 U10038 ( .A1(n8271), .A2(n8270), .ZN(n15162) );
  NAND2_X1 U10039 ( .A1(n8639), .A2(n12759), .ZN(n8640) );
  AND2_X1 U10040 ( .A1(n9141), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12759) );
  NOR2_X1 U10041 ( .A1(n8494), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12764) );
  INV_X1 U10042 ( .A(SI_17_), .ZN(n15257) );
  INV_X1 U10043 ( .A(SI_12_), .ZN(n15232) );
  INV_X1 U10044 ( .A(n9177), .ZN(n9319) );
  INV_X1 U10045 ( .A(n12875), .ZN(n12865) );
  INV_X1 U10046 ( .A(n13006), .ZN(n13035) );
  INV_X1 U10047 ( .A(n14790), .ZN(n9395) );
  INV_X1 U10048 ( .A(n14791), .ZN(n14733) );
  AND2_X1 U10049 ( .A1(n9730), .A2(n9418), .ZN(n9755) );
  INV_X1 U10050 ( .A(n14908), .ZN(n14905) );
  INV_X1 U10051 ( .A(n14887), .ZN(n14886) );
  NAND2_X1 U10052 ( .A1(n14805), .A2(n14800), .ZN(n14801) );
  INV_X1 U10053 ( .A(n14805), .ZN(n14803) );
  INV_X1 U10054 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13367) );
  INV_X1 U10055 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8786) );
  AND2_X1 U10056 ( .A1(n8792), .A2(n8760), .ZN(n14517) );
  OR2_X1 U10057 ( .A1(n13462), .A2(n14615), .ZN(n14426) );
  INV_X1 U10058 ( .A(n14415), .ZN(n14423) );
  NAND2_X1 U10059 ( .A1(n9607), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14436) );
  OR3_X1 U10060 ( .A1(n11363), .A2(n11362), .A3(n11361), .ZN(n13894) );
  INV_X1 U10061 ( .A(n14124), .ZN(n13994) );
  OR2_X1 U10062 ( .A1(n14499), .A2(n9126), .ZN(n14553) );
  OR2_X1 U10063 ( .A1(n14499), .A2(n7231), .ZN(n14538) );
  OR2_X1 U10064 ( .A1(n14499), .A2(n8802), .ZN(n14536) );
  NAND2_X1 U10065 ( .A1(n14730), .A2(n14701), .ZN(n14155) );
  OR2_X1 U10066 ( .A1(n10145), .A2(n10144), .ZN(n14727) );
  AND3_X1 U10067 ( .A1(n14712), .A2(n14711), .A3(n14710), .ZN(n14729) );
  XNOR2_X1 U10068 ( .A(n8443), .B(n8754), .ZN(n10747) );
  INV_X1 U10069 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9221) );
  AND2_X1 U10070 ( .A1(n12759), .A2(n8450), .ZN(P3_U3897) );
  OAI211_X1 U10071 ( .C1(n12214), .C2(n8397), .A(n8396), .B(n8395), .ZN(
        P3_U3165) );
  NOR2_X1 U10072 ( .A1(n8920), .A2(n8422), .ZN(P2_U3947) );
  INV_X2 U10073 ( .A(n13721), .ZN(P1_U4016) );
  INV_X1 U10074 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8272) );
  NOR2_X1 U10075 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7851) );
  NAND2_X1 U10076 ( .A1(n7851), .A2(n7852), .ZN(n7868) );
  INV_X1 U10077 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7694) );
  INV_X1 U10078 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7696) );
  INV_X1 U10079 ( .A(n8150), .ZN(n7698) );
  INV_X1 U10080 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15209) );
  INV_X1 U10081 ( .A(n8179), .ZN(n7699) );
  INV_X1 U10082 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15324) );
  NAND2_X1 U10083 ( .A1(n7699), .A2(n15324), .ZN(n8181) );
  NAND2_X1 U10084 ( .A1(n8181), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U10085 ( .A1(n8195), .A2(n7700), .ZN(n12428) );
  NAND4_X1 U10086 ( .A1(n7710), .A2(n7709), .A3(n7708), .A4(n7993), .ZN(n8201)
         );
  NAND2_X1 U10087 ( .A1(n7718), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7719) );
  MUX2_X1 U10088 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7719), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7720) );
  INV_X1 U10089 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n7727) );
  AND2_X2 U10090 ( .A1(n7724), .A2(n12048), .ZN(n7805) );
  NAND2_X1 U10091 ( .A1(n6482), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U10092 ( .A1(n7806), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7725) );
  OAI211_X1 U10093 ( .C1(n8142), .C2(n7727), .A(n7726), .B(n7725), .ZN(n7728)
         );
  INV_X1 U10094 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U10095 ( .A1(n8966), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U10096 ( .A1(n7730), .A2(n7729), .ZN(n7813) );
  NAND2_X1 U10097 ( .A1(n8976), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7732) );
  INV_X1 U10098 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U10099 ( .A1(n9282), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10100 ( .A1(n8559), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7734) );
  INV_X1 U10101 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U10102 ( .A1(n8499), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U10103 ( .A1(n9326), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7736) );
  INV_X1 U10104 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U10105 ( .A1(n9595), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U10106 ( .A1(n8574), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10107 ( .A1(n9770), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10108 ( .A1(n7859), .A2(n7858), .ZN(n7861) );
  NAND2_X1 U10109 ( .A1(n7861), .A2(n7738), .ZN(n7876) );
  NAND2_X1 U10110 ( .A1(n8523), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U10111 ( .A1(n7876), .A2(n7739), .ZN(n7741) );
  NAND2_X1 U10112 ( .A1(n8562), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U10113 ( .A1(n7002), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U10114 ( .A1(n8567), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7742) );
  INV_X1 U10115 ( .A(n7886), .ZN(n7743) );
  NAND2_X1 U10116 ( .A1(n8593), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U10117 ( .A1(n8590), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7745) );
  NAND2_X1 U10118 ( .A1(n7909), .A2(n7746), .ZN(n7921) );
  NAND2_X1 U10119 ( .A1(n8605), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U10120 ( .A1(n8610), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U10121 ( .A1(n7921), .A2(n7920), .ZN(n7923) );
  NAND2_X1 U10122 ( .A1(n7923), .A2(n7748), .ZN(n7933) );
  NAND2_X1 U10123 ( .A1(n8681), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U10124 ( .A1(n8677), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U10125 ( .A1(n7933), .A2(n7932), .ZN(n7935) );
  NAND2_X1 U10126 ( .A1(n8697), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7751) );
  XNOR2_X1 U10127 ( .A(n8786), .B(P2_DATAO_REG_12__SCAN_IN), .ZN(n7960) );
  INV_X1 U10128 ( .A(n7960), .ZN(n7752) );
  NAND2_X1 U10129 ( .A1(n8790), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7753) );
  NAND2_X1 U10130 ( .A1(n7976), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7757) );
  NAND2_X1 U10131 ( .A1(n7755), .A2(n10697), .ZN(n7756) );
  NAND2_X1 U10132 ( .A1(n9022), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U10133 ( .A1(n9221), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7761) );
  NAND2_X1 U10134 ( .A1(n9214), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7760) );
  NAND2_X1 U10135 ( .A1(n7761), .A2(n7760), .ZN(n8004) );
  NAND2_X1 U10136 ( .A1(n9013), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7763) );
  INV_X1 U10137 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U10138 ( .A1(n9019), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U10139 ( .A1(n9199), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7765) );
  INV_X1 U10140 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U10141 ( .A1(n9203), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7764) );
  INV_X1 U10142 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U10143 ( .A1(n9475), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7767) );
  INV_X1 U10144 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9480) );
  NAND2_X1 U10145 ( .A1(n9480), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7766) );
  INV_X1 U10146 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U10147 ( .A1(n9527), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n7769) );
  INV_X1 U10148 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U10149 ( .A1(n9525), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7768) );
  INV_X1 U10150 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11316) );
  NAND2_X1 U10151 ( .A1(n11316), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7772) );
  INV_X1 U10152 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11530) );
  NAND2_X1 U10153 ( .A1(n11530), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7771) );
  AND2_X1 U10154 ( .A1(n7772), .A2(n7771), .ZN(n8092) );
  INV_X1 U10155 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11543) );
  XNOR2_X1 U10156 ( .A(n11543), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10157 ( .A1(n11543), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7773) );
  XNOR2_X1 U10158 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8118) );
  INV_X1 U10159 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11576) );
  INV_X1 U10160 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U10161 ( .A1(n7774), .A2(n11664), .ZN(n7775) );
  NAND2_X1 U10162 ( .A1(n7776), .A2(n7775), .ZN(n8132) );
  INV_X1 U10163 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11672) );
  NAND2_X1 U10164 ( .A1(n11672), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7777) );
  INV_X1 U10165 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11395) );
  NAND2_X1 U10166 ( .A1(n11395), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7778) );
  INV_X1 U10167 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11419) );
  AND2_X1 U10168 ( .A1(n11419), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7779) );
  INV_X1 U10169 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11689) );
  NAND2_X1 U10170 ( .A1(n11689), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7780) );
  AND2_X1 U10171 ( .A1(n13367), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7781) );
  INV_X1 U10172 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14222) );
  NAND2_X1 U10173 ( .A1(n14222), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7782) );
  INV_X1 U10174 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n11722) );
  XNOR2_X1 U10175 ( .A(n11722), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n7784) );
  XNOR2_X1 U10176 ( .A(n8191), .B(n7784), .ZN(n11182) );
  NAND2_X1 U10177 ( .A1(n7785), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10178 ( .A1(n11182), .A2(n11108), .ZN(n7788) );
  INV_X1 U10179 ( .A(SI_28_), .ZN(n15243) );
  OR2_X1 U10180 ( .A1(n11100), .A2(n15243), .ZN(n7787) );
  NAND2_X1 U10181 ( .A1(n7797), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U10182 ( .A1(n7806), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U10183 ( .A1(n6478), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7789) );
  INV_X1 U10184 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7793) );
  INV_X1 U10185 ( .A(SI_1_), .ZN(n8460) );
  XNOR2_X1 U10186 ( .A(n7794), .B(n7803), .ZN(n8459) );
  NAND2_X1 U10187 ( .A1(n7797), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U10188 ( .A1(n7805), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10189 ( .A1(n7806), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U10190 ( .A1(n6479), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7798) );
  INV_X1 U10191 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U10192 ( .A1(n9061), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7802) );
  AND2_X1 U10193 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  NAND2_X1 U10194 ( .A1(n8494), .A2(SI_0_), .ZN(n8912) );
  OAI21_X1 U10195 ( .B1(n11332), .B2(n7804), .A(n8912), .ZN(n12772) );
  NAND2_X1 U10196 ( .A1(n15094), .A2(n9700), .ZN(n15089) );
  NAND2_X1 U10197 ( .A1(n7018), .A2(n7430), .ZN(n15073) );
  NAND2_X1 U10198 ( .A1(n6481), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U10199 ( .A1(n7797), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7810) );
  NAND2_X1 U10200 ( .A1(n7806), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7809) );
  NAND2_X1 U10201 ( .A1(n6478), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7808) );
  XNOR2_X1 U10202 ( .A(n7812), .B(n7813), .ZN(n8463) );
  OR2_X1 U10203 ( .A1(n8096), .A2(n8463), .ZN(n7816) );
  OR2_X1 U10204 ( .A1(n9140), .A2(n9177), .ZN(n7815) );
  NAND2_X1 U10205 ( .A1(n15097), .A2(n15082), .ZN(n7819) );
  NAND2_X1 U10206 ( .A1(n6482), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7823) );
  INV_X1 U10207 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15360) );
  NAND2_X1 U10208 ( .A1(n7797), .A2(n15360), .ZN(n7822) );
  NAND2_X1 U10209 ( .A1(n7806), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7821) );
  NAND2_X1 U10210 ( .A1(n6479), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7820) );
  AND4_X2 U10211 ( .A1(n7823), .A2(n7822), .A3(n7821), .A4(n7820), .ZN(n15071)
         );
  OR2_X1 U10212 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  NAND2_X1 U10213 ( .A1(n7827), .A2(n7826), .ZN(n8471) );
  OR2_X1 U10214 ( .A1(n8096), .A2(n8471), .ZN(n7831) );
  NAND2_X1 U10215 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n7828), .ZN(n7829) );
  XNOR2_X1 U10216 ( .A(n7829), .B(P3_IR_REG_3__SCAN_IN), .ZN(n14924) );
  OR2_X1 U10217 ( .A1(n9140), .A2(n14924), .ZN(n7830) );
  NAND2_X1 U10218 ( .A1(n12232), .A2(n9898), .ZN(n7834) );
  AND2_X1 U10219 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7835) );
  OR2_X1 U10220 ( .A1(n7835), .A2(n7851), .ZN(n10084) );
  NAND2_X1 U10221 ( .A1(n7797), .A2(n10084), .ZN(n7839) );
  NAND2_X1 U10222 ( .A1(n6481), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10223 ( .A1(n7806), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10224 ( .A1(n6479), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7836) );
  OR2_X1 U10225 ( .A1(n11100), .A2(SI_4_), .ZN(n7848) );
  XNOR2_X1 U10226 ( .A(n7841), .B(n7840), .ZN(n8469) );
  OR2_X1 U10227 ( .A1(n8096), .A2(n8469), .ZN(n7847) );
  NAND2_X1 U10228 ( .A1(n7842), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7843) );
  MUX2_X1 U10229 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7843), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7845) );
  AND2_X1 U10230 ( .A1(n7845), .A2(n7844), .ZN(n9172) );
  OR2_X1 U10231 ( .A1(n9140), .A2(n9172), .ZN(n7846) );
  NAND2_X1 U10232 ( .A1(n10247), .A2(n10083), .ZN(n10983) );
  INV_X1 U10233 ( .A(n10083), .ZN(n7849) );
  NAND2_X1 U10234 ( .A1(n12231), .A2(n7849), .ZN(n10984) );
  NAND2_X1 U10235 ( .A1(n10983), .A2(n10984), .ZN(n10075) );
  NAND2_X1 U10236 ( .A1(n12231), .A2(n10083), .ZN(n7850) );
  OR2_X1 U10237 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  NAND2_X1 U10238 ( .A1(n7868), .A2(n7853), .ZN(n10250) );
  NAND2_X1 U10239 ( .A1(n7797), .A2(n10250), .ZN(n7857) );
  NAND2_X1 U10240 ( .A1(n6482), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U10241 ( .A1(n7806), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U10242 ( .A1(n6479), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7854) );
  OR2_X1 U10243 ( .A1(n11100), .A2(SI_5_), .ZN(n7865) );
  OR2_X1 U10244 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  NAND2_X1 U10245 ( .A1(n7861), .A2(n7860), .ZN(n8474) );
  OR2_X1 U10246 ( .A1(n8096), .A2(n8474), .ZN(n7864) );
  NAND2_X1 U10247 ( .A1(n7844), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7862) );
  OR2_X1 U10248 ( .A1(n9140), .A2(n14940), .ZN(n7863) );
  NAND2_X1 U10249 ( .A1(n15055), .A2(n10249), .ZN(n10988) );
  INV_X1 U10250 ( .A(n15055), .ZN(n12230) );
  INV_X1 U10251 ( .A(n10249), .ZN(n15132) );
  NAND2_X1 U10252 ( .A1(n15055), .A2(n15132), .ZN(n7867) );
  NAND2_X1 U10253 ( .A1(n6482), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U10254 ( .A1(n7868), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U10255 ( .A1(n7880), .A2(n7869), .ZN(n15060) );
  NAND2_X1 U10256 ( .A1(n8045), .A2(n15060), .ZN(n7872) );
  NAND2_X1 U10257 ( .A1(n7806), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10258 ( .A1(n6479), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7870) );
  NOR2_X1 U10259 ( .A1(n7844), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7889) );
  OR2_X1 U10260 ( .A1(n7889), .A2(n8021), .ZN(n7874) );
  XNOR2_X1 U10261 ( .A(n7874), .B(n7888), .ZN(n9880) );
  INV_X1 U10262 ( .A(SI_6_), .ZN(n8465) );
  OR2_X1 U10263 ( .A1(n11100), .A2(n8465), .ZN(n7878) );
  XNOR2_X1 U10264 ( .A(n8562), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7875) );
  XNOR2_X1 U10265 ( .A(n7876), .B(n7875), .ZN(n8466) );
  OR2_X1 U10266 ( .A1(n8096), .A2(n8466), .ZN(n7877) );
  OAI211_X1 U10267 ( .C1(n9140), .C2(n9880), .A(n7878), .B(n7877), .ZN(n10276)
         );
  NAND2_X1 U10268 ( .A1(n10401), .A2(n10276), .ZN(n10995) );
  INV_X1 U10269 ( .A(n10401), .ZN(n12229) );
  INV_X1 U10270 ( .A(n10276), .ZN(n15063) );
  NAND2_X1 U10271 ( .A1(n12229), .A2(n15063), .ZN(n10994) );
  NAND2_X1 U10272 ( .A1(n10995), .A2(n10994), .ZN(n11134) );
  NAND2_X1 U10273 ( .A1(n12229), .A2(n10276), .ZN(n7879) );
  AND2_X1 U10274 ( .A1(n7880), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7881) );
  OR2_X1 U10275 ( .A1(n7881), .A2(n7895), .ZN(n12070) );
  NAND2_X1 U10276 ( .A1(n8045), .A2(n12070), .ZN(n7885) );
  NAND2_X1 U10277 ( .A1(n6481), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U10278 ( .A1(n7806), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7883) );
  NAND2_X1 U10279 ( .A1(n6479), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7882) );
  XNOR2_X1 U10280 ( .A(n7887), .B(n7886), .ZN(n8467) );
  OR2_X1 U10281 ( .A1(n8096), .A2(n8467), .ZN(n7893) );
  OR2_X1 U10282 ( .A1(n7010), .A2(SI_7_), .ZN(n7892) );
  NAND2_X1 U10283 ( .A1(n7889), .A2(n7888), .ZN(n7901) );
  NAND2_X1 U10284 ( .A1(n7901), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7890) );
  OR2_X1 U10285 ( .A1(n9140), .A2(n14956), .ZN(n7891) );
  NAND2_X1 U10286 ( .A1(n15056), .A2(n12069), .ZN(n10998) );
  INV_X1 U10287 ( .A(n12069), .ZN(n10406) );
  NAND2_X1 U10288 ( .A1(n12228), .A2(n10406), .ZN(n10999) );
  NAND2_X1 U10289 ( .A1(n10998), .A2(n10999), .ZN(n8224) );
  NAND2_X1 U10290 ( .A1(n12228), .A2(n12069), .ZN(n7894) );
  NAND2_X1 U10291 ( .A1(n6482), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7900) );
  NOR2_X1 U10292 ( .A1(n7895), .A2(n15348), .ZN(n7896) );
  OR2_X1 U10293 ( .A1(n7913), .A2(n7896), .ZN(n12093) );
  NAND2_X1 U10294 ( .A1(n8045), .A2(n12093), .ZN(n7899) );
  NAND2_X1 U10295 ( .A1(n7806), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7898) );
  NAND2_X1 U10296 ( .A1(n6479), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7897) );
  NAND4_X1 U10297 ( .A1(n7900), .A2(n7899), .A3(n7898), .A4(n7897), .ZN(n15044) );
  INV_X1 U10298 ( .A(n7937), .ZN(n7905) );
  NAND2_X1 U10299 ( .A1(n7902), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7903) );
  MUX2_X1 U10300 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7903), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n7904) );
  OR2_X1 U10301 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  NAND2_X1 U10302 ( .A1(n7909), .A2(n7908), .ZN(n8462) );
  OR2_X1 U10303 ( .A1(n8096), .A2(n8462), .ZN(n7911) );
  INV_X1 U10304 ( .A(SI_8_), .ZN(n8461) );
  OR2_X1 U10305 ( .A1(n11100), .A2(n8461), .ZN(n7910) );
  OAI211_X1 U10306 ( .C1(n9140), .C2(n10234), .A(n7911), .B(n7910), .ZN(n12092) );
  AND2_X1 U10307 ( .A1(n15044), .A2(n12092), .ZN(n15036) );
  NAND2_X1 U10308 ( .A1(n6481), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7918) );
  OR2_X1 U10309 ( .A1(n7913), .A2(n7912), .ZN(n7914) );
  AND2_X1 U10310 ( .A1(n7926), .A2(n7914), .ZN(n15054) );
  INV_X1 U10311 ( .A(n15054), .ZN(n10662) );
  NAND2_X1 U10312 ( .A1(n8045), .A2(n10662), .ZN(n7917) );
  NAND2_X1 U10313 ( .A1(n7806), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10314 ( .A1(n6479), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7915) );
  OR2_X1 U10315 ( .A1(n7937), .A2(n8021), .ZN(n7919) );
  XNOR2_X1 U10316 ( .A(n7919), .B(P3_IR_REG_9__SCAN_IN), .ZN(n10571) );
  OR2_X1 U10317 ( .A1(n11100), .A2(SI_9_), .ZN(n7925) );
  OR2_X1 U10318 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  AND2_X1 U10319 ( .A1(n7923), .A2(n7922), .ZN(n8476) );
  OR2_X1 U10320 ( .A1(n8096), .A2(n8476), .ZN(n7924) );
  OAI211_X1 U10321 ( .C1(n10571), .C2(n9140), .A(n7925), .B(n7924), .ZN(n15048) );
  INV_X1 U10322 ( .A(n15048), .ZN(n15152) );
  AND2_X1 U10323 ( .A1(n15024), .A2(n15152), .ZN(n7943) );
  OR2_X1 U10324 ( .A1(n15036), .A2(n7943), .ZN(n15017) );
  NAND2_X1 U10325 ( .A1(n7926), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U10326 ( .A1(n7945), .A2(n7927), .ZN(n15028) );
  NAND2_X1 U10327 ( .A1(n8045), .A2(n15028), .ZN(n7931) );
  NAND2_X1 U10328 ( .A1(n6482), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10329 ( .A1(n7806), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10330 ( .A1(n6479), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7928) );
  OR2_X1 U10331 ( .A1(n7933), .A2(n7932), .ZN(n7934) );
  AND2_X1 U10332 ( .A1(n7935), .A2(n7934), .ZN(n8478) );
  OR2_X1 U10333 ( .A1(n8478), .A2(n8096), .ZN(n7941) );
  OR2_X1 U10334 ( .A1(n11100), .A2(SI_10_), .ZN(n7940) );
  INV_X1 U10335 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10336 ( .A1(n7937), .A2(n7936), .ZN(n7953) );
  NAND2_X1 U10337 ( .A1(n7953), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7938) );
  XNOR2_X1 U10338 ( .A(n7938), .B(P3_IR_REG_10__SCAN_IN), .ZN(n14982) );
  OR2_X1 U10339 ( .A1(n9140), .A2(n14982), .ZN(n7939) );
  AND2_X1 U10340 ( .A1(n8302), .A2(n10785), .ZN(n7944) );
  OR2_X1 U10341 ( .A1(n15017), .A2(n7944), .ZN(n7942) );
  INV_X1 U10342 ( .A(n12092), .ZN(n10432) );
  NAND2_X1 U10343 ( .A1(n10659), .A2(n10432), .ZN(n15038) );
  XNOR2_X1 U10344 ( .A(n15024), .B(n15048), .ZN(n15042) );
  AND2_X1 U10345 ( .A1(n15038), .A2(n15042), .ZN(n15039) );
  OR2_X1 U10346 ( .A1(n7943), .A2(n15039), .ZN(n15018) );
  NAND2_X1 U10347 ( .A1(n12179), .A2(n10785), .ZN(n11012) );
  INV_X1 U10348 ( .A(n10785), .ZN(n15029) );
  NAND2_X1 U10349 ( .A1(n8302), .A2(n15029), .ZN(n11011) );
  NAND2_X1 U10350 ( .A1(n11012), .A2(n11011), .ZN(n15022) );
  NAND2_X1 U10351 ( .A1(n6482), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10352 ( .A1(n7945), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U10353 ( .A1(n7968), .A2(n7946), .ZN(n12175) );
  NAND2_X1 U10354 ( .A1(n8045), .A2(n12175), .ZN(n7949) );
  NAND2_X1 U10355 ( .A1(n7806), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U10356 ( .A1(n6479), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7947) );
  XNOR2_X1 U10357 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7951) );
  XNOR2_X1 U10358 ( .A(n7952), .B(n7951), .ZN(n8481) );
  NAND2_X1 U10359 ( .A1(n8481), .A2(n11108), .ZN(n7956) );
  OAI21_X1 U10360 ( .B1(n7953), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7954) );
  XNOR2_X1 U10361 ( .A(n7954), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12251) );
  INV_X1 U10362 ( .A(n12251), .ZN(n10578) );
  AOI22_X1 U10363 ( .A1(n8070), .A2(n8688), .B1(n8136), .B2(n10578), .ZN(n7955) );
  NAND2_X1 U10364 ( .A1(n7956), .A2(n7955), .ZN(n10874) );
  NAND2_X1 U10365 ( .A1(n12173), .A2(n10874), .ZN(n7957) );
  NAND2_X1 U10366 ( .A1(n10666), .A2(n7957), .ZN(n7959) );
  INV_X1 U10367 ( .A(n10874), .ZN(n12181) );
  NAND2_X1 U10368 ( .A1(n15025), .A2(n12181), .ZN(n7958) );
  XNOR2_X1 U10369 ( .A(n7961), .B(n7960), .ZN(n8575) );
  NAND2_X1 U10370 ( .A1(n8575), .A2(n11108), .ZN(n7967) );
  NOR2_X1 U10371 ( .A1(n7962), .A2(n8021), .ZN(n7963) );
  MUX2_X1 U10372 ( .A(n8021), .B(n7963), .S(P3_IR_REG_12__SCAN_IN), .Z(n7965)
         );
  OR2_X1 U10373 ( .A1(n7965), .A2(n7964), .ZN(n14992) );
  INV_X1 U10374 ( .A(n14992), .ZN(n12253) );
  AOI22_X1 U10375 ( .A1(n8070), .A2(SI_12_), .B1(n8136), .B2(n12253), .ZN(
        n7966) );
  NAND2_X1 U10376 ( .A1(n7968), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10377 ( .A1(n7983), .A2(n7969), .ZN(n12111) );
  NAND2_X1 U10378 ( .A1(n8045), .A2(n12111), .ZN(n7973) );
  NAND2_X1 U10379 ( .A1(n6481), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U10380 ( .A1(n7806), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U10381 ( .A1(n6479), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7970) );
  NAND4_X1 U10382 ( .A1(n7973), .A2(n7972), .A3(n7971), .A4(n7970), .ZN(n12227) );
  NAND2_X1 U10383 ( .A1(n14366), .A2(n12227), .ZN(n11015) );
  INV_X1 U10384 ( .A(n14366), .ZN(n7974) );
  NAND2_X1 U10385 ( .A1(n14356), .A2(n7974), .ZN(n10956) );
  NAND2_X1 U10386 ( .A1(n11015), .A2(n10956), .ZN(n11140) );
  NAND2_X1 U10387 ( .A1(n7974), .A2(n12227), .ZN(n7975) );
  XNOR2_X1 U10388 ( .A(n7976), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U10389 ( .A1(n8641), .A2(n11108), .ZN(n7982) );
  NOR2_X1 U10390 ( .A1(n7964), .A2(n8021), .ZN(n7977) );
  MUX2_X1 U10391 ( .A(n8021), .B(n7977), .S(P3_IR_REG_13__SCAN_IN), .Z(n7980)
         );
  AOI22_X1 U10392 ( .A1(n8070), .A2(n8999), .B1(n8136), .B2(n12280), .ZN(n7981) );
  NAND2_X1 U10393 ( .A1(n7982), .A2(n7981), .ZN(n14357) );
  NAND2_X1 U10394 ( .A1(n6482), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10395 ( .A1(n7983), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U10396 ( .A1(n7997), .A2(n7984), .ZN(n14358) );
  NAND2_X1 U10397 ( .A1(n8045), .A2(n14358), .ZN(n7987) );
  NAND2_X1 U10398 ( .A1(n7806), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10399 ( .A1(n6479), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7985) );
  NOR2_X1 U10400 ( .A1(n14357), .A2(n12619), .ZN(n7990) );
  NAND2_X1 U10401 ( .A1(n14357), .A2(n12619), .ZN(n7989) );
  XNOR2_X1 U10402 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n7991) );
  XNOR2_X1 U10403 ( .A(n7992), .B(n7991), .ZN(n8711) );
  NAND2_X1 U10404 ( .A1(n8711), .A2(n11108), .ZN(n7996) );
  XNOR2_X1 U10405 ( .A(n7994), .B(n7993), .ZN(n12289) );
  AOI22_X1 U10406 ( .A1(n8070), .A2(n15322), .B1(n8136), .B2(n12289), .ZN(
        n7995) );
  NAND2_X1 U10407 ( .A1(n7996), .A2(n7995), .ZN(n12756) );
  NAND2_X1 U10408 ( .A1(n6481), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U10409 ( .A1(n7997), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U10410 ( .A1(n8011), .A2(n7998), .ZN(n11218) );
  NAND2_X1 U10411 ( .A1(n8045), .A2(n11218), .ZN(n8001) );
  NAND2_X1 U10412 ( .A1(n7806), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10413 ( .A1(n6479), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7999) );
  NAND4_X1 U10414 ( .A1(n8002), .A2(n8001), .A3(n8000), .A4(n7999), .ZN(n12225) );
  OR2_X1 U10415 ( .A1(n12756), .A2(n12225), .ZN(n11027) );
  NAND2_X1 U10416 ( .A1(n12756), .A2(n12225), .ZN(n11023) );
  OR2_X1 U10417 ( .A1(n12756), .A2(n14355), .ZN(n8003) );
  NAND2_X1 U10418 ( .A1(n8005), .A2(n8004), .ZN(n8006) );
  NAND2_X1 U10419 ( .A1(n8007), .A2(n8006), .ZN(n8761) );
  NAND2_X1 U10420 ( .A1(n8761), .A2(n11108), .ZN(n8010) );
  NAND2_X1 U10421 ( .A1(n6512), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8008) );
  XNOR2_X1 U10422 ( .A(n8008), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12331) );
  INV_X1 U10423 ( .A(n12331), .ZN(n12305) );
  AOI22_X1 U10424 ( .A1(n8070), .A2(n9208), .B1(n8136), .B2(n12305), .ZN(n8009) );
  NAND2_X1 U10425 ( .A1(n6481), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10426 ( .A1(n7806), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U10427 ( .A1(n8011), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10428 ( .A1(n8028), .A2(n8012), .ZN(n12613) );
  NAND2_X1 U10429 ( .A1(n8045), .A2(n12613), .ZN(n8014) );
  NAND2_X1 U10430 ( .A1(n6479), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8013) );
  OR2_X1 U10431 ( .A1(n8018), .A2(n8017), .ZN(n8019) );
  NAND2_X1 U10432 ( .A1(n8020), .A2(n8019), .ZN(n8816) );
  OR2_X1 U10433 ( .A1(n8816), .A2(n8096), .ZN(n8027) );
  OR2_X1 U10434 ( .A1(n8024), .A2(n8021), .ZN(n8022) );
  INV_X1 U10435 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8023) );
  MUX2_X1 U10436 ( .A(n8022), .B(P3_IR_REG_31__SCAN_IN), .S(n8023), .Z(n8025)
         );
  AOI22_X1 U10437 ( .A1(n8070), .A2(SI_16_), .B1(n8136), .B2(n12333), .ZN(
        n8026) );
  NAND2_X1 U10438 ( .A1(n8027), .A2(n8026), .ZN(n12127) );
  NAND2_X1 U10439 ( .A1(n6482), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10440 ( .A1(n8028), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10441 ( .A1(n8043), .A2(n8029), .ZN(n12602) );
  NAND2_X1 U10442 ( .A1(n8045), .A2(n12602), .ZN(n8032) );
  NAND2_X1 U10443 ( .A1(n7806), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10444 ( .A1(n6479), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8030) );
  NAND4_X1 U10445 ( .A1(n8033), .A2(n8032), .A3(n8031), .A4(n8030), .ZN(n12583) );
  AND2_X1 U10446 ( .A1(n12127), .A2(n12583), .ZN(n8034) );
  OR2_X1 U10447 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  NAND2_X1 U10448 ( .A1(n8038), .A2(n8037), .ZN(n8869) );
  NAND2_X1 U10449 ( .A1(n8869), .A2(n11108), .ZN(n8042) );
  MUX2_X1 U10450 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8039), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8040) );
  NAND2_X1 U10451 ( .A1(n8040), .A2(n7683), .ZN(n12371) );
  AOI22_X1 U10452 ( .A1(n8070), .A2(n15257), .B1(n8136), .B2(n12371), .ZN(
        n8041) );
  NAND2_X1 U10453 ( .A1(n6481), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10454 ( .A1(n8043), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8044) );
  NAND2_X1 U10455 ( .A1(n8058), .A2(n8044), .ZN(n12591) );
  NAND2_X1 U10456 ( .A1(n8045), .A2(n12591), .ZN(n8048) );
  NAND2_X1 U10457 ( .A1(n7806), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10458 ( .A1(n6479), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8046) );
  NAND4_X1 U10459 ( .A1(n8049), .A2(n8048), .A3(n8047), .A4(n8046), .ZN(n12570) );
  NAND2_X1 U10460 ( .A1(n12689), .A2(n12570), .ZN(n11041) );
  INV_X1 U10461 ( .A(n12570), .ZN(n12598) );
  OR2_X1 U10462 ( .A1(n12689), .A2(n12598), .ZN(n8050) );
  OR2_X1 U10463 ( .A1(n8052), .A2(n8051), .ZN(n8053) );
  NAND2_X1 U10464 ( .A1(n8054), .A2(n8053), .ZN(n9020) );
  OR2_X1 U10465 ( .A1(n9020), .A2(n8096), .ZN(n8057) );
  NAND2_X1 U10466 ( .A1(n7683), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8055) );
  XNOR2_X1 U10467 ( .A(n8055), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U10468 ( .A1(n8070), .A2(SI_18_), .B1(n8136), .B2(n12395), .ZN(
        n8056) );
  NAND2_X1 U10469 ( .A1(n6481), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U10470 ( .A1(n7806), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8062) );
  NAND2_X1 U10471 ( .A1(n8058), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10472 ( .A1(n8073), .A2(n8059), .ZN(n12186) );
  NAND2_X1 U10473 ( .A1(n8045), .A2(n12186), .ZN(n8061) );
  NAND2_X1 U10474 ( .A1(n6479), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10475 ( .A1(n12681), .A2(n8322), .ZN(n11044) );
  OR2_X1 U10476 ( .A1(n12681), .A2(n12584), .ZN(n8064) );
  NAND2_X1 U10477 ( .A1(n12568), .A2(n8064), .ZN(n12547) );
  OR2_X1 U10478 ( .A1(n8066), .A2(n8065), .ZN(n8067) );
  NAND2_X1 U10479 ( .A1(n8068), .A2(n8067), .ZN(n9246) );
  OR2_X1 U10480 ( .A1(n9246), .A2(n8096), .ZN(n8072) );
  AOI22_X1 U10481 ( .A1(n8070), .A2(SI_19_), .B1(n6480), .B2(n8136), .ZN(n8071) );
  NAND2_X1 U10482 ( .A1(n8073), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10483 ( .A1(n8085), .A2(n8074), .ZN(n12554) );
  NAND2_X1 U10484 ( .A1(n12554), .A2(n8045), .ZN(n8078) );
  NAND2_X1 U10485 ( .A1(n6482), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10486 ( .A1(n7806), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10487 ( .A1(n6479), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8075) );
  NAND4_X1 U10488 ( .A1(n8078), .A2(n8077), .A3(n8076), .A4(n8075), .ZN(n12571) );
  NOR2_X1 U10489 ( .A1(n12677), .A2(n12571), .ZN(n8079) );
  INV_X1 U10490 ( .A(n12677), .ZN(n12556) );
  NAND2_X1 U10491 ( .A1(n8080), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U10492 ( .A1(n8082), .A2(n8081), .ZN(n9451) );
  OR2_X1 U10493 ( .A1(n9451), .A2(n8096), .ZN(n8084) );
  OR2_X1 U10494 ( .A1(n11100), .A2(n15325), .ZN(n8083) );
  NAND2_X1 U10495 ( .A1(n8085), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8086) );
  NAND2_X1 U10496 ( .A1(n8099), .A2(n8086), .ZN(n12542) );
  NAND2_X1 U10497 ( .A1(n12542), .A2(n8045), .ZN(n8089) );
  AOI22_X1 U10498 ( .A1(n6482), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n7806), .B2(
        P3_REG0_REG_20__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10499 ( .A1(n6479), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10500 ( .A1(n12536), .A2(n12522), .ZN(n11057) );
  NAND2_X1 U10501 ( .A1(n11056), .A2(n11057), .ZN(n12538) );
  NAND2_X1 U10502 ( .A1(n12536), .A2(n12548), .ZN(n8090) );
  OR2_X1 U10503 ( .A1(n8093), .A2(n8092), .ZN(n8094) );
  NAND2_X1 U10504 ( .A1(n8095), .A2(n8094), .ZN(n9633) );
  INV_X1 U10505 ( .A(SI_21_), .ZN(n15361) );
  NAND2_X1 U10506 ( .A1(n8099), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U10507 ( .A1(n8109), .A2(n8100), .ZN(n12527) );
  NAND2_X1 U10508 ( .A1(n12527), .A2(n8045), .ZN(n8103) );
  AOI22_X1 U10509 ( .A1(n6482), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n7806), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U10510 ( .A1(n6479), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8101) );
  OR2_X1 U10511 ( .A1(n12526), .A2(n12535), .ZN(n11061) );
  NAND2_X1 U10512 ( .A1(n12526), .A2(n12535), .ZN(n11060) );
  INV_X1 U10513 ( .A(n12535), .ZN(n12508) );
  OR2_X1 U10514 ( .A1(n12526), .A2(n12508), .ZN(n8104) );
  XNOR2_X1 U10515 ( .A(n8106), .B(n8105), .ZN(n9721) );
  NAND2_X1 U10516 ( .A1(n9721), .A2(n11108), .ZN(n8108) );
  INV_X1 U10517 ( .A(SI_22_), .ZN(n15228) );
  OR2_X1 U10518 ( .A1(n11100), .A2(n15228), .ZN(n8107) );
  NAND2_X1 U10519 ( .A1(n8109), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U10520 ( .A1(n8122), .A2(n8110), .ZN(n12513) );
  NAND2_X1 U10521 ( .A1(n12513), .A2(n8045), .ZN(n8116) );
  INV_X1 U10522 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10523 ( .A1(n6481), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U10524 ( .A1(n7806), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8111) );
  OAI211_X1 U10525 ( .C1(n8113), .C2(n8142), .A(n8112), .B(n8111), .ZN(n8114)
         );
  INV_X1 U10526 ( .A(n8114), .ZN(n8115) );
  NAND2_X1 U10527 ( .A1(n12665), .A2(n12496), .ZN(n8117) );
  XNOR2_X1 U10528 ( .A(n8119), .B(n8118), .ZN(n9966) );
  NAND2_X1 U10529 ( .A1(n9966), .A2(n11108), .ZN(n8121) );
  INV_X1 U10530 ( .A(SI_23_), .ZN(n9968) );
  OR2_X1 U10531 ( .A1(n7010), .A2(n9968), .ZN(n8120) );
  NAND2_X1 U10532 ( .A1(n8122), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10533 ( .A1(n8137), .A2(n8123), .ZN(n12502) );
  NAND2_X1 U10534 ( .A1(n12502), .A2(n8045), .ZN(n8129) );
  INV_X1 U10535 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U10536 ( .A1(n6481), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8125) );
  NAND2_X1 U10537 ( .A1(n7806), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8124) );
  OAI211_X1 U10538 ( .C1(n8126), .C2(n8142), .A(n8125), .B(n8124), .ZN(n8127)
         );
  INV_X1 U10539 ( .A(n8127), .ZN(n8128) );
  XNOR2_X1 U10540 ( .A(n12501), .B(n12509), .ZN(n12499) );
  NAND2_X1 U10541 ( .A1(n12501), .A2(n12509), .ZN(n8131) );
  NAND2_X1 U10542 ( .A1(n8132), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10543 ( .A1(n8134), .A2(n8133), .ZN(n8135) );
  NAND2_X1 U10544 ( .A1(n8137), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U10545 ( .A1(n8150), .A2(n8138), .ZN(n12490) );
  NAND2_X1 U10546 ( .A1(n12490), .A2(n8045), .ZN(n8145) );
  INV_X1 U10547 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U10548 ( .A1(n6482), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10549 ( .A1(n7806), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8139) );
  OAI211_X1 U10550 ( .C1(n8142), .C2(n8141), .A(n8140), .B(n8139), .ZN(n8143)
         );
  INV_X1 U10551 ( .A(n8143), .ZN(n8144) );
  XNOR2_X1 U10552 ( .A(n11672), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8146) );
  XNOR2_X1 U10553 ( .A(n8147), .B(n8146), .ZN(n10493) );
  NAND2_X1 U10554 ( .A1(n10493), .A2(n11108), .ZN(n8149) );
  INV_X1 U10555 ( .A(SI_25_), .ZN(n10536) );
  OR2_X1 U10556 ( .A1(n11100), .A2(n10536), .ZN(n8148) );
  NAND2_X1 U10557 ( .A1(n8150), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10558 ( .A1(n8164), .A2(n8151), .ZN(n12473) );
  NAND2_X1 U10559 ( .A1(n12473), .A2(n8045), .ZN(n8157) );
  INV_X1 U10560 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U10561 ( .A1(n6481), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10562 ( .A1(n7806), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8152) );
  OAI211_X1 U10563 ( .C1(n8154), .C2(n8142), .A(n8153), .B(n8152), .ZN(n8155)
         );
  INV_X1 U10564 ( .A(n8155), .ZN(n8156) );
  NAND2_X1 U10565 ( .A1(n12653), .A2(n12480), .ZN(n11075) );
  NAND2_X1 U10566 ( .A1(n11080), .A2(n11075), .ZN(n12467) );
  AND2_X1 U10567 ( .A1(n12486), .A2(n12467), .ZN(n8158) );
  INV_X1 U10568 ( .A(n12467), .ZN(n11074) );
  INV_X1 U10569 ( .A(n12725), .ZN(n8231) );
  NAND2_X1 U10570 ( .A1(n8231), .A2(n12469), .ZN(n12465) );
  NAND2_X1 U10571 ( .A1(n12653), .A2(n12224), .ZN(n8159) );
  XNOR2_X1 U10572 ( .A(n11689), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8160) );
  XNOR2_X1 U10573 ( .A(n8161), .B(n8160), .ZN(n10630) );
  NAND2_X1 U10574 ( .A1(n10630), .A2(n11108), .ZN(n8163) );
  INV_X1 U10575 ( .A(SI_26_), .ZN(n15358) );
  NAND2_X1 U10576 ( .A1(n8164), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10577 ( .A1(n8179), .A2(n8165), .ZN(n12459) );
  NAND2_X1 U10578 ( .A1(n12459), .A2(n8045), .ZN(n8171) );
  INV_X1 U10579 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10580 ( .A1(n6482), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U10581 ( .A1(n7806), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8166) );
  OAI211_X1 U10582 ( .C1(n8168), .C2(n8142), .A(n8167), .B(n8166), .ZN(n8169)
         );
  INV_X1 U10583 ( .A(n8169), .ZN(n8170) );
  OR2_X1 U10584 ( .A1(n12648), .A2(n12223), .ZN(n8172) );
  NAND2_X1 U10585 ( .A1(n12450), .A2(n8172), .ZN(n8174) );
  NAND2_X1 U10586 ( .A1(n12648), .A2(n12223), .ZN(n8173) );
  XNOR2_X1 U10587 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8175) );
  XNOR2_X1 U10588 ( .A(n8176), .B(n8175), .ZN(n11753) );
  NAND2_X1 U10589 ( .A1(n11753), .A2(n11108), .ZN(n8178) );
  INV_X1 U10590 ( .A(SI_27_), .ZN(n15347) );
  NAND2_X1 U10591 ( .A1(n8179), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U10592 ( .A1(n8181), .A2(n8180), .ZN(n12443) );
  NAND2_X1 U10593 ( .A1(n12443), .A2(n8045), .ZN(n8187) );
  INV_X1 U10594 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10595 ( .A1(n6481), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U10596 ( .A1(n7806), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8182) );
  OAI211_X1 U10597 ( .C1(n8184), .C2(n8142), .A(n8183), .B(n8182), .ZN(n8185)
         );
  INV_X1 U10598 ( .A(n8185), .ZN(n8186) );
  XNOR2_X1 U10599 ( .A(n12444), .B(n12425), .ZN(n12433) );
  OR2_X1 U10600 ( .A1(n12444), .A2(n12425), .ZN(n8188) );
  NAND2_X1 U10601 ( .A1(n12061), .A2(n12440), .ZN(n8232) );
  NOR2_X1 U10602 ( .A1(n11722), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10603 ( .A1(n11722), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8192) );
  XNOR2_X1 U10604 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n11097) );
  XNOR2_X1 U10605 ( .A(n11099), .B(n11097), .ZN(n12767) );
  NAND2_X1 U10606 ( .A1(n12767), .A2(n11108), .ZN(n8194) );
  INV_X1 U10607 ( .A(SI_29_), .ZN(n15364) );
  OR2_X1 U10608 ( .A1(n7010), .A2(n15364), .ZN(n8193) );
  NAND2_X1 U10609 ( .A1(n12408), .A2(n8045), .ZN(n11115) );
  INV_X1 U10610 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12415) );
  NAND2_X1 U10611 ( .A1(n6481), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8197) );
  NAND2_X1 U10612 ( .A1(n7806), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8196) );
  OAI211_X1 U10613 ( .C1(n8142), .C2(n12415), .A(n8197), .B(n8196), .ZN(n8198)
         );
  INV_X1 U10614 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U10615 ( .A1(n12417), .A2(n12427), .ZN(n11123) );
  XNOR2_X1 U10616 ( .A(n8200), .B(n11147), .ZN(n8211) );
  NAND2_X1 U10617 ( .A1(n8263), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8205) );
  INV_X2 U10618 ( .A(n10853), .ZN(n11160) );
  NAND2_X1 U10619 ( .A1(n6480), .A2(n11160), .ZN(n8268) );
  NAND2_X1 U10620 ( .A1(n8209), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8206) );
  MUX2_X1 U10621 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8206), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8207) );
  NAND2_X1 U10622 ( .A1(n6534), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8208) );
  MUX2_X1 U10623 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8208), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8210) );
  INV_X1 U10624 ( .A(n9452), .ZN(n10852) );
  NAND2_X1 U10625 ( .A1(n10960), .A2(n10852), .ZN(n11154) );
  NAND2_X1 U10626 ( .A1(n8211), .A2(n15099), .ZN(n8222) );
  INV_X1 U10627 ( .A(n8212), .ZN(n11157) );
  NAND2_X1 U10628 ( .A1(n11157), .A2(n6812), .ZN(n9142) );
  NAND2_X1 U10629 ( .A1(n9140), .A2(n9142), .ZN(n8363) );
  INV_X1 U10630 ( .A(n8363), .ZN(n8214) );
  INV_X4 U10631 ( .A(n6475), .ZN(n11093) );
  INV_X1 U10632 ( .A(n12440), .ZN(n12222) );
  INV_X1 U10633 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8217) );
  NAND2_X1 U10634 ( .A1(n6482), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10635 ( .A1(n7806), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8215) );
  OAI211_X1 U10636 ( .C1(n8217), .C2(n8142), .A(n8216), .B(n8215), .ZN(n8218)
         );
  INV_X1 U10637 ( .A(n8218), .ZN(n8219) );
  NAND2_X1 U10638 ( .A1(n11115), .A2(n8219), .ZN(n12221) );
  AND2_X1 U10639 ( .A1(n11157), .A2(P3_B_REG_SCAN_IN), .ZN(n8220) );
  NOR2_X1 U10640 ( .A1(n15096), .A2(n8220), .ZN(n12406) );
  AOI22_X1 U10641 ( .A1(n15093), .A2(n12222), .B1(n12221), .B2(n12406), .ZN(
        n8221) );
  INV_X1 U10642 ( .A(n9700), .ZN(n12707) );
  NAND2_X1 U10643 ( .A1(n15088), .A2(n10969), .ZN(n8280) );
  NAND2_X1 U10644 ( .A1(n8280), .A2(n10968), .ZN(n15070) );
  NAND2_X1 U10645 ( .A1(n10062), .A2(n11133), .ZN(n10064) );
  INV_X1 U10646 ( .A(n10075), .ZN(n11131) );
  NAND2_X1 U10647 ( .A1(n10076), .A2(n11131), .ZN(n8223) );
  INV_X1 U10648 ( .A(n11134), .ZN(n15061) );
  NAND2_X1 U10649 ( .A1(n10397), .A2(n10998), .ZN(n10428) );
  NAND2_X1 U10650 ( .A1(n10659), .A2(n12092), .ZN(n11002) );
  NAND2_X1 U10651 ( .A1(n15044), .A2(n10432), .ZN(n11003) );
  NAND2_X1 U10652 ( .A1(n10428), .A2(n11129), .ZN(n8225) );
  NAND2_X1 U10653 ( .A1(n12173), .A2(n12181), .ZN(n10955) );
  NAND2_X1 U10654 ( .A1(n15025), .A2(n10874), .ZN(n11014) );
  INV_X1 U10655 ( .A(n11140), .ZN(n10753) );
  NAND2_X1 U10656 ( .A1(n10752), .A2(n10956), .ZN(n14351) );
  NOR2_X1 U10657 ( .A1(n14357), .A2(n12226), .ZN(n10957) );
  NAND2_X1 U10658 ( .A1(n14357), .A2(n12226), .ZN(n10951) );
  INV_X1 U10659 ( .A(n11023), .ZN(n8226) );
  NAND2_X1 U10660 ( .A1(n12752), .A2(n8315), .ZN(n11024) );
  INV_X1 U10661 ( .A(n12583), .ZN(n12610) );
  OR2_X1 U10662 ( .A1(n12127), .A2(n12610), .ZN(n11036) );
  NAND2_X1 U10663 ( .A1(n12127), .A2(n12610), .ZN(n11035) );
  NAND2_X1 U10664 ( .A1(n12601), .A2(n12600), .ZN(n12599) );
  INV_X1 U10665 ( .A(n12560), .ZN(n11043) );
  NOR2_X1 U10666 ( .A1(n12561), .A2(n11043), .ZN(n8227) );
  OR2_X1 U10667 ( .A1(n12677), .A2(n12534), .ZN(n11052) );
  NAND2_X1 U10668 ( .A1(n12677), .A2(n12534), .ZN(n12537) );
  NAND2_X1 U10669 ( .A1(n11052), .A2(n12537), .ZN(n12552) );
  INV_X1 U10670 ( .A(n12537), .ZN(n8229) );
  NOR2_X1 U10671 ( .A1(n12538), .A2(n8229), .ZN(n8230) );
  NAND2_X1 U10672 ( .A1(n12550), .A2(n8230), .ZN(n12540) );
  NAND2_X1 U10673 ( .A1(n12540), .A2(n11056), .ZN(n12525) );
  NAND2_X1 U10674 ( .A1(n12665), .A2(n12523), .ZN(n11064) );
  NAND2_X1 U10675 ( .A1(n12500), .A2(n12499), .ZN(n12485) );
  INV_X1 U10676 ( .A(n12509), .ZN(n12479) );
  OR2_X1 U10677 ( .A1(n12501), .A2(n12479), .ZN(n12484) );
  AND2_X1 U10678 ( .A1(n11065), .A2(n12484), .ZN(n11068) );
  NAND2_X1 U10679 ( .A1(n8231), .A2(n7366), .ZN(n11071) );
  NAND2_X1 U10680 ( .A1(n12648), .A2(n12472), .ZN(n11082) );
  INV_X1 U10681 ( .A(n12425), .ZN(n12454) );
  NAND2_X1 U10682 ( .A1(n12444), .A2(n12454), .ZN(n12420) );
  AND2_X1 U10683 ( .A1(n8232), .A2(n12420), .ZN(n11089) );
  NAND2_X1 U10684 ( .A1(n12436), .A2(n11089), .ZN(n8233) );
  NAND2_X1 U10685 ( .A1(n8233), .A2(n11091), .ZN(n11122) );
  INV_X1 U10686 ( .A(n11147), .ZN(n8234) );
  XNOR2_X1 U10687 ( .A(n11122), .B(n8234), .ZN(n12412) );
  NAND2_X1 U10688 ( .A1(n11160), .A2(n9452), .ZN(n8235) );
  NAND2_X1 U10689 ( .A1(n6480), .A2(n8235), .ZN(n8236) );
  NAND2_X1 U10690 ( .A1(n8236), .A2(n10965), .ZN(n8239) );
  NAND2_X1 U10691 ( .A1(n10965), .A2(n9452), .ZN(n8237) );
  NAND2_X1 U10692 ( .A1(n8237), .A2(n10853), .ZN(n8238) );
  NAND2_X1 U10693 ( .A1(n8239), .A2(n8238), .ZN(n8365) );
  INV_X1 U10694 ( .A(n6480), .ZN(n9247) );
  NAND2_X1 U10695 ( .A1(n9247), .A2(n9452), .ZN(n10854) );
  INV_X1 U10696 ( .A(n10854), .ZN(n11155) );
  NAND3_X1 U10697 ( .A1(n8365), .A2(n11155), .A3(n15131), .ZN(n8240) );
  OR3_X1 U10698 ( .A1(n6480), .A2(n9452), .A3(n10853), .ZN(n9690) );
  AND2_X1 U10699 ( .A1(n12412), .A2(n15160), .ZN(n8241) );
  MUX2_X1 U10700 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8242), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8244) );
  XNOR2_X1 U10701 ( .A(n10372), .B(P3_B_REG_SCAN_IN), .ZN(n8247) );
  NAND2_X1 U10702 ( .A1(n8243), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8245) );
  MUX2_X1 U10703 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8245), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8246) );
  NAND2_X1 U10704 ( .A1(n8246), .A2(n8248), .ZN(n10495) );
  INV_X1 U10705 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U10706 ( .A1(n10632), .A2(n10495), .ZN(n8250) );
  NAND2_X1 U10707 ( .A1(n8251), .A2(n8250), .ZN(n10858) );
  INV_X1 U10708 ( .A(n10858), .ZN(n10860) );
  NAND2_X1 U10709 ( .A1(n12760), .A2(n10860), .ZN(n10863) );
  NOR2_X1 U10710 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8255) );
  NOR4_X1 U10711 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8254) );
  NOR4_X1 U10712 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8253) );
  NOR4_X1 U10713 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8252) );
  NAND4_X1 U10714 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n8261)
         );
  NOR4_X1 U10715 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8259) );
  NOR4_X1 U10716 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8258) );
  NOR4_X1 U10717 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8257) );
  NOR4_X1 U10718 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8256) );
  NAND4_X1 U10719 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n8260)
         );
  NOR2_X1 U10720 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  NOR2_X1 U10721 ( .A1(n10863), .A2(n9694), .ZN(n8372) );
  NOR2_X1 U10722 ( .A1(n10854), .A2(n6476), .ZN(n9687) );
  NOR2_X1 U10723 ( .A1(n10495), .A2(n10372), .ZN(n8266) );
  NAND2_X1 U10724 ( .A1(n8267), .A2(n8266), .ZN(n8449) );
  NAND2_X1 U10725 ( .A1(n9687), .A2(n8355), .ZN(n8374) );
  NAND2_X1 U10726 ( .A1(n10965), .A2(n10852), .ZN(n11153) );
  NOR2_X1 U10727 ( .A1(n8268), .A2(n11153), .ZN(n8367) );
  NAND2_X1 U10728 ( .A1(n8367), .A2(n8355), .ZN(n8356) );
  NAND2_X1 U10729 ( .A1(n8374), .A2(n8356), .ZN(n8269) );
  NAND2_X1 U10730 ( .A1(n8372), .A2(n8269), .ZN(n8271) );
  NAND2_X1 U10731 ( .A1(n9691), .A2(n10858), .ZN(n9695) );
  NOR2_X1 U10732 ( .A1(n9695), .A2(n9694), .ZN(n8375) );
  NAND3_X1 U10733 ( .A1(n8375), .A2(n8355), .A3(n8365), .ZN(n8270) );
  INV_X1 U10734 ( .A(n12757), .ZN(n8273) );
  NAND2_X1 U10735 ( .A1(n12417), .A2(n8273), .ZN(n8274) );
  INV_X2 U10736 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U10737 ( .A(n11153), .ZN(n8275) );
  NAND2_X1 U10738 ( .A1(n12402), .A2(n10965), .ZN(n8276) );
  XNOR2_X1 U10739 ( .A(n12444), .B(n12051), .ZN(n12057) );
  NOR2_X1 U10740 ( .A1(n12057), .A2(n12425), .ZN(n12053) );
  AOI21_X1 U10741 ( .B1(n12057), .B2(n12425), .A(n12053), .ZN(n8354) );
  XNOR2_X1 U10742 ( .A(n14357), .B(n6474), .ZN(n12157) );
  INV_X1 U10743 ( .A(n12157), .ZN(n8312) );
  XNOR2_X1 U10744 ( .A(n15063), .B(n6474), .ZN(n8289) );
  INV_X1 U10745 ( .A(n8286), .ZN(n8287) );
  XNOR2_X1 U10746 ( .A(n9898), .B(n6474), .ZN(n8285) );
  INV_X1 U10747 ( .A(n15089), .ZN(n9404) );
  NAND2_X1 U10748 ( .A1(n8278), .A2(n7018), .ZN(n8281) );
  INV_X1 U10749 ( .A(n8281), .ZN(n8282) );
  NOR2_X1 U10750 ( .A1(n9401), .A2(n8282), .ZN(n9510) );
  XNOR2_X1 U10751 ( .A(n15097), .B(n8283), .ZN(n9511) );
  INV_X1 U10752 ( .A(n8283), .ZN(n8284) );
  XNOR2_X1 U10753 ( .A(n15071), .B(n8285), .ZN(n9895) );
  XNOR2_X1 U10754 ( .A(n10249), .B(n6474), .ZN(n8288) );
  XNOR2_X1 U10755 ( .A(n12230), .B(n8288), .ZN(n10245) );
  XNOR2_X1 U10756 ( .A(n8289), .B(n10401), .ZN(n10272) );
  NAND2_X1 U10757 ( .A1(n10273), .A2(n10272), .ZN(n10271) );
  XNOR2_X1 U10758 ( .A(n12069), .B(n6474), .ZN(n8290) );
  XNOR2_X1 U10759 ( .A(n12228), .B(n8290), .ZN(n12067) );
  INV_X1 U10760 ( .A(n8290), .ZN(n8291) );
  NAND2_X1 U10761 ( .A1(n12228), .A2(n8291), .ZN(n8292) );
  XNOR2_X1 U10762 ( .A(n12092), .B(n6474), .ZN(n8293) );
  XNOR2_X1 U10763 ( .A(n8293), .B(n15044), .ZN(n12089) );
  INV_X1 U10764 ( .A(n8293), .ZN(n8294) );
  NAND2_X1 U10765 ( .A1(n15044), .A2(n8294), .ZN(n8295) );
  XNOR2_X1 U10766 ( .A(n15048), .B(n6474), .ZN(n8296) );
  XNOR2_X1 U10767 ( .A(n8296), .B(n15024), .ZN(n10658) );
  INV_X1 U10768 ( .A(n8296), .ZN(n8298) );
  INV_X1 U10769 ( .A(n10780), .ZN(n8300) );
  XNOR2_X1 U10770 ( .A(n10785), .B(n6474), .ZN(n8301) );
  XNOR2_X1 U10771 ( .A(n12179), .B(n8301), .ZN(n10779) );
  NAND2_X1 U10772 ( .A1(n8300), .A2(n8299), .ZN(n10781) );
  INV_X1 U10773 ( .A(n8301), .ZN(n8303) );
  NAND2_X1 U10774 ( .A1(n10781), .A2(n8304), .ZN(n12105) );
  XNOR2_X1 U10775 ( .A(n10874), .B(n6474), .ZN(n12106) );
  INV_X1 U10776 ( .A(n12106), .ZN(n8305) );
  XNOR2_X1 U10777 ( .A(n14366), .B(n6474), .ZN(n12107) );
  NAND2_X1 U10778 ( .A1(n12107), .A2(n12227), .ZN(n8308) );
  OAI21_X1 U10779 ( .B1(n12173), .B2(n8305), .A(n8308), .ZN(n8310) );
  NOR2_X1 U10780 ( .A1(n15025), .A2(n12106), .ZN(n8307) );
  INV_X1 U10781 ( .A(n12107), .ZN(n8306) );
  AOI22_X1 U10782 ( .A1(n8308), .A2(n8307), .B1(n14356), .B2(n8306), .ZN(n8309) );
  NOR2_X1 U10783 ( .A1(n12157), .A2(n12226), .ZN(n8311) );
  XNOR2_X1 U10784 ( .A(n12756), .B(n12051), .ZN(n8313) );
  NAND2_X1 U10785 ( .A1(n8313), .A2(n14355), .ZN(n8314) );
  OAI21_X1 U10786 ( .B1(n8313), .B2(n14355), .A(n8314), .ZN(n11217) );
  XNOR2_X1 U10787 ( .A(n12752), .B(n12051), .ZN(n12120) );
  INV_X1 U10788 ( .A(n12120), .ZN(n12209) );
  XNOR2_X1 U10789 ( .A(n12127), .B(n12051), .ZN(n8318) );
  NAND2_X1 U10790 ( .A1(n8318), .A2(n12583), .ZN(n12121) );
  NOR2_X1 U10791 ( .A1(n8318), .A2(n12583), .ZN(n12123) );
  AOI21_X1 U10792 ( .B1(n8319), .B2(n12121), .A(n12123), .ZN(n12133) );
  XNOR2_X1 U10793 ( .A(n12689), .B(n6474), .ZN(n8320) );
  XNOR2_X1 U10794 ( .A(n8320), .B(n12598), .ZN(n12132) );
  XNOR2_X1 U10795 ( .A(n12681), .B(n6474), .ZN(n8321) );
  XNOR2_X1 U10796 ( .A(n8321), .B(n8322), .ZN(n12184) );
  OAI22_X1 U10797 ( .A1(n12185), .A2(n12184), .B1(n8322), .B2(n8321), .ZN(
        n12081) );
  XNOR2_X1 U10798 ( .A(n12677), .B(n6474), .ZN(n8323) );
  XNOR2_X1 U10799 ( .A(n8323), .B(n12571), .ZN(n12082) );
  NAND2_X1 U10800 ( .A1(n12081), .A2(n12082), .ZN(n8326) );
  NAND2_X1 U10801 ( .A1(n8326), .A2(n8325), .ZN(n12151) );
  XNOR2_X1 U10802 ( .A(n12536), .B(n6474), .ZN(n8327) );
  XNOR2_X1 U10803 ( .A(n8327), .B(n12548), .ZN(n12150) );
  INV_X1 U10804 ( .A(n8327), .ZN(n8328) );
  NAND2_X1 U10805 ( .A1(n8328), .A2(n12548), .ZN(n8329) );
  XNOR2_X1 U10806 ( .A(n12526), .B(n6474), .ZN(n8330) );
  NAND2_X1 U10807 ( .A1(n8330), .A2(n12535), .ZN(n8332) );
  OAI21_X1 U10808 ( .B1(n8330), .B2(n12535), .A(n8332), .ZN(n12099) );
  INV_X1 U10809 ( .A(n12099), .ZN(n8331) );
  XNOR2_X1 U10810 ( .A(n12665), .B(n6474), .ZN(n8333) );
  NAND2_X1 U10811 ( .A1(n8334), .A2(n8333), .ZN(n8335) );
  XNOR2_X1 U10812 ( .A(n12501), .B(n6474), .ZN(n8336) );
  XNOR2_X1 U10813 ( .A(n12725), .B(n12051), .ZN(n8338) );
  NAND2_X1 U10814 ( .A1(n8338), .A2(n7366), .ZN(n8391) );
  INV_X1 U10815 ( .A(n8338), .ZN(n8339) );
  NAND2_X1 U10816 ( .A1(n8339), .A2(n12469), .ZN(n8340) );
  AND2_X1 U10817 ( .A1(n8391), .A2(n8340), .ZN(n12140) );
  XNOR2_X1 U10818 ( .A(n12653), .B(n6474), .ZN(n8342) );
  NAND2_X1 U10819 ( .A1(n8342), .A2(n12480), .ZN(n8348) );
  INV_X1 U10820 ( .A(n8342), .ZN(n8343) );
  NAND2_X1 U10821 ( .A1(n8343), .A2(n12224), .ZN(n8344) );
  AND2_X1 U10822 ( .A1(n8348), .A2(n8344), .ZN(n8347) );
  XNOR2_X1 U10823 ( .A(n12648), .B(n12051), .ZN(n8345) );
  NOR2_X1 U10824 ( .A1(n8345), .A2(n12223), .ZN(n8350) );
  AOI21_X1 U10825 ( .B1(n8345), .B2(n12223), .A(n8350), .ZN(n12202) );
  AND2_X1 U10826 ( .A1(n8387), .A2(n12202), .ZN(n8346) );
  NAND2_X1 U10827 ( .A1(n8389), .A2(n8346), .ZN(n12199) );
  INV_X1 U10828 ( .A(n12202), .ZN(n8349) );
  INV_X1 U10829 ( .A(n8347), .ZN(n8390) );
  OR2_X1 U10830 ( .A1(n8390), .A2(n8391), .ZN(n8388) );
  AND2_X1 U10831 ( .A1(n8388), .A2(n8348), .ZN(n12196) );
  INV_X1 U10832 ( .A(n8350), .ZN(n8351) );
  AND2_X1 U10833 ( .A1(n12198), .A2(n8351), .ZN(n8352) );
  NAND2_X1 U10834 ( .A1(n12199), .A2(n8352), .ZN(n8353) );
  OAI21_X1 U10835 ( .B1(n8354), .B2(n8353), .A(n12064), .ZN(n8360) );
  NAND4_X1 U10836 ( .A1(n8372), .A2(n8355), .A3(n15131), .A4(n8365), .ZN(n8359) );
  INV_X1 U10837 ( .A(n8356), .ZN(n8357) );
  NAND2_X1 U10838 ( .A1(n8375), .A2(n8357), .ZN(n8358) );
  NAND2_X1 U10839 ( .A1(n8360), .A2(n12203), .ZN(n8383) );
  OR2_X1 U10840 ( .A1(n8372), .A2(n11121), .ZN(n8361) );
  NOR2_X1 U10841 ( .A1(n9693), .A2(n15131), .ZN(n9686) );
  NAND2_X1 U10842 ( .A1(n8361), .A2(n9686), .ZN(n12214) );
  INV_X1 U10843 ( .A(n8374), .ZN(n11158) );
  NAND2_X1 U10844 ( .A1(n8375), .A2(n11158), .ZN(n8364) );
  INV_X1 U10845 ( .A(n8364), .ZN(n8362) );
  INV_X1 U10846 ( .A(n8365), .ZN(n8371) );
  NAND2_X1 U10847 ( .A1(n8449), .A2(n9141), .ZN(n8366) );
  NOR2_X1 U10848 ( .A1(n10857), .A2(n8366), .ZN(n8370) );
  INV_X1 U10849 ( .A(n8367), .ZN(n8368) );
  OR2_X1 U10850 ( .A1(n8375), .A2(n8368), .ZN(n8369) );
  OAI211_X1 U10851 ( .C1(n8372), .C2(n8371), .A(n8370), .B(n8369), .ZN(n8373)
         );
  NAND2_X1 U10852 ( .A1(n8373), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8377) );
  OR2_X1 U10853 ( .A1(n8375), .A2(n8374), .ZN(n8376) );
  AOI22_X1 U10854 ( .A1(n12443), .A2(n12217), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8378) );
  OAI21_X1 U10855 ( .B1(n12472), .B2(n12213), .A(n8378), .ZN(n8379) );
  AOI21_X1 U10856 ( .B1(n12222), .B2(n12211), .A(n8379), .ZN(n8380) );
  INV_X1 U10857 ( .A(n8381), .ZN(n8382) );
  NAND2_X1 U10858 ( .A1(n8383), .A2(n8382), .ZN(P3_U3154) );
  INV_X1 U10859 ( .A(n12653), .ZN(n8397) );
  INV_X1 U10860 ( .A(n12211), .ZN(n12187) );
  AOI22_X1 U10861 ( .A1(n12469), .A2(n12189), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8385) );
  NAND2_X1 U10862 ( .A1(n12473), .A2(n12217), .ZN(n8384) );
  OAI211_X1 U10863 ( .C1(n12472), .C2(n12187), .A(n8385), .B(n8384), .ZN(n8386) );
  INV_X1 U10864 ( .A(n8386), .ZN(n8396) );
  NAND2_X1 U10865 ( .A1(n8389), .A2(n8387), .ZN(n12197) );
  AND2_X1 U10866 ( .A1(n12197), .A2(n8388), .ZN(n8393) );
  NAND2_X1 U10867 ( .A1(n8389), .A2(n12140), .ZN(n12142) );
  NAND3_X1 U10868 ( .A1(n12142), .A2(n8391), .A3(n8390), .ZN(n8392) );
  AOI21_X1 U10869 ( .B1(n8393), .B2(n8392), .A(n12219), .ZN(n8394) );
  INV_X1 U10870 ( .A(n8394), .ZN(n8395) );
  NOR2_X1 U10871 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .ZN(n8403) );
  NOR2_X1 U10872 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n8402) );
  INV_X1 U10873 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10874 ( .A1(n8611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10875 ( .A1(n6635), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U10876 ( .A(n8417), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U10877 ( .A1(n8887), .A2(n8886), .ZN(n8418) );
  INV_X1 U10878 ( .A(n8891), .ZN(n8422) );
  INV_X1 U10879 ( .A(n8712), .ZN(n8426) );
  NOR2_X1 U10880 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8425) );
  NOR2_X1 U10881 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8424) );
  INV_X2 U10882 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8715) );
  INV_X2 U10883 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8825) );
  NAND2_X1 U10884 ( .A1(n6569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10885 ( .A1(n6513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8446) );
  MUX2_X1 U10886 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8446), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n8448) );
  NAND2_X1 U10887 ( .A1(n8448), .A2(n8447), .ZN(n9120) );
  NAND2_X1 U10888 ( .A1(n9120), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10949) );
  INV_X1 U10889 ( .A(n8449), .ZN(n8450) );
  NAND2_X2 U10890 ( .A1(n11332), .A2(P1_U3086), .ZN(n14223) );
  NOR2_X1 U10891 ( .A1(n11332), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14215) );
  INV_X2 U10892 ( .A(n14215), .ZN(n14221) );
  INV_X1 U10893 ( .A(n8912), .ZN(n8451) );
  NAND2_X1 U10894 ( .A1(n8451), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8914) );
  AND2_X1 U10895 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8452) );
  NAND2_X1 U10896 ( .A1(n8945), .A2(n8452), .ZN(n9064) );
  NAND2_X1 U10897 ( .A1(n8914), .A2(n9064), .ZN(n8482) );
  XNOR2_X1 U10898 ( .A(n8483), .B(n8482), .ZN(n9079) );
  NAND2_X1 U10899 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8453) );
  MUX2_X1 U10900 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8453), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8455) );
  INV_X1 U10901 ( .A(n8454), .ZN(n8487) );
  NAND2_X1 U10902 ( .A1(n8455), .A2(n8487), .ZN(n13736) );
  OAI222_X1 U10903 ( .A1(n14223), .A2(n7611), .B1(n14221), .B2(n9079), .C1(
        P1_U3086), .C2(n13736), .ZN(P1_U3354) );
  NOR2_X1 U10904 ( .A1(n11332), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13361) );
  INV_X2 U10905 ( .A(n13361), .ZN(n13368) );
  INV_X2 U10906 ( .A(n10257), .ZN(n13366) );
  NAND2_X1 U10907 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8457) );
  INV_X1 U10908 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8456) );
  MUX2_X1 U10909 ( .A(n8457), .B(P2_IR_REG_31__SCAN_IN), .S(n8456), .Z(n8458)
         );
  OAI222_X1 U10910 ( .A1(n13368), .A2(n8966), .B1(n13366), .B2(n9079), .C1(
        P2_U3088), .C2(n8967), .ZN(P2_U3326) );
  NAND2_X2 U10911 ( .A1(n8494), .A2(P3_U3151), .ZN(n12771) );
  INV_X1 U10912 ( .A(n12764), .ZN(n12770) );
  OAI222_X1 U10913 ( .A1(P3_U3151), .A2(n9365), .B1(n12771), .B2(n8460), .C1(
        n12770), .C2(n8459), .ZN(P3_U3294) );
  OAI222_X1 U10914 ( .A1(n12770), .A2(n8462), .B1(n12771), .B2(n8461), .C1(
        n10234), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U10915 ( .A(n8463), .ZN(n8464) );
  INV_X1 U10916 ( .A(SI_2_), .ZN(n15258) );
  OAI222_X1 U10917 ( .A1(n12770), .A2(n8464), .B1(n12771), .B2(n15258), .C1(
        n9319), .C2(P3_U3151), .ZN(P3_U3293) );
  OAI222_X1 U10918 ( .A1(n9880), .A2(P3_U3151), .B1(n12770), .B2(n8466), .C1(
        n8465), .C2(n12771), .ZN(P3_U3289) );
  INV_X1 U10919 ( .A(n12771), .ZN(n8473) );
  AOI222_X1 U10920 ( .A1(n8467), .A2(n12764), .B1(SI_7_), .B2(n8473), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n14956), .ZN(n8468) );
  INV_X1 U10921 ( .A(n8468), .ZN(P3_U3288) );
  AOI222_X1 U10922 ( .A1(n8469), .A2(n12764), .B1(SI_4_), .B2(n8473), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n9172), .ZN(n8470) );
  INV_X1 U10923 ( .A(n8470), .ZN(P3_U3291) );
  AOI222_X1 U10924 ( .A1(n8471), .A2(n12764), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14924), .C1(SI_3_), .C2(n8473), .ZN(n8472) );
  INV_X1 U10925 ( .A(n8472), .ZN(P3_U3292) );
  AOI222_X1 U10926 ( .A1(n8474), .A2(n12764), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14940), .C1(SI_5_), .C2(n8473), .ZN(n8475) );
  INV_X1 U10927 ( .A(n8475), .ZN(P3_U3290) );
  INV_X1 U10928 ( .A(n8476), .ZN(n8477) );
  INV_X1 U10929 ( .A(SI_9_), .ZN(n15335) );
  OAI222_X1 U10930 ( .A1(n12770), .A2(n8477), .B1(n12771), .B2(n15335), .C1(
        n7055), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U10931 ( .A(n8478), .ZN(n8480) );
  INV_X1 U10932 ( .A(SI_10_), .ZN(n8479) );
  INV_X1 U10933 ( .A(n14982), .ZN(n10579) );
  OAI222_X1 U10934 ( .A1(n12770), .A2(n8480), .B1(n12771), .B2(n8479), .C1(
        n10579), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U10935 ( .A1(n12770), .A2(n8481), .B1(n12771), .B2(n8688), .C1(
        n10578), .C2(P3_U3151), .ZN(P3_U3284) );
  NAND2_X1 U10936 ( .A1(n8484), .A2(SI_1_), .ZN(n8485) );
  XNOR2_X1 U10937 ( .A(n8504), .B(SI_2_), .ZN(n8490) );
  MUX2_X1 U10938 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8494), .Z(n8505) );
  XNOR2_X1 U10939 ( .A(n8505), .B(n8490), .ZN(n9281) );
  INV_X1 U10940 ( .A(n9281), .ZN(n8548) );
  NAND2_X1 U10941 ( .A1(n8487), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8488) );
  MUX2_X1 U10942 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8488), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n8489) );
  NAND2_X1 U10943 ( .A1(n8489), .A2(n8520), .ZN(n9285) );
  OAI222_X1 U10944 ( .A1(n14223), .A2(n9282), .B1(n14221), .B2(n8548), .C1(
        P1_U3086), .C2(n9285), .ZN(P1_U3353) );
  INV_X1 U10945 ( .A(n8490), .ZN(n8491) );
  NAND2_X1 U10946 ( .A1(n8491), .A2(n8505), .ZN(n8493) );
  NAND2_X1 U10947 ( .A1(n8504), .A2(SI_2_), .ZN(n8492) );
  NAND2_X1 U10948 ( .A1(n8493), .A2(n8492), .ZN(n8496) );
  XNOR2_X1 U10949 ( .A(n8507), .B(SI_3_), .ZN(n8495) );
  INV_X1 U10950 ( .A(n9574), .ZN(n8558) );
  NAND2_X1 U10951 ( .A1(n8520), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8497) );
  XNOR2_X1 U10952 ( .A(n8497), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13747) );
  INV_X1 U10953 ( .A(n13747), .ZN(n8498) );
  OAI222_X1 U10954 ( .A1(n14223), .A2(n8499), .B1(n14221), .B2(n8558), .C1(
        P1_U3086), .C2(n8498), .ZN(P1_U3352) );
  INV_X1 U10955 ( .A(SI_3_), .ZN(n8500) );
  NAND2_X1 U10956 ( .A1(n8501), .A2(n8500), .ZN(n8508) );
  OAI21_X1 U10957 ( .B1(SI_2_), .B2(n8505), .A(n8508), .ZN(n8502) );
  INV_X1 U10958 ( .A(n8502), .ZN(n8503) );
  NAND2_X1 U10959 ( .A1(n8504), .A2(n8503), .ZN(n8511) );
  INV_X1 U10960 ( .A(n8505), .ZN(n8506) );
  NOR2_X1 U10961 ( .A1(n8506), .A2(n15258), .ZN(n8509) );
  AOI22_X1 U10962 ( .A1(n8509), .A2(n8508), .B1(n8507), .B2(SI_3_), .ZN(n8510)
         );
  MUX2_X1 U10963 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8494), .Z(n8513) );
  XNOR2_X1 U10964 ( .A(n8513), .B(SI_4_), .ZN(n8529) );
  INV_X1 U10965 ( .A(n8529), .ZN(n8512) );
  NAND2_X1 U10966 ( .A1(n8530), .A2(n8512), .ZN(n8515) );
  NAND2_X1 U10967 ( .A1(n8513), .A2(SI_4_), .ZN(n8514) );
  NAND2_X1 U10968 ( .A1(n8525), .A2(n8516), .ZN(n8519) );
  NAND2_X1 U10969 ( .A1(n8517), .A2(SI_5_), .ZN(n8518) );
  XNOR2_X1 U10970 ( .A(n8537), .B(n8535), .ZN(n9822) );
  INV_X1 U10971 ( .A(n9822), .ZN(n8561) );
  OR2_X1 U10972 ( .A1(n8520), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8531) );
  INV_X1 U10973 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8521) );
  INV_X1 U10974 ( .A(n8540), .ZN(n8527) );
  NAND2_X1 U10975 ( .A1(n8527), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8522) );
  XNOR2_X1 U10976 ( .A(n8522), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9823) );
  INV_X1 U10977 ( .A(n9823), .ZN(n8868) );
  OAI222_X1 U10978 ( .A1(n14223), .A2(n8523), .B1(n14221), .B2(n8561), .C1(
        P1_U3086), .C2(n8868), .ZN(P1_U3349) );
  XNOR2_X1 U10979 ( .A(n8525), .B(n8524), .ZN(n9769) );
  INV_X1 U10980 ( .A(n9769), .ZN(n8573) );
  INV_X1 U10981 ( .A(n9216), .ZN(n8533) );
  NAND2_X1 U10982 ( .A1(n8533), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8526) );
  MUX2_X1 U10983 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8526), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n8528) );
  NAND2_X1 U10984 ( .A1(n8528), .A2(n8527), .ZN(n13769) );
  OAI222_X1 U10985 ( .A1(n14223), .A2(n9770), .B1(n14221), .B2(n8573), .C1(
        P1_U3086), .C2(n13769), .ZN(P1_U3350) );
  XNOR2_X1 U10986 ( .A(n8530), .B(n8529), .ZN(n9594) );
  INV_X1 U10987 ( .A(n9594), .ZN(n8553) );
  NAND2_X1 U10988 ( .A1(n8531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8532) );
  MUX2_X1 U10989 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8532), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n8534) );
  NAND2_X1 U10990 ( .A1(n8534), .A2(n8533), .ZN(n9598) );
  OAI222_X1 U10991 ( .A1(n14223), .A2(n9595), .B1(n14221), .B2(n8553), .C1(
        P1_U3086), .C2(n9598), .ZN(P1_U3351) );
  INV_X1 U10992 ( .A(n8535), .ZN(n8536) );
  XNOR2_X1 U10993 ( .A(n8582), .B(SI_7_), .ZN(n8579) );
  XNOR2_X1 U10994 ( .A(n8581), .B(n8579), .ZN(n9970) );
  INV_X1 U10995 ( .A(n9970), .ZN(n8566) );
  INV_X1 U10996 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10997 ( .A1(n8540), .A2(n8539), .ZN(n8542) );
  NAND2_X1 U10998 ( .A1(n8542), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8541) );
  MUX2_X1 U10999 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8541), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n8543) );
  AND2_X1 U11000 ( .A1(n8543), .A2(n8591), .ZN(n9971) );
  INV_X1 U11001 ( .A(n9971), .ZN(n8837) );
  OAI222_X1 U11002 ( .A1(n14223), .A2(n7002), .B1(n14221), .B2(n8566), .C1(
        P1_U3086), .C2(n8837), .ZN(P1_U3348) );
  NAND2_X1 U11003 ( .A1(n8546), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8545) );
  INV_X1 U11004 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8544) );
  MUX2_X1 U11005 ( .A(n8545), .B(P2_IR_REG_31__SCAN_IN), .S(n8544), .Z(n8547)
         );
  NOR2_X1 U11006 ( .A1(n8546), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U11007 ( .A1(n8547), .A2(n8554), .ZN(n8660) );
  OAI222_X1 U11008 ( .A1(n13368), .A2(n8976), .B1(n13366), .B2(n8548), .C1(
        P2_U3088), .C2(n8660), .ZN(P2_U3325) );
  INV_X1 U11009 ( .A(n8556), .ZN(n8549) );
  NAND2_X1 U11010 ( .A1(n8549), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8550) );
  MUX2_X1 U11011 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8550), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8552) );
  NAND2_X1 U11012 ( .A1(n8556), .A2(n8551), .ZN(n8568) );
  AND2_X1 U11013 ( .A1(n8552), .A2(n8568), .ZN(n9323) );
  INV_X1 U11014 ( .A(n9323), .ZN(n8746) );
  OAI222_X1 U11015 ( .A1(n13368), .A2(n9326), .B1(n13366), .B2(n8553), .C1(
        P2_U3088), .C2(n8746), .ZN(P2_U3323) );
  NOR2_X1 U11016 ( .A1(n8557), .A2(n8556), .ZN(n12905) );
  INV_X1 U11017 ( .A(n12905), .ZN(n8662) );
  OAI222_X1 U11018 ( .A1(n13368), .A2(n8559), .B1(n13366), .B2(n8558), .C1(
        P2_U3088), .C2(n8662), .ZN(P2_U3324) );
  NAND2_X1 U11019 ( .A1(n8571), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8560) );
  XNOR2_X1 U11020 ( .A(n8560), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9528) );
  INV_X1 U11021 ( .A(n9528), .ZN(n8733) );
  OAI222_X1 U11022 ( .A1(n13368), .A2(n8562), .B1(n13366), .B2(n8561), .C1(
        P2_U3088), .C2(n8733), .ZN(P2_U3321) );
  INV_X1 U11023 ( .A(n8571), .ZN(n8564) );
  INV_X1 U11024 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U11025 ( .A1(n8564), .A2(n8563), .ZN(n8583) );
  NAND2_X1 U11026 ( .A1(n8583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8565) );
  XNOR2_X1 U11027 ( .A(n8565), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9635) );
  INV_X1 U11028 ( .A(n9635), .ZN(n8710) );
  OAI222_X1 U11029 ( .A1(n13368), .A2(n8567), .B1(n13366), .B2(n8566), .C1(
        P2_U3088), .C2(n8710), .ZN(P2_U3320) );
  NAND2_X1 U11030 ( .A1(n8568), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8570) );
  MUX2_X1 U11031 ( .A(n8570), .B(P2_IR_REG_31__SCAN_IN), .S(n8569), .Z(n8572)
         );
  AND2_X1 U11032 ( .A1(n8572), .A2(n8571), .ZN(n9556) );
  INV_X1 U11033 ( .A(n9556), .ZN(n8669) );
  OAI222_X1 U11034 ( .A1(n13368), .A2(n8574), .B1(n13366), .B2(n8573), .C1(
        P2_U3088), .C2(n8669), .ZN(P2_U3322) );
  INV_X1 U11035 ( .A(n8575), .ZN(n8576) );
  OAI222_X1 U11036 ( .A1(n12770), .A2(n8576), .B1(n12771), .B2(n15232), .C1(
        n14992), .C2(P3_U3151), .ZN(P3_U3283) );
  NAND2_X1 U11037 ( .A1(n10860), .A2(n12759), .ZN(n8577) );
  OAI21_X1 U11038 ( .B1(n12759), .B2(n8578), .A(n8577), .ZN(P3_U3377) );
  INV_X1 U11039 ( .A(n8579), .ZN(n8580) );
  MUX2_X1 U11040 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11332), .Z(n8597) );
  XNOR2_X1 U11041 ( .A(n8597), .B(SI_8_), .ZN(n8594) );
  XNOR2_X1 U11042 ( .A(n8596), .B(n8594), .ZN(n9976) );
  INV_X1 U11043 ( .A(n9976), .ZN(n8592) );
  INV_X1 U11044 ( .A(n8583), .ZN(n8585) );
  INV_X1 U11045 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U11046 ( .A1(n8585), .A2(n8584), .ZN(n8587) );
  AND2_X1 U11047 ( .A1(n8587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8586) );
  MUX2_X1 U11048 ( .A(n7012), .B(n8586), .S(P2_IR_REG_8__SCAN_IN), .Z(n8588)
         );
  NOR2_X1 U11049 ( .A1(n8588), .A2(n8675), .ZN(n9643) );
  INV_X1 U11050 ( .A(n9643), .ZN(n8589) );
  OAI222_X1 U11051 ( .A1(n13368), .A2(n8590), .B1(n13366), .B2(n8592), .C1(
        P2_U3088), .C2(n8589), .ZN(P2_U3319) );
  NAND2_X1 U11052 ( .A1(n8591), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8600) );
  XNOR2_X1 U11053 ( .A(n8600), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9977) );
  INV_X1 U11054 ( .A(n9977), .ZN(n8829) );
  OAI222_X1 U11055 ( .A1(n14223), .A2(n8593), .B1(n14221), .B2(n8592), .C1(
        P1_U3086), .C2(n8829), .ZN(P1_U3347) );
  INV_X1 U11056 ( .A(n8594), .ZN(n8595) );
  NAND2_X1 U11057 ( .A1(n8597), .A2(SI_8_), .ZN(n8598) );
  MUX2_X1 U11058 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n11332), .Z(n8673) );
  XNOR2_X1 U11059 ( .A(n8673), .B(SI_9_), .ZN(n8670) );
  XNOR2_X1 U11060 ( .A(n8672), .B(n8670), .ZN(n10329) );
  INV_X1 U11061 ( .A(n10329), .ZN(n8609) );
  NAND2_X1 U11062 ( .A1(n8600), .A2(n8599), .ZN(n8601) );
  NAND2_X1 U11063 ( .A1(n8601), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11064 ( .A1(n8714), .A2(n8602), .ZN(n8678) );
  OR2_X1 U11065 ( .A1(n8714), .A2(n8602), .ZN(n8603) );
  INV_X1 U11066 ( .A(n10330), .ZN(n8604) );
  OAI222_X1 U11067 ( .A1(n14223), .A2(n8605), .B1(n14221), .B2(n8609), .C1(
        P1_U3086), .C2(n8604), .ZN(P1_U3346) );
  INV_X1 U11068 ( .A(n8675), .ZN(n8606) );
  NAND2_X1 U11069 ( .A1(n8606), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U11070 ( .A(n8607), .B(P2_IR_REG_9__SCAN_IN), .ZN(n12926) );
  INV_X1 U11071 ( .A(n12926), .ZN(n8608) );
  OAI222_X1 U11072 ( .A1(n13368), .A2(n8610), .B1(n13366), .B2(n8609), .C1(
        P2_U3088), .C2(n8608), .ZN(P2_U3318) );
  INV_X1 U11073 ( .A(n10258), .ZN(n8621) );
  XNOR2_X2 U11074 ( .A(n8615), .B(n8614), .ZN(n8622) );
  NAND2_X1 U11075 ( .A1(n8617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11076 ( .A1(n8960), .A2(n10258), .ZN(n8619) );
  NAND2_X1 U11077 ( .A1(n8968), .A2(n8619), .ZN(n8620) );
  OAI21_X1 U11078 ( .B1(n8920), .B2(n8621), .A(n8620), .ZN(n8624) );
  AND2_X1 U11079 ( .A1(n8624), .A2(n8622), .ZN(n14751) );
  AND2_X1 U11080 ( .A1(n14751), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14790) );
  OR2_X1 U11081 ( .A1(n8624), .A2(P2_U3088), .ZN(n9257) );
  INV_X1 U11082 ( .A(n9257), .ZN(n14784) );
  INV_X1 U11083 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U11084 ( .A1(n10041), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8628) );
  INV_X1 U11085 ( .A(n8967), .ZN(n8649) );
  INV_X1 U11086 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n14889) );
  MUX2_X1 U11087 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n14889), .S(n8967), .Z(n8645) );
  INV_X1 U11088 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8623) );
  NOR3_X1 U11089 ( .A1(n8645), .A2(n8623), .A3(n7612), .ZN(n8644) );
  AOI21_X1 U11090 ( .B1(n8649), .B2(P2_REG1_REG_1__SCAN_IN), .A(n8644), .ZN(
        n8626) );
  INV_X1 U11091 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n14891) );
  MUX2_X1 U11092 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n14891), .S(n8660), .Z(n8625) );
  NOR2_X1 U11093 ( .A1(n8626), .A2(n8625), .ZN(n12912) );
  NOR2_X1 U11094 ( .A1(n8622), .A2(P2_U3088), .ZN(n13360) );
  NAND2_X1 U11095 ( .A1(n8624), .A2(n13360), .ZN(n8632) );
  INV_X1 U11096 ( .A(n13365), .ZN(n12039) );
  AOI211_X1 U11097 ( .C1(n8626), .C2(n8625), .A(n12912), .B(n14742), .ZN(n8627) );
  AOI211_X1 U11098 ( .C1(n14784), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n8628), .B(
        n8627), .ZN(n8638) );
  INV_X1 U11099 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8629) );
  MUX2_X1 U11100 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n8629), .S(n8967), .Z(n8642)
         );
  INV_X1 U11101 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8905) );
  NOR3_X1 U11102 ( .A1(n8642), .A2(n8905), .A3(n7612), .ZN(n8652) );
  INV_X1 U11103 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10042) );
  MUX2_X1 U11104 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10042), .S(n8660), .Z(n8631) );
  NOR2_X1 U11105 ( .A1(n8967), .A2(n8629), .ZN(n8635) );
  INV_X1 U11106 ( .A(n8635), .ZN(n8630) );
  NAND2_X1 U11107 ( .A1(n8631), .A2(n8630), .ZN(n8636) );
  INV_X1 U11108 ( .A(n8632), .ZN(n8633) );
  AND2_X1 U11109 ( .A1(n8633), .A2(n12039), .ZN(n14791) );
  MUX2_X1 U11110 ( .A(n10042), .B(P2_REG2_REG_2__SCAN_IN), .S(n8660), .Z(n8634) );
  OAI21_X1 U11111 ( .B1(n8652), .B2(n8635), .A(n8634), .ZN(n12901) );
  OAI211_X1 U11112 ( .C1(n8652), .C2(n8636), .A(n14791), .B(n12901), .ZN(n8637) );
  OAI211_X1 U11113 ( .C1(n9395), .C2(n8660), .A(n8638), .B(n8637), .ZN(
        P2_U3216) );
  AND2_X1 U11114 ( .A1(n8640), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11115 ( .A1(n8640), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11116 ( .A1(n8640), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11117 ( .A1(n8640), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11118 ( .A1(n8640), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11119 ( .A1(n8640), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11120 ( .A1(n8640), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11121 ( .A1(n8640), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11122 ( .A1(n8640), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11123 ( .A1(n8640), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U11124 ( .A1(n8640), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11125 ( .A1(n8640), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11126 ( .A1(n8640), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11127 ( .A1(n8640), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11128 ( .A1(n8640), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11129 ( .A1(n8640), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11130 ( .A1(n8640), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11131 ( .A1(n8640), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11132 ( .A1(n8640), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11133 ( .A1(n8640), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11134 ( .A1(n8640), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11135 ( .A1(n8640), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11136 ( .A1(n8640), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11137 ( .A1(n8640), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11138 ( .A1(n8640), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U11139 ( .A1(n8640), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11140 ( .A1(n8640), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11141 ( .A1(n8640), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11142 ( .A1(n8640), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11143 ( .A1(n8640), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  OAI222_X1 U11144 ( .A1(n12770), .A2(n8641), .B1(n12771), .B2(n8999), .C1(
        n12280), .C2(P3_U3151), .ZN(P3_U3282) );
  NAND2_X1 U11145 ( .A1(n14791), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n14731) );
  OAI22_X1 U11146 ( .A1(n7612), .A2(n14731), .B1(n14733), .B2(n8642), .ZN(
        n8643) );
  INV_X1 U11147 ( .A(n8643), .ZN(n8651) );
  INV_X1 U11148 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8924) );
  OAI22_X1 U11149 ( .A1(n9257), .A2(n6738), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8924), .ZN(n8648) );
  OR2_X1 U11150 ( .A1(n7612), .A2(n8623), .ZN(n8646) );
  AOI211_X1 U11151 ( .C1(n8646), .C2(n8645), .A(n8644), .B(n14742), .ZN(n8647)
         );
  AOI211_X1 U11152 ( .C1(n14790), .C2(n8649), .A(n8648), .B(n8647), .ZN(n8650)
         );
  OAI21_X1 U11153 ( .B1(n8652), .B2(n8651), .A(n8650), .ZN(P2_U3215) );
  INV_X1 U11154 ( .A(n8660), .ZN(n8974) );
  NAND2_X1 U11155 ( .A1(n8974), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n12900) );
  INV_X1 U11156 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8653) );
  MUX2_X1 U11157 ( .A(n8653), .B(P2_REG2_REG_3__SCAN_IN), .S(n12905), .Z(
        n12899) );
  AOI21_X1 U11158 ( .B1(n12905), .B2(P2_REG2_REG_3__SCAN_IN), .A(n12903), .ZN(
        n8736) );
  INV_X1 U11159 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8654) );
  MUX2_X1 U11160 ( .A(n8654), .B(P2_REG2_REG_4__SCAN_IN), .S(n9323), .Z(n8735)
         );
  MUX2_X1 U11161 ( .A(n9819), .B(P2_REG2_REG_5__SCAN_IN), .S(n9556), .Z(n8656)
         );
  NOR2_X1 U11162 ( .A1(n8746), .A2(n8654), .ZN(n8658) );
  INV_X1 U11163 ( .A(n8658), .ZN(n8655) );
  NAND2_X1 U11164 ( .A1(n8656), .A2(n8655), .ZN(n8659) );
  INV_X1 U11165 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9819) );
  MUX2_X1 U11166 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9819), .S(n9556), .Z(n8657)
         );
  OAI21_X1 U11167 ( .B1(n8734), .B2(n8658), .A(n8657), .ZN(n8728) );
  OAI211_X1 U11168 ( .C1(n8734), .C2(n8659), .A(n8728), .B(n14791), .ZN(n8668)
         );
  NAND2_X1 U11169 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n12819) );
  INV_X1 U11170 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14893) );
  INV_X1 U11171 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n12906) );
  NOR2_X1 U11172 ( .A1(n8660), .A2(n14891), .ZN(n12907) );
  MUX2_X1 U11173 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n12906), .S(n12905), .Z(
        n8661) );
  OAI21_X1 U11174 ( .B1(n12912), .B2(n12907), .A(n8661), .ZN(n12910) );
  OAI21_X1 U11175 ( .B1(n12906), .B2(n8662), .A(n12910), .ZN(n8740) );
  MUX2_X1 U11176 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n14893), .S(n9323), .Z(n8739) );
  NAND2_X1 U11177 ( .A1(n8740), .A2(n8739), .ZN(n8738) );
  OAI21_X1 U11178 ( .B1(n14893), .B2(n8746), .A(n8738), .ZN(n8664) );
  INV_X1 U11179 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9333) );
  MUX2_X1 U11180 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9333), .S(n9556), .Z(n8663)
         );
  NAND2_X1 U11181 ( .A1(n8664), .A2(n8663), .ZN(n8720) );
  OAI211_X1 U11182 ( .C1(n8664), .C2(n8663), .A(n14785), .B(n8720), .ZN(n8665)
         );
  NAND2_X1 U11183 ( .A1(n12819), .A2(n8665), .ZN(n8666) );
  AOI21_X1 U11184 ( .B1(n14784), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8666), .ZN(
        n8667) );
  OAI211_X1 U11185 ( .C1(n9395), .C2(n8669), .A(n8668), .B(n8667), .ZN(
        P2_U3219) );
  INV_X1 U11186 ( .A(n8670), .ZN(n8671) );
  MUX2_X1 U11187 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n11332), .Z(n8685) );
  XNOR2_X1 U11188 ( .A(n8685), .B(SI_10_), .ZN(n8682) );
  XNOR2_X1 U11189 ( .A(n8684), .B(n8682), .ZN(n10335) );
  INV_X1 U11190 ( .A(n10335), .ZN(n8680) );
  INV_X1 U11191 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U11192 ( .A1(n8675), .A2(n8674), .ZN(n8695) );
  NAND2_X1 U11193 ( .A1(n8695), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8676) );
  XNOR2_X1 U11194 ( .A(n8676), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10172) );
  INV_X1 U11195 ( .A(n10172), .ZN(n9037) );
  OAI222_X1 U11196 ( .A1(n13368), .A2(n8677), .B1(n13366), .B2(n8680), .C1(
        P2_U3088), .C2(n9037), .ZN(P2_U3317) );
  NAND2_X1 U11197 ( .A1(n8678), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8679) );
  XNOR2_X1 U11198 ( .A(n8679), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10336) );
  INV_X1 U11199 ( .A(n10336), .ZN(n9442) );
  OAI222_X1 U11200 ( .A1(n14223), .A2(n8681), .B1(n14221), .B2(n8680), .C1(
        P1_U3086), .C2(n9442), .ZN(P1_U3345) );
  INV_X1 U11201 ( .A(n8682), .ZN(n8683) );
  NAND2_X1 U11202 ( .A1(n8685), .A2(SI_10_), .ZN(n8686) );
  MUX2_X1 U11203 ( .A(n8717), .B(n8697), .S(n11332), .Z(n8689) );
  NAND2_X1 U11204 ( .A1(n8689), .A2(n8688), .ZN(n8775) );
  INV_X1 U11205 ( .A(n8689), .ZN(n8690) );
  NAND2_X1 U11206 ( .A1(n8690), .A2(SI_11_), .ZN(n8691) );
  NAND2_X1 U11207 ( .A1(n8775), .A2(n8691), .ZN(n8692) );
  NAND2_X1 U11208 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  NAND2_X1 U11209 ( .A1(n8776), .A2(n8694), .ZN(n10547) );
  INV_X1 U11210 ( .A(n10547), .ZN(n8716) );
  OAI21_X1 U11211 ( .B1(n8695), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8696) );
  XNOR2_X1 U11212 ( .A(n8696), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10178) );
  INV_X1 U11213 ( .A(n10178), .ZN(n9381) );
  OAI222_X1 U11214 ( .A1(n13368), .A2(n8697), .B1(n13366), .B2(n8716), .C1(
        P2_U3088), .C2(n9381), .ZN(P2_U3316) );
  NAND2_X1 U11215 ( .A1(n9556), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8727) );
  INV_X1 U11216 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8698) );
  MUX2_X1 U11217 ( .A(n8698), .B(P2_REG2_REG_6__SCAN_IN), .S(n9528), .Z(n8726)
         );
  NOR2_X1 U11218 ( .A1(n8733), .A2(n8698), .ZN(n8701) );
  INV_X1 U11219 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9945) );
  MUX2_X1 U11220 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9945), .S(n9635), .Z(n8700)
         );
  NOR3_X1 U11221 ( .A1(n8725), .A2(n8701), .A3(n8700), .ZN(n8699) );
  NOR2_X1 U11222 ( .A1(n8699), .A2(n14733), .ZN(n8706) );
  NAND2_X1 U11223 ( .A1(n9556), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8719) );
  INV_X1 U11224 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14896) );
  MUX2_X1 U11225 ( .A(n14896), .B(P2_REG1_REG_6__SCAN_IN), .S(n9528), .Z(n8718) );
  AOI21_X1 U11226 ( .B1(n8720), .B2(n8719), .A(n8718), .ZN(n8722) );
  NOR2_X1 U11227 ( .A1(n8733), .A2(n14896), .ZN(n8704) );
  INV_X1 U11228 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9531) );
  MUX2_X1 U11229 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9531), .S(n9635), .Z(n8703)
         );
  NOR3_X1 U11230 ( .A1(n8722), .A2(n8704), .A3(n8703), .ZN(n8702) );
  NOR2_X1 U11231 ( .A1(n8702), .A2(n14742), .ZN(n8705) );
  OAI21_X1 U11232 ( .B1(n8722), .B2(n8704), .A(n8703), .ZN(n8769) );
  AOI22_X1 U11233 ( .A1(n8706), .A2(n8765), .B1(n8705), .B2(n8769), .ZN(n8709)
         );
  NAND2_X1 U11234 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9704) );
  INV_X1 U11235 ( .A(n9704), .ZN(n8707) );
  AOI21_X1 U11236 ( .B1(n14784), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8707), .ZN(
        n8708) );
  OAI211_X1 U11237 ( .C1(n8710), .C2(n9395), .A(n8709), .B(n8708), .ZN(
        P2_U3221) );
  OAI222_X1 U11238 ( .A1(n12770), .A2(n8711), .B1(n12771), .B2(n15322), .C1(
        n12289), .C2(P3_U3151), .ZN(P3_U3281) );
  NAND2_X1 U11239 ( .A1(n8712), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U11240 ( .A1(n8714), .A2(n8713), .ZN(n8787) );
  XNOR2_X1 U11241 ( .A(n8787), .B(n8715), .ZN(n13783) );
  INV_X1 U11242 ( .A(n13783), .ZN(n9443) );
  OAI222_X1 U11243 ( .A1(n8717), .A2(n14223), .B1(P1_U3086), .B2(n9443), .C1(
        n14221), .C2(n8716), .ZN(P1_U3344) );
  NAND2_X1 U11244 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9546) );
  INV_X1 U11245 ( .A(n9546), .ZN(n8724) );
  AND3_X1 U11246 ( .A1(n8720), .A2(n8719), .A3(n8718), .ZN(n8721) );
  NOR3_X1 U11247 ( .A1(n8722), .A2(n8721), .A3(n14742), .ZN(n8723) );
  AOI211_X1 U11248 ( .C1(n14784), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n8724), .B(
        n8723), .ZN(n8732) );
  INV_X1 U11249 ( .A(n8725), .ZN(n8730) );
  NAND3_X1 U11250 ( .A1(n8728), .A2(n8727), .A3(n8726), .ZN(n8729) );
  NAND3_X1 U11251 ( .A1(n8730), .A2(n14791), .A3(n8729), .ZN(n8731) );
  OAI211_X1 U11252 ( .C1(n9395), .C2(n8733), .A(n8732), .B(n8731), .ZN(
        P2_U3220) );
  AOI211_X1 U11253 ( .C1(n8736), .C2(n8735), .A(n8734), .B(n14733), .ZN(n8737)
         );
  INV_X1 U11254 ( .A(n8737), .ZN(n8742) );
  OAI211_X1 U11255 ( .C1(n8740), .C2(n8739), .A(n14785), .B(n8738), .ZN(n8741)
         );
  NAND2_X1 U11256 ( .A1(n8742), .A2(n8741), .ZN(n8744) );
  NAND2_X1 U11257 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n9346) );
  INV_X1 U11258 ( .A(n9346), .ZN(n8743) );
  AOI211_X1 U11259 ( .C1(n14784), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n8744), .B(
        n8743), .ZN(n8745) );
  OAI21_X1 U11260 ( .B1(n9395), .B2(n8746), .A(n8745), .ZN(P2_U3218) );
  INV_X1 U11261 ( .A(n10949), .ZN(n8747) );
  INV_X1 U11262 ( .A(n10947), .ZN(n8749) );
  INV_X1 U11263 ( .A(n9120), .ZN(n8748) );
  NAND2_X1 U11264 ( .A1(n8748), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13714) );
  NAND2_X1 U11265 ( .A1(n8749), .A2(n13714), .ZN(n8792) );
  NAND2_X1 U11266 ( .A1(n8750), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U11267 ( .A1(n8752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11268 ( .A1(n14225), .A2(n13645), .ZN(n13659) );
  NAND2_X1 U11269 ( .A1(n9127), .A2(n9120), .ZN(n8759) );
  NAND2_X1 U11270 ( .A1(n8757), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8758) );
  XNOR2_X2 U11271 ( .A(n8758), .B(n8755), .ZN(n14496) );
  AND2_X1 U11272 ( .A1(n8759), .A2(n11335), .ZN(n8791) );
  INV_X1 U11273 ( .A(n8791), .ZN(n8760) );
  NOR2_X1 U11274 ( .A1(n14517), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U11275 ( .A1(n12770), .A2(n8761), .B1(n12771), .B2(n9208), .C1(
        n12305), .C2(P3_U3151), .ZN(P3_U3280) );
  NAND2_X1 U11276 ( .A1(n9635), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8764) );
  INV_X1 U11277 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8762) );
  MUX2_X1 U11278 ( .A(n8762), .B(P2_REG2_REG_8__SCAN_IN), .S(n9643), .Z(n8763)
         );
  NAND3_X1 U11279 ( .A1(n8765), .A2(n8764), .A3(n8763), .ZN(n8766) );
  NAND2_X1 U11280 ( .A1(n8766), .A2(n14791), .ZN(n8774) );
  NAND2_X1 U11281 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9761) );
  OAI21_X1 U11282 ( .B1(n9257), .B2(n6724), .A(n9761), .ZN(n8772) );
  NAND2_X1 U11283 ( .A1(n9635), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8768) );
  INV_X1 U11284 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14899) );
  MUX2_X1 U11285 ( .A(n14899), .B(P2_REG1_REG_8__SCAN_IN), .S(n9643), .Z(n8767) );
  AOI21_X1 U11286 ( .B1(n8769), .B2(n8768), .A(n8767), .ZN(n9032) );
  AND3_X1 U11287 ( .A1(n8769), .A2(n8768), .A3(n8767), .ZN(n8770) );
  NOR3_X1 U11288 ( .A1(n9032), .A2(n8770), .A3(n14742), .ZN(n8771) );
  AOI211_X1 U11289 ( .C1(n14790), .C2(n9643), .A(n8772), .B(n8771), .ZN(n8773)
         );
  OAI21_X1 U11290 ( .B1(n9027), .B2(n8774), .A(n8773), .ZN(P2_U3222) );
  MUX2_X1 U11291 ( .A(n8790), .B(n8786), .S(n11332), .Z(n8777) );
  NAND2_X1 U11292 ( .A1(n8777), .A2(n15232), .ZN(n8819) );
  INV_X1 U11293 ( .A(n8777), .ZN(n8778) );
  NAND2_X1 U11294 ( .A1(n8778), .A2(SI_12_), .ZN(n8779) );
  INV_X1 U11295 ( .A(n10607), .ZN(n8789) );
  NAND3_X1 U11296 ( .A1(n8782), .A2(n8781), .A3(n8780), .ZN(n8784) );
  NAND2_X1 U11297 ( .A1(n8784), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8783) );
  MUX2_X1 U11298 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8783), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8785) );
  INV_X1 U11299 ( .A(n12948), .ZN(n12933) );
  OAI222_X1 U11300 ( .A1(n13368), .A2(n8786), .B1(n13366), .B2(n8789), .C1(
        n12933), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U11301 ( .A1(n8788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8823) );
  XNOR2_X1 U11302 ( .A(n8823), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10608) );
  INV_X1 U11303 ( .A(n10608), .ZN(n14510) );
  OAI222_X1 U11304 ( .A1(n14223), .A2(n8790), .B1(n14221), .B2(n8789), .C1(
        n14510), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U11305 ( .A1(n8792), .A2(n8791), .ZN(n14499) );
  INV_X1 U11306 ( .A(n11594), .ZN(n9126) );
  INV_X1 U11307 ( .A(n13769), .ZN(n13763) );
  INV_X1 U11308 ( .A(n9598), .ZN(n8798) );
  INV_X1 U11309 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9074) );
  MUX2_X1 U11310 ( .A(n9074), .B(P1_REG1_REG_1__SCAN_IN), .S(n13736), .Z(n8794) );
  AND2_X1 U11311 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n8793) );
  NAND2_X1 U11312 ( .A1(n8794), .A2(n8793), .ZN(n13740) );
  INV_X1 U11313 ( .A(n13736), .ZN(n13741) );
  NAND2_X1 U11314 ( .A1(n13741), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U11315 ( .A1(n13740), .A2(n8795), .ZN(n9238) );
  INV_X1 U11316 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9128) );
  MUX2_X1 U11317 ( .A(n9128), .B(P1_REG1_REG_2__SCAN_IN), .S(n9285), .Z(n9239)
         );
  NAND2_X1 U11318 ( .A1(n9238), .A2(n9239), .ZN(n13750) );
  INV_X1 U11319 ( .A(n9285), .ZN(n9240) );
  NAND2_X1 U11320 ( .A1(n9240), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U11321 ( .A1(n13750), .A2(n13749), .ZN(n8797) );
  INV_X1 U11322 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9297) );
  MUX2_X1 U11323 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9297), .S(n13747), .Z(n8796) );
  NAND2_X1 U11324 ( .A1(n8797), .A2(n8796), .ZN(n13752) );
  NAND2_X1 U11325 ( .A1(n13747), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9272) );
  INV_X1 U11326 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14719) );
  MUX2_X1 U11327 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n14719), .S(n9598), .Z(n9273) );
  AOI21_X1 U11328 ( .B1(n13752), .B2(n9272), .A(n9273), .ZN(n9271) );
  AOI21_X1 U11329 ( .B1(n8798), .B2(P1_REG1_REG_4__SCAN_IN), .A(n9271), .ZN(
        n13765) );
  INV_X1 U11330 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14721) );
  MUX2_X1 U11331 ( .A(n14721), .B(P1_REG1_REG_5__SCAN_IN), .S(n13769), .Z(
        n13766) );
  NAND2_X1 U11332 ( .A1(n13765), .A2(n13766), .ZN(n13764) );
  OAI21_X1 U11333 ( .B1(n13763), .B2(P1_REG1_REG_5__SCAN_IN), .A(n13764), .ZN(
        n8859) );
  INV_X1 U11334 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10146) );
  MUX2_X1 U11335 ( .A(n10146), .B(P1_REG1_REG_6__SCAN_IN), .S(n9823), .Z(n8858) );
  NOR2_X1 U11336 ( .A1(n8859), .A2(n8858), .ZN(n8857) );
  NOR2_X1 U11337 ( .A1(n8868), .A2(n10146), .ZN(n8801) );
  INV_X1 U11338 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9849) );
  MUX2_X1 U11339 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9849), .S(n9971), .Z(n8800)
         );
  NOR3_X1 U11340 ( .A1(n8857), .A2(n8801), .A3(n8800), .ZN(n8799) );
  NOR2_X1 U11341 ( .A1(n14538), .A2(n8799), .ZN(n8813) );
  OAI21_X1 U11342 ( .B1(n8857), .B2(n8801), .A(n8800), .ZN(n8836) );
  OR2_X1 U11343 ( .A1(n11594), .A2(n14496), .ZN(n8802) );
  INV_X1 U11344 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10119) );
  MUX2_X1 U11345 ( .A(n10119), .B(P1_REG2_REG_1__SCAN_IN), .S(n13736), .Z(
        n13734) );
  AND2_X1 U11346 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13735) );
  NAND2_X1 U11347 ( .A1(n13734), .A2(n13735), .ZN(n13733) );
  NAND2_X1 U11348 ( .A1(n13741), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U11349 ( .A1(n13733), .A2(n8803), .ZN(n9236) );
  INV_X1 U11350 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9129) );
  MUX2_X1 U11351 ( .A(n9129), .B(P1_REG2_REG_2__SCAN_IN), .S(n9285), .Z(n9237)
         );
  NAND2_X1 U11352 ( .A1(n9236), .A2(n9237), .ZN(n13755) );
  NAND2_X1 U11353 ( .A1(n9240), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13754) );
  INV_X1 U11354 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n8804) );
  MUX2_X1 U11355 ( .A(n8804), .B(P1_REG2_REG_3__SCAN_IN), .S(n13747), .Z(
        n13753) );
  AOI21_X1 U11356 ( .B1(n13755), .B2(n13754), .A(n13753), .ZN(n8805) );
  INV_X1 U11357 ( .A(n8805), .ZN(n13757) );
  NAND2_X1 U11358 ( .A1(n13747), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9268) );
  INV_X1 U11359 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8806) );
  MUX2_X1 U11360 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n8806), .S(n9598), .Z(n9267)
         );
  AOI21_X1 U11361 ( .B1(n13757), .B2(n9268), .A(n9267), .ZN(n9266) );
  NOR2_X1 U11362 ( .A1(n9598), .A2(n8806), .ZN(n13768) );
  MUX2_X1 U11363 ( .A(n13770), .B(P1_REG2_REG_5__SCAN_IN), .S(n13769), .Z(
        n8807) );
  OAI21_X1 U11364 ( .B1(n9266), .B2(n13768), .A(n8807), .ZN(n13775) );
  NAND2_X1 U11365 ( .A1(n13763), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8861) );
  INV_X1 U11366 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9858) );
  MUX2_X1 U11367 ( .A(n9858), .B(P1_REG2_REG_6__SCAN_IN), .S(n9823), .Z(n8860)
         );
  AOI21_X1 U11368 ( .B1(n13775), .B2(n8861), .A(n8860), .ZN(n8863) );
  NOR2_X1 U11369 ( .A1(n8868), .A2(n9858), .ZN(n8809) );
  INV_X1 U11370 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9847) );
  MUX2_X1 U11371 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n9847), .S(n9971), .Z(n8808)
         );
  OAI21_X1 U11372 ( .B1(n8863), .B2(n8809), .A(n8808), .ZN(n8851) );
  INV_X1 U11373 ( .A(n8851), .ZN(n8811) );
  NOR3_X1 U11374 ( .A1(n8863), .A2(n8809), .A3(n8808), .ZN(n8810) );
  NOR3_X1 U11375 ( .A1(n14536), .A2(n8811), .A3(n8810), .ZN(n8812) );
  AOI21_X1 U11376 ( .B1(n8813), .B2(n8836), .A(n8812), .ZN(n8815) );
  AND2_X1 U11377 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10164) );
  AOI21_X1 U11378 ( .B1(n14517), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10164), .ZN(
        n8814) );
  OAI211_X1 U11379 ( .C1(n8837), .C2(n14553), .A(n8815), .B(n8814), .ZN(
        P1_U3250) );
  INV_X1 U11380 ( .A(n12333), .ZN(n12347) );
  OAI222_X1 U11381 ( .A1(n12770), .A2(n8816), .B1(n12347), .B2(P3_U3151), .C1(
        n15336), .C2(n12771), .ZN(P3_U3279) );
  NAND2_X1 U11382 ( .A1(n8817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8818) );
  XNOR2_X1 U11383 ( .A(n8818), .B(P2_IR_REG_13__SCAN_IN), .ZN(n14746) );
  INV_X1 U11384 ( .A(n14746), .ZN(n12935) );
  MUX2_X1 U11385 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n11332), .Z(n8998) );
  XNOR2_X1 U11386 ( .A(n8998), .B(n8999), .ZN(n8820) );
  XNOR2_X1 U11387 ( .A(n8997), .B(n8820), .ZN(n10696) );
  INV_X1 U11388 ( .A(n10696), .ZN(n8828) );
  INV_X1 U11389 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n8821) );
  OAI222_X1 U11390 ( .A1(P2_U3088), .A2(n12935), .B1(n13366), .B2(n8828), .C1(
        n8821), .C2(n13368), .ZN(P2_U3314) );
  NAND2_X1 U11391 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  NAND2_X1 U11392 ( .A1(n8824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8826) );
  NAND2_X1 U11393 ( .A1(n8826), .A2(n8825), .ZN(n9023) );
  OR2_X1 U11394 ( .A1(n8826), .A2(n8825), .ZN(n8827) );
  NAND2_X1 U11395 ( .A1(n9023), .A2(n8827), .ZN(n14520) );
  OAI222_X1 U11396 ( .A1(n14223), .A2(n10697), .B1(n14221), .B2(n8828), .C1(
        n14520), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U11397 ( .A(n14553), .ZN(n13797) );
  INV_X1 U11398 ( .A(n14517), .ZN(n14557) );
  INV_X1 U11399 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14251) );
  NAND2_X1 U11400 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10515) );
  OAI21_X1 U11401 ( .B1(n14557), .B2(n14251), .A(n10515), .ZN(n8835) );
  NAND2_X1 U11402 ( .A1(n9971), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8850) );
  INV_X1 U11403 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10001) );
  MUX2_X1 U11404 ( .A(n10001), .B(P1_REG2_REG_8__SCAN_IN), .S(n9977), .Z(n8849) );
  AOI21_X1 U11405 ( .B1(n8851), .B2(n8850), .A(n8849), .ZN(n8848) );
  NOR2_X1 U11406 ( .A1(n8829), .A2(n10001), .ZN(n8831) );
  INV_X1 U11407 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9989) );
  MUX2_X1 U11408 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9989), .S(n10330), .Z(n8830) );
  OAI21_X1 U11409 ( .B1(n8848), .B2(n8831), .A(n8830), .ZN(n8934) );
  INV_X1 U11410 ( .A(n8934), .ZN(n8833) );
  NOR3_X1 U11411 ( .A1(n8848), .A2(n8831), .A3(n8830), .ZN(n8832) );
  NOR3_X1 U11412 ( .A1(n8833), .A2(n8832), .A3(n14536), .ZN(n8834) );
  AOI211_X1 U11413 ( .C1(n13797), .C2(n10330), .A(n8835), .B(n8834), .ZN(n8843) );
  OAI21_X1 U11414 ( .B1(n9849), .B2(n8837), .A(n8836), .ZN(n8845) );
  INV_X1 U11415 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9984) );
  MUX2_X1 U11416 ( .A(n9984), .B(P1_REG1_REG_8__SCAN_IN), .S(n9977), .Z(n8846)
         );
  NOR2_X1 U11417 ( .A1(n8845), .A2(n8846), .ZN(n8844) );
  NOR2_X1 U11418 ( .A1(n9977), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8838) );
  INV_X1 U11419 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14725) );
  MUX2_X1 U11420 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14725), .S(n10330), .Z(
        n8839) );
  OAI21_X1 U11421 ( .B1(n8844), .B2(n8838), .A(n8839), .ZN(n8937) );
  INV_X1 U11422 ( .A(n8937), .ZN(n8841) );
  NOR3_X1 U11423 ( .A1(n8844), .A2(n8839), .A3(n8838), .ZN(n8840) );
  OAI21_X1 U11424 ( .B1(n8841), .B2(n8840), .A(n14545), .ZN(n8842) );
  NAND2_X1 U11425 ( .A1(n8843), .A2(n8842), .ZN(P1_U3252) );
  AOI21_X1 U11426 ( .B1(n8846), .B2(n8845), .A(n8844), .ZN(n8856) );
  NAND2_X1 U11427 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10388) );
  OAI21_X1 U11428 ( .B1(n14557), .B2(n14249), .A(n10388), .ZN(n8847) );
  AOI21_X1 U11429 ( .B1(n9977), .B2(n13797), .A(n8847), .ZN(n8855) );
  INV_X1 U11430 ( .A(n8848), .ZN(n8853) );
  NAND3_X1 U11431 ( .A1(n8851), .A2(n8850), .A3(n8849), .ZN(n8852) );
  NAND3_X1 U11432 ( .A1(n8853), .A2(n14548), .A3(n8852), .ZN(n8854) );
  OAI211_X1 U11433 ( .C1(n8856), .C2(n14538), .A(n8855), .B(n8854), .ZN(
        P1_U3251) );
  AOI211_X1 U11434 ( .C1(n8859), .C2(n8858), .A(n8857), .B(n14538), .ZN(n8865)
         );
  AND3_X1 U11435 ( .A1(n13775), .A2(n8861), .A3(n8860), .ZN(n8862) );
  NOR3_X1 U11436 ( .A1(n14536), .A2(n8863), .A3(n8862), .ZN(n8864) );
  NOR2_X1 U11437 ( .A1(n8865), .A2(n8864), .ZN(n8867) );
  AND2_X1 U11438 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9914) );
  AOI21_X1 U11439 ( .B1(n14517), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9914), .ZN(
        n8866) );
  OAI211_X1 U11440 ( .C1(n8868), .C2(n14553), .A(n8867), .B(n8866), .ZN(
        P1_U3249) );
  OAI222_X1 U11441 ( .A1(n12770), .A2(n8869), .B1(n12771), .B2(n15257), .C1(
        n12371), .C2(P3_U3151), .ZN(P3_U3278) );
  NOR4_X1 U11442 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8873) );
  NOR4_X1 U11443 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8872) );
  NOR4_X1 U11444 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8871) );
  NOR4_X1 U11445 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8870) );
  NAND4_X1 U11446 ( .A1(n8873), .A2(n8872), .A3(n8871), .A4(n8870), .ZN(n8881)
         );
  NOR2_X1 U11447 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8877) );
  NOR4_X1 U11448 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8876) );
  NOR4_X1 U11449 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8875) );
  NOR4_X1 U11450 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8874) );
  NAND4_X1 U11451 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(n8880)
         );
  INV_X1 U11452 ( .A(n8886), .ZN(n10540) );
  XNOR2_X1 U11453 ( .A(n10442), .B(P2_B_REG_SCAN_IN), .ZN(n8878) );
  NAND2_X1 U11454 ( .A1(n10540), .A2(n8878), .ZN(n8879) );
  OAI21_X1 U11455 ( .B1(n8881), .B2(n8880), .A(n14799), .ZN(n9409) );
  INV_X1 U11456 ( .A(n8887), .ZN(n10749) );
  NAND2_X1 U11457 ( .A1(n10442), .A2(n10749), .ZN(n8884) );
  INV_X1 U11458 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U11459 ( .A1(n14799), .A2(n8882), .ZN(n8883) );
  NAND2_X1 U11460 ( .A1(n8884), .A2(n8883), .ZN(n14802) );
  INV_X1 U11461 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U11462 ( .A1(n14799), .A2(n8885), .ZN(n8889) );
  OR2_X1 U11463 ( .A1(n8887), .A2(n8886), .ZN(n8888) );
  NAND2_X1 U11464 ( .A1(n8889), .A2(n8888), .ZN(n14804) );
  NOR2_X1 U11465 ( .A1(n14802), .A2(n14804), .ZN(n8890) );
  NAND2_X1 U11466 ( .A1(n9409), .A2(n8890), .ZN(n8919) );
  NOR2_X2 U11467 ( .A1(n9212), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U11468 ( .A1(n9014), .A2(n8893), .ZN(n9200) );
  INV_X1 U11469 ( .A(n8916), .ZN(n8963) );
  NAND2_X1 U11470 ( .A1(n8894), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8896) );
  INV_X1 U11471 ( .A(n9463), .ZN(n8897) );
  INV_X1 U11472 ( .A(n8960), .ZN(n8898) );
  INV_X1 U11473 ( .A(n12877), .ZN(n12808) );
  INV_X1 U11474 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8903) );
  INV_X1 U11475 ( .A(n11726), .ZN(n8906) );
  NAND2_X1 U11476 ( .A1(n8906), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U11477 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  AND2_X1 U11478 ( .A1(n8914), .A2(n8913), .ZN(n13369) );
  INV_X1 U11479 ( .A(n9685), .ZN(n12003) );
  INV_X1 U11480 ( .A(n9668), .ZN(n11702) );
  NAND2_X1 U11481 ( .A1(n8915), .A2(n9668), .ZN(n8969) );
  NOR2_X1 U11482 ( .A1(n9463), .A2(n9685), .ZN(n9736) );
  NAND2_X1 U11483 ( .A1(n8923), .A2(n9736), .ZN(n8918) );
  OR2_X1 U11484 ( .A1(n9463), .A2(n9459), .ZN(n9410) );
  INV_X1 U11485 ( .A(n9410), .ZN(n8917) );
  AOI21_X1 U11486 ( .B1(n12808), .B2(n8969), .A(n12875), .ZN(n8931) );
  INV_X1 U11487 ( .A(n13244), .ZN(n9464) );
  NAND2_X1 U11488 ( .A1(n8919), .A2(n9410), .ZN(n8922) );
  NAND2_X1 U11489 ( .A1(n11993), .A2(n8960), .ZN(n9455) );
  AND3_X1 U11490 ( .A1(n9455), .A2(n8920), .A3(n10258), .ZN(n8921) );
  NAND2_X1 U11491 ( .A1(n8922), .A2(n8921), .ZN(n8947) );
  NOR2_X1 U11492 ( .A1(n8947), .A2(P2_U3088), .ZN(n9371) );
  INV_X1 U11493 ( .A(n9371), .ZN(n9225) );
  INV_X1 U11494 ( .A(n11993), .ZN(n12038) );
  INV_X1 U11495 ( .A(n12897), .ZN(n8928) );
  NAND2_X1 U11496 ( .A1(n8960), .A2(n8622), .ZN(n12988) );
  NOR2_X1 U11497 ( .A1(n8928), .A2(n12988), .ZN(n9461) );
  AOI22_X1 U11498 ( .A1(n9225), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n12871), .B2(
        n9461), .ZN(n8930) );
  INV_X1 U11499 ( .A(n12828), .ZN(n11651) );
  NAND3_X1 U11500 ( .A1(n11651), .A2(n12898), .A3(n13241), .ZN(n8929) );
  OAI211_X1 U11501 ( .C1(n8931), .C2(n9464), .A(n8930), .B(n8929), .ZN(
        P2_U3204) );
  NAND2_X1 U11502 ( .A1(n10330), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8933) );
  INV_X1 U11503 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10364) );
  MUX2_X1 U11504 ( .A(n10364), .B(P1_REG2_REG_10__SCAN_IN), .S(n10336), .Z(
        n8932) );
  AOI21_X1 U11505 ( .B1(n8934), .B2(n8933), .A(n8932), .ZN(n13786) );
  INV_X1 U11506 ( .A(n13786), .ZN(n8936) );
  NAND3_X1 U11507 ( .A1(n8934), .A2(n8933), .A3(n8932), .ZN(n8935) );
  NAND3_X1 U11508 ( .A1(n8936), .A2(n14548), .A3(n8935), .ZN(n8944) );
  NAND2_X1 U11509 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10650)
         );
  INV_X1 U11510 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14728) );
  MUX2_X1 U11511 ( .A(n14728), .B(P1_REG1_REG_10__SCAN_IN), .S(n10336), .Z(
        n8939) );
  OAI21_X1 U11512 ( .B1(n10330), .B2(P1_REG1_REG_9__SCAN_IN), .A(n8937), .ZN(
        n8938) );
  NOR2_X1 U11513 ( .A1(n8938), .A2(n8939), .ZN(n9435) );
  AOI211_X1 U11514 ( .C1(n8939), .C2(n8938), .A(n9435), .B(n14538), .ZN(n8940)
         );
  INV_X1 U11515 ( .A(n8940), .ZN(n8941) );
  NAND2_X1 U11516 ( .A1(n10650), .A2(n8941), .ZN(n8942) );
  AOI21_X1 U11517 ( .B1(n14517), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n8942), .ZN(
        n8943) );
  OAI211_X1 U11518 ( .C1(n14553), .C2(n9442), .A(n8944), .B(n8943), .ZN(
        P1_U3253) );
  INV_X4 U11519 ( .A(n11953), .ZN(n11507) );
  INV_X2 U11520 ( .A(n8968), .ZN(n11506) );
  INV_X1 U11521 ( .A(n11786), .ZN(n11790) );
  INV_X1 U11522 ( .A(n12873), .ZN(n12861) );
  INV_X1 U11523 ( .A(n12871), .ZN(n12859) );
  NAND2_X1 U11524 ( .A1(n11959), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8954) );
  OR2_X1 U11525 ( .A1(n11962), .A2(n8654), .ZN(n8953) );
  OR2_X1 U11526 ( .A1(n6950), .A2(n14893), .ZN(n8952) );
  INV_X1 U11527 ( .A(n9334), .ZN(n9336) );
  INV_X1 U11528 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9748) );
  INV_X1 U11529 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U11530 ( .A1(n9748), .A2(n8949), .ZN(n8950) );
  NAND2_X1 U11531 ( .A1(n9336), .A2(n8950), .ZN(n9345) );
  OR2_X1 U11532 ( .A1(n8956), .A2(n9345), .ZN(n8951) );
  INV_X1 U11533 ( .A(n12894), .ZN(n12827) );
  INV_X1 U11534 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8957) );
  INV_X1 U11535 ( .A(n8622), .ZN(n8959) );
  INV_X1 U11536 ( .A(n13020), .ZN(n12775) );
  OAI22_X1 U11537 ( .A1(n12827), .A2(n12988), .B1(n9224), .B2(n12775), .ZN(
        n9426) );
  INV_X1 U11538 ( .A(n9426), .ZN(n8961) );
  NAND2_X1 U11539 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n12915) );
  OAI21_X1 U11540 ( .B1(n12859), .B2(n8961), .A(n12915), .ZN(n8962) );
  AOI21_X1 U11541 ( .B1(n12861), .B2(n9748), .A(n8962), .ZN(n8995) );
  NAND2_X1 U11542 ( .A1(n12897), .A2(n9668), .ZN(n8972) );
  INV_X1 U11543 ( .A(n12042), .ZN(n11956) );
  XNOR2_X1 U11544 ( .A(n11956), .B(n11762), .ZN(n8964) );
  NAND2_X2 U11545 ( .A1(n8964), .A2(n8963), .ZN(n14871) );
  NAND2_X1 U11546 ( .A1(n9464), .A2(n11579), .ZN(n9223) );
  INV_X1 U11547 ( .A(n9372), .ZN(n8971) );
  NAND2_X1 U11548 ( .A1(n8972), .A2(n8971), .ZN(n8973) );
  NAND2_X1 U11549 ( .A1(n9373), .A2(n8973), .ZN(n8977) );
  NAND2_X1 U11550 ( .A1(n12896), .A2(n9668), .ZN(n8980) );
  NAND2_X1 U11551 ( .A1(n9281), .A2(n6486), .ZN(n8975) );
  XNOR2_X1 U11552 ( .A(n11781), .B(n9327), .ZN(n8978) );
  XNOR2_X1 U11553 ( .A(n8980), .B(n8978), .ZN(n9374) );
  NAND2_X1 U11554 ( .A1(n8977), .A2(n9374), .ZN(n9380) );
  INV_X1 U11555 ( .A(n8978), .ZN(n8979) );
  NAND2_X1 U11556 ( .A1(n8980), .A2(n8979), .ZN(n8981) );
  NAND2_X1 U11557 ( .A1(n8982), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8987) );
  OR2_X1 U11558 ( .A1(n6950), .A2(n12906), .ZN(n8986) );
  INV_X1 U11559 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8983) );
  OR2_X1 U11560 ( .A1(n11743), .A2(n8983), .ZN(n8984) );
  NAND2_X1 U11561 ( .A1(n12895), .A2(n9668), .ZN(n8988) );
  OR2_X1 U11562 ( .A1(n9332), .A2(n8988), .ZN(n9328) );
  NAND2_X1 U11563 ( .A1(n9332), .A2(n8988), .ZN(n8989) );
  NAND2_X1 U11564 ( .A1(n9328), .A2(n8989), .ZN(n8991) );
  AOI21_X1 U11565 ( .B1(n8990), .B2(n8991), .A(n12877), .ZN(n8993) );
  NAND2_X1 U11566 ( .A1(n8993), .A2(n9329), .ZN(n8994) );
  OAI211_X1 U11567 ( .C1(n11790), .C2(n12865), .A(n8995), .B(n8994), .ZN(
        P2_U3190) );
  NAND2_X1 U11568 ( .A1(n8998), .A2(SI_13_), .ZN(n8996) );
  INV_X1 U11569 ( .A(n8998), .ZN(n9000) );
  NAND2_X1 U11570 ( .A1(n9000), .A2(n8999), .ZN(n9001) );
  MUX2_X1 U11571 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n11332), .Z(n9206) );
  INV_X1 U11572 ( .A(n9206), .ZN(n9003) );
  MUX2_X1 U11573 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n11332), .Z(n9209) );
  NAND2_X1 U11574 ( .A1(n9209), .A2(SI_15_), .ZN(n9007) );
  OAI21_X1 U11575 ( .B1(n9003), .B2(n15322), .A(n9007), .ZN(n9004) );
  INV_X1 U11576 ( .A(n9004), .ZN(n9005) );
  NOR2_X1 U11577 ( .A1(n9206), .A2(SI_14_), .ZN(n9008) );
  INV_X1 U11578 ( .A(n9209), .ZN(n9006) );
  AOI22_X1 U11579 ( .A1(n9008), .A2(n9007), .B1(n9006), .B2(n9208), .ZN(n9009)
         );
  MUX2_X1 U11580 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n11332), .Z(n9192) );
  XNOR2_X1 U11581 ( .A(n9192), .B(n15336), .ZN(n9190) );
  XNOR2_X1 U11582 ( .A(n9191), .B(n9190), .ZN(n11258) );
  INV_X1 U11583 ( .A(n11258), .ZN(n9018) );
  NAND2_X1 U11584 ( .A1(n9010), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9011) );
  MUX2_X1 U11585 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9011), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9012) );
  AND2_X1 U11586 ( .A1(n9012), .A2(n9197), .ZN(n13796) );
  INV_X1 U11587 ( .A(n13796), .ZN(n10419) );
  OAI222_X1 U11588 ( .A1(n14223), .A2(n9013), .B1(n14221), .B2(n9018), .C1(
        n10419), .C2(P1_U3086), .ZN(P1_U3339) );
  NOR2_X1 U11589 ( .A1(n9014), .A2(n7012), .ZN(n9015) );
  MUX2_X1 U11590 ( .A(n7012), .B(n9015), .S(P2_IR_REG_16__SCAN_IN), .Z(n9017)
         );
  INV_X1 U11591 ( .A(n9200), .ZN(n9016) );
  NOR2_X1 U11592 ( .A1(n9017), .A2(n9016), .ZN(n14773) );
  INV_X1 U11593 ( .A(n14773), .ZN(n12953) );
  OAI222_X1 U11594 ( .A1(n13368), .A2(n9019), .B1(n13366), .B2(n9018), .C1(
        n12953), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U11595 ( .A(n12395), .ZN(n12378) );
  OAI222_X1 U11596 ( .A1(n12770), .A2(n9020), .B1(n12771), .B2(n15344), .C1(
        n12378), .C2(P3_U3151), .ZN(P3_U3277) );
  XNOR2_X1 U11597 ( .A(n9204), .B(n15322), .ZN(n9207) );
  XNOR2_X1 U11598 ( .A(n9207), .B(n9206), .ZN(n10704) );
  INV_X1 U11599 ( .A(n10704), .ZN(n9025) );
  XNOR2_X1 U11600 ( .A(n9021), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12949) );
  INV_X1 U11601 ( .A(n12949), .ZN(n14752) );
  OAI222_X1 U11602 ( .A1(n13368), .A2(n9022), .B1(n13366), .B2(n9025), .C1(
        n14752), .C2(P2_U3088), .ZN(P2_U3313) );
  NAND2_X1 U11603 ( .A1(n9023), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9024) );
  XNOR2_X1 U11604 ( .A(n9024), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10705) );
  INV_X1 U11605 ( .A(n10705), .ZN(n10416) );
  OAI222_X1 U11606 ( .A1(n14223), .A2(n9026), .B1(n14221), .B2(n9025), .C1(
        n10416), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U11607 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9028) );
  MUX2_X1 U11608 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9028), .S(n12926), .Z(
        n12918) );
  NAND2_X1 U11609 ( .A1(n12919), .A2(n12918), .ZN(n12917) );
  OAI21_X1 U11610 ( .B1(n12926), .B2(P2_REG2_REG_9__SCAN_IN), .A(n12917), .ZN(
        n9031) );
  INV_X1 U11611 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9029) );
  MUX2_X1 U11612 ( .A(n9029), .B(P2_REG2_REG_10__SCAN_IN), .S(n10172), .Z(
        n9030) );
  AOI211_X1 U11613 ( .C1(n9031), .C2(n9030), .A(n14733), .B(n9248), .ZN(n9040)
         );
  AOI21_X1 U11614 ( .B1(n9643), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9032), .ZN(
        n12924) );
  INV_X1 U11615 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n14901) );
  MUX2_X1 U11616 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14901), .S(n12926), .Z(
        n12923) );
  NAND2_X1 U11617 ( .A1(n12924), .A2(n12923), .ZN(n12922) );
  OAI21_X1 U11618 ( .B1(n12926), .B2(P2_REG1_REG_9__SCAN_IN), .A(n12922), .ZN(
        n9035) );
  INV_X1 U11619 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14903) );
  MUX2_X1 U11620 ( .A(n14903), .B(P2_REG1_REG_10__SCAN_IN), .S(n10172), .Z(
        n9034) );
  INV_X1 U11621 ( .A(n9260), .ZN(n9033) );
  AOI211_X1 U11622 ( .C1(n9035), .C2(n9034), .A(n14742), .B(n9033), .ZN(n9039)
         );
  NAND2_X1 U11623 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10263)
         );
  NAND2_X1 U11624 ( .A1(n14784), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n9036) );
  OAI211_X1 U11625 ( .C1(n9395), .C2(n9037), .A(n10263), .B(n9036), .ZN(n9038)
         );
  OR3_X1 U11626 ( .A1(n9040), .A2(n9039), .A3(n9038), .ZN(P2_U3224) );
  NAND2_X1 U11627 ( .A1(n9041), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9043) );
  AND2_X2 U11628 ( .A1(n9122), .A2(n9838), .ZN(n9068) );
  INV_X1 U11629 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14210) );
  NAND2_X1 U11630 ( .A1(n9047), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9049) );
  XNOR2_X1 U11631 ( .A(n9049), .B(n9048), .ZN(n9051) );
  NAND2_X1 U11632 ( .A1(n11632), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9060) );
  INV_X2 U11633 ( .A(n9054), .ZN(n9055) );
  NAND2_X4 U11634 ( .A1(n9055), .A2(n9053), .ZN(n9585) );
  INV_X1 U11635 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9052) );
  OR2_X1 U11636 ( .A1(n9585), .A2(n9052), .ZN(n9059) );
  INV_X1 U11637 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14495) );
  OR2_X1 U11638 ( .A1(n6463), .A2(n14495), .ZN(n9058) );
  INV_X1 U11639 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9056) );
  OR2_X1 U11640 ( .A1(n13638), .A2(n9056), .ZN(n9057) );
  NAND2_X1 U11641 ( .A1(n11367), .A2(n13732), .ZN(n9067) );
  INV_X1 U11642 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13738) );
  INV_X1 U11643 ( .A(SI_0_), .ZN(n9062) );
  OAI21_X1 U11644 ( .B1(n11332), .B2(n9062), .A(n9061), .ZN(n9063) );
  NAND2_X1 U11645 ( .A1(n9064), .A2(n9063), .ZN(n14226) );
  MUX2_X1 U11646 ( .A(n13738), .B(n14226), .S(n11335), .Z(n14618) );
  INV_X1 U11647 ( .A(n14618), .ZN(n14632) );
  INV_X1 U11648 ( .A(n9122), .ZN(n9065) );
  AOI22_X1 U11649 ( .A1(n11436), .A2(n14632), .B1(n9065), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9066) );
  NAND2_X1 U11650 ( .A1(n13732), .A2(n11234), .ZN(n9071) );
  OAI22_X1 U11651 ( .A1(n11476), .A2(n14618), .B1(n14495), .B2(n9122), .ZN(
        n9069) );
  INV_X1 U11652 ( .A(n9069), .ZN(n9070) );
  NAND2_X1 U11653 ( .A1(n9071), .A2(n9070), .ZN(n9186) );
  NAND2_X1 U11654 ( .A1(n9187), .A2(n9186), .ZN(n9185) );
  OR2_X1 U11655 ( .A1(n9186), .A2(n11410), .ZN(n9073) );
  NAND2_X1 U11656 ( .A1(n11632), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9078) );
  INV_X1 U11657 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10109) );
  OR2_X1 U11658 ( .A1(n9585), .A2(n10109), .ZN(n9077) );
  OR2_X1 U11659 ( .A1(n6463), .A2(n9074), .ZN(n9076) );
  NAND4_X2 U11660 ( .A1(n9078), .A2(n9077), .A3(n9076), .A4(n9075), .ZN(n13731) );
  NAND2_X1 U11661 ( .A1(n11367), .A2(n13731), .ZN(n9083) );
  NAND2_X4 U11662 ( .A1(n11335), .A2(n11332), .ZN(n13653) );
  OR2_X1 U11663 ( .A1(n13653), .A2(n7611), .ZN(n9080) );
  NAND2_X1 U11664 ( .A1(n6668), .A2(n11234), .ZN(n9082) );
  INV_X1 U11665 ( .A(n9087), .ZN(n9086) );
  NAND2_X1 U11666 ( .A1(n13731), .A2(n11234), .ZN(n9084) );
  INV_X1 U11667 ( .A(n9088), .ZN(n9085) );
  NAND2_X1 U11668 ( .A1(n9086), .A2(n9085), .ZN(n9089) );
  NAND2_X1 U11669 ( .A1(n9088), .A2(n9087), .ZN(n9292) );
  NAND2_X1 U11670 ( .A1(n9089), .A2(n9292), .ZN(n9093) );
  INV_X1 U11671 ( .A(n9094), .ZN(n9091) );
  INV_X1 U11672 ( .A(n9093), .ZN(n9090) );
  NAND2_X1 U11673 ( .A1(n9091), .A2(n9090), .ZN(n9293) );
  INV_X1 U11674 ( .A(n9293), .ZN(n9092) );
  AOI21_X1 U11675 ( .B1(n9094), .B2(n9093), .A(n9092), .ZN(n9136) );
  INV_X1 U11676 ( .A(n10747), .ZN(n10948) );
  AND2_X1 U11677 ( .A1(n9096), .A2(n10948), .ZN(n9099) );
  NAND3_X1 U11678 ( .A1(n9097), .A2(P1_B_REG_SCAN_IN), .A3(n9095), .ZN(n9098)
         );
  NAND2_X1 U11679 ( .A1(n9095), .A2(n10747), .ZN(n9100) );
  NAND2_X1 U11680 ( .A1(n9101), .A2(n9100), .ZN(n9833) );
  NOR4_X1 U11681 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9110) );
  NOR4_X1 U11682 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9109) );
  NOR4_X1 U11683 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9105) );
  NOR4_X1 U11684 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9104) );
  NOR4_X1 U11685 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9103) );
  NOR4_X1 U11686 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9102) );
  NAND4_X1 U11687 ( .A1(n9105), .A2(n9104), .A3(n9103), .A4(n9102), .ZN(n9106)
         );
  NOR4_X1 U11688 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9107), .A4(n9106), .ZN(n9108) );
  AND3_X1 U11689 ( .A1(n9110), .A2(n9109), .A3(n9108), .ZN(n9111) );
  NOR2_X1 U11690 ( .A1(n10946), .A2(n9111), .ZN(n9834) );
  OR2_X1 U11691 ( .A1(n10946), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U11692 ( .A1(n9097), .A2(n10747), .ZN(n9112) );
  OR2_X1 U11693 ( .A1(n10145), .A2(n11638), .ZN(n9118) );
  INV_X1 U11694 ( .A(n9118), .ZN(n9114) );
  NAND2_X1 U11695 ( .A1(n9114), .A2(n10947), .ZN(n9125) );
  NAND2_X1 U11696 ( .A1(n14633), .A2(n13664), .ZN(n9857) );
  NAND2_X1 U11697 ( .A1(n14633), .A2(n13489), .ZN(n9115) );
  NAND2_X1 U11698 ( .A1(n9857), .A2(n9115), .ZN(n14701) );
  OR2_X1 U11699 ( .A1(n9125), .A2(n9857), .ZN(n9117) );
  NAND2_X1 U11700 ( .A1(n9118), .A2(n10143), .ZN(n9606) );
  NAND2_X1 U11701 ( .A1(n14614), .A2(n13656), .ZN(n9119) );
  NAND2_X1 U11702 ( .A1(n9127), .A2(n9119), .ZN(n9123) );
  AND2_X1 U11703 ( .A1(n9123), .A2(n9120), .ZN(n9121) );
  NAND2_X1 U11704 ( .A1(n9122), .A2(n9121), .ZN(n9604) );
  NAND2_X1 U11705 ( .A1(n9606), .A2(n13711), .ZN(n9303) );
  AOI22_X1 U11706 ( .A1(n14415), .A2(n6668), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9303), .ZN(n9135) );
  INV_X1 U11707 ( .A(n9123), .ZN(n9124) );
  AND2_X2 U11708 ( .A1(n9127), .A2(n9126), .ZN(n14683) );
  INV_X1 U11709 ( .A(n14683), .ZN(n14704) );
  INV_X1 U11710 ( .A(n14427), .ZN(n13442) );
  INV_X1 U11711 ( .A(n14635), .ZN(n14615) );
  INV_X1 U11712 ( .A(n14426), .ZN(n9799) );
  NAND2_X1 U11713 ( .A1(n11632), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9133) );
  INV_X1 U11714 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10123) );
  OR2_X1 U11715 ( .A1(n9585), .A2(n10123), .ZN(n9132) );
  OR2_X1 U11716 ( .A1(n9589), .A2(n9128), .ZN(n9131) );
  OR2_X1 U11717 ( .A1(n13638), .A2(n9129), .ZN(n9130) );
  AOI22_X1 U11718 ( .A1(n13442), .A2(n13732), .B1(n9799), .B2(n14636), .ZN(
        n9134) );
  OAI211_X1 U11719 ( .C1(n9136), .C2(n14410), .A(n9135), .B(n9134), .ZN(
        P1_U3222) );
  AND2_X1 U11720 ( .A1(n15094), .A2(n12707), .ZN(n10959) );
  NOR2_X1 U11721 ( .A1(n15088), .A2(n10959), .ZN(n11127) );
  INV_X1 U11722 ( .A(n12214), .ZN(n12193) );
  AOI22_X1 U11723 ( .A1(n12234), .A2(n12211), .B1(n12193), .B2(n9700), .ZN(
        n9138) );
  NAND2_X1 U11724 ( .A1(n12191), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9514) );
  NAND2_X1 U11725 ( .A1(n9514), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9137) );
  OAI211_X1 U11726 ( .C1(n11127), .C2(n12219), .A(n9138), .B(n9137), .ZN(
        P3_U3172) );
  NAND2_X1 U11727 ( .A1(n11093), .A2(n9141), .ZN(n9139) );
  AND2_X1 U11728 ( .A1(n9140), .A2(n9139), .ZN(n9166) );
  OR2_X1 U11729 ( .A1(n9141), .A2(P3_U3151), .ZN(n11162) );
  NAND2_X1 U11730 ( .A1(n9693), .A2(n11162), .ZN(n9165) );
  AND2_X1 U11731 ( .A1(n9166), .A2(n9165), .ZN(n9164) );
  MUX2_X1 U11732 ( .A(P3_U3897), .B(n9164), .S(n8212), .Z(n14983) );
  INV_X1 U11733 ( .A(n9172), .ZN(n9498) );
  INV_X1 U11734 ( .A(n9142), .ZN(n9143) );
  INV_X1 U11735 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15087) );
  INV_X1 U11736 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U11737 ( .A1(n9145), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9146) );
  INV_X1 U11738 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15109) );
  NAND2_X1 U11739 ( .A1(n9319), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9147) );
  INV_X1 U11740 ( .A(n14924), .ZN(n9173) );
  INV_X1 U11741 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n14929) );
  NOR2_X1 U11742 ( .A1(n9149), .A2(n14930), .ZN(n9151) );
  INV_X1 U11743 ( .A(n9151), .ZN(n9153) );
  INV_X1 U11744 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10081) );
  MUX2_X1 U11745 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10081), .S(n9172), .Z(n9150) );
  INV_X1 U11746 ( .A(n9150), .ZN(n9152) );
  OAI21_X1 U11747 ( .B1(n9153), .B2(n9152), .A(n9482), .ZN(n9171) );
  INV_X1 U11748 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15167) );
  MUX2_X1 U11749 ( .A(n15167), .B(P3_REG1_REG_2__SCAN_IN), .S(n9177), .Z(n9310) );
  NAND2_X1 U11750 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n14915), .ZN(n9156) );
  NAND2_X1 U11751 ( .A1(n9365), .A2(n9156), .ZN(n9155) );
  INV_X1 U11752 ( .A(n9156), .ZN(n14910) );
  NAND2_X1 U11753 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n14910), .ZN(n9154) );
  NAND2_X1 U11754 ( .A1(n9155), .A2(n9154), .ZN(n9355) );
  NAND2_X1 U11755 ( .A1(n9355), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9354) );
  OR2_X1 U11756 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9156), .ZN(n9157) );
  NAND2_X1 U11757 ( .A1(n9354), .A2(n9157), .ZN(n9309) );
  NAND2_X1 U11758 ( .A1(n9319), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9158) );
  INV_X1 U11759 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15169) );
  INV_X1 U11760 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9161) );
  MUX2_X1 U11761 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n9161), .S(n9172), .Z(n9162)
         );
  AOI21_X1 U11762 ( .B1(n9163), .B2(n9162), .A(n9497), .ZN(n9169) );
  INV_X2 U11763 ( .A(n6812), .ZN(n12369) );
  NAND2_X1 U11764 ( .A1(n9164), .A2(n12369), .ZN(n14977) );
  INV_X1 U11765 ( .A(n9165), .ZN(n9167) );
  INV_X1 U11766 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15230) );
  NOR2_X1 U11767 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15230), .ZN(n10014) );
  AOI21_X1 U11768 ( .B1(n14996), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10014), .ZN(
        n9168) );
  OAI21_X1 U11769 ( .B1(n9169), .B2(n14977), .A(n9168), .ZN(n9170) );
  AOI21_X1 U11770 ( .B1(n14997), .B2(n9171), .A(n9170), .ZN(n9184) );
  MUX2_X1 U11771 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12369), .Z(n9488) );
  XNOR2_X1 U11772 ( .A(n9488), .B(n9172), .ZN(n9181) );
  MUX2_X1 U11773 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12369), .Z(n9174) );
  OR2_X1 U11774 ( .A1(n9174), .A2(n9173), .ZN(n9179) );
  XNOR2_X1 U11775 ( .A(n9174), .B(n14924), .ZN(n14922) );
  INV_X1 U11776 ( .A(n9365), .ZN(n9176) );
  MUX2_X1 U11777 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12369), .Z(n9178) );
  XOR2_X1 U11778 ( .A(n9177), .B(n9178), .Z(n9306) );
  OAI21_X1 U11779 ( .B1(n9181), .B2(n9180), .A(n9489), .ZN(n9182) );
  NAND2_X1 U11780 ( .A1(P3_U3897), .A2(n8212), .ZN(n14911) );
  NAND2_X1 U11781 ( .A1(n9182), .A2(n15007), .ZN(n9183) );
  OAI211_X1 U11782 ( .C1(n14993), .C2(n9498), .A(n9184), .B(n9183), .ZN(
        P3_U3186) );
  INV_X1 U11783 ( .A(n13731), .ZN(n14616) );
  OAI21_X1 U11784 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(n9232) );
  AOI22_X1 U11785 ( .A1(n14431), .A2(n9232), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9303), .ZN(n9189) );
  NAND2_X1 U11786 ( .A1(n14415), .A2(n14632), .ZN(n9188) );
  OAI211_X1 U11787 ( .C1(n14616), .C2(n14426), .A(n9189), .B(n9188), .ZN(
        P1_U3232) );
  INV_X1 U11788 ( .A(n9192), .ZN(n9193) );
  NAND2_X1 U11789 ( .A1(n9193), .A2(n15336), .ZN(n9194) );
  MUX2_X1 U11790 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n11332), .Z(n9468) );
  XNOR2_X1 U11791 ( .A(n9468), .B(n15257), .ZN(n9196) );
  XNOR2_X1 U11792 ( .A(n9469), .B(n9196), .ZN(n11268) );
  INV_X1 U11793 ( .A(n11268), .ZN(n9202) );
  NAND2_X1 U11794 ( .A1(n9197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9198) );
  XNOR2_X1 U11795 ( .A(n9198), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11269) );
  INV_X1 U11796 ( .A(n11269), .ZN(n10790) );
  OAI222_X1 U11797 ( .A1(n14223), .A2(n9199), .B1(n14221), .B2(n9202), .C1(
        n10790), .C2(P1_U3086), .ZN(P1_U3338) );
  NAND2_X1 U11798 ( .A1(n9200), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9201) );
  XNOR2_X1 U11799 ( .A(n9201), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14789) );
  INV_X1 U11800 ( .A(n14789), .ZN(n12956) );
  OAI222_X1 U11801 ( .A1(n13368), .A2(n9203), .B1(n13366), .B2(n9202), .C1(
        n12956), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U11802 ( .A(n9204), .ZN(n9205) );
  OAI22_X1 U11803 ( .A1(n9207), .A2(n9206), .B1(n9205), .B2(SI_14_), .ZN(n9211) );
  XNOR2_X1 U11804 ( .A(n9209), .B(n9208), .ZN(n9210) );
  XNOR2_X1 U11805 ( .A(n9211), .B(n9210), .ZN(n10926) );
  INV_X1 U11806 ( .A(n10926), .ZN(n9220) );
  NAND2_X1 U11807 ( .A1(n9212), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9213) );
  XNOR2_X1 U11808 ( .A(n9213), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14764) );
  INV_X1 U11809 ( .A(n14764), .ZN(n12940) );
  OAI222_X1 U11810 ( .A1(n13368), .A2(n9214), .B1(n13366), .B2(n9220), .C1(
        n12940), .C2(P2_U3088), .ZN(P2_U3312) );
  NAND2_X1 U11811 ( .A1(n9216), .A2(n9215), .ZN(n9217) );
  NAND2_X1 U11812 ( .A1(n9217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9218) );
  MUX2_X1 U11813 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9218), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9219) );
  AND2_X1 U11814 ( .A1(n9219), .A2(n9010), .ZN(n10927) );
  INV_X1 U11815 ( .A(n10927), .ZN(n14539) );
  OAI222_X1 U11816 ( .A1(n14223), .A2(n9221), .B1(n14221), .B2(n9220), .C1(
        n14539), .C2(P1_U3086), .ZN(P1_U3340) );
  OAI21_X1 U11817 ( .B1(n9223), .B2(n9222), .A(n9373), .ZN(n9229) );
  NOR3_X1 U11818 ( .A1(n12828), .A2(n9222), .A3(n13241), .ZN(n9228) );
  INV_X1 U11819 ( .A(n14814), .ZN(n9420) );
  OAI22_X1 U11820 ( .A1(n6906), .A2(n12775), .B1(n9224), .B2(n12988), .ZN(
        n13250) );
  AOI22_X1 U11821 ( .A1(n9225), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n12871), .B2(
        n13250), .ZN(n9226) );
  OAI21_X1 U11822 ( .B1(n9420), .B2(n12865), .A(n9226), .ZN(n9227) );
  AOI211_X1 U11823 ( .C1(n12808), .C2(n9229), .A(n9228), .B(n9227), .ZN(n9230)
         );
  INV_X1 U11824 ( .A(n9230), .ZN(P2_U3194) );
  NOR2_X1 U11825 ( .A1(n14496), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9231) );
  OR2_X1 U11826 ( .A1(n11594), .A2(n9231), .ZN(n14494) );
  INV_X1 U11827 ( .A(n13735), .ZN(n9233) );
  MUX2_X1 U11828 ( .A(n9233), .B(n9232), .S(n14496), .Z(n9234) );
  NOR2_X1 U11829 ( .A1(n9234), .A2(n11594), .ZN(n9235) );
  AOI211_X1 U11830 ( .C1(n13738), .C2(n14494), .A(n13721), .B(n9235), .ZN(
        n9279) );
  AOI22_X1 U11831 ( .A1(n14517), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9244) );
  OAI211_X1 U11832 ( .C1(n9237), .C2(n9236), .A(n14548), .B(n13755), .ZN(n9243) );
  OAI211_X1 U11833 ( .C1(n9239), .C2(n9238), .A(n14545), .B(n13750), .ZN(n9242) );
  NAND2_X1 U11834 ( .A1(n13797), .A2(n9240), .ZN(n9241) );
  NAND4_X1 U11835 ( .A1(n9244), .A2(n9243), .A3(n9242), .A4(n9241), .ZN(n9245)
         );
  OR2_X1 U11836 ( .A1(n9279), .A2(n9245), .ZN(P1_U3245) );
  OAI222_X1 U11837 ( .A1(P3_U3151), .A2(n9247), .B1(n12771), .B2(n15267), .C1(
        n12770), .C2(n9246), .ZN(P3_U3276) );
  INV_X1 U11838 ( .A(n9251), .ZN(n9254) );
  INV_X1 U11839 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9249) );
  MUX2_X1 U11840 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n9249), .S(n10178), .Z(
        n9250) );
  INV_X1 U11841 ( .A(n9250), .ZN(n9253) );
  INV_X1 U11842 ( .A(n9387), .ZN(n9252) );
  AOI21_X1 U11843 ( .B1(n9254), .B2(n9253), .A(n9252), .ZN(n9265) );
  INV_X1 U11844 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9256) );
  INV_X1 U11845 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9255) );
  OAI22_X1 U11846 ( .A1(n9257), .A2(n9256), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9255), .ZN(n9263) );
  NAND2_X1 U11847 ( .A1(n10172), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9259) );
  INV_X1 U11848 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14906) );
  MUX2_X1 U11849 ( .A(n14906), .B(P2_REG1_REG_11__SCAN_IN), .S(n10178), .Z(
        n9258) );
  AOI21_X1 U11850 ( .B1(n9260), .B2(n9259), .A(n9258), .ZN(n9389) );
  AND3_X1 U11851 ( .A1(n9260), .A2(n9259), .A3(n9258), .ZN(n9261) );
  NOR3_X1 U11852 ( .A1(n9389), .A2(n9261), .A3(n14742), .ZN(n9262) );
  AOI211_X1 U11853 ( .C1(n14790), .C2(n10178), .A(n9263), .B(n9262), .ZN(n9264) );
  OAI21_X1 U11854 ( .B1(n9265), .B2(n14733), .A(n9264), .ZN(P2_U3225) );
  INV_X1 U11855 ( .A(n9266), .ZN(n13773) );
  NAND3_X1 U11856 ( .A1(n13757), .A2(n9268), .A3(n9267), .ZN(n9269) );
  NAND3_X1 U11857 ( .A1(n14548), .A2(n13773), .A3(n9269), .ZN(n9270) );
  NAND2_X1 U11858 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9619) );
  OAI211_X1 U11859 ( .C1(n14237), .C2(n14557), .A(n9270), .B(n9619), .ZN(n9278) );
  INV_X1 U11860 ( .A(n9271), .ZN(n9275) );
  NAND3_X1 U11861 ( .A1(n9273), .A2(n13752), .A3(n9272), .ZN(n9274) );
  NAND2_X1 U11862 ( .A1(n9275), .A2(n9274), .ZN(n9276) );
  OAI22_X1 U11863 ( .A1(n9598), .A2(n14553), .B1(n14538), .B2(n9276), .ZN(
        n9277) );
  OR3_X1 U11864 ( .A1(n9279), .A2(n9278), .A3(n9277), .ZN(P1_U3247) );
  NAND2_X1 U11865 ( .A1(n10703), .A2(n9281), .ZN(n9284) );
  OR2_X1 U11866 ( .A1(n13653), .A2(n9282), .ZN(n9283) );
  INV_X1 U11867 ( .A(n13498), .ZN(n14649) );
  NAND2_X1 U11868 ( .A1(n14636), .A2(n11459), .ZN(n9287) );
  INV_X2 U11869 ( .A(n11476), .ZN(n11422) );
  NAND2_X1 U11870 ( .A1(n11422), .A2(n13498), .ZN(n9286) );
  NAND2_X1 U11871 ( .A1(n9287), .A2(n9286), .ZN(n9288) );
  XNOR2_X1 U11872 ( .A(n9288), .B(n11410), .ZN(n9571) );
  NAND2_X1 U11873 ( .A1(n11367), .A2(n14636), .ZN(n9291) );
  NAND2_X1 U11874 ( .A1(n11459), .A2(n13498), .ZN(n9290) );
  NAND2_X1 U11875 ( .A1(n9291), .A2(n9290), .ZN(n9569) );
  XNOR2_X1 U11876 ( .A(n9571), .B(n9569), .ZN(n9295) );
  NAND2_X1 U11877 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  NAND2_X1 U11878 ( .A1(n9294), .A2(n9295), .ZN(n9573) );
  OAI21_X1 U11879 ( .B1(n9295), .B2(n9294), .A(n9573), .ZN(n9296) );
  NAND2_X1 U11880 ( .A1(n9296), .A2(n14431), .ZN(n9305) );
  NAND2_X1 U11881 ( .A1(n11632), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9301) );
  OR2_X1 U11882 ( .A1(n9585), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9300) );
  OR2_X1 U11883 ( .A1(n13638), .A2(n8804), .ZN(n9299) );
  OR2_X1 U11884 ( .A1(n6463), .A2(n9297), .ZN(n9298) );
  NAND4_X1 U11885 ( .A1(n9301), .A2(n9300), .A3(n9299), .A4(n9298), .ZN(n13730) );
  INV_X1 U11886 ( .A(n13730), .ZN(n9302) );
  OAI22_X1 U11887 ( .A1(n14616), .A2(n14704), .B1(n9302), .B2(n14615), .ZN(
        n10129) );
  AOI22_X1 U11888 ( .A1(n14387), .A2(n10129), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n9303), .ZN(n9304) );
  OAI211_X1 U11889 ( .C1(n14649), .C2(n14423), .A(n9305), .B(n9304), .ZN(
        P1_U3237) );
  XNOR2_X1 U11890 ( .A(n9307), .B(n9306), .ZN(n9321) );
  INV_X1 U11891 ( .A(n14977), .ZN(n15005) );
  OAI21_X1 U11892 ( .B1(n9310), .B2(n9309), .A(n9308), .ZN(n9312) );
  INV_X1 U11893 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15253) );
  OAI22_X1 U11894 ( .A1(n14974), .A2(n14233), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15253), .ZN(n9311) );
  AOI21_X1 U11895 ( .B1(n15005), .B2(n9312), .A(n9311), .ZN(n9318) );
  OAI21_X1 U11896 ( .B1(n9315), .B2(n9314), .A(n9313), .ZN(n9316) );
  NAND2_X1 U11897 ( .A1(n14997), .A2(n9316), .ZN(n9317) );
  OAI211_X1 U11898 ( .C1(n14993), .C2(n9319), .A(n9318), .B(n9317), .ZN(n9320)
         );
  AOI21_X1 U11899 ( .B1(n9321), .B2(n15007), .A(n9320), .ZN(n9322) );
  INV_X1 U11900 ( .A(n9322), .ZN(P3_U3184) );
  NAND2_X1 U11901 ( .A1(n12894), .A2(n9668), .ZN(n9554) );
  NAND2_X1 U11902 ( .A1(n11506), .A2(n9323), .ZN(n9324) );
  OAI211_X1 U11903 ( .C1(n11953), .C2(n9326), .A(n9325), .B(n9324), .ZN(n11801) );
  OAI21_X1 U11904 ( .B1(n9330), .B2(n9329), .A(n12832), .ZN(n9351) );
  INV_X1 U11905 ( .A(n12895), .ZN(n9331) );
  NOR4_X1 U11906 ( .A1(n12828), .A2(n9332), .A3(n9331), .A4(n9330), .ZN(n9350)
         );
  NAND2_X1 U11907 ( .A1(n8982), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9342) );
  OR2_X1 U11908 ( .A1(n6950), .A2(n9333), .ZN(n9341) );
  INV_X1 U11909 ( .A(n9532), .ZN(n9542) );
  INV_X1 U11910 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U11911 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  NAND2_X1 U11912 ( .A1(n9542), .A2(n9337), .ZN(n12822) );
  OR2_X1 U11913 ( .A1(n11741), .A2(n12822), .ZN(n9340) );
  INV_X1 U11914 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9338) );
  OR2_X1 U11915 ( .A1(n11743), .A2(n9338), .ZN(n9339) );
  NAND2_X1 U11916 ( .A1(n12893), .A2(n12858), .ZN(n9344) );
  NAND2_X1 U11917 ( .A1(n12895), .A2(n13020), .ZN(n9343) );
  NAND2_X1 U11918 ( .A1(n9344), .A2(n9343), .ZN(n9727) );
  INV_X1 U11919 ( .A(n9727), .ZN(n9348) );
  INV_X1 U11920 ( .A(n9345), .ZN(n9740) );
  AOI22_X1 U11921 ( .A1(n11801), .A2(n12875), .B1(n12861), .B2(n9740), .ZN(
        n9347) );
  OAI211_X1 U11922 ( .C1(n9348), .C2(n12859), .A(n9347), .B(n9346), .ZN(n9349)
         );
  AOI211_X1 U11923 ( .C1(n12808), .C2(n9351), .A(n9350), .B(n9349), .ZN(n9352)
         );
  INV_X1 U11924 ( .A(n9352), .ZN(P2_U3202) );
  XNOR2_X1 U11925 ( .A(n9353), .B(n14912), .ZN(n9367) );
  OAI21_X1 U11926 ( .B1(n9355), .B2(P3_REG1_REG_1__SCAN_IN), .A(n9354), .ZN(
        n9358) );
  INV_X1 U11927 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n9356) );
  OAI22_X1 U11928 ( .A1(n14974), .A2(n14232), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9356), .ZN(n9357) );
  AOI21_X1 U11929 ( .B1(n15005), .B2(n9358), .A(n9357), .ZN(n9364) );
  NAND2_X1 U11930 ( .A1(n9359), .A2(n15109), .ZN(n9360) );
  NAND2_X1 U11931 ( .A1(n9361), .A2(n9360), .ZN(n9362) );
  NAND2_X1 U11932 ( .A1(n14997), .A2(n9362), .ZN(n9363) );
  OAI211_X1 U11933 ( .C1(n14993), .C2(n9365), .A(n9364), .B(n9363), .ZN(n9366)
         );
  AOI21_X1 U11934 ( .B1(n15007), .B2(n9367), .A(n9366), .ZN(n9368) );
  INV_X1 U11935 ( .A(n9368), .ZN(P3_U3183) );
  NAND2_X1 U11936 ( .A1(n12895), .A2(n12858), .ZN(n9370) );
  NAND2_X1 U11937 ( .A1(n12897), .A2(n13020), .ZN(n9369) );
  AND2_X1 U11938 ( .A1(n9370), .A2(n9369), .ZN(n10033) );
  OAI22_X1 U11939 ( .A1(n12859), .A2(n10033), .B1(n9371), .B2(n10041), .ZN(
        n9378) );
  AOI22_X1 U11940 ( .A1(n11651), .A2(n12897), .B1(n12808), .B2(n9372), .ZN(
        n9376) );
  INV_X1 U11941 ( .A(n9373), .ZN(n9375) );
  NOR3_X1 U11942 ( .A1(n9376), .A2(n9375), .A3(n9374), .ZN(n9377) );
  AOI211_X1 U11943 ( .C1(n11781), .C2(n12875), .A(n9378), .B(n9377), .ZN(n9379) );
  OAI21_X1 U11944 ( .B1(n9380), .B2(n12877), .A(n9379), .ZN(P2_U3209) );
  NAND2_X1 U11945 ( .A1(n9381), .A2(n9249), .ZN(n9386) );
  INV_X1 U11946 ( .A(n9386), .ZN(n9383) );
  INV_X1 U11947 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U11948 ( .A1(n12948), .A2(n12932), .ZN(n9382) );
  OAI21_X1 U11949 ( .B1(n12948), .B2(n12932), .A(n9382), .ZN(n9384) );
  NOR2_X1 U11950 ( .A1(n9383), .A2(n9384), .ZN(n9388) );
  INV_X1 U11951 ( .A(n9384), .ZN(n9385) );
  AOI21_X1 U11952 ( .B1(n9388), .B2(n9387), .A(n12931), .ZN(n9400) );
  INV_X1 U11953 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10501) );
  NOR2_X1 U11954 ( .A1(n12948), .A2(n10501), .ZN(n9390) );
  AOI21_X1 U11955 ( .B1(n10178), .B2(P2_REG1_REG_11__SCAN_IN), .A(n9389), .ZN(
        n9392) );
  AOI211_X1 U11956 ( .C1(n10501), .C2(n12948), .A(n9390), .B(n9392), .ZN(n9394) );
  NAND2_X1 U11957 ( .A1(n12948), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9391) );
  OAI211_X1 U11958 ( .C1(n12948), .C2(P2_REG1_REG_12__SCAN_IN), .A(n9392), .B(
        n9391), .ZN(n12947) );
  INV_X1 U11959 ( .A(n12947), .ZN(n9393) );
  OAI21_X1 U11960 ( .B1(n9394), .B2(n9393), .A(n14785), .ZN(n9399) );
  NOR2_X1 U11961 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10193), .ZN(n9397) );
  NOR2_X1 U11962 ( .A1(n9395), .A2(n12933), .ZN(n9396) );
  AOI211_X1 U11963 ( .C1(n14784), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n9397), .B(
        n9396), .ZN(n9398) );
  OAI211_X1 U11964 ( .C1(n9400), .C2(n14733), .A(n9399), .B(n9398), .ZN(
        P2_U3226) );
  INV_X1 U11965 ( .A(n15090), .ZN(n11132) );
  NOR3_X1 U11966 ( .A1(n11132), .A2(n15088), .A3(n12051), .ZN(n9402) );
  AOI211_X1 U11967 ( .C1(n9404), .C2(n9403), .A(n9402), .B(n9401), .ZN(n9408)
         );
  OAI22_X1 U11968 ( .A1(n12187), .A2(n15097), .B1(n7430), .B2(n12214), .ZN(
        n9405) );
  AOI21_X1 U11969 ( .B1(n12189), .B2(n15094), .A(n9405), .ZN(n9407) );
  NAND2_X1 U11970 ( .A1(n9514), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9406) );
  OAI211_X1 U11971 ( .C1(n9408), .C2(n12219), .A(n9407), .B(n9406), .ZN(
        P3_U3162) );
  NAND2_X1 U11972 ( .A1(n9409), .A2(n14805), .ZN(n9458) );
  NAND3_X1 U11973 ( .A1(n9410), .A2(n14804), .A3(n9455), .ZN(n9411) );
  NOR2_X1 U11974 ( .A1(n9458), .A2(n9411), .ZN(n9432) );
  OR2_X1 U11975 ( .A1(n12897), .A2(n14814), .ZN(n9412) );
  NAND2_X1 U11976 ( .A1(n12896), .A2(n14822), .ZN(n9414) );
  NAND2_X1 U11977 ( .A1(n10037), .A2(n7021), .ZN(n10036) );
  OR2_X1 U11978 ( .A1(n12896), .A2(n11781), .ZN(n9415) );
  INV_X1 U11979 ( .A(n12008), .ZN(n9416) );
  OR2_X1 U11980 ( .A1(n9417), .A2(n9416), .ZN(n9418) );
  NAND2_X1 U11981 ( .A1(n9417), .A2(n9416), .ZN(n9730) );
  NAND2_X1 U11982 ( .A1(n8916), .A2(n12042), .ZN(n9419) );
  NAND2_X1 U11983 ( .A1(n11957), .A2(n12003), .ZN(n11997) );
  OR2_X1 U11984 ( .A1(n11768), .A2(n9420), .ZN(n9421) );
  NAND2_X1 U11985 ( .A1(n10030), .A2(n9423), .ZN(n9424) );
  OAI21_X1 U11986 ( .B1(n9424), .B2(n12008), .A(n9725), .ZN(n9427) );
  NOR2_X1 U11987 ( .A1(n9755), .A2(n14871), .ZN(n9425) );
  AOI211_X1 U11988 ( .C1(n13251), .C2(n9427), .A(n9426), .B(n9425), .ZN(n9746)
         );
  AOI21_X1 U11989 ( .B1(n10040), .B2(n11786), .A(n13243), .ZN(n9428) );
  AND2_X1 U11990 ( .A1(n9428), .A2(n9737), .ZN(n9747) );
  AOI21_X1 U11991 ( .B1(n14879), .B2(n11786), .A(n9747), .ZN(n9429) );
  OAI211_X1 U11992 ( .C1(n9755), .C2(n14881), .A(n9746), .B(n9429), .ZN(n9433)
         );
  NAND2_X1 U11993 ( .A1(n9433), .A2(n14887), .ZN(n9430) );
  OAI21_X1 U11994 ( .B1(n14887), .B2(n8983), .A(n9430), .ZN(P2_U3439) );
  INV_X1 U11995 ( .A(n14802), .ZN(n9431) );
  NAND2_X1 U11996 ( .A1(n9433), .A2(n14908), .ZN(n9434) );
  OAI21_X1 U11997 ( .B1(n14908), .B2(n12906), .A(n9434), .ZN(P2_U3502) );
  INV_X1 U11998 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U11999 ( .A1(n10705), .A2(n14455), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10416), .ZN(n9437) );
  INV_X1 U12000 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10829) );
  INV_X1 U12001 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10817) );
  AOI21_X1 U12002 ( .B1(n10336), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9435), .ZN(
        n13779) );
  INV_X1 U12003 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14461) );
  MUX2_X1 U12004 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14461), .S(n13783), .Z(
        n13780) );
  NAND2_X1 U12005 ( .A1(n13779), .A2(n13780), .ZN(n14504) );
  NAND2_X1 U12006 ( .A1(n9443), .A2(n14461), .ZN(n14502) );
  MUX2_X1 U12007 ( .A(n10817), .B(P1_REG1_REG_12__SCAN_IN), .S(n10608), .Z(
        n14503) );
  AOI21_X1 U12008 ( .B1(n14504), .B2(n14502), .A(n14503), .ZN(n14501) );
  AOI21_X1 U12009 ( .B1(n10817), .B2(n14510), .A(n14501), .ZN(n14524) );
  MUX2_X1 U12010 ( .A(n10829), .B(P1_REG1_REG_13__SCAN_IN), .S(n14520), .Z(
        n14523) );
  NAND2_X1 U12011 ( .A1(n14524), .A2(n14523), .ZN(n14522) );
  OAI21_X1 U12012 ( .B1(n10829), .B2(n14520), .A(n14522), .ZN(n9436) );
  NOR2_X1 U12013 ( .A1(n9437), .A2(n9436), .ZN(n10415) );
  AOI21_X1 U12014 ( .B1(n9437), .B2(n9436), .A(n10415), .ZN(n9450) );
  NAND2_X1 U12015 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14382)
         );
  NAND2_X1 U12016 ( .A1(n14517), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9438) );
  OAI211_X1 U12017 ( .C1(n14553), .C2(n10416), .A(n14382), .B(n9438), .ZN(
        n9439) );
  INV_X1 U12018 ( .A(n9439), .ZN(n9449) );
  INV_X1 U12019 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9440) );
  MUX2_X1 U12020 ( .A(n9440), .B(P1_REG2_REG_14__SCAN_IN), .S(n10705), .Z(
        n9441) );
  INV_X1 U12021 ( .A(n9441), .ZN(n9447) );
  INV_X1 U12022 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9445) );
  MUX2_X1 U12023 ( .A(n9445), .B(P1_REG2_REG_13__SCAN_IN), .S(n14520), .Z(
        n14526) );
  INV_X1 U12024 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9444) );
  AOI22_X1 U12025 ( .A1(n10608), .A2(n9444), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14510), .ZN(n14508) );
  INV_X1 U12026 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10556) );
  NOR2_X1 U12027 ( .A1(n9442), .A2(n10364), .ZN(n13785) );
  MUX2_X1 U12028 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10556), .S(n13783), .Z(
        n13784) );
  OAI21_X1 U12029 ( .B1(n13786), .B2(n13785), .A(n13784), .ZN(n13788) );
  OAI21_X1 U12030 ( .B1(n9443), .B2(n10556), .A(n13788), .ZN(n14509) );
  NOR2_X1 U12031 ( .A1(n14508), .A2(n14509), .ZN(n14507) );
  AOI21_X1 U12032 ( .B1(n14510), .B2(n9444), .A(n14507), .ZN(n14527) );
  NAND2_X1 U12033 ( .A1(n14526), .A2(n14527), .ZN(n14525) );
  OAI21_X1 U12034 ( .B1(n14520), .B2(n9445), .A(n14525), .ZN(n9446) );
  NAND2_X1 U12035 ( .A1(n9447), .A2(n9446), .ZN(n10411) );
  OAI211_X1 U12036 ( .C1(n9447), .C2(n9446), .A(n14548), .B(n10411), .ZN(n9448) );
  OAI211_X1 U12037 ( .C1(n9450), .C2(n14538), .A(n9449), .B(n9448), .ZN(
        P1_U3257) );
  OAI222_X1 U12038 ( .A1(P3_U3151), .A2(n9452), .B1(n12771), .B2(n15325), .C1(
        n12770), .C2(n9451), .ZN(P3_U3275) );
  NAND2_X1 U12039 ( .A1(n12898), .A2(n9464), .ZN(n9453) );
  AND2_X1 U12040 ( .A1(n9454), .A2(n9453), .ZN(n14806) );
  INV_X1 U12041 ( .A(n14804), .ZN(n9456) );
  NAND3_X1 U12042 ( .A1(n14802), .A2(n9456), .A3(n9455), .ZN(n9457) );
  INV_X1 U12043 ( .A(n11957), .ZN(n12031) );
  OR2_X1 U12044 ( .A1(n9459), .A2(n12031), .ZN(n11757) );
  INV_X1 U12045 ( .A(n11757), .ZN(n9460) );
  NAND2_X1 U12046 ( .A1(n13228), .A2(n9460), .ZN(n9754) );
  AOI21_X1 U12047 ( .B1(n13226), .B2(n14871), .A(n14806), .ZN(n9462) );
  NOR2_X1 U12048 ( .A1(n9462), .A2(n9461), .ZN(n14807) );
  NOR2_X1 U12049 ( .A1(n9464), .A2(n9463), .ZN(n14809) );
  INV_X1 U12050 ( .A(n13232), .ZN(n13247) );
  AOI22_X1 U12051 ( .A1(n14809), .A2(n9459), .B1(n13247), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n9465) );
  AOI21_X1 U12052 ( .B1(n14807), .B2(n9465), .A(n6466), .ZN(n9466) );
  AOI21_X1 U12053 ( .B1(n6466), .B2(P2_REG2_REG_0__SCAN_IN), .A(n9466), .ZN(
        n9467) );
  OAI21_X1 U12054 ( .B1(n14806), .B2(n9754), .A(n9467), .ZN(P2_U3265) );
  XNOR2_X1 U12055 ( .A(n9626), .B(SI_18_), .ZN(n9517) );
  MUX2_X1 U12056 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n11332), .Z(n9627) );
  XNOR2_X1 U12057 ( .A(n9517), .B(n9627), .ZN(n11495) );
  INV_X1 U12058 ( .A(n11495), .ZN(n9479) );
  INV_X1 U12059 ( .A(n9470), .ZN(n9471) );
  NAND2_X1 U12060 ( .A1(n9471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9472) );
  MUX2_X1 U12061 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9472), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n9474) );
  NAND2_X1 U12062 ( .A1(n9474), .A2(n9473), .ZN(n14552) );
  OAI222_X1 U12063 ( .A1(n14223), .A2(n9475), .B1(n14221), .B2(n9479), .C1(
        P1_U3086), .C2(n14552), .ZN(P1_U3337) );
  INV_X1 U12064 ( .A(n9476), .ZN(n9477) );
  NAND2_X1 U12065 ( .A1(n9477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9478) );
  XNOR2_X1 U12066 ( .A(n9478), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12972) );
  INV_X1 U12067 ( .A(n12972), .ZN(n12958) );
  OAI222_X1 U12068 ( .A1(n13368), .A2(n9480), .B1(n13366), .B2(n9479), .C1(
        P2_U3088), .C2(n12958), .ZN(P2_U3309) );
  NAND2_X1 U12069 ( .A1(n9498), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9481) );
  INV_X1 U12070 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14942) );
  INV_X1 U12071 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9485) );
  MUX2_X1 U12072 ( .A(n9485), .B(P3_REG2_REG_6__SCAN_IN), .S(n9880), .Z(n9484)
         );
  INV_X1 U12073 ( .A(n9864), .ZN(n9483) );
  AOI21_X1 U12074 ( .B1(n6641), .B2(n9484), .A(n9483), .ZN(n9509) );
  INV_X1 U12075 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9501) );
  MUX2_X1 U12076 ( .A(n9485), .B(n9501), .S(n12369), .Z(n9872) );
  XNOR2_X1 U12077 ( .A(n9872), .B(n9880), .ZN(n9493) );
  MUX2_X1 U12078 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12369), .Z(n9487) );
  INV_X1 U12079 ( .A(n9487), .ZN(n9486) );
  NAND2_X1 U12080 ( .A1(n14940), .A2(n9486), .ZN(n9491) );
  XNOR2_X1 U12081 ( .A(n9487), .B(n14940), .ZN(n14938) );
  OR2_X1 U12082 ( .A1(n9488), .A2(n9498), .ZN(n9490) );
  NAND2_X1 U12083 ( .A1(n9490), .A2(n9489), .ZN(n14937) );
  OAI21_X1 U12084 ( .B1(n9493), .B2(n9492), .A(n9874), .ZN(n9507) );
  INV_X1 U12085 ( .A(n9880), .ZN(n9873) );
  NAND2_X1 U12086 ( .A1(n14983), .A2(n9873), .ZN(n9496) );
  INV_X1 U12087 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n9494) );
  NOR2_X1 U12088 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9494), .ZN(n10275) );
  AOI21_X1 U12089 ( .B1(n14996), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10275), .ZN(
        n9495) );
  NAND2_X1 U12090 ( .A1(n9496), .A2(n9495), .ZN(n9506) );
  NOR2_X1 U12091 ( .A1(n14940), .A2(n9499), .ZN(n9500) );
  INV_X1 U12092 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15172) );
  XNOR2_X1 U12093 ( .A(n9499), .B(n14940), .ZN(n14945) );
  NOR2_X1 U12094 ( .A1(n15172), .A2(n14945), .ZN(n14944) );
  NOR2_X1 U12095 ( .A1(n9500), .A2(n14944), .ZN(n9503) );
  MUX2_X1 U12096 ( .A(n9501), .B(P3_REG1_REG_6__SCAN_IN), .S(n9880), .Z(n9502)
         );
  NAND2_X1 U12097 ( .A1(n9503), .A2(n9502), .ZN(n9504) );
  AOI21_X1 U12098 ( .B1(n9882), .B2(n9504), .A(n14977), .ZN(n9505) );
  AOI211_X1 U12099 ( .C1(n15007), .C2(n9507), .A(n9506), .B(n9505), .ZN(n9508)
         );
  OAI21_X1 U12100 ( .B1(n9509), .B2(n14990), .A(n9508), .ZN(P3_U3188) );
  XOR2_X1 U12101 ( .A(n9511), .B(n9510), .Z(n9516) );
  OAI21_X1 U12102 ( .B1(n7018), .B2(n12213), .A(n9512), .ZN(n9513) );
  AOI21_X1 U12103 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n9514), .A(n9513), .ZN(
        n9515) );
  OAI21_X1 U12104 ( .B1(n9516), .B2(n12219), .A(n9515), .ZN(P3_U3177) );
  INV_X1 U12105 ( .A(n9517), .ZN(n9518) );
  NAND2_X1 U12106 ( .A1(n9518), .A2(n9627), .ZN(n9520) );
  NAND2_X1 U12107 ( .A1(n9626), .A2(SI_18_), .ZN(n9519) );
  NAND2_X1 U12108 ( .A1(n9520), .A2(n9519), .ZN(n9524) );
  MUX2_X1 U12109 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n11332), .Z(n9521) );
  NAND2_X1 U12110 ( .A1(n9521), .A2(SI_19_), .ZN(n9630) );
  INV_X1 U12111 ( .A(n9521), .ZN(n9522) );
  NAND2_X1 U12112 ( .A1(n9522), .A2(n15267), .ZN(n9628) );
  NAND2_X1 U12113 ( .A1(n9630), .A2(n9628), .ZN(n9523) );
  INV_X1 U12114 ( .A(n11505), .ZN(n9526) );
  OAI222_X1 U12115 ( .A1(n13368), .A2(n9525), .B1(n13366), .B2(n9526), .C1(
        n8963), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U12116 ( .A1(n14223), .A2(n9527), .B1(n14221), .B2(n9526), .C1(
        P1_U3086), .C2(n14614), .ZN(P1_U3336) );
  AOI22_X1 U12117 ( .A1(n11507), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11506), 
        .B2(n9528), .ZN(n9529) );
  NAND2_X1 U12118 ( .A1(n9530), .A2(n9529), .ZN(n11812) );
  NAND2_X1 U12119 ( .A1(n8982), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9537) );
  OR2_X1 U12120 ( .A1(n6950), .A2(n9531), .ZN(n9536) );
  NAND2_X1 U12121 ( .A1(n9540), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9647) );
  OAI21_X1 U12122 ( .B1(n9540), .B2(P2_REG3_REG_7__SCAN_IN), .A(n9647), .ZN(
        n9948) );
  OR2_X1 U12123 ( .A1(n11741), .A2(n9948), .ZN(n9535) );
  INV_X1 U12124 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9533) );
  OR2_X1 U12125 ( .A1(n11743), .A2(n9533), .ZN(n9534) );
  NAND4_X1 U12126 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), .ZN(n12891) );
  NAND2_X1 U12127 ( .A1(n12891), .A2(n12858), .ZN(n9539) );
  NAND2_X1 U12128 ( .A1(n12893), .A2(n13020), .ZN(n9538) );
  AND2_X1 U12129 ( .A1(n9539), .A2(n9538), .ZN(n9927) );
  INV_X1 U12130 ( .A(n9540), .ZN(n9544) );
  INV_X1 U12131 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U12132 ( .A1(n9542), .A2(n9541), .ZN(n9543) );
  NAND2_X1 U12133 ( .A1(n9544), .A2(n9543), .ZN(n9931) );
  INV_X1 U12134 ( .A(n9931), .ZN(n9545) );
  NAND2_X1 U12135 ( .A1(n12861), .A2(n9545), .ZN(n9547) );
  OAI211_X1 U12136 ( .C1(n12859), .C2(n9927), .A(n9547), .B(n9546), .ZN(n9567)
         );
  XNOR2_X1 U12137 ( .A(n11812), .B(n11736), .ZN(n9706) );
  NAND2_X1 U12138 ( .A1(n8906), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9552) );
  OR2_X1 U12139 ( .A1(n11962), .A2(n8698), .ZN(n9551) );
  OR2_X1 U12140 ( .A1(n11741), .A2(n9931), .ZN(n9550) );
  INV_X1 U12141 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9548) );
  OR2_X1 U12142 ( .A1(n11743), .A2(n9548), .ZN(n9549) );
  AND2_X1 U12143 ( .A1(n12892), .A2(n9668), .ZN(n9553) );
  NAND2_X1 U12144 ( .A1(n9706), .A2(n9553), .ZN(n9634) );
  OAI21_X1 U12145 ( .B1(n9706), .B2(n9553), .A(n9634), .ZN(n9565) );
  INV_X1 U12146 ( .A(n9554), .ZN(n9555) );
  NOR2_X1 U12147 ( .A1(n9555), .A2(n12825), .ZN(n9559) );
  AOI22_X1 U12148 ( .A1(n11507), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11506), 
        .B2(n9556), .ZN(n9558) );
  NAND2_X1 U12149 ( .A1(n9558), .A2(n9557), .ZN(n12824) );
  XNOR2_X1 U12150 ( .A(n12824), .B(n11736), .ZN(n9562) );
  NAND2_X1 U12151 ( .A1(n12893), .A2(n9668), .ZN(n9561) );
  XNOR2_X1 U12152 ( .A(n9562), .B(n9561), .ZN(n12829) );
  INV_X1 U12153 ( .A(n9561), .ZN(n9563) );
  AOI211_X1 U12154 ( .C1(n9565), .C2(n9564), .A(n12877), .B(n6508), .ZN(n9566)
         );
  AOI211_X1 U12155 ( .C1(n11812), .C2(n12875), .A(n9567), .B(n9566), .ZN(n9568) );
  INV_X1 U12156 ( .A(n9568), .ZN(P2_U3211) );
  INV_X1 U12157 ( .A(n9569), .ZN(n9570) );
  NAND2_X1 U12158 ( .A1(n9571), .A2(n9570), .ZN(n9572) );
  NAND2_X1 U12159 ( .A1(n13730), .A2(n11459), .ZN(n9578) );
  INV_X2 U12160 ( .A(n13653), .ZN(n11284) );
  AOI22_X1 U12161 ( .A1(n11284), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n11283), 
        .B2(n13747), .ZN(n9576) );
  NAND2_X1 U12162 ( .A1(n9574), .A2(n6468), .ZN(n9575) );
  NAND2_X1 U12163 ( .A1(n11422), .A2(n14602), .ZN(n9577) );
  NAND2_X1 U12164 ( .A1(n9578), .A2(n9577), .ZN(n9579) );
  XNOR2_X1 U12165 ( .A(n9579), .B(n11477), .ZN(n9583) );
  NAND2_X1 U12166 ( .A1(n11367), .A2(n13730), .ZN(n9581) );
  NAND2_X1 U12167 ( .A1(n11459), .A2(n14602), .ZN(n9580) );
  NAND2_X1 U12168 ( .A1(n9581), .A2(n9580), .ZN(n9582) );
  XNOR2_X1 U12169 ( .A(n9583), .B(n9582), .ZN(n13387) );
  NAND2_X1 U12170 ( .A1(n9583), .A2(n9582), .ZN(n9584) );
  NAND2_X1 U12171 ( .A1(n11632), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9593) );
  OR2_X1 U12172 ( .A1(n13638), .A2(n8806), .ZN(n9592) );
  INV_X1 U12173 ( .A(n9609), .ZN(n9611) );
  INV_X1 U12174 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9587) );
  INV_X1 U12175 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9586) );
  NAND2_X1 U12176 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  NAND2_X1 U12177 ( .A1(n9611), .A2(n9588), .ZN(n10022) );
  OR2_X1 U12178 ( .A1(n9585), .A2(n10022), .ZN(n9591) );
  OR2_X1 U12179 ( .A1(n9589), .A2(n14719), .ZN(n9590) );
  NAND4_X1 U12180 ( .A1(n9593), .A2(n9592), .A3(n9591), .A4(n9590), .ZN(n13729) );
  NAND2_X1 U12181 ( .A1(n11367), .A2(n13729), .ZN(n9600) );
  NAND2_X1 U12182 ( .A1(n6468), .A2(n9594), .ZN(n9597) );
  OR2_X1 U12183 ( .A1(n13653), .A2(n9595), .ZN(n9596) );
  OAI211_X1 U12184 ( .C1(n11335), .C2(n9598), .A(n9597), .B(n9596), .ZN(n14662) );
  NAND2_X1 U12185 ( .A1(n11459), .A2(n14662), .ZN(n9599) );
  AND2_X1 U12186 ( .A1(n9600), .A2(n9599), .ZN(n9784) );
  NAND2_X1 U12187 ( .A1(n13729), .A2(n11459), .ZN(n9602) );
  NAND2_X1 U12188 ( .A1(n11422), .A2(n14662), .ZN(n9601) );
  NAND2_X1 U12189 ( .A1(n9602), .A2(n9601), .ZN(n9603) );
  XNOR2_X1 U12190 ( .A(n9603), .B(n11477), .ZN(n9782) );
  XNOR2_X1 U12191 ( .A(n9783), .B(n9782), .ZN(n9623) );
  INV_X1 U12192 ( .A(n9604), .ZN(n9605) );
  NAND2_X1 U12193 ( .A1(n9606), .A2(n9605), .ZN(n9607) );
  NOR2_X1 U12194 ( .A1(n14436), .A2(n10022), .ZN(n9621) );
  NAND2_X1 U12195 ( .A1(n11483), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9616) );
  INV_X1 U12196 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9608) );
  OR2_X1 U12197 ( .A1(n13639), .A2(n9608), .ZN(n9615) );
  INV_X1 U12198 ( .A(n9790), .ZN(n9792) );
  INV_X1 U12199 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9610) );
  NAND2_X1 U12200 ( .A1(n9611), .A2(n9610), .ZN(n9612) );
  NAND2_X1 U12201 ( .A1(n9792), .A2(n9612), .ZN(n10090) );
  OR2_X1 U12202 ( .A1(n9585), .A2(n10090), .ZN(n9614) );
  OR2_X1 U12203 ( .A1(n6463), .A2(n14721), .ZN(n9613) );
  NAND2_X1 U12204 ( .A1(n13728), .A2(n14635), .ZN(n9618) );
  NAND2_X1 U12205 ( .A1(n13730), .A2(n14683), .ZN(n9617) );
  AND2_X1 U12206 ( .A1(n9618), .A2(n9617), .ZN(n14665) );
  OAI21_X1 U12207 ( .B1(n13462), .B2(n14665), .A(n9619), .ZN(n9620) );
  AOI211_X1 U12208 ( .C1(n14662), .C2(n14415), .A(n9621), .B(n9620), .ZN(n9622) );
  OAI21_X1 U12209 ( .B1(n9623), .B2(n14410), .A(n9622), .ZN(P1_U3230) );
  INV_X1 U12210 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11302) );
  INV_X1 U12211 ( .A(n9627), .ZN(n9624) );
  OAI21_X1 U12212 ( .B1(n15344), .B2(n9624), .A(n9630), .ZN(n9625) );
  NOR2_X1 U12213 ( .A1(n9627), .A2(SI_18_), .ZN(n9631) );
  INV_X1 U12214 ( .A(n9628), .ZN(n9629) );
  INV_X1 U12215 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11519) );
  MUX2_X1 U12216 ( .A(n11302), .B(n11519), .S(n11332), .Z(n9714) );
  XNOR2_X1 U12217 ( .A(n9716), .B(n9714), .ZN(n11518) );
  INV_X1 U12218 ( .A(n11518), .ZN(n9684) );
  OAI222_X1 U12219 ( .A1(n14223), .A2(n11302), .B1(n14221), .B2(n9684), .C1(
        n13656), .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U12220 ( .A1(P3_U3151), .A2(n10965), .B1(n12771), .B2(n15361), 
        .C1(n12770), .C2(n9633), .ZN(P3_U3274) );
  INV_X1 U12221 ( .A(n9634), .ZN(n9642) );
  AOI22_X1 U12222 ( .A1(n11507), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11506), 
        .B2(n9635), .ZN(n9636) );
  NAND2_X1 U12223 ( .A1(n9637), .A2(n9636), .ZN(n11820) );
  XNOR2_X1 U12224 ( .A(n11820), .B(n11736), .ZN(n9638) );
  AND2_X1 U12225 ( .A1(n12891), .A2(n9668), .ZN(n9639) );
  NAND2_X1 U12226 ( .A1(n9638), .A2(n9639), .ZN(n9654) );
  INV_X1 U12227 ( .A(n9638), .ZN(n9756) );
  INV_X1 U12228 ( .A(n9639), .ZN(n9640) );
  NAND2_X1 U12229 ( .A1(n9756), .A2(n9640), .ZN(n9641) );
  AND2_X1 U12230 ( .A1(n9654), .A2(n9641), .ZN(n9707) );
  AOI22_X1 U12231 ( .A1(n11507), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9643), 
        .B2(n11506), .ZN(n9644) );
  XNOR2_X1 U12232 ( .A(n11826), .B(n11736), .ZN(n9678) );
  NAND2_X1 U12233 ( .A1(n8982), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9653) );
  OR2_X1 U12234 ( .A1(n6950), .A2(n14899), .ZN(n9652) );
  AND2_X1 U12235 ( .A1(n9647), .A2(n9646), .ZN(n9648) );
  OR2_X1 U12236 ( .A1(n9648), .A2(n9662), .ZN(n10057) );
  OR2_X1 U12237 ( .A1(n11741), .A2(n10057), .ZN(n9651) );
  INV_X1 U12238 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9649) );
  OR2_X1 U12239 ( .A1(n11743), .A2(n9649), .ZN(n9650) );
  NAND4_X1 U12240 ( .A1(n9653), .A2(n9652), .A3(n9651), .A4(n9650), .ZN(n12890) );
  NAND2_X1 U12241 ( .A1(n12890), .A2(n9668), .ZN(n9656) );
  XNOR2_X1 U12242 ( .A(n9678), .B(n9656), .ZN(n9767) );
  AND2_X1 U12243 ( .A1(n9767), .A2(n9654), .ZN(n9655) );
  NAND2_X1 U12244 ( .A1(n9708), .A2(n9655), .ZN(n9763) );
  INV_X1 U12245 ( .A(n9656), .ZN(n9657) );
  AOI22_X1 U12246 ( .A1(n11507), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n11506), 
        .B2(n12926), .ZN(n9659) );
  XNOR2_X1 U12247 ( .A(n14860), .B(n11736), .ZN(n10169) );
  NAND2_X1 U12248 ( .A1(n11958), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9667) );
  INV_X1 U12249 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9661) );
  OR2_X1 U12250 ( .A1(n11743), .A2(n9661), .ZN(n9666) );
  NAND2_X1 U12251 ( .A1(n9662), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10184) );
  OR2_X1 U12252 ( .A1(n9662), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U12253 ( .A1(n10184), .A2(n9663), .ZN(n9961) );
  OR2_X1 U12254 ( .A1(n11741), .A2(n9961), .ZN(n9665) );
  OR2_X1 U12255 ( .A1(n11962), .A2(n9028), .ZN(n9664) );
  NAND4_X1 U12256 ( .A1(n9667), .A2(n9666), .A3(n9665), .A4(n9664), .ZN(n12889) );
  NAND2_X1 U12257 ( .A1(n12889), .A2(n9668), .ZN(n10167) );
  XNOR2_X1 U12258 ( .A(n10169), .B(n10167), .ZN(n9677) );
  NAND2_X1 U12259 ( .A1(n8982), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9673) );
  OR2_X1 U12260 ( .A1(n6950), .A2(n14903), .ZN(n9672) );
  INV_X1 U12261 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10182) );
  XNOR2_X1 U12262 ( .A(n10184), .B(n10182), .ZN(n10289) );
  OR2_X1 U12263 ( .A1(n11741), .A2(n10289), .ZN(n9671) );
  INV_X1 U12264 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9669) );
  OR2_X1 U12265 ( .A1(n11743), .A2(n9669), .ZN(n9670) );
  NAND4_X1 U12266 ( .A1(n9673), .A2(n9672), .A3(n9671), .A4(n9670), .ZN(n12888) );
  AOI22_X1 U12267 ( .A1(n13020), .A2(n12890), .B1(n12888), .B2(n12858), .ZN(
        n9959) );
  INV_X1 U12268 ( .A(n9959), .ZN(n9674) );
  AOI22_X1 U12269 ( .A1(n12871), .A2(n9674), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3088), .ZN(n9675) );
  OAI21_X1 U12270 ( .B1(n9961), .B2(n12873), .A(n9675), .ZN(n9676) );
  AOI21_X1 U12271 ( .B1(n14860), .B2(n12875), .A(n9676), .ZN(n9683) );
  INV_X1 U12272 ( .A(n9677), .ZN(n9681) );
  INV_X1 U12273 ( .A(n9678), .ZN(n9679) );
  OAI22_X1 U12274 ( .A1(n12828), .A2(n9958), .B1(n9679), .B2(n12877), .ZN(
        n9680) );
  NAND3_X1 U12275 ( .A1(n9763), .A2(n9681), .A3(n9680), .ZN(n9682) );
  OAI211_X1 U12276 ( .C1(n10171), .C2(n12877), .A(n9683), .B(n9682), .ZN(
        P2_U3203) );
  OAI222_X1 U12277 ( .A1(n13368), .A2(n11519), .B1(P2_U3088), .B2(n9685), .C1(
        n13366), .C2(n9684), .ZN(P2_U3307) );
  INV_X2 U12278 ( .A(n15053), .ZN(n15102) );
  INV_X1 U12279 ( .A(n15096), .ZN(n15045) );
  NOR3_X1 U12280 ( .A1(n11127), .A2(n9687), .A3(n15151), .ZN(n9688) );
  AOI21_X1 U12281 ( .B1(n15045), .B2(n12234), .A(n9688), .ZN(n12706) );
  INV_X1 U12282 ( .A(n12706), .ZN(n9689) );
  AOI21_X1 U12283 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15102), .A(n9689), .ZN(
        n9702) );
  NAND2_X1 U12284 ( .A1(n9691), .A2(n10861), .ZN(n9692) );
  OAI21_X1 U12285 ( .B1(n10860), .B2(n10861), .A(n9692), .ZN(n9698) );
  NOR2_X1 U12286 ( .A1(n9694), .A2(n9693), .ZN(n9696) );
  INV_X1 U12287 ( .A(n10857), .ZN(n9697) );
  NAND3_X1 U12288 ( .A1(n9698), .A2(n10864), .A3(n9697), .ZN(n9699) );
  OR2_X1 U12289 ( .A1(n9699), .A2(n11121), .ZN(n10082) );
  AOI22_X1 U12290 ( .A1(n12627), .A2(n9700), .B1(n15068), .B2(
        P3_REG2_REG_0__SCAN_IN), .ZN(n9701) );
  OAI21_X1 U12291 ( .B1(n9702), .B2(n15068), .A(n9701), .ZN(P3_U3233) );
  AOI22_X1 U12292 ( .A1(n12858), .A2(n12890), .B1(n12892), .B2(n13020), .ZN(
        n9942) );
  INV_X1 U12293 ( .A(n9948), .ZN(n9703) );
  NAND2_X1 U12294 ( .A1(n12861), .A2(n9703), .ZN(n9705) );
  OAI211_X1 U12295 ( .C1(n12859), .C2(n9942), .A(n9705), .B(n9704), .ZN(n9712)
         );
  NAND3_X1 U12296 ( .A1(n11651), .A2(n9706), .A3(n12892), .ZN(n9710) );
  OAI21_X1 U12297 ( .B1(n6508), .B2(n9707), .A(n12808), .ZN(n9709) );
  INV_X1 U12298 ( .A(n9708), .ZN(n9758) );
  AOI21_X1 U12299 ( .B1(n9710), .B2(n9709), .A(n9758), .ZN(n9711) );
  AOI211_X1 U12300 ( .C1(n11820), .C2(n12875), .A(n9712), .B(n9711), .ZN(n9713) );
  INV_X1 U12301 ( .A(n9713), .ZN(P2_U3185) );
  INV_X1 U12302 ( .A(n9714), .ZN(n9715) );
  MUX2_X1 U12303 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n11332), .Z(n10104) );
  XNOR2_X1 U12304 ( .A(n10104), .B(SI_21_), .ZN(n10101) );
  XNOR2_X1 U12305 ( .A(n10103), .B(n10101), .ZN(n11529) );
  INV_X1 U12306 ( .A(n11529), .ZN(n9720) );
  INV_X1 U12307 ( .A(n13645), .ZN(n13665) );
  OAI222_X1 U12308 ( .A1(n14223), .A2(n11316), .B1(n14221), .B2(n9720), .C1(
        P1_U3086), .C2(n13665), .ZN(P1_U3334) );
  OAI222_X1 U12309 ( .A1(n13368), .A2(n11530), .B1(n13366), .B2(n9720), .C1(
        n12031), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U12310 ( .A(n9721), .ZN(n9723) );
  OAI22_X1 U12311 ( .A1(n11160), .A2(P3_U3151), .B1(SI_22_), .B2(n12771), .ZN(
        n9722) );
  AOI21_X1 U12312 ( .B1(n9723), .B2(n12764), .A(n9722), .ZN(P3_U3273) );
  OR2_X1 U12313 ( .A1(n12895), .A2(n11790), .ZN(n9724) );
  INV_X1 U12314 ( .A(n11801), .ZN(n14829) );
  NAND3_X1 U12315 ( .A1(n9725), .A2(n12006), .A3(n9724), .ZN(n9726) );
  NAND2_X1 U12316 ( .A1(n9812), .A2(n9726), .ZN(n9728) );
  AOI21_X1 U12317 ( .B1(n9728), .B2(n13251), .A(n9727), .ZN(n9734) );
  OR2_X1 U12318 ( .A1(n12895), .A2(n11786), .ZN(n9729) );
  OR2_X1 U12319 ( .A1(n9731), .A2(n12006), .ZN(n9732) );
  NAND2_X1 U12320 ( .A1(n9805), .A2(n9732), .ZN(n14832) );
  INV_X1 U12321 ( .A(n14871), .ZN(n14885) );
  NAND2_X1 U12322 ( .A1(n14832), .A2(n14885), .ZN(n9733) );
  NAND2_X1 U12323 ( .A1(n9734), .A2(n9733), .ZN(n14830) );
  MUX2_X1 U12324 ( .A(n14830), .B(P2_REG2_REG_4__SCAN_IN), .S(n6466), .Z(n9735) );
  INV_X1 U12325 ( .A(n9735), .ZN(n9745) );
  INV_X1 U12326 ( .A(n9754), .ZN(n10046) );
  NAND2_X1 U12327 ( .A1(n9737), .A2(n11801), .ZN(n9738) );
  NAND2_X1 U12328 ( .A1(n9738), .A2(n13332), .ZN(n9739) );
  NOR2_X1 U12329 ( .A1(n9809), .A2(n9739), .ZN(n14827) );
  NAND2_X1 U12330 ( .A1(n13245), .A2(n14827), .ZN(n9742) );
  NAND2_X1 U12331 ( .A1(n13247), .A2(n9740), .ZN(n9741) );
  OAI211_X1 U12332 ( .C1(n14829), .C2(n13231), .A(n9742), .B(n9741), .ZN(n9743) );
  AOI21_X1 U12333 ( .B1(n14832), .B2(n10046), .A(n9743), .ZN(n9744) );
  NAND2_X1 U12334 ( .A1(n9745), .A2(n9744), .ZN(P2_U3261) );
  MUX2_X1 U12335 ( .A(n8653), .B(n9746), .S(n13228), .Z(n9753) );
  NAND2_X1 U12336 ( .A1(n13245), .A2(n9747), .ZN(n9750) );
  NAND2_X1 U12337 ( .A1(n13247), .A2(n9748), .ZN(n9749) );
  OAI211_X1 U12338 ( .C1(n11790), .C2(n13231), .A(n9750), .B(n9749), .ZN(n9751) );
  INV_X1 U12339 ( .A(n9751), .ZN(n9752) );
  OAI211_X1 U12340 ( .C1(n9755), .C2(n9754), .A(n9753), .B(n9752), .ZN(
        P2_U3262) );
  INV_X1 U12341 ( .A(n12891), .ZN(n11822) );
  NOR3_X1 U12342 ( .A1(n12828), .A2(n9756), .A3(n11822), .ZN(n9757) );
  AOI21_X1 U12343 ( .B1(n9758), .B2(n12808), .A(n9757), .ZN(n9768) );
  NAND2_X1 U12344 ( .A1(n12889), .A2(n12858), .ZN(n9760) );
  NAND2_X1 U12345 ( .A1(n12891), .A2(n13020), .ZN(n9759) );
  NAND2_X1 U12346 ( .A1(n9760), .A2(n9759), .ZN(n10050) );
  NAND2_X1 U12347 ( .A1(n12871), .A2(n10050), .ZN(n9762) );
  OAI211_X1 U12348 ( .C1(n12873), .C2(n10057), .A(n9762), .B(n9761), .ZN(n9765) );
  NOR2_X1 U12349 ( .A1(n9763), .A2(n12877), .ZN(n9764) );
  AOI211_X1 U12350 ( .C1(n11826), .C2(n12875), .A(n9765), .B(n9764), .ZN(n9766) );
  OAI21_X1 U12351 ( .B1(n9768), .B2(n9767), .A(n9766), .ZN(P2_U3193) );
  NAND2_X1 U12352 ( .A1(n13728), .A2(n11459), .ZN(n9774) );
  NAND2_X1 U12353 ( .A1(n9769), .A2(n6468), .ZN(n9772) );
  OR2_X1 U12354 ( .A1(n13653), .A2(n9770), .ZN(n9771) );
  OAI211_X1 U12355 ( .C1(n11335), .C2(n13769), .A(n9772), .B(n9771), .ZN(
        n13511) );
  NAND2_X1 U12356 ( .A1(n11422), .A2(n13511), .ZN(n9773) );
  NAND2_X1 U12357 ( .A1(n9774), .A2(n9773), .ZN(n9775) );
  XNOR2_X1 U12358 ( .A(n9775), .B(n11410), .ZN(n9778) );
  NAND2_X1 U12359 ( .A1(n11367), .A2(n13728), .ZN(n9777) );
  NAND2_X1 U12360 ( .A1(n11459), .A2(n13511), .ZN(n9776) );
  AND2_X1 U12361 ( .A1(n9777), .A2(n9776), .ZN(n9779) );
  NAND2_X1 U12362 ( .A1(n9778), .A2(n9779), .ZN(n9901) );
  INV_X1 U12363 ( .A(n9778), .ZN(n9781) );
  INV_X1 U12364 ( .A(n9779), .ZN(n9780) );
  NAND2_X1 U12365 ( .A1(n9781), .A2(n9780), .ZN(n9903) );
  NAND2_X1 U12366 ( .A1(n9901), .A2(n9903), .ZN(n9789) );
  INV_X1 U12367 ( .A(n9784), .ZN(n9785) );
  NAND2_X1 U12368 ( .A1(n9786), .A2(n9785), .ZN(n9787) );
  XOR2_X1 U12369 ( .A(n9789), .B(n9902), .Z(n9803) );
  NAND2_X1 U12370 ( .A1(n11632), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9798) );
  OR2_X1 U12371 ( .A1(n9589), .A2(n10146), .ZN(n9797) );
  INV_X1 U12372 ( .A(n9848), .ZN(n9794) );
  INV_X1 U12373 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U12374 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  NAND2_X1 U12375 ( .A1(n9794), .A2(n9793), .ZN(n9911) );
  OR2_X1 U12376 ( .A1(n9585), .A2(n9911), .ZN(n9796) );
  OR2_X1 U12377 ( .A1(n13638), .A2(n9858), .ZN(n9795) );
  NAND4_X1 U12378 ( .A1(n9798), .A2(n9797), .A3(n9796), .A4(n9795), .ZN(n13727) );
  AOI22_X1 U12379 ( .A1(n9799), .A2(n13727), .B1(n13442), .B2(n13729), .ZN(
        n9802) );
  NAND2_X1 U12380 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13761) );
  OAI21_X1 U12381 ( .B1(n14436), .B2(n10090), .A(n13761), .ZN(n9800) );
  AOI21_X1 U12382 ( .B1(n13511), .B2(n14415), .A(n9800), .ZN(n9801) );
  OAI211_X1 U12383 ( .C1(n9803), .C2(n14410), .A(n9802), .B(n9801), .ZN(
        P1_U3227) );
  OR2_X1 U12384 ( .A1(n12894), .A2(n11801), .ZN(n9804) );
  OR2_X1 U12385 ( .A1(n12893), .A2(n14836), .ZN(n9924) );
  NAND2_X1 U12386 ( .A1(n12893), .A2(n14836), .ZN(n9806) );
  XNOR2_X1 U12387 ( .A(n9919), .B(n12005), .ZN(n14838) );
  NAND2_X1 U12388 ( .A1(n11757), .A2(n14871), .ZN(n9807) );
  INV_X1 U12389 ( .A(n9930), .ZN(n9808) );
  OAI211_X1 U12390 ( .C1(n14836), .C2(n9809), .A(n9808), .B(n13332), .ZN(
        n14834) );
  NOR2_X1 U12391 ( .A1(n13159), .A2(n14834), .ZN(n9811) );
  OAI22_X1 U12392 ( .A1(n13231), .A2(n14836), .B1(n13232), .B2(n12822), .ZN(
        n9810) );
  AOI211_X1 U12393 ( .C1(n14838), .C2(n13246), .A(n9811), .B(n9810), .ZN(n9821) );
  OR2_X1 U12394 ( .A1(n12894), .A2(n14829), .ZN(n9814) );
  INV_X1 U12395 ( .A(n12005), .ZN(n9813) );
  NAND3_X1 U12396 ( .A1(n9812), .A2(n12005), .A3(n9814), .ZN(n9815) );
  NAND2_X1 U12397 ( .A1(n9923), .A2(n9815), .ZN(n9818) );
  NAND2_X1 U12398 ( .A1(n12892), .A2(n12858), .ZN(n9817) );
  NAND2_X1 U12399 ( .A1(n12894), .A2(n13020), .ZN(n9816) );
  NAND2_X1 U12400 ( .A1(n9817), .A2(n9816), .ZN(n12821) );
  AOI21_X1 U12401 ( .B1(n9818), .B2(n13251), .A(n12821), .ZN(n14835) );
  MUX2_X1 U12402 ( .A(n9819), .B(n14835), .S(n13228), .Z(n9820) );
  NAND2_X1 U12403 ( .A1(n9821), .A2(n9820), .ZN(P2_U3260) );
  NAND2_X1 U12404 ( .A1(n9822), .A2(n6468), .ZN(n9825) );
  AOI22_X1 U12405 ( .A1(n11284), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11283), 
        .B2(n9823), .ZN(n9824) );
  NAND2_X1 U12406 ( .A1(n9825), .A2(n9824), .ZN(n13515) );
  XNOR2_X1 U12407 ( .A(n13727), .B(n10147), .ZN(n13676) );
  NAND2_X1 U12408 ( .A1(n13731), .A2(n10110), .ZN(n13493) );
  AND2_X1 U12409 ( .A1(n13494), .A2(n13493), .ZN(n13675) );
  AND2_X1 U12410 ( .A1(n13732), .A2(n14632), .ZN(n10108) );
  INV_X1 U12411 ( .A(n13496), .ZN(n13678) );
  NAND2_X1 U12412 ( .A1(n10122), .A2(n13678), .ZN(n9827) );
  OR2_X1 U12413 ( .A1(n14636), .A2(n13498), .ZN(n9826) );
  NAND2_X1 U12414 ( .A1(n9827), .A2(n9826), .ZN(n14592) );
  XNOR2_X1 U12415 ( .A(n13730), .B(n14602), .ZN(n13502) );
  NAND2_X1 U12416 ( .A1(n14592), .A2(n14593), .ZN(n9829) );
  OR2_X1 U12417 ( .A1(n13730), .A2(n14602), .ZN(n9828) );
  NAND2_X1 U12418 ( .A1(n9829), .A2(n9828), .ZN(n10020) );
  XNOR2_X1 U12419 ( .A(n13729), .B(n14662), .ZN(n13673) );
  INV_X1 U12420 ( .A(n13673), .ZN(n10019) );
  NAND2_X1 U12421 ( .A1(n10020), .A2(n10019), .ZN(n9831) );
  OR2_X1 U12422 ( .A1(n13729), .A2(n14662), .ZN(n9830) );
  XNOR2_X1 U12423 ( .A(n13728), .B(n13511), .ZN(n13674) );
  OR2_X1 U12424 ( .A1(n13728), .A2(n13511), .ZN(n9832) );
  XOR2_X1 U12425 ( .A(n13676), .B(n9969), .Z(n10134) );
  INV_X1 U12426 ( .A(n13711), .ZN(n9836) );
  INV_X1 U12427 ( .A(n9833), .ZN(n9835) );
  OR2_X1 U12428 ( .A1(n14614), .A2(n9838), .ZN(n13660) );
  NOR2_X1 U12429 ( .A1(n14016), .A2(n13660), .ZN(n14610) );
  INV_X1 U12430 ( .A(n14610), .ZN(n13910) );
  OAI21_X1 U12431 ( .B1(n13490), .B2(n9838), .A(n11477), .ZN(n9839) );
  OR2_X2 U12432 ( .A1(n13732), .A2(n14618), .ZN(n13672) );
  NAND2_X1 U12433 ( .A1(n13494), .A2(n13672), .ZN(n9840) );
  NAND2_X1 U12434 ( .A1(n10128), .A2(n13496), .ZN(n9842) );
  OR2_X1 U12435 ( .A1(n14636), .A2(n14649), .ZN(n9841) );
  NAND2_X1 U12436 ( .A1(n14594), .A2(n13502), .ZN(n9844) );
  INV_X1 U12437 ( .A(n14602), .ZN(n14655) );
  OR2_X1 U12438 ( .A1(n13730), .A2(n14655), .ZN(n9843) );
  NAND2_X1 U12439 ( .A1(n9844), .A2(n9843), .ZN(n10018) );
  INV_X1 U12440 ( .A(n14662), .ZN(n10021) );
  OR2_X1 U12441 ( .A1(n13729), .A2(n10021), .ZN(n9845) );
  INV_X1 U12442 ( .A(n13511), .ZN(n14671) );
  XOR2_X1 U12443 ( .A(n9997), .B(n13676), .Z(n9855) );
  NAND2_X1 U12444 ( .A1(n13489), .A2(n14225), .ZN(n9846) );
  NAND2_X1 U12445 ( .A1(n13645), .A2(n13664), .ZN(n13647) );
  NAND2_X1 U12446 ( .A1(n11632), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9853) );
  OR2_X1 U12447 ( .A1(n13638), .A2(n9847), .ZN(n9852) );
  NAND2_X1 U12448 ( .A1(n9848), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9982) );
  OAI21_X1 U12449 ( .B1(n9848), .B2(P1_REG3_REG_7__SCAN_IN), .A(n9982), .ZN(
        n14583) );
  OR2_X1 U12450 ( .A1(n9585), .A2(n14583), .ZN(n9851) );
  OR2_X1 U12451 ( .A1(n9589), .A2(n9849), .ZN(n9850) );
  NAND4_X1 U12452 ( .A1(n9853), .A2(n9852), .A3(n9851), .A4(n9850), .ZN(n14682) );
  INV_X1 U12453 ( .A(n14682), .ZN(n10390) );
  INV_X1 U12454 ( .A(n13728), .ZN(n9912) );
  OAI22_X1 U12455 ( .A1(n10390), .A2(n14615), .B1(n9912), .B2(n14704), .ZN(
        n9854) );
  AOI21_X1 U12456 ( .B1(n9855), .B2(n14699), .A(n9854), .ZN(n9856) );
  OAI21_X1 U12457 ( .B1(n10134), .B2(n14647), .A(n9856), .ZN(n10136) );
  NAND2_X1 U12458 ( .A1(n10136), .A2(n6464), .ZN(n9862) );
  NAND2_X1 U12459 ( .A1(n10110), .A2(n14618), .ZN(n10124) );
  AOI211_X1 U12460 ( .C1(n13515), .C2(n10089), .A(n13980), .B(n14588), .ZN(
        n10137) );
  INV_X1 U12461 ( .A(n9857), .ZN(n14613) );
  NOR2_X1 U12462 ( .A1(n13982), .A2(n10147), .ZN(n9860) );
  OAI22_X1 U12463 ( .A1(n6464), .A2(n9858), .B1(n9911), .B2(n14599), .ZN(n9859) );
  AOI211_X1 U12464 ( .C1(n10137), .C2(n14609), .A(n9860), .B(n9859), .ZN(n9861) );
  OAI211_X1 U12465 ( .C1(n10134), .C2(n13910), .A(n9862), .B(n9861), .ZN(
        P1_U3287) );
  NAND2_X1 U12466 ( .A1(n9880), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9863) );
  NOR2_X1 U12467 ( .A1(n14956), .A2(n9865), .ZN(n9866) );
  INV_X1 U12468 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n14961) );
  XNOR2_X1 U12469 ( .A(n14956), .B(n9865), .ZN(n14960) );
  INV_X1 U12470 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10434) );
  MUX2_X1 U12471 ( .A(n10434), .B(P3_REG2_REG_8__SCAN_IN), .S(n10234), .Z(
        n9868) );
  INV_X1 U12472 ( .A(n10223), .ZN(n9867) );
  AOI21_X1 U12473 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9892) );
  INV_X1 U12474 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9884) );
  MUX2_X1 U12475 ( .A(n10434), .B(n9884), .S(n12369), .Z(n10227) );
  XNOR2_X1 U12476 ( .A(n10227), .B(n10234), .ZN(n9878) );
  MUX2_X1 U12477 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12369), .Z(n9871) );
  INV_X1 U12478 ( .A(n9871), .ZN(n9870) );
  NAND2_X1 U12479 ( .A1(n14956), .A2(n9870), .ZN(n9876) );
  XNOR2_X1 U12480 ( .A(n9871), .B(n14956), .ZN(n14954) );
  NAND2_X1 U12481 ( .A1(n9873), .A2(n9872), .ZN(n9875) );
  OAI21_X1 U12482 ( .B1(n9878), .B2(n9877), .A(n10225), .ZN(n9890) );
  NOR2_X1 U12483 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15348), .ZN(n12091) );
  AOI21_X1 U12484 ( .B1(n14996), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12091), .ZN(
        n9879) );
  OAI21_X1 U12485 ( .B1(n14993), .B2(n10234), .A(n9879), .ZN(n9889) );
  NAND2_X1 U12486 ( .A1(n9880), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9881) );
  INV_X1 U12487 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15175) );
  MUX2_X1 U12488 ( .A(n9884), .B(P3_REG1_REG_8__SCAN_IN), .S(n10234), .Z(n9885) );
  NAND2_X1 U12489 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  AOI21_X1 U12490 ( .B1(n10236), .B2(n9887), .A(n14977), .ZN(n9888) );
  AOI211_X1 U12491 ( .C1(n15007), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9891)
         );
  OAI21_X1 U12492 ( .B1(n9892), .B2(n14990), .A(n9891), .ZN(P3_U3190) );
  AOI211_X1 U12493 ( .C1(n9895), .C2(n9894), .A(n12219), .B(n9893), .ZN(n9896)
         );
  INV_X1 U12494 ( .A(n9896), .ZN(n9900) );
  NOR2_X1 U12495 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15360), .ZN(n14920) );
  OAI22_X1 U12496 ( .A1(n12187), .A2(n10247), .B1(n15097), .B2(n12213), .ZN(
        n9897) );
  AOI211_X1 U12497 ( .C1(n12193), .C2(n9898), .A(n14920), .B(n9897), .ZN(n9899) );
  OAI211_X1 U12498 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12191), .A(n9900), .B(
        n9899), .ZN(P3_U3158) );
  NAND2_X1 U12499 ( .A1(n13727), .A2(n11459), .ZN(n9905) );
  NAND2_X1 U12500 ( .A1(n13515), .A2(n11422), .ZN(n9904) );
  NAND2_X1 U12501 ( .A1(n9905), .A2(n9904), .ZN(n9906) );
  XNOR2_X1 U12502 ( .A(n9906), .B(n11410), .ZN(n10151) );
  NAND2_X1 U12503 ( .A1(n11367), .A2(n13727), .ZN(n9908) );
  NAND2_X1 U12504 ( .A1(n13515), .A2(n11234), .ZN(n9907) );
  NAND2_X1 U12505 ( .A1(n9908), .A2(n9907), .ZN(n10152) );
  XNOR2_X1 U12506 ( .A(n10151), .B(n10152), .ZN(n9909) );
  OAI211_X1 U12507 ( .C1(n9910), .C2(n9909), .A(n10155), .B(n14431), .ZN(n9917) );
  INV_X1 U12508 ( .A(n14436), .ZN(n13474) );
  INV_X1 U12509 ( .A(n9911), .ZN(n9915) );
  OAI22_X1 U12510 ( .A1(n10390), .A2(n14426), .B1(n14427), .B2(n9912), .ZN(
        n9913) );
  AOI211_X1 U12511 ( .C1(n13474), .C2(n9915), .A(n9914), .B(n9913), .ZN(n9916)
         );
  OAI211_X1 U12512 ( .C1(n10147), .C2(n14423), .A(n9917), .B(n9916), .ZN(
        P1_U3239) );
  INV_X1 U12513 ( .A(n12893), .ZN(n9918) );
  XNOR2_X1 U12514 ( .A(n11812), .B(n12892), .ZN(n12007) );
  NAND2_X1 U12515 ( .A1(n9921), .A2(n12007), .ZN(n9922) );
  NAND2_X1 U12516 ( .A1(n9937), .A2(n9922), .ZN(n14839) );
  NOR2_X1 U12517 ( .A1(n12007), .A2(n6897), .ZN(n9925) );
  AND2_X1 U12518 ( .A1(n9923), .A2(n9925), .ZN(n9926) );
  OAI21_X1 U12519 ( .B1(n9940), .B2(n9926), .A(n13251), .ZN(n9928) );
  NAND2_X1 U12520 ( .A1(n9928), .A2(n9927), .ZN(n14843) );
  INV_X1 U12521 ( .A(n14843), .ZN(n9929) );
  MUX2_X1 U12522 ( .A(n8698), .B(n9929), .S(n13228), .Z(n9935) );
  NAND2_X1 U12523 ( .A1(n9930), .A2(n14841), .ZN(n9946) );
  OAI211_X1 U12524 ( .C1(n9930), .C2(n14841), .A(n13332), .B(n9946), .ZN(
        n14840) );
  INV_X1 U12525 ( .A(n14840), .ZN(n9933) );
  OAI22_X1 U12526 ( .A1(n13231), .A2(n14841), .B1(n13232), .B2(n9931), .ZN(
        n9932) );
  AOI21_X1 U12527 ( .B1(n13245), .B2(n9933), .A(n9932), .ZN(n9934) );
  OAI211_X1 U12528 ( .C1(n13239), .C2(n14839), .A(n9935), .B(n9934), .ZN(
        P2_U3259) );
  INV_X1 U12529 ( .A(n12892), .ZN(n9941) );
  NAND2_X1 U12530 ( .A1(n9937), .A2(n9936), .ZN(n9939) );
  XNOR2_X1 U12531 ( .A(n11820), .B(n12891), .ZN(n12009) );
  INV_X1 U12532 ( .A(n12009), .ZN(n9938) );
  OAI21_X1 U12533 ( .B1(n9939), .B2(n9938), .A(n9954), .ZN(n14845) );
  XNOR2_X1 U12534 ( .A(n9957), .B(n12009), .ZN(n9943) );
  OAI21_X1 U12535 ( .B1(n9943), .B2(n13226), .A(n9942), .ZN(n14848) );
  INV_X1 U12536 ( .A(n14848), .ZN(n9944) );
  MUX2_X1 U12537 ( .A(n9945), .B(n9944), .S(n13228), .Z(n9952) );
  AOI21_X1 U12538 ( .B1(n9946), .B2(n11820), .A(n13243), .ZN(n9947) );
  NAND2_X1 U12539 ( .A1(n9947), .A2(n10054), .ZN(n14846) );
  INV_X1 U12540 ( .A(n14846), .ZN(n9950) );
  INV_X1 U12541 ( .A(n11820), .ZN(n14847) );
  OAI22_X1 U12542 ( .A1(n13231), .A2(n14847), .B1(n13232), .B2(n9948), .ZN(
        n9949) );
  AOI21_X1 U12543 ( .B1(n9950), .B2(n13245), .A(n9949), .ZN(n9951) );
  OAI211_X1 U12544 ( .C1(n13239), .C2(n14845), .A(n9952), .B(n9951), .ZN(
        P2_U3258) );
  NAND2_X1 U12545 ( .A1(n9954), .A2(n9953), .ZN(n10053) );
  XNOR2_X1 U12546 ( .A(n11826), .B(n9958), .ZN(n12012) );
  INV_X1 U12547 ( .A(n11826), .ZN(n14853) );
  NAND2_X1 U12548 ( .A1(n11826), .A2(n12890), .ZN(n9955) );
  INV_X1 U12549 ( .A(n12889), .ZN(n10283) );
  XNOR2_X1 U12550 ( .A(n14860), .B(n10283), .ZN(n12013) );
  NAND2_X1 U12551 ( .A1(n9956), .A2(n12013), .ZN(n10285) );
  OAI21_X1 U12552 ( .B1(n9956), .B2(n12013), .A(n10285), .ZN(n14862) );
  INV_X1 U12553 ( .A(n12012), .ZN(n10048) );
  XOR2_X1 U12554 ( .A(n10280), .B(n12013), .Z(n9960) );
  OAI21_X1 U12555 ( .B1(n9960), .B2(n13226), .A(n9959), .ZN(n14863) );
  NAND2_X1 U12556 ( .A1(n14863), .A2(n13228), .ZN(n9965) );
  AOI211_X1 U12557 ( .C1(n14860), .C2(n10055), .A(n13243), .B(n10288), .ZN(
        n14859) );
  INV_X1 U12558 ( .A(n14860), .ZN(n10284) );
  NOR2_X1 U12559 ( .A1(n13231), .A2(n10284), .ZN(n9963) );
  OAI22_X1 U12560 ( .A1(n13155), .A2(n9028), .B1(n9961), .B2(n13232), .ZN(
        n9962) );
  AOI211_X1 U12561 ( .C1(n14859), .C2(n13245), .A(n9963), .B(n9962), .ZN(n9964) );
  OAI211_X1 U12562 ( .C1(n13239), .C2(n14862), .A(n9965), .B(n9964), .ZN(
        P2_U3256) );
  NAND2_X1 U12563 ( .A1(n9966), .A2(n12764), .ZN(n9967) );
  OAI211_X1 U12564 ( .C1(n9968), .C2(n12771), .A(n9967), .B(n11162), .ZN(
        P3_U3272) );
  INV_X1 U12565 ( .A(n14647), .ZN(n14598) );
  AOI21_X1 U12566 ( .B1(n14598), .B2(n6464), .A(n14610), .ZN(n14004) );
  INV_X1 U12567 ( .A(n14004), .ZN(n14624) );
  NAND2_X1 U12568 ( .A1(n9970), .A2(n6468), .ZN(n9973) );
  AOI22_X1 U12569 ( .A1(n11284), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11283), 
        .B2(n9971), .ZN(n9972) );
  NAND2_X1 U12570 ( .A1(n9973), .A2(n9972), .ZN(n14585) );
  XNOR2_X1 U12571 ( .A(n14585), .B(n14682), .ZN(n14578) );
  NAND2_X1 U12572 ( .A1(n14577), .A2(n14576), .ZN(n9975) );
  OR2_X1 U12573 ( .A1(n14585), .A2(n14682), .ZN(n9974) );
  NAND2_X1 U12574 ( .A1(n9975), .A2(n9974), .ZN(n10326) );
  NAND2_X1 U12575 ( .A1(n9976), .A2(n6468), .ZN(n9979) );
  AOI22_X1 U12576 ( .A1(n11284), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11283), 
        .B2(n9977), .ZN(n9978) );
  NAND2_X1 U12577 ( .A1(n9979), .A2(n9978), .ZN(n14684) );
  NAND2_X1 U12578 ( .A1(n11483), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9988) );
  INV_X1 U12579 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9980) );
  OR2_X1 U12580 ( .A1(n13639), .A2(n9980), .ZN(n9987) );
  AND2_X1 U12581 ( .A1(n9982), .A2(n9981), .ZN(n9983) );
  OR2_X1 U12582 ( .A1(n9983), .A2(n9990), .ZN(n10389) );
  OR2_X1 U12583 ( .A1(n9585), .A2(n10389), .ZN(n9986) );
  OR2_X1 U12584 ( .A1(n6463), .A2(n9984), .ZN(n9985) );
  NAND4_X1 U12585 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n13726) );
  XNOR2_X1 U12586 ( .A(n14684), .B(n13726), .ZN(n13679) );
  INV_X1 U12587 ( .A(n13679), .ZN(n10325) );
  XNOR2_X1 U12588 ( .A(n10326), .B(n10325), .ZN(n14689) );
  INV_X1 U12589 ( .A(n14689), .ZN(n10008) );
  NAND2_X1 U12590 ( .A1(n11632), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9995) );
  OR2_X1 U12591 ( .A1(n13638), .A2(n9989), .ZN(n9994) );
  NAND2_X1 U12592 ( .A1(n9990), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10341) );
  OR2_X1 U12593 ( .A1(n9990), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U12594 ( .A1(n10341), .A2(n9991), .ZN(n14566) );
  OR2_X1 U12595 ( .A1(n9585), .A2(n14566), .ZN(n9993) );
  OR2_X1 U12596 ( .A1(n9589), .A2(n14725), .ZN(n9992) );
  NAND4_X1 U12597 ( .A1(n9995), .A2(n9994), .A3(n9993), .A4(n9992), .ZN(n13725) );
  INV_X1 U12598 ( .A(n13725), .ZN(n14705) );
  NOR2_X1 U12599 ( .A1(n10147), .A2(n13727), .ZN(n9996) );
  NAND2_X1 U12600 ( .A1(n10147), .A2(n13727), .ZN(n9998) );
  NAND2_X1 U12601 ( .A1(n9999), .A2(n9998), .ZN(n14579) );
  OAI211_X1 U12602 ( .C1(n6638), .C2(n13679), .A(n10349), .B(n14699), .ZN(
        n10000) );
  OAI21_X1 U12603 ( .B1(n14705), .B2(n14615), .A(n10000), .ZN(n14687) );
  INV_X1 U12604 ( .A(n14585), .ZN(n14676) );
  INV_X1 U12605 ( .A(n14684), .ZN(n10003) );
  OAI211_X1 U12606 ( .C1(n14586), .C2(n10003), .A(n14604), .B(n14569), .ZN(
        n14686) );
  NAND2_X1 U12607 ( .A1(n6464), .A2(n14683), .ZN(n14029) );
  INV_X1 U12608 ( .A(n14029), .ZN(n10366) );
  OAI22_X1 U12609 ( .A1(n6464), .A2(n10001), .B1(n10389), .B2(n14599), .ZN(
        n10002) );
  AOI21_X1 U12610 ( .B1(n10366), .B2(n14682), .A(n10002), .ZN(n10005) );
  OR2_X1 U12611 ( .A1(n13982), .A2(n10003), .ZN(n10004) );
  OAI211_X1 U12612 ( .C1(n14686), .C2(n14035), .A(n10005), .B(n10004), .ZN(
        n10006) );
  AOI21_X1 U12613 ( .B1(n14687), .B2(n6464), .A(n10006), .ZN(n10007) );
  OAI21_X1 U12614 ( .B1(n14004), .B2(n10008), .A(n10007), .ZN(P1_U3285) );
  INV_X1 U12615 ( .A(n10084), .ZN(n10017) );
  OAI21_X1 U12616 ( .B1(n10011), .B2(n10010), .A(n10009), .ZN(n10012) );
  NAND2_X1 U12617 ( .A1(n10012), .A2(n12203), .ZN(n10016) );
  OAI22_X1 U12618 ( .A1(n12187), .A2(n15055), .B1(n15071), .B2(n12213), .ZN(
        n10013) );
  AOI211_X1 U12619 ( .C1(n12193), .C2(n10083), .A(n10014), .B(n10013), .ZN(
        n10015) );
  OAI211_X1 U12620 ( .C1(n10017), .C2(n12191), .A(n10016), .B(n10015), .ZN(
        P3_U3170) );
  XNOR2_X1 U12621 ( .A(n10018), .B(n13673), .ZN(n14668) );
  INV_X1 U12622 ( .A(n14668), .ZN(n10028) );
  INV_X1 U12623 ( .A(n14623), .ZN(n14038) );
  XNOR2_X1 U12624 ( .A(n10020), .B(n10019), .ZN(n14661) );
  OAI211_X1 U12625 ( .C1(n14606), .C2(n10021), .A(n14604), .B(n10088), .ZN(
        n14664) );
  INV_X1 U12626 ( .A(n10022), .ZN(n10023) );
  INV_X1 U12627 ( .A(n14599), .ZN(n14621) );
  AOI22_X1 U12628 ( .A1(n14601), .A2(n14662), .B1(n10023), .B2(n14621), .ZN(
        n10025) );
  MUX2_X1 U12629 ( .A(n8806), .B(n14665), .S(n6464), .Z(n10024) );
  OAI211_X1 U12630 ( .C1(n14664), .C2(n14035), .A(n10025), .B(n10024), .ZN(
        n10026) );
  AOI21_X1 U12631 ( .B1(n14661), .B2(n14624), .A(n10026), .ZN(n10027) );
  OAI21_X1 U12632 ( .B1(n10028), .B2(n14038), .A(n10027), .ZN(P1_U3289) );
  NAND2_X1 U12633 ( .A1(n12235), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10029) );
  OAI21_X1 U12634 ( .B1(n12427), .B2(n12235), .A(n10029), .ZN(P3_U3520) );
  OAI21_X1 U12635 ( .B1(n10032), .B2(n10031), .A(n10030), .ZN(n10035) );
  INV_X1 U12636 ( .A(n10033), .ZN(n10034) );
  AOI21_X1 U12637 ( .B1(n10035), .B2(n13251), .A(n10034), .ZN(n10039) );
  OAI21_X1 U12638 ( .B1(n10037), .B2(n7021), .A(n10036), .ZN(n14824) );
  NAND2_X1 U12639 ( .A1(n14824), .A2(n14885), .ZN(n10038) );
  AND2_X1 U12640 ( .A1(n10039), .A2(n10038), .ZN(n14826) );
  OAI211_X1 U12641 ( .C1(n13242), .C2(n14822), .A(n13332), .B(n10040), .ZN(
        n14821) );
  OAI22_X1 U12642 ( .A1(n13155), .A2(n10042), .B1(n10041), .B2(n13232), .ZN(
        n10043) );
  AOI21_X1 U12643 ( .B1(n13248), .B2(n11781), .A(n10043), .ZN(n10044) );
  OAI21_X1 U12644 ( .B1(n13159), .B2(n14821), .A(n10044), .ZN(n10045) );
  AOI21_X1 U12645 ( .B1(n10046), .B2(n14824), .A(n10045), .ZN(n10047) );
  OAI21_X1 U12646 ( .B1(n6466), .B2(n14826), .A(n10047), .ZN(P2_U3263) );
  XNOR2_X1 U12647 ( .A(n10049), .B(n10048), .ZN(n10051) );
  AOI21_X1 U12648 ( .B1(n10051), .B2(n13251), .A(n10050), .ZN(n14854) );
  OAI21_X1 U12649 ( .B1(n10053), .B2(n12012), .A(n10052), .ZN(n14855) );
  INV_X1 U12650 ( .A(n14855), .ZN(n14858) );
  AOI21_X1 U12651 ( .B1(n10054), .B2(n11826), .A(n13243), .ZN(n10056) );
  NAND2_X1 U12652 ( .A1(n10056), .A2(n10055), .ZN(n14852) );
  OAI22_X1 U12653 ( .A1(n13155), .A2(n8762), .B1(n10057), .B2(n13232), .ZN(
        n10058) );
  AOI21_X1 U12654 ( .B1(n13248), .B2(n11826), .A(n10058), .ZN(n10059) );
  OAI21_X1 U12655 ( .B1(n14852), .B2(n13159), .A(n10059), .ZN(n10060) );
  AOI21_X1 U12656 ( .B1(n14858), .B2(n13246), .A(n10060), .ZN(n10061) );
  OAI21_X1 U12657 ( .B1(n14854), .B2(n6466), .A(n10061), .ZN(P2_U3257) );
  AND2_X1 U12658 ( .A1(n11121), .A2(n10960), .ZN(n15083) );
  NAND2_X1 U12659 ( .A1(n15107), .A2(n15083), .ZN(n12447) );
  INV_X1 U12660 ( .A(n12447), .ZN(n15030) );
  OR2_X1 U12661 ( .A1(n10062), .A2(n11133), .ZN(n10063) );
  NAND2_X1 U12662 ( .A1(n10064), .A2(n10063), .ZN(n15123) );
  OAI22_X1 U12663 ( .A1(n15049), .A2(n15120), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15053), .ZN(n10073) );
  NAND2_X1 U12664 ( .A1(n15123), .A2(n15080), .ZN(n10071) );
  NAND2_X1 U12665 ( .A1(n10065), .A2(n11133), .ZN(n10066) );
  NAND3_X1 U12666 ( .A1(n10067), .A2(n15099), .A3(n10066), .ZN(n10070) );
  OAI22_X1 U12667 ( .A1(n10247), .A2(n15096), .B1(n15097), .B2(n15072), .ZN(
        n10068) );
  INV_X1 U12668 ( .A(n10068), .ZN(n10069) );
  NAND3_X1 U12669 ( .A1(n10071), .A2(n10070), .A3(n10069), .ZN(n15121) );
  MUX2_X1 U12670 ( .A(n15121), .B(P3_REG2_REG_3__SCAN_IN), .S(n15068), .Z(
        n10072) );
  AOI211_X1 U12671 ( .C1(n15030), .C2(n15123), .A(n10073), .B(n10072), .ZN(
        n10074) );
  INV_X1 U12672 ( .A(n10074), .ZN(P3_U3230) );
  XNOR2_X1 U12673 ( .A(n10076), .B(n10075), .ZN(n15125) );
  XNOR2_X1 U12674 ( .A(n10077), .B(n11131), .ZN(n10080) );
  OAI22_X1 U12675 ( .A1(n15071), .A2(n15072), .B1(n15055), .B2(n15096), .ZN(
        n10079) );
  INV_X1 U12676 ( .A(n15080), .ZN(n12453) );
  NOR2_X1 U12677 ( .A1(n15125), .A2(n12453), .ZN(n10078) );
  AOI211_X1 U12678 ( .C1(n10080), .C2(n15099), .A(n10079), .B(n10078), .ZN(
        n15126) );
  MUX2_X1 U12679 ( .A(n10081), .B(n15126), .S(n15107), .Z(n10086) );
  INV_X1 U12680 ( .A(n10082), .ZN(n15064) );
  AND2_X1 U12681 ( .A1(n10083), .A2(n15151), .ZN(n15128) );
  AOI22_X1 U12682 ( .A1(n15064), .A2(n15128), .B1(n15102), .B2(n10084), .ZN(
        n10085) );
  OAI211_X1 U12683 ( .C1(n15125), .C2(n12447), .A(n10086), .B(n10085), .ZN(
        P3_U3229) );
  XNOR2_X1 U12684 ( .A(n10087), .B(n10093), .ZN(n14674) );
  OAI211_X1 U12685 ( .C1(n7197), .C2(n14671), .A(n14604), .B(n10089), .ZN(
        n14670) );
  INV_X1 U12686 ( .A(n10090), .ZN(n10091) );
  AOI22_X1 U12687 ( .A1(n14601), .A2(n13511), .B1(n14621), .B2(n10091), .ZN(
        n10092) );
  OAI21_X1 U12688 ( .B1(n14035), .B2(n14670), .A(n10092), .ZN(n10099) );
  INV_X1 U12689 ( .A(n14699), .ZN(n14629) );
  XNOR2_X1 U12690 ( .A(n10094), .B(n10093), .ZN(n10097) );
  NAND2_X1 U12691 ( .A1(n14674), .A2(n14598), .ZN(n10096) );
  AOI22_X1 U12692 ( .A1(n14635), .A2(n13727), .B1(n13729), .B2(n14683), .ZN(
        n10095) );
  OAI211_X1 U12693 ( .C1(n14629), .C2(n10097), .A(n10096), .B(n10095), .ZN(
        n14672) );
  MUX2_X1 U12694 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n14672), .S(n6464), .Z(
        n10098) );
  AOI211_X1 U12695 ( .C1(n14674), .C2(n14610), .A(n10099), .B(n10098), .ZN(
        n10100) );
  INV_X1 U12696 ( .A(n10100), .ZN(P1_U3288) );
  INV_X1 U12697 ( .A(n10101), .ZN(n10102) );
  NAND2_X1 U12698 ( .A1(n10104), .A2(SI_21_), .ZN(n10105) );
  MUX2_X1 U12699 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n11332), .Z(n10254) );
  XNOR2_X1 U12700 ( .A(n11333), .B(n10254), .ZN(n11542) );
  INV_X1 U12701 ( .A(n11542), .ZN(n10107) );
  OAI222_X1 U12702 ( .A1(n13368), .A2(n11543), .B1(n13366), .B2(n10107), .C1(
        n11956), .C2(P2_U3088), .ZN(P2_U3305) );
  XOR2_X1 U12703 ( .A(n13675), .B(n10108), .Z(n14640) );
  AND2_X1 U12704 ( .A1(n6464), .A2(n14635), .ZN(n14032) );
  OAI22_X1 U12705 ( .A1(n13982), .A2(n10110), .B1(n10109), .B2(n14599), .ZN(
        n10113) );
  INV_X1 U12706 ( .A(n10124), .ZN(n10111) );
  AOI21_X1 U12707 ( .B1(n14632), .B2(n6668), .A(n10111), .ZN(n10114) );
  NAND2_X1 U12708 ( .A1(n10114), .A2(n14604), .ZN(n14637) );
  NOR2_X1 U12709 ( .A1(n14035), .A2(n14637), .ZN(n10112) );
  AOI211_X1 U12710 ( .C1(n14032), .C2(n14636), .A(n10113), .B(n10112), .ZN(
        n10121) );
  AOI21_X1 U12711 ( .B1(n13675), .B2(n13732), .A(n14629), .ZN(n10118) );
  INV_X1 U12712 ( .A(n10114), .ZN(n10115) );
  XNOR2_X1 U12713 ( .A(n14616), .B(n10115), .ZN(n10116) );
  NOR2_X1 U12714 ( .A1(n10116), .A2(n14629), .ZN(n10117) );
  OAI22_X1 U12715 ( .A1(n14683), .A2(n10118), .B1(n10117), .B2(n13732), .ZN(
        n14641) );
  MUX2_X1 U12716 ( .A(n10119), .B(n14641), .S(n6464), .Z(n10120) );
  OAI211_X1 U12717 ( .C1(n14004), .C2(n14640), .A(n10121), .B(n10120), .ZN(
        P1_U3292) );
  XNOR2_X1 U12718 ( .A(n10122), .B(n13496), .ZN(n14645) );
  OAI22_X1 U12719 ( .A1(n6464), .A2(n9129), .B1(n10123), .B2(n14599), .ZN(
        n10127) );
  AOI21_X1 U12720 ( .B1(n10124), .B2(n13498), .A(n13980), .ZN(n10125) );
  NAND2_X1 U12721 ( .A1(n10125), .A2(n14603), .ZN(n14648) );
  NOR2_X1 U12722 ( .A1(n14035), .A2(n14648), .ZN(n10126) );
  AOI211_X1 U12723 ( .C1(n14601), .C2(n13498), .A(n10127), .B(n10126), .ZN(
        n10133) );
  XNOR2_X1 U12724 ( .A(n13678), .B(n10128), .ZN(n10131) );
  INV_X1 U12725 ( .A(n10129), .ZN(n10130) );
  OAI21_X1 U12726 ( .B1(n10131), .B2(n14629), .A(n10130), .ZN(n14651) );
  NAND2_X1 U12727 ( .A1(n14651), .A2(n6464), .ZN(n10132) );
  OAI211_X1 U12728 ( .C1(n14004), .C2(n14645), .A(n10133), .B(n10132), .ZN(
        P1_U3291) );
  INV_X1 U12729 ( .A(n10134), .ZN(n10138) );
  NOR2_X1 U12730 ( .A1(n14614), .A2(n13664), .ZN(n10135) );
  INV_X1 U12731 ( .A(n14225), .ZN(n13657) );
  NAND2_X1 U12732 ( .A1(n10135), .A2(n13657), .ZN(n14646) );
  AOI211_X1 U12733 ( .C1(n10138), .C2(n14697), .A(n10137), .B(n10136), .ZN(
        n10150) );
  NAND2_X1 U12734 ( .A1(n11638), .A2(n10143), .ZN(n10139) );
  NAND2_X1 U12735 ( .A1(n14714), .A2(n14701), .ZN(n14209) );
  INV_X1 U12736 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10140) );
  OAI22_X1 U12737 ( .A1(n14209), .A2(n10147), .B1(n14714), .B2(n10140), .ZN(
        n10141) );
  INV_X1 U12738 ( .A(n10141), .ZN(n10142) );
  OAI21_X1 U12739 ( .B1(n10150), .B2(n14713), .A(n10142), .ZN(P1_U3477) );
  NAND3_X1 U12740 ( .A1(n13711), .A2(n11638), .A3(n10143), .ZN(n10144) );
  OAI22_X1 U12741 ( .A1(n14155), .A2(n10147), .B1(n14730), .B2(n10146), .ZN(
        n10148) );
  INV_X1 U12742 ( .A(n10148), .ZN(n10149) );
  OAI21_X1 U12743 ( .B1(n10150), .B2(n14727), .A(n10149), .ZN(P1_U3534) );
  INV_X1 U12744 ( .A(n10151), .ZN(n10153) );
  NAND2_X1 U12745 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  NAND2_X1 U12746 ( .A1(n10155), .A2(n10154), .ZN(n10160) );
  NAND2_X1 U12747 ( .A1(n14585), .A2(n11422), .ZN(n10157) );
  NAND2_X1 U12748 ( .A1(n14682), .A2(n11234), .ZN(n10156) );
  NAND2_X1 U12749 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  XNOR2_X1 U12750 ( .A(n10158), .B(n11477), .ZN(n10380) );
  AOI22_X1 U12751 ( .A1(n14585), .A2(n11436), .B1(n11367), .B2(n14682), .ZN(
        n10381) );
  XNOR2_X1 U12752 ( .A(n10380), .B(n10381), .ZN(n10159) );
  OAI211_X1 U12753 ( .C1(n10160), .C2(n10159), .A(n10384), .B(n14431), .ZN(
        n10166) );
  NAND2_X1 U12754 ( .A1(n13726), .A2(n14635), .ZN(n10162) );
  NAND2_X1 U12755 ( .A1(n13727), .A2(n14683), .ZN(n10161) );
  NAND2_X1 U12756 ( .A1(n10162), .A2(n10161), .ZN(n14582) );
  NOR2_X1 U12757 ( .A1(n14436), .A2(n14583), .ZN(n10163) );
  AOI211_X1 U12758 ( .C1(n14387), .C2(n14582), .A(n10164), .B(n10163), .ZN(
        n10165) );
  OAI211_X1 U12759 ( .C1(n14676), .C2(n14423), .A(n10166), .B(n10165), .ZN(
        P1_U3213) );
  INV_X1 U12760 ( .A(n10167), .ZN(n10168) );
  OR2_X1 U12761 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  AOI22_X1 U12762 ( .A1(n10172), .A2(n11506), .B1(n11507), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n10173) );
  XNOR2_X1 U12763 ( .A(n11837), .B(n11736), .ZN(n10176) );
  AND2_X1 U12764 ( .A1(n12888), .A2(n9668), .ZN(n10175) );
  NAND2_X1 U12765 ( .A1(n10176), .A2(n10175), .ZN(n10190) );
  OAI21_X1 U12766 ( .B1(n10176), .B2(n10175), .A(n10190), .ZN(n10267) );
  INV_X1 U12767 ( .A(n12888), .ZN(n11839) );
  NOR2_X1 U12768 ( .A1(n12828), .A2(n11839), .ZN(n10177) );
  AOI22_X1 U12769 ( .A1(n10265), .A2(n12808), .B1(n10177), .B2(n10176), .ZN(
        n10207) );
  AOI22_X1 U12770 ( .A1(n10178), .A2(n11506), .B1(n11507), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n10179) );
  XNOR2_X1 U12771 ( .A(n14878), .B(n11579), .ZN(n10305) );
  NAND2_X1 U12772 ( .A1(n11958), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10189) );
  INV_X1 U12773 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10181) );
  OR2_X1 U12774 ( .A1(n11743), .A2(n10181), .ZN(n10188) );
  OAI21_X1 U12775 ( .B1(n10184), .B2(n10182), .A(n9255), .ZN(n10185) );
  NAND2_X1 U12776 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n10183) );
  NAND2_X1 U12777 ( .A1(n10185), .A2(n10194), .ZN(n10300) );
  OR2_X1 U12778 ( .A1(n11741), .A2(n10300), .ZN(n10187) );
  OR2_X1 U12779 ( .A1(n11962), .A2(n9249), .ZN(n10186) );
  NAND4_X1 U12780 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n12887) );
  NAND2_X1 U12781 ( .A1(n12887), .A2(n9668), .ZN(n10306) );
  XNOR2_X1 U12782 ( .A(n10305), .B(n10306), .ZN(n10191) );
  INV_X1 U12783 ( .A(n10191), .ZN(n10206) );
  INV_X1 U12784 ( .A(n10190), .ZN(n10192) );
  NAND2_X1 U12785 ( .A1(n14878), .A2(n12875), .ZN(n10203) );
  NAND2_X1 U12786 ( .A1(n11958), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10200) );
  OR2_X1 U12787 ( .A1(n11962), .A2(n12932), .ZN(n10199) );
  NAND2_X1 U12788 ( .A1(n10194), .A2(n10193), .ZN(n10195) );
  NAND2_X1 U12789 ( .A1(n10469), .A2(n10195), .ZN(n10446) );
  OR2_X1 U12790 ( .A1(n11741), .A2(n10446), .ZN(n10198) );
  INV_X1 U12791 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10196) );
  OR2_X1 U12792 ( .A1(n11743), .A2(n10196), .ZN(n10197) );
  NAND4_X1 U12793 ( .A1(n10200), .A2(n10199), .A3(n10198), .A4(n10197), .ZN(
        n12886) );
  AOI22_X1 U12794 ( .A1(n13020), .A2(n12888), .B1(n12886), .B2(n12858), .ZN(
        n10296) );
  INV_X1 U12795 ( .A(n10296), .ZN(n10201) );
  AOI22_X1 U12796 ( .A1(n12871), .A2(n10201), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10202) );
  OAI211_X1 U12797 ( .C1(n12873), .C2(n10300), .A(n10203), .B(n10202), .ZN(
        n10204) );
  AOI21_X1 U12798 ( .B1(n10321), .B2(n12808), .A(n10204), .ZN(n10205) );
  OAI21_X1 U12799 ( .B1(n10207), .B2(n10206), .A(n10205), .ZN(P2_U3208) );
  OR2_X1 U12800 ( .A1(n10208), .A2(n11130), .ZN(n10209) );
  NAND2_X1 U12801 ( .A1(n10210), .A2(n10209), .ZN(n15135) );
  INV_X1 U12802 ( .A(n15135), .ZN(n10221) );
  OAI22_X1 U12803 ( .A1(n10247), .A2(n15072), .B1(n10401), .B2(n15096), .ZN(
        n10211) );
  AOI21_X1 U12804 ( .B1(n15135), .B2(n15080), .A(n10211), .ZN(n10217) );
  NAND2_X1 U12805 ( .A1(n10212), .A2(n11130), .ZN(n10213) );
  NAND2_X1 U12806 ( .A1(n10214), .A2(n10213), .ZN(n10215) );
  NAND2_X1 U12807 ( .A1(n10215), .A2(n15099), .ZN(n10216) );
  NAND2_X1 U12808 ( .A1(n10217), .A2(n10216), .ZN(n15133) );
  MUX2_X1 U12809 ( .A(n15133), .B(P3_REG2_REG_5__SCAN_IN), .S(n15068), .Z(
        n10218) );
  INV_X1 U12810 ( .A(n10218), .ZN(n10220) );
  AOI22_X1 U12811 ( .A1(n12627), .A2(n10249), .B1(n15102), .B2(n10250), .ZN(
        n10219) );
  OAI211_X1 U12812 ( .C1(n10221), .C2(n12447), .A(n10220), .B(n10219), .ZN(
        P3_U3228) );
  INV_X1 U12813 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U12814 ( .A1(n10234), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10222) );
  AOI21_X1 U12815 ( .B1(n10228), .B2(n10224), .A(n10563), .ZN(n10244) );
  INV_X1 U12816 ( .A(n10234), .ZN(n10226) );
  INV_X1 U12817 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10238) );
  MUX2_X1 U12818 ( .A(n10228), .B(n10238), .S(n12369), .Z(n10229) );
  NAND2_X1 U12819 ( .A1(n10229), .A2(n10571), .ZN(n10582) );
  INV_X1 U12820 ( .A(n10229), .ZN(n10230) );
  NAND2_X1 U12821 ( .A1(n10230), .A2(n7055), .ZN(n10581) );
  NAND2_X1 U12822 ( .A1(n10582), .A2(n10581), .ZN(n10231) );
  XNOR2_X1 U12823 ( .A(n10583), .B(n10231), .ZN(n10242) );
  NAND2_X1 U12824 ( .A1(n14983), .A2(n10571), .ZN(n10233) );
  NOR2_X1 U12825 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7912), .ZN(n10661) );
  AOI21_X1 U12826 ( .B1(n14996), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10661), .ZN(
        n10232) );
  NAND2_X1 U12827 ( .A1(n10233), .A2(n10232), .ZN(n10241) );
  NAND2_X1 U12828 ( .A1(n10234), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10235) );
  AOI21_X1 U12829 ( .B1(n10238), .B2(n10237), .A(n10572), .ZN(n10239) );
  NOR2_X1 U12830 ( .A1(n10239), .A2(n14977), .ZN(n10240) );
  AOI211_X1 U12831 ( .C1(n15007), .C2(n10242), .A(n10241), .B(n10240), .ZN(
        n10243) );
  OAI21_X1 U12832 ( .B1(n10244), .B2(n14990), .A(n10243), .ZN(P3_U3191) );
  XOR2_X1 U12833 ( .A(n10246), .B(n10245), .Z(n10253) );
  NOR2_X1 U12834 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7852), .ZN(n14935) );
  OAI22_X1 U12835 ( .A1(n12187), .A2(n10401), .B1(n10247), .B2(n12213), .ZN(
        n10248) );
  AOI211_X1 U12836 ( .C1(n12193), .C2(n10249), .A(n14935), .B(n10248), .ZN(
        n10252) );
  NAND2_X1 U12837 ( .A1(n12217), .A2(n10250), .ZN(n10251) );
  OAI211_X1 U12838 ( .C1(n10253), .C2(n12219), .A(n10252), .B(n10251), .ZN(
        P3_U3167) );
  NAND2_X1 U12839 ( .A1(n10255), .A2(SI_22_), .ZN(n10256) );
  MUX2_X1 U12840 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n11332), .Z(n10441) );
  XNOR2_X1 U12841 ( .A(n10441), .B(SI_23_), .ZN(n10438) );
  XNOR2_X1 U12842 ( .A(n10440), .B(n10438), .ZN(n11575) );
  NAND2_X1 U12843 ( .A1(n11575), .A2(n10257), .ZN(n10259) );
  OR2_X1 U12844 ( .A1(n10258), .A2(P2_U3088), .ZN(n12041) );
  OAI211_X1 U12845 ( .C1(n11576), .C2(n13368), .A(n10259), .B(n12041), .ZN(
        P2_U3304) );
  INV_X1 U12846 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11352) );
  NAND2_X1 U12847 ( .A1(n11575), .A2(n14215), .ZN(n10260) );
  OAI211_X1 U12848 ( .C1(n11352), .C2(n14223), .A(n10260), .B(n13714), .ZN(
        P1_U3332) );
  NAND2_X1 U12849 ( .A1(n12887), .A2(n12858), .ZN(n10262) );
  NAND2_X1 U12850 ( .A1(n12889), .A2(n13020), .ZN(n10261) );
  NAND2_X1 U12851 ( .A1(n10262), .A2(n10261), .ZN(n10281) );
  NAND2_X1 U12852 ( .A1(n12871), .A2(n10281), .ZN(n10264) );
  OAI211_X1 U12853 ( .C1(n12873), .C2(n10289), .A(n10264), .B(n10263), .ZN(
        n10269) );
  AOI211_X1 U12854 ( .C1(n10267), .C2(n10266), .A(n12877), .B(n10265), .ZN(
        n10268) );
  AOI211_X1 U12855 ( .C1(n11837), .C2(n12875), .A(n10269), .B(n10268), .ZN(
        n10270) );
  INV_X1 U12856 ( .A(n10270), .ZN(P2_U3189) );
  INV_X1 U12857 ( .A(n15060), .ZN(n10279) );
  OAI211_X1 U12858 ( .C1(n10273), .C2(n10272), .A(n10271), .B(n12203), .ZN(
        n10278) );
  OAI22_X1 U12859 ( .A1(n12187), .A2(n15056), .B1(n15055), .B2(n12213), .ZN(
        n10274) );
  AOI211_X1 U12860 ( .C1(n12193), .C2(n10276), .A(n10275), .B(n10274), .ZN(
        n10277) );
  OAI211_X1 U12861 ( .C1(n10279), .C2(n12191), .A(n10278), .B(n10277), .ZN(
        P3_U3179) );
  XNOR2_X1 U12862 ( .A(n11837), .B(n12888), .ZN(n12015) );
  XNOR2_X1 U12863 ( .A(n10295), .B(n12015), .ZN(n10282) );
  AOI21_X1 U12864 ( .B1(n10282), .B2(n13251), .A(n10281), .ZN(n14869) );
  INV_X1 U12865 ( .A(n12015), .ZN(n10286) );
  OAI21_X1 U12866 ( .B1(n10287), .B2(n10286), .A(n10294), .ZN(n14870) );
  INV_X1 U12867 ( .A(n14870), .ZN(n14874) );
  OAI211_X1 U12868 ( .C1(n10288), .C2(n14868), .A(n10299), .B(n13332), .ZN(
        n14866) );
  OAI22_X1 U12869 ( .A1(n13155), .A2(n9029), .B1(n10289), .B2(n13232), .ZN(
        n10290) );
  AOI21_X1 U12870 ( .B1(n13248), .B2(n11837), .A(n10290), .ZN(n10291) );
  OAI21_X1 U12871 ( .B1(n14866), .B2(n13159), .A(n10291), .ZN(n10292) );
  AOI21_X1 U12872 ( .B1(n14874), .B2(n13246), .A(n10292), .ZN(n10293) );
  OAI21_X1 U12873 ( .B1(n14869), .B2(n6466), .A(n10293), .ZN(P2_U3255) );
  XOR2_X1 U12874 ( .A(n12887), .B(n14878), .Z(n12014) );
  XNOR2_X1 U12875 ( .A(n10444), .B(n12014), .ZN(n14882) );
  XOR2_X1 U12876 ( .A(n10450), .B(n12014), .Z(n10297) );
  OAI21_X1 U12877 ( .B1(n10297), .B2(n13226), .A(n10296), .ZN(n14876) );
  NAND2_X1 U12878 ( .A1(n14876), .A2(n13228), .ZN(n10304) );
  INV_X1 U12879 ( .A(n10445), .ZN(n10298) );
  AOI211_X1 U12880 ( .C1(n14878), .C2(n10299), .A(n13243), .B(n10298), .ZN(
        n14877) );
  INV_X1 U12881 ( .A(n14878), .ZN(n10449) );
  NOR2_X1 U12882 ( .A1(n10449), .A2(n13231), .ZN(n10302) );
  OAI22_X1 U12883 ( .A1(n13155), .A2(n9249), .B1(n10300), .B2(n13232), .ZN(
        n10301) );
  AOI211_X1 U12884 ( .C1(n14877), .C2(n13245), .A(n10302), .B(n10301), .ZN(
        n10303) );
  OAI211_X1 U12885 ( .C1(n13239), .C2(n14882), .A(n10304), .B(n10303), .ZN(
        P2_U3254) );
  INV_X1 U12886 ( .A(n10305), .ZN(n10318) );
  INV_X1 U12887 ( .A(n10306), .ZN(n10307) );
  NOR2_X1 U12888 ( .A1(n10318), .A2(n10307), .ZN(n10309) );
  AOI22_X1 U12889 ( .A1(n11507), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11506), 
        .B2(n12948), .ZN(n10308) );
  XNOR2_X1 U12890 ( .A(n11851), .B(n11736), .ZN(n10458) );
  NAND2_X1 U12891 ( .A1(n12886), .A2(n9668), .ZN(n10456) );
  NAND2_X1 U12892 ( .A1(n11959), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10314) );
  INV_X1 U12893 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10310) );
  OR2_X1 U12894 ( .A1(n6950), .A2(n10310), .ZN(n10313) );
  INV_X1 U12895 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10527) );
  OR2_X1 U12896 ( .A1(n11962), .A2(n10527), .ZN(n10312) );
  INV_X1 U12897 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10599) );
  XNOR2_X1 U12898 ( .A(n10469), .B(n10599), .ZN(n10598) );
  OR2_X1 U12899 ( .A1(n11741), .A2(n10598), .ZN(n10311) );
  NAND4_X1 U12900 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n12885) );
  NAND2_X1 U12901 ( .A1(n12885), .A2(n12858), .ZN(n10316) );
  NAND2_X1 U12902 ( .A1(n12887), .A2(n13020), .ZN(n10315) );
  NAND2_X1 U12903 ( .A1(n10316), .A2(n10315), .ZN(n10451) );
  AOI22_X1 U12904 ( .A1(n12871), .A2(n10451), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10317) );
  OAI21_X1 U12905 ( .B1(n10446), .B2(n12873), .A(n10317), .ZN(n10323) );
  AOI22_X1 U12906 ( .A1(n10318), .A2(n12808), .B1(n11651), .B2(n12887), .ZN(
        n10320) );
  NOR3_X1 U12907 ( .A1(n10321), .A2(n10320), .A3(n10319), .ZN(n10322) );
  AOI211_X1 U12908 ( .C1(n11851), .C2(n12875), .A(n10323), .B(n10322), .ZN(
        n10324) );
  OAI21_X1 U12909 ( .B1(n10457), .B2(n12877), .A(n10324), .ZN(P2_U3196) );
  NAND2_X1 U12910 ( .A1(n10326), .A2(n10325), .ZN(n10328) );
  OR2_X1 U12911 ( .A1(n14684), .A2(n13726), .ZN(n10327) );
  NAND2_X1 U12912 ( .A1(n10329), .A2(n6468), .ZN(n10332) );
  AOI22_X1 U12913 ( .A1(n11284), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11283), 
        .B2(n10330), .ZN(n10331) );
  XNOR2_X1 U12914 ( .A(n14570), .B(n13725), .ZN(n14561) );
  INV_X1 U12915 ( .A(n14561), .ZN(n10333) );
  OR2_X1 U12916 ( .A1(n14570), .A2(n13725), .ZN(n10334) );
  NAND2_X1 U12917 ( .A1(n10335), .A2(n6468), .ZN(n10338) );
  AOI22_X1 U12918 ( .A1(n11284), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10336), 
        .B2(n11283), .ZN(n10337) );
  NAND2_X1 U12919 ( .A1(n11483), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10346) );
  INV_X1 U12920 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10339) );
  OR2_X1 U12921 ( .A1(n13639), .A2(n10339), .ZN(n10345) );
  NAND2_X1 U12922 ( .A1(n10341), .A2(n10340), .ZN(n10342) );
  NAND2_X1 U12923 ( .A1(n10356), .A2(n10342), .ZN(n10648) );
  OR2_X1 U12924 ( .A1(n9585), .A2(n10648), .ZN(n10344) );
  OR2_X1 U12925 ( .A1(n9589), .A2(n14728), .ZN(n10343) );
  NAND4_X1 U12926 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n13724) );
  XNOR2_X1 U12927 ( .A(n14702), .B(n14404), .ZN(n13683) );
  XNOR2_X1 U12928 ( .A(n10553), .B(n13683), .ZN(n14709) );
  INV_X1 U12929 ( .A(n14709), .ZN(n10371) );
  INV_X1 U12930 ( .A(n13726), .ZN(n10347) );
  OR2_X1 U12931 ( .A1(n14684), .A2(n10347), .ZN(n10348) );
  NAND2_X1 U12932 ( .A1(n14560), .A2(n14561), .ZN(n14559) );
  NAND2_X1 U12933 ( .A1(n14570), .A2(n14705), .ZN(n10350) );
  OR2_X1 U12934 ( .A1(n10351), .A2(n7220), .ZN(n10352) );
  AND2_X1 U12935 ( .A1(n10352), .A2(n10551), .ZN(n14700) );
  INV_X1 U12936 ( .A(n14702), .ZN(n10656) );
  NAND2_X1 U12937 ( .A1(n14571), .A2(n14702), .ZN(n10353) );
  NAND2_X1 U12938 ( .A1(n10353), .A2(n14604), .ZN(n10354) );
  OR2_X1 U12939 ( .A1(n6628), .A2(n10354), .ZN(n10363) );
  NAND2_X1 U12940 ( .A1(n11632), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10361) );
  AND2_X1 U12941 ( .A1(n10356), .A2(n10355), .ZN(n10357) );
  OR2_X1 U12942 ( .A1(n10357), .A2(n10541), .ZN(n14419) );
  OR2_X1 U12943 ( .A1(n9585), .A2(n14419), .ZN(n10360) );
  OR2_X1 U12944 ( .A1(n13638), .A2(n10556), .ZN(n10359) );
  OR2_X1 U12945 ( .A1(n6463), .A2(n14461), .ZN(n10358) );
  NAND4_X1 U12946 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n13723) );
  NAND2_X1 U12947 ( .A1(n13723), .A2(n14635), .ZN(n10362) );
  NAND2_X1 U12948 ( .A1(n10363), .A2(n10362), .ZN(n14707) );
  NAND2_X1 U12949 ( .A1(n14707), .A2(n14609), .ZN(n10368) );
  OAI22_X1 U12950 ( .A1(n6464), .A2(n10364), .B1(n10648), .B2(n14599), .ZN(
        n10365) );
  AOI21_X1 U12951 ( .B1(n10366), .B2(n13725), .A(n10365), .ZN(n10367) );
  OAI211_X1 U12952 ( .C1(n10656), .C2(n13982), .A(n10368), .B(n10367), .ZN(
        n10369) );
  AOI21_X1 U12953 ( .B1(n14700), .B2(n14623), .A(n10369), .ZN(n10370) );
  OAI21_X1 U12954 ( .B1(n14004), .B2(n10371), .A(n10370), .ZN(P1_U3283) );
  INV_X1 U12955 ( .A(n10372), .ZN(n10373) );
  NAND2_X1 U12956 ( .A1(n10373), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10374) );
  OAI21_X1 U12957 ( .B1(n10375), .B2(P3_STATE_REG_SCAN_IN), .A(n10374), .ZN(
        P3_U3271) );
  NAND2_X1 U12958 ( .A1(n14684), .A2(n11422), .ZN(n10377) );
  NAND2_X1 U12959 ( .A1(n13726), .A2(n11234), .ZN(n10376) );
  NAND2_X1 U12960 ( .A1(n10377), .A2(n10376), .ZN(n10378) );
  XNOR2_X1 U12961 ( .A(n10378), .B(n11410), .ZN(n10505) );
  AND2_X1 U12962 ( .A1(n11367), .A2(n13726), .ZN(n10379) );
  AOI21_X1 U12963 ( .B1(n14684), .B2(n11436), .A(n10379), .ZN(n10504) );
  XNOR2_X1 U12964 ( .A(n10505), .B(n10504), .ZN(n10387) );
  INV_X1 U12965 ( .A(n10380), .ZN(n10382) );
  OR2_X1 U12966 ( .A1(n10382), .A2(n10381), .ZN(n10383) );
  INV_X1 U12967 ( .A(n10507), .ZN(n10385) );
  AOI21_X1 U12968 ( .B1(n10387), .B2(n10386), .A(n10385), .ZN(n10394) );
  OAI21_X1 U12969 ( .B1(n14436), .B2(n10389), .A(n10388), .ZN(n10392) );
  OAI22_X1 U12970 ( .A1(n14705), .A2(n14426), .B1(n14427), .B2(n10390), .ZN(
        n10391) );
  AOI211_X1 U12971 ( .C1(n14684), .C2(n14415), .A(n10392), .B(n10391), .ZN(
        n10393) );
  OAI21_X1 U12972 ( .B1(n10394), .B2(n14410), .A(n10393), .ZN(P1_U3221) );
  OR2_X1 U12973 ( .A1(n10395), .A2(n11128), .ZN(n10396) );
  NAND2_X1 U12974 ( .A1(n10397), .A2(n10396), .ZN(n15144) );
  INV_X1 U12975 ( .A(n15144), .ZN(n10409) );
  XNOR2_X1 U12976 ( .A(n10398), .B(n11128), .ZN(n10399) );
  NAND2_X1 U12977 ( .A1(n10399), .A2(n15099), .ZN(n10404) );
  NAND2_X1 U12978 ( .A1(n15044), .A2(n15045), .ZN(n10400) );
  OAI21_X1 U12979 ( .B1(n10401), .B2(n15072), .A(n10400), .ZN(n10402) );
  AOI21_X1 U12980 ( .B1(n15144), .B2(n15080), .A(n10402), .ZN(n10403) );
  NAND2_X1 U12981 ( .A1(n10404), .A2(n10403), .ZN(n15142) );
  MUX2_X1 U12982 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n15142), .S(n15107), .Z(
        n10405) );
  INV_X1 U12983 ( .A(n10405), .ZN(n10408) );
  NOR2_X1 U12984 ( .A1(n10406), .A2(n15131), .ZN(n15143) );
  AOI22_X1 U12985 ( .A1(n15143), .A2(n15064), .B1(n15102), .B2(n12070), .ZN(
        n10407) );
  OAI211_X1 U12986 ( .C1(n10409), .C2(n12447), .A(n10408), .B(n10407), .ZN(
        P3_U3226) );
  INV_X1 U12987 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10410) );
  MUX2_X1 U12988 ( .A(n10410), .B(P1_REG2_REG_17__SCAN_IN), .S(n11269), .Z(
        n10794) );
  INV_X1 U12989 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U12990 ( .A1(n10705), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U12991 ( .A1(n10412), .A2(n10411), .ZN(n10413) );
  NOR2_X1 U12992 ( .A1(n10927), .A2(n10413), .ZN(n10414) );
  XNOR2_X1 U12993 ( .A(n10413), .B(n10927), .ZN(n14534) );
  NOR2_X1 U12994 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14534), .ZN(n14533) );
  NOR2_X1 U12995 ( .A1(n10414), .A2(n14533), .ZN(n13800) );
  MUX2_X1 U12996 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n14028), .S(n13796), .Z(
        n13799) );
  NAND2_X1 U12997 ( .A1(n13800), .A2(n13799), .ZN(n13798) );
  OAI21_X1 U12998 ( .B1(n14028), .B2(n10419), .A(n13798), .ZN(n10796) );
  XOR2_X1 U12999 ( .A(n10794), .B(n10796), .Z(n10427) );
  NOR2_X1 U13000 ( .A1(n14553), .A2(n10790), .ZN(n10425) );
  NAND2_X1 U13001 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3086), .ZN(n14401)
         );
  INV_X1 U13002 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14143) );
  AOI21_X1 U13003 ( .B1(n10416), .B2(n14455), .A(n10415), .ZN(n10417) );
  NOR2_X1 U13004 ( .A1(n10927), .A2(n10417), .ZN(n10418) );
  XNOR2_X1 U13005 ( .A(n10927), .B(n10417), .ZN(n14532) );
  NOR2_X1 U13006 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14532), .ZN(n14531) );
  NOR2_X1 U13007 ( .A1(n10418), .A2(n14531), .ZN(n13794) );
  MUX2_X1 U13008 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14143), .S(n13796), .Z(
        n13793) );
  NAND2_X1 U13009 ( .A1(n13794), .A2(n13793), .ZN(n13792) );
  OAI21_X1 U13010 ( .B1(n14143), .B2(n10419), .A(n13792), .ZN(n10422) );
  NOR2_X1 U13011 ( .A1(n11269), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n10420) );
  AOI21_X1 U13012 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n11269), .A(n10420), 
        .ZN(n10421) );
  NAND2_X1 U13013 ( .A1(n10422), .A2(n10421), .ZN(n10789) );
  OAI211_X1 U13014 ( .C1(n10422), .C2(n10421), .A(n10789), .B(n14545), .ZN(
        n10423) );
  NAND2_X1 U13015 ( .A1(n14401), .A2(n10423), .ZN(n10424) );
  AOI211_X1 U13016 ( .C1(n14517), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n10425), 
        .B(n10424), .ZN(n10426) );
  OAI21_X1 U13017 ( .B1(n10427), .B2(n14536), .A(n10426), .ZN(P1_U3260) );
  XOR2_X1 U13018 ( .A(n11129), .B(n15037), .Z(n10431) );
  AOI22_X1 U13019 ( .A1(n12228), .A2(n15093), .B1(n15045), .B2(n15024), .ZN(
        n10430) );
  XNOR2_X1 U13020 ( .A(n10428), .B(n11129), .ZN(n15149) );
  NAND2_X1 U13021 ( .A1(n15149), .A2(n15080), .ZN(n10429) );
  OAI211_X1 U13022 ( .C1(n10431), .C2(n15075), .A(n10430), .B(n10429), .ZN(
        n15146) );
  INV_X1 U13023 ( .A(n15146), .ZN(n10437) );
  NOR2_X1 U13024 ( .A1(n10432), .A2(n15131), .ZN(n15147) );
  AOI22_X1 U13025 ( .A1(n15064), .A2(n15147), .B1(n15102), .B2(n12093), .ZN(
        n10433) );
  OAI21_X1 U13026 ( .B1(n10434), .B2(n15107), .A(n10433), .ZN(n10435) );
  AOI21_X1 U13027 ( .B1(n15149), .B2(n15030), .A(n10435), .ZN(n10436) );
  OAI21_X1 U13028 ( .B1(n10437), .B2(n15068), .A(n10436), .ZN(P3_U3225) );
  INV_X1 U13029 ( .A(n10438), .ZN(n10439) );
  MUX2_X1 U13030 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n11332), .Z(n10533) );
  INV_X1 U13031 ( .A(n11663), .ZN(n10945) );
  OAI222_X1 U13032 ( .A1(n13368), .A2(n11664), .B1(n13366), .B2(n10945), .C1(
        P2_U3088), .C2(n10442), .ZN(P2_U3303) );
  NAND2_X1 U13033 ( .A1(n10449), .A2(n7527), .ZN(n10443) );
  XNOR2_X1 U13034 ( .A(n11851), .B(n12886), .ZN(n12016) );
  XNOR2_X1 U13035 ( .A(n10520), .B(n12016), .ZN(n10499) );
  AOI211_X1 U13036 ( .C1(n11851), .C2(n10445), .A(n13243), .B(n10525), .ZN(
        n10496) );
  INV_X1 U13037 ( .A(n11851), .ZN(n10523) );
  INV_X1 U13038 ( .A(n10446), .ZN(n10447) );
  AOI22_X1 U13039 ( .A1(n6466), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n10447), 
        .B2(n13247), .ZN(n10448) );
  OAI21_X1 U13040 ( .B1(n10523), .B2(n13231), .A(n10448), .ZN(n10454) );
  XNOR2_X1 U13041 ( .A(n10522), .B(n12016), .ZN(n10452) );
  AOI21_X1 U13042 ( .B1(n10452), .B2(n13251), .A(n10451), .ZN(n10498) );
  NOR2_X1 U13043 ( .A1(n10498), .A2(n6466), .ZN(n10453) );
  AOI211_X1 U13044 ( .C1(n10496), .C2(n13245), .A(n10454), .B(n10453), .ZN(
        n10455) );
  OAI21_X1 U13045 ( .B1(n10499), .B2(n13239), .A(n10455), .ZN(P2_U3253) );
  INV_X1 U13046 ( .A(n10456), .ZN(n10459) );
  AOI22_X1 U13047 ( .A1(n11507), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11506), 
        .B2(n14746), .ZN(n10460) );
  XNOR2_X1 U13048 ( .A(n11860), .B(n11736), .ZN(n10463) );
  AND2_X1 U13049 ( .A1(n12885), .A2(n9668), .ZN(n10462) );
  NAND2_X1 U13050 ( .A1(n10463), .A2(n10462), .ZN(n10477) );
  OAI21_X1 U13051 ( .B1(n10463), .B2(n10462), .A(n10477), .ZN(n10596) );
  INV_X1 U13052 ( .A(n12885), .ZN(n10684) );
  NOR2_X1 U13053 ( .A1(n12828), .A2(n10684), .ZN(n10464) );
  AOI22_X1 U13054 ( .A1(n10594), .A2(n12808), .B1(n10464), .B2(n10463), .ZN(
        n10492) );
  AOI22_X1 U13055 ( .A1(n11507), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n11506), 
        .B2(n12949), .ZN(n10465) );
  XNOR2_X1 U13056 ( .A(n11866), .B(n11579), .ZN(n11185) );
  NAND2_X1 U13057 ( .A1(n11958), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10476) );
  INV_X1 U13058 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10679) );
  OR2_X1 U13059 ( .A1(n11962), .A2(n10679), .ZN(n10475) );
  NAND2_X1 U13060 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n10467) );
  INV_X1 U13061 ( .A(n10481), .ZN(n10471) );
  INV_X1 U13062 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10468) );
  OAI21_X1 U13063 ( .B1(n10469), .B2(n10599), .A(n10468), .ZN(n10470) );
  NAND2_X1 U13064 ( .A1(n10471), .A2(n10470), .ZN(n10678) );
  OR2_X1 U13065 ( .A1(n11741), .A2(n10678), .ZN(n10474) );
  INV_X1 U13066 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10472) );
  OR2_X1 U13067 ( .A1(n11743), .A2(n10472), .ZN(n10473) );
  NAND4_X1 U13068 ( .A1(n10476), .A2(n10475), .A3(n10474), .A4(n10473), .ZN(
        n12884) );
  NAND2_X1 U13069 ( .A1(n12884), .A2(n9668), .ZN(n11184) );
  XNOR2_X1 U13070 ( .A(n11185), .B(n11184), .ZN(n10479) );
  INV_X1 U13071 ( .A(n10479), .ZN(n10491) );
  INV_X1 U13072 ( .A(n10477), .ZN(n10478) );
  NAND2_X1 U13073 ( .A1(n11186), .A2(n12808), .ZN(n10490) );
  NAND2_X1 U13074 ( .A1(n11959), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n10486) );
  INV_X1 U13075 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10835) );
  OR2_X1 U13076 ( .A1(n11962), .A2(n10835), .ZN(n10485) );
  INV_X1 U13077 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10480) );
  OR2_X1 U13078 ( .A1(n6950), .A2(n10480), .ZN(n10484) );
  OR2_X1 U13079 ( .A1(n10481), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U13080 ( .A1(n10887), .A2(n10482), .ZN(n11655) );
  OR2_X1 U13081 ( .A1(n11741), .A2(n11655), .ZN(n10483) );
  NAND4_X1 U13082 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n12883) );
  INV_X1 U13083 ( .A(n12883), .ZN(n11187) );
  OAI22_X1 U13084 ( .A1(n11187), .A2(n12988), .B1(n10684), .B2(n12775), .ZN(
        n10676) );
  AOI22_X1 U13085 ( .A1(n12871), .A2(n10676), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10487) );
  OAI21_X1 U13086 ( .B1(n10678), .B2(n12873), .A(n10487), .ZN(n10488) );
  AOI21_X1 U13087 ( .B1(n11866), .B2(n12875), .A(n10488), .ZN(n10489) );
  OAI211_X1 U13088 ( .C1(n10492), .C2(n10491), .A(n10490), .B(n10489), .ZN(
        P2_U3187) );
  INV_X1 U13089 ( .A(n10493), .ZN(n10494) );
  OAI222_X1 U13090 ( .A1(n10495), .A2(P3_U3151), .B1(n12771), .B2(n10536), 
        .C1(n12770), .C2(n10494), .ZN(P3_U3270) );
  AOI21_X1 U13091 ( .B1(n14879), .B2(n11851), .A(n10496), .ZN(n10497) );
  OAI211_X1 U13092 ( .C1(n13337), .C2(n10499), .A(n10498), .B(n10497), .ZN(
        n10502) );
  NAND2_X1 U13093 ( .A1(n10502), .A2(n14908), .ZN(n10500) );
  OAI21_X1 U13094 ( .B1(n14908), .B2(n10501), .A(n10500), .ZN(P2_U3511) );
  NAND2_X1 U13095 ( .A1(n10502), .A2(n14887), .ZN(n10503) );
  OAI21_X1 U13096 ( .B1(n14887), .B2(n10196), .A(n10503), .ZN(P2_U3466) );
  NAND2_X1 U13097 ( .A1(n10505), .A2(n10504), .ZN(n10506) );
  NAND2_X1 U13098 ( .A1(n14570), .A2(n11436), .ZN(n10509) );
  NAND2_X1 U13099 ( .A1(n11367), .A2(n13725), .ZN(n10508) );
  INV_X1 U13100 ( .A(n10639), .ZN(n10643) );
  XNOR2_X1 U13101 ( .A(n10641), .B(n10643), .ZN(n10633) );
  NAND2_X1 U13102 ( .A1(n14570), .A2(n11422), .ZN(n10511) );
  NAND2_X1 U13103 ( .A1(n13725), .A2(n11436), .ZN(n10510) );
  NAND2_X1 U13104 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  XNOR2_X1 U13105 ( .A(n10512), .B(n11410), .ZN(n10638) );
  INV_X1 U13106 ( .A(n10638), .ZN(n10642) );
  XNOR2_X1 U13107 ( .A(n10633), .B(n10642), .ZN(n10519) );
  NAND2_X1 U13108 ( .A1(n13724), .A2(n14635), .ZN(n10514) );
  NAND2_X1 U13109 ( .A1(n13726), .A2(n14683), .ZN(n10513) );
  NAND2_X1 U13110 ( .A1(n10514), .A2(n10513), .ZN(n14564) );
  NAND2_X1 U13111 ( .A1(n14387), .A2(n14564), .ZN(n10516) );
  OAI211_X1 U13112 ( .C1(n14436), .C2(n14566), .A(n10516), .B(n10515), .ZN(
        n10517) );
  AOI21_X1 U13113 ( .B1(n14570), .B2(n14415), .A(n10517), .ZN(n10518) );
  OAI21_X1 U13114 ( .B1(n10519), .B2(n14410), .A(n10518), .ZN(P1_U3231) );
  INV_X1 U13115 ( .A(n12886), .ZN(n11853) );
  NOR2_X1 U13116 ( .A1(n10685), .A2(n12885), .ZN(n10674) );
  NOR2_X1 U13117 ( .A1(n11860), .A2(n10684), .ZN(n10673) );
  NOR2_X1 U13118 ( .A1(n10674), .A2(n10673), .ZN(n12018) );
  XNOR2_X1 U13119 ( .A(n10683), .B(n12018), .ZN(n10691) );
  XOR2_X1 U13120 ( .A(n12018), .B(n10675), .Z(n10524) );
  AOI22_X1 U13121 ( .A1(n13020), .A2(n12886), .B1(n12884), .B2(n12858), .ZN(
        n10600) );
  OAI21_X1 U13122 ( .B1(n10524), .B2(n13226), .A(n10600), .ZN(n10688) );
  NAND2_X1 U13123 ( .A1(n10688), .A2(n13228), .ZN(n10531) );
  INV_X1 U13124 ( .A(n10525), .ZN(n10526) );
  AOI211_X1 U13125 ( .C1(n11860), .C2(n10526), .A(n13243), .B(n10680), .ZN(
        n10689) );
  NOR2_X1 U13126 ( .A1(n10685), .A2(n13231), .ZN(n10529) );
  OAI22_X1 U13127 ( .A1(n13155), .A2(n10527), .B1(n10598), .B2(n13232), .ZN(
        n10528) );
  AOI211_X1 U13128 ( .C1(n10689), .C2(n13245), .A(n10529), .B(n10528), .ZN(
        n10530) );
  OAI211_X1 U13129 ( .C1(n10691), .C2(n13239), .A(n10531), .B(n10530), .ZN(
        P2_U3252) );
  NAND2_X1 U13130 ( .A1(n10534), .A2(SI_24_), .ZN(n10535) );
  MUX2_X1 U13131 ( .A(n11395), .B(n11672), .S(n11332), .Z(n10537) );
  NAND2_X1 U13132 ( .A1(n10537), .A2(n10536), .ZN(n10746) );
  INV_X1 U13133 ( .A(n10537), .ZN(n10538) );
  NAND2_X1 U13134 ( .A1(n10538), .A2(SI_25_), .ZN(n10539) );
  NAND2_X1 U13135 ( .A1(n10746), .A2(n10539), .ZN(n10744) );
  XNOR2_X1 U13136 ( .A(n10745), .B(n10744), .ZN(n11671) );
  INV_X1 U13137 ( .A(n11671), .ZN(n11164) );
  OAI222_X1 U13138 ( .A1(n13368), .A2(n11672), .B1(n13366), .B2(n11164), .C1(
        P2_U3088), .C2(n10540), .ZN(P2_U3302) );
  NAND2_X1 U13139 ( .A1(n11632), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10546) );
  OR2_X1 U13140 ( .A1(n13638), .A2(n9444), .ZN(n10545) );
  NOR2_X1 U13141 ( .A1(n10541), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10542) );
  OR2_X1 U13142 ( .A1(n10612), .A2(n10542), .ZN(n10901) );
  OR2_X1 U13143 ( .A1(n9585), .A2(n10901), .ZN(n10544) );
  OR2_X1 U13144 ( .A1(n6463), .A2(n10817), .ZN(n10543) );
  NAND4_X1 U13145 ( .A1(n10546), .A2(n10545), .A3(n10544), .A4(n10543), .ZN(
        n13722) );
  NAND2_X1 U13146 ( .A1(n10547), .A2(n6468), .ZN(n10549) );
  AOI22_X1 U13147 ( .A1(n11284), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n13783), 
        .B2(n11283), .ZN(n10548) );
  XNOR2_X1 U13148 ( .A(n14416), .B(n10649), .ZN(n13682) );
  OR2_X1 U13149 ( .A1(n14702), .A2(n14404), .ZN(n10550) );
  XOR2_X1 U13150 ( .A(n13682), .B(n10606), .Z(n10552) );
  OAI222_X1 U13151 ( .A1(n14704), .A2(n14404), .B1(n14615), .B2(n14405), .C1(
        n10552), .C2(n14629), .ZN(n14458) );
  INV_X1 U13152 ( .A(n14458), .ZN(n10561) );
  OR2_X1 U13153 ( .A1(n14702), .A2(n13724), .ZN(n10554) );
  XNOR2_X1 U13154 ( .A(n10622), .B(n13682), .ZN(n14460) );
  INV_X1 U13155 ( .A(n14416), .ZN(n14457) );
  INV_X1 U13156 ( .A(n10625), .ZN(n10555) );
  OAI211_X1 U13157 ( .C1(n14457), .C2(n6628), .A(n10555), .B(n14604), .ZN(
        n14456) );
  OAI22_X1 U13158 ( .A1(n6464), .A2(n10556), .B1(n14419), .B2(n14599), .ZN(
        n10557) );
  AOI21_X1 U13159 ( .B1(n14416), .B2(n14601), .A(n10557), .ZN(n10558) );
  OAI21_X1 U13160 ( .B1(n14456), .B2(n14035), .A(n10558), .ZN(n10559) );
  AOI21_X1 U13161 ( .B1(n14460), .B2(n14624), .A(n10559), .ZN(n10560) );
  OAI21_X1 U13162 ( .B1(n10561), .B2(n14016), .A(n10560), .ZN(P1_U3282) );
  INV_X1 U13163 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n10569) );
  NOR2_X1 U13164 ( .A1(n10571), .A2(n10562), .ZN(n10564) );
  NOR2_X1 U13165 ( .A1(n10564), .A2(n10563), .ZN(n14970) );
  INV_X1 U13166 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10565) );
  OR2_X1 U13167 ( .A1(n14982), .A2(n10565), .ZN(n10567) );
  NAND2_X1 U13168 ( .A1(n14982), .A2(n10565), .ZN(n10566) );
  NAND2_X1 U13169 ( .A1(n10567), .A2(n10566), .ZN(n14969) );
  AOI21_X1 U13170 ( .B1(n10569), .B2(n10568), .A(n12236), .ZN(n10593) );
  INV_X1 U13171 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n10869) );
  INV_X1 U13172 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10573) );
  OR2_X1 U13173 ( .A1(n14982), .A2(n10573), .ZN(n10575) );
  NAND2_X1 U13174 ( .A1(n14982), .A2(n10573), .ZN(n10574) );
  NAND2_X1 U13175 ( .A1(n10575), .A2(n10574), .ZN(n14975) );
  AOI21_X1 U13176 ( .B1(n10869), .B2(n10576), .A(n12242), .ZN(n10577) );
  NOR2_X1 U13177 ( .A1(n10577), .A2(n14977), .ZN(n10591) );
  MUX2_X1 U13178 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12369), .Z(n12249) );
  XNOR2_X1 U13179 ( .A(n12249), .B(n10578), .ZN(n10586) );
  MUX2_X1 U13180 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12369), .Z(n10580) );
  NOR2_X1 U13181 ( .A1(n10580), .A2(n10579), .ZN(n10584) );
  AOI21_X1 U13182 ( .B1(n10580), .B2(n10579), .A(n10584), .ZN(n14985) );
  AOI21_X1 U13183 ( .B1(n10586), .B2(n10585), .A(n12250), .ZN(n10589) );
  NAND2_X1 U13184 ( .A1(n14983), .A2(n12251), .ZN(n10588) );
  INV_X1 U13185 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15345) );
  NOR2_X1 U13186 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15345), .ZN(n12176) );
  AOI21_X1 U13187 ( .B1(n14996), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12176), 
        .ZN(n10587) );
  OAI211_X1 U13188 ( .C1(n10589), .C2(n14911), .A(n10588), .B(n10587), .ZN(
        n10590) );
  NOR2_X1 U13189 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  OAI21_X1 U13190 ( .B1(n10593), .B2(n14990), .A(n10592), .ZN(P3_U3193) );
  AOI211_X1 U13191 ( .C1(n10596), .C2(n10595), .A(n12877), .B(n10594), .ZN(
        n10597) );
  INV_X1 U13192 ( .A(n10597), .ZN(n10604) );
  INV_X1 U13193 ( .A(n10598), .ZN(n10602) );
  OAI22_X1 U13194 ( .A1(n12859), .A2(n10600), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10599), .ZN(n10601) );
  AOI21_X1 U13195 ( .B1(n10602), .B2(n12861), .A(n10601), .ZN(n10603) );
  OAI211_X1 U13196 ( .C1(n10685), .C2(n12865), .A(n10604), .B(n10603), .ZN(
        P2_U3206) );
  NOR2_X1 U13197 ( .A1(n14416), .A2(n10649), .ZN(n10605) );
  NAND2_X1 U13198 ( .A1(n10607), .A2(n6468), .ZN(n10610) );
  AOI22_X1 U13199 ( .A1(n10608), .A2(n11283), .B1(n11284), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n10609) );
  XNOR2_X1 U13200 ( .A(n13538), .B(n14405), .ZN(n13684) );
  OAI211_X1 U13201 ( .C1(n10611), .C2(n10717), .A(n10771), .B(n14699), .ZN(
        n10620) );
  NAND2_X1 U13202 ( .A1(n11632), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10617) );
  OR2_X1 U13203 ( .A1(n10612), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10613) );
  NAND2_X1 U13204 ( .A1(n10709), .A2(n10613), .ZN(n13448) );
  OR2_X1 U13205 ( .A1(n9585), .A2(n13448), .ZN(n10616) );
  OR2_X1 U13206 ( .A1(n9589), .A2(n10829), .ZN(n10615) );
  OR2_X1 U13207 ( .A1(n13638), .A2(n9445), .ZN(n10614) );
  NAND4_X1 U13208 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n14446) );
  NAND2_X1 U13209 ( .A1(n14446), .A2(n14635), .ZN(n10619) );
  NAND2_X1 U13210 ( .A1(n13723), .A2(n14683), .ZN(n10618) );
  AND2_X1 U13211 ( .A1(n10619), .A2(n10618), .ZN(n10904) );
  AND2_X1 U13212 ( .A1(n10620), .A2(n10904), .ZN(n10813) );
  NOR2_X1 U13213 ( .A1(n14416), .A2(n13723), .ZN(n10621) );
  NAND2_X1 U13214 ( .A1(n14416), .A2(n13723), .ZN(n10623) );
  NAND2_X1 U13215 ( .A1(n10624), .A2(n10623), .ZN(n10718) );
  XNOR2_X1 U13216 ( .A(n10718), .B(n10717), .ZN(n10810) );
  NAND2_X1 U13217 ( .A1(n10625), .A2(n10819), .ZN(n10763) );
  OAI211_X1 U13218 ( .C1(n10625), .C2(n10819), .A(n14604), .B(n10763), .ZN(
        n10811) );
  OAI22_X1 U13219 ( .A1(n6464), .A2(n9444), .B1(n10901), .B2(n14599), .ZN(
        n10626) );
  AOI21_X1 U13220 ( .B1(n13538), .B2(n14601), .A(n10626), .ZN(n10627) );
  OAI21_X1 U13221 ( .B1(n10811), .B2(n14035), .A(n10627), .ZN(n10628) );
  AOI21_X1 U13222 ( .B1(n10810), .B2(n14624), .A(n10628), .ZN(n10629) );
  OAI21_X1 U13223 ( .B1(n10813), .B2(n14016), .A(n10629), .ZN(P1_U3281) );
  INV_X1 U13224 ( .A(n10630), .ZN(n10631) );
  OAI222_X1 U13225 ( .A1(n10632), .A2(P3_U3151), .B1(n12771), .B2(n15358), 
        .C1(n12770), .C2(n10631), .ZN(P3_U3269) );
  AOI22_X1 U13226 ( .A1(n10633), .A2(n10638), .B1(n10639), .B2(n10641), .ZN(
        n10647) );
  NAND2_X1 U13227 ( .A1(n14702), .A2(n11422), .ZN(n10635) );
  NAND2_X1 U13228 ( .A1(n13724), .A2(n11459), .ZN(n10634) );
  NAND2_X1 U13229 ( .A1(n10635), .A2(n10634), .ZN(n10636) );
  XNOR2_X1 U13230 ( .A(n10636), .B(n11477), .ZN(n10916) );
  AND2_X1 U13231 ( .A1(n11367), .A2(n13724), .ZN(n10637) );
  AOI21_X1 U13232 ( .B1(n14702), .B2(n11436), .A(n10637), .ZN(n10914) );
  XNOR2_X1 U13233 ( .A(n10916), .B(n10914), .ZN(n10646) );
  NAND2_X1 U13234 ( .A1(n10642), .A2(n10643), .ZN(n10640) );
  AND2_X1 U13235 ( .A1(n10646), .A2(n10644), .ZN(n10645) );
  OAI211_X1 U13236 ( .C1(n10647), .C2(n10646), .A(n14431), .B(n14408), .ZN(
        n10655) );
  INV_X1 U13237 ( .A(n10648), .ZN(n10653) );
  OAI22_X1 U13238 ( .A1(n10649), .A2(n14426), .B1(n14427), .B2(n14705), .ZN(
        n10652) );
  INV_X1 U13239 ( .A(n10650), .ZN(n10651) );
  AOI211_X1 U13240 ( .C1(n10653), .C2(n13474), .A(n10652), .B(n10651), .ZN(
        n10654) );
  OAI211_X1 U13241 ( .C1(n10656), .C2(n14423), .A(n10655), .B(n10654), .ZN(
        P1_U3217) );
  AOI21_X1 U13242 ( .B1(n10658), .B2(n10657), .A(n6633), .ZN(n10665) );
  OAI22_X1 U13243 ( .A1(n12187), .A2(n12179), .B1(n10659), .B2(n12213), .ZN(
        n10660) );
  AOI211_X1 U13244 ( .C1(n12193), .C2(n15152), .A(n10661), .B(n10660), .ZN(
        n10664) );
  NAND2_X1 U13245 ( .A1(n12217), .A2(n10662), .ZN(n10663) );
  OAI211_X1 U13246 ( .C1(n10665), .C2(n12219), .A(n10664), .B(n10663), .ZN(
        P3_U3171) );
  XOR2_X1 U13247 ( .A(n10666), .B(n11137), .Z(n10667) );
  OAI222_X1 U13248 ( .A1(n15096), .A2(n14356), .B1(n15072), .B2(n12179), .C1(
        n10667), .C2(n15075), .ZN(n10867) );
  INV_X1 U13249 ( .A(n10867), .ZN(n10672) );
  XNOR2_X1 U13250 ( .A(n10668), .B(n11137), .ZN(n10868) );
  NAND2_X1 U13251 ( .A1(n15107), .A2(n15034), .ZN(n12579) );
  AOI22_X1 U13252 ( .A1(n15068), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15102), 
        .B2(n12175), .ZN(n10669) );
  OAI21_X1 U13253 ( .B1(n15049), .B2(n10874), .A(n10669), .ZN(n10670) );
  AOI21_X1 U13254 ( .B1(n10868), .B2(n15065), .A(n10670), .ZN(n10671) );
  OAI21_X1 U13255 ( .B1(n10672), .B2(n15068), .A(n10671), .ZN(P3_U3222) );
  INV_X1 U13256 ( .A(n12884), .ZN(n11868) );
  XNOR2_X1 U13257 ( .A(n11866), .B(n11868), .ZN(n12021) );
  XNOR2_X1 U13258 ( .A(n10837), .B(n12021), .ZN(n10677) );
  AOI21_X1 U13259 ( .B1(n10677), .B2(n13251), .A(n10676), .ZN(n10738) );
  OAI22_X1 U13260 ( .A1(n13155), .A2(n10679), .B1(n10678), .B2(n13232), .ZN(
        n10682) );
  NAND2_X1 U13261 ( .A1(n10836), .A2(n10680), .ZN(n10847) );
  OAI211_X1 U13262 ( .C1(n10836), .C2(n10680), .A(n13332), .B(n10847), .ZN(
        n10737) );
  NOR2_X1 U13263 ( .A1(n10737), .A2(n13159), .ZN(n10681) );
  AOI211_X1 U13264 ( .C1(n13248), .C2(n11866), .A(n10682), .B(n10681), .ZN(
        n10687) );
  XNOR2_X1 U13265 ( .A(n6624), .B(n12021), .ZN(n10740) );
  NAND2_X1 U13266 ( .A1(n10740), .A2(n13246), .ZN(n10686) );
  OAI211_X1 U13267 ( .C1(n10738), .C2(n6466), .A(n10687), .B(n10686), .ZN(
        P2_U3251) );
  AOI211_X1 U13268 ( .C1(n14879), .C2(n11860), .A(n10689), .B(n10688), .ZN(
        n10690) );
  OAI21_X1 U13269 ( .B1(n13337), .B2(n10691), .A(n10690), .ZN(n10693) );
  NAND2_X1 U13270 ( .A1(n10693), .A2(n14908), .ZN(n10692) );
  OAI21_X1 U13271 ( .B1(n14908), .B2(n10310), .A(n10692), .ZN(P2_U3512) );
  INV_X1 U13272 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10695) );
  NAND2_X1 U13273 ( .A1(n10693), .A2(n14887), .ZN(n10694) );
  OAI21_X1 U13274 ( .B1(n14887), .B2(n10695), .A(n10694), .ZN(P2_U3469) );
  OR2_X1 U13275 ( .A1(n13538), .A2(n14405), .ZN(n10768) );
  NAND2_X1 U13276 ( .A1(n10771), .A2(n10768), .ZN(n10701) );
  NAND2_X1 U13277 ( .A1(n10696), .A2(n6468), .ZN(n10700) );
  OAI22_X1 U13278 ( .A1(n14520), .A2(n11335), .B1(n13653), .B2(n10697), .ZN(
        n10698) );
  INV_X1 U13279 ( .A(n10698), .ZN(n10699) );
  XNOR2_X1 U13280 ( .A(n13550), .B(n14446), .ZN(n13685) );
  INV_X1 U13281 ( .A(n14446), .ZN(n14375) );
  OR2_X1 U13282 ( .A1(n13550), .A2(n14375), .ZN(n10702) );
  NAND2_X1 U13283 ( .A1(n10704), .A2(n6468), .ZN(n10707) );
  AOI22_X1 U13284 ( .A1(n10705), .A2(n11283), .B1(n11284), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10706) );
  NAND2_X1 U13285 ( .A1(n11632), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n10714) );
  NAND2_X1 U13286 ( .A1(n10709), .A2(n10708), .ZN(n10710) );
  NAND2_X1 U13287 ( .A1(n10722), .A2(n10710), .ZN(n14384) );
  OR2_X1 U13288 ( .A1(n9585), .A2(n14384), .ZN(n10713) );
  OR2_X1 U13289 ( .A1(n6463), .A2(n14455), .ZN(n10712) );
  OR2_X1 U13290 ( .A1(n13638), .A2(n9440), .ZN(n10711) );
  INV_X1 U13291 ( .A(n14428), .ZN(n14147) );
  XNOR2_X1 U13292 ( .A(n14445), .B(n14147), .ZN(n13559) );
  XNOR2_X1 U13293 ( .A(n10924), .B(n13689), .ZN(n10715) );
  NAND2_X1 U13294 ( .A1(n10715), .A2(n14699), .ZN(n14451) );
  OR2_X1 U13295 ( .A1(n13538), .A2(n13722), .ZN(n10716) );
  INV_X1 U13296 ( .A(n13685), .ZN(n10759) );
  OR2_X1 U13297 ( .A1(n13550), .A2(n14446), .ZN(n10719) );
  XNOR2_X1 U13298 ( .A(n10930), .B(n13689), .ZN(n14454) );
  OR2_X2 U13299 ( .A1(n10763), .A2(n13550), .ZN(n10764) );
  AOI21_X1 U13300 ( .B1(n10764), .B2(n14445), .A(n13980), .ZN(n10720) );
  NAND2_X1 U13301 ( .A1(n10720), .A2(n6616), .ZN(n14449) );
  INV_X1 U13302 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10721) );
  NAND2_X1 U13303 ( .A1(n10722), .A2(n10721), .ZN(n10723) );
  NAND2_X1 U13304 ( .A1(n10934), .A2(n10723), .ZN(n14435) );
  INV_X1 U13305 ( .A(n14435), .ZN(n10724) );
  INV_X1 U13306 ( .A(n9585), .ZN(n11227) );
  NAND2_X1 U13307 ( .A1(n10724), .A2(n11227), .ZN(n10730) );
  NAND2_X1 U13308 ( .A1(n11632), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n10729) );
  INV_X1 U13309 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10725) );
  OR2_X1 U13310 ( .A1(n9589), .A2(n10725), .ZN(n10728) );
  INV_X1 U13311 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10726) );
  OR2_X1 U13312 ( .A1(n13638), .A2(n10726), .ZN(n10727) );
  NAND4_X1 U13313 ( .A1(n10730), .A2(n10729), .A3(n10728), .A4(n10727), .ZN(
        n14447) );
  OAI22_X1 U13314 ( .A1(n6464), .A2(n9440), .B1(n14384), .B2(n14599), .ZN(
        n10731) );
  AOI21_X1 U13315 ( .B1(n14032), .B2(n14447), .A(n10731), .ZN(n10732) );
  OAI21_X1 U13316 ( .B1(n14375), .B2(n14029), .A(n10732), .ZN(n10733) );
  AOI21_X1 U13317 ( .B1(n14445), .B2(n14601), .A(n10733), .ZN(n10734) );
  OAI21_X1 U13318 ( .B1(n14449), .B2(n14035), .A(n10734), .ZN(n10735) );
  AOI21_X1 U13319 ( .B1(n14454), .B2(n14624), .A(n10735), .ZN(n10736) );
  OAI21_X1 U13320 ( .B1(n14451), .B2(n14016), .A(n10736), .ZN(P1_U3279) );
  OAI211_X1 U13321 ( .C1(n10836), .C2(n14867), .A(n10738), .B(n10737), .ZN(
        n10739) );
  AOI21_X1 U13322 ( .B1(n14850), .B2(n10740), .A(n10739), .ZN(n10743) );
  NAND2_X1 U13323 ( .A1(n14905), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10741) );
  OAI21_X1 U13324 ( .B1(n10743), .B2(n14905), .A(n10741), .ZN(P2_U3513) );
  NAND2_X1 U13325 ( .A1(n14886), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10742) );
  OAI21_X1 U13326 ( .B1(n10743), .B2(n14886), .A(n10742), .ZN(P2_U3472) );
  MUX2_X1 U13327 ( .A(n11419), .B(n11689), .S(n11332), .Z(n11170) );
  XNOR2_X1 U13328 ( .A(n11170), .B(SI_26_), .ZN(n11167) );
  XNOR2_X1 U13329 ( .A(n11169), .B(n11167), .ZN(n11688) );
  INV_X1 U13330 ( .A(n11688), .ZN(n10748) );
  OAI222_X1 U13331 ( .A1(n10747), .A2(P1_U3086), .B1(n14221), .B2(n10748), 
        .C1(n11419), .C2(n14223), .ZN(P1_U3329) );
  OAI222_X1 U13332 ( .A1(P2_U3088), .A2(n10749), .B1(n13366), .B2(n10748), 
        .C1(n11689), .C2(n13368), .ZN(P2_U3301) );
  XNOR2_X1 U13333 ( .A(n10750), .B(n11140), .ZN(n10751) );
  OAI222_X1 U13334 ( .A1(n15096), .A2(n12619), .B1(n15072), .B2(n12173), .C1(
        n10751), .C2(n15075), .ZN(n14367) );
  INV_X1 U13335 ( .A(n14367), .ZN(n10758) );
  OAI21_X1 U13336 ( .B1(n10754), .B2(n10753), .A(n10752), .ZN(n14369) );
  AOI22_X1 U13337 ( .A1(n15068), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n15102), 
        .B2(n12111), .ZN(n10755) );
  OAI21_X1 U13338 ( .B1(n15049), .B2(n14366), .A(n10755), .ZN(n10756) );
  AOI21_X1 U13339 ( .B1(n14369), .B2(n15065), .A(n10756), .ZN(n10757) );
  OAI21_X1 U13340 ( .B1(n10758), .B2(n15068), .A(n10757), .ZN(P3_U3221) );
  OR2_X1 U13341 ( .A1(n10760), .A2(n10759), .ZN(n10761) );
  NAND2_X1 U13342 ( .A1(n10762), .A2(n10761), .ZN(n10823) );
  AOI21_X1 U13343 ( .B1(n10763), .B2(n13550), .A(n13980), .ZN(n10765) );
  NAND2_X1 U13344 ( .A1(n10765), .A2(n10764), .ZN(n10821) );
  OAI22_X1 U13345 ( .A1(n6464), .A2(n9445), .B1(n13448), .B2(n14599), .ZN(
        n10766) );
  AOI21_X1 U13346 ( .B1(n13550), .B2(n14601), .A(n10766), .ZN(n10767) );
  OAI21_X1 U13347 ( .B1(n10821), .B2(n14035), .A(n10767), .ZN(n10777) );
  INV_X1 U13348 ( .A(n10768), .ZN(n10769) );
  NOR2_X1 U13349 ( .A1(n13685), .A2(n10769), .ZN(n10770) );
  AOI21_X1 U13350 ( .B1(n10771), .B2(n10770), .A(n14629), .ZN(n10772) );
  NAND2_X1 U13351 ( .A1(n10773), .A2(n10772), .ZN(n10825) );
  OR2_X1 U13352 ( .A1(n14428), .A2(n14615), .ZN(n10775) );
  NAND2_X1 U13353 ( .A1(n13722), .A2(n14683), .ZN(n10774) );
  NAND2_X1 U13354 ( .A1(n10775), .A2(n10774), .ZN(n13446) );
  INV_X1 U13355 ( .A(n13446), .ZN(n10820) );
  AOI21_X1 U13356 ( .B1(n10825), .B2(n10820), .A(n14016), .ZN(n10776) );
  AOI211_X1 U13357 ( .C1(n14624), .C2(n10823), .A(n10777), .B(n10776), .ZN(
        n10778) );
  INV_X1 U13358 ( .A(n10778), .ZN(P1_U3280) );
  INV_X1 U13359 ( .A(n15028), .ZN(n10788) );
  AOI21_X1 U13360 ( .B1(n10780), .B2(n10779), .A(n12219), .ZN(n10782) );
  NAND2_X1 U13361 ( .A1(n10782), .A2(n10781), .ZN(n10787) );
  INV_X1 U13362 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15363) );
  NOR2_X1 U13363 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15363), .ZN(n14971) );
  AOI21_X1 U13364 ( .B1(n12189), .B2(n15024), .A(n14971), .ZN(n10783) );
  OAI21_X1 U13365 ( .B1(n12187), .B2(n12173), .A(n10783), .ZN(n10784) );
  AOI21_X1 U13366 ( .B1(n10785), .B2(n12193), .A(n10784), .ZN(n10786) );
  OAI211_X1 U13367 ( .C1(n10788), .C2(n12191), .A(n10787), .B(n10786), .ZN(
        P3_U3157) );
  INV_X1 U13368 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14444) );
  OAI21_X1 U13369 ( .B1(n14444), .B2(n10790), .A(n10789), .ZN(n10791) );
  XNOR2_X1 U13370 ( .A(n10791), .B(n14552), .ZN(n14546) );
  NAND2_X1 U13371 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14546), .ZN(n14544) );
  INV_X1 U13372 ( .A(n14552), .ZN(n11282) );
  NAND2_X1 U13373 ( .A1(n10791), .A2(n11282), .ZN(n10792) );
  NAND2_X1 U13374 ( .A1(n14544), .A2(n10792), .ZN(n10793) );
  INV_X1 U13375 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n11230) );
  XNOR2_X1 U13376 ( .A(n10793), .B(n11230), .ZN(n10805) );
  INV_X1 U13377 ( .A(n10805), .ZN(n10803) );
  NAND2_X1 U13378 ( .A1(n11269), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10798) );
  INV_X1 U13379 ( .A(n10794), .ZN(n10795) );
  NAND2_X1 U13380 ( .A1(n10796), .A2(n10795), .ZN(n10797) );
  NAND2_X1 U13381 ( .A1(n10798), .A2(n10797), .ZN(n10799) );
  XNOR2_X1 U13382 ( .A(n10799), .B(n14552), .ZN(n14549) );
  NAND2_X1 U13383 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14549), .ZN(n14547) );
  NAND2_X1 U13384 ( .A1(n10799), .A2(n11282), .ZN(n10800) );
  NAND2_X1 U13385 ( .A1(n14547), .A2(n10800), .ZN(n10801) );
  XOR2_X1 U13386 ( .A(n10801), .B(P1_REG2_REG_19__SCAN_IN), .Z(n10804) );
  OAI21_X1 U13387 ( .B1(n10804), .B2(n14536), .A(n14553), .ZN(n10802) );
  AOI21_X1 U13388 ( .B1(n10803), .B2(n14545), .A(n10802), .ZN(n10807) );
  AOI22_X1 U13389 ( .A1(n10805), .A2(n14545), .B1(n14548), .B2(n10804), .ZN(
        n10806) );
  MUX2_X1 U13390 ( .A(n10807), .B(n10806), .S(n14614), .Z(n10808) );
  NAND2_X1 U13391 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13401)
         );
  OAI211_X1 U13392 ( .C1(n10809), .C2(n14557), .A(n10808), .B(n13401), .ZN(
        P1_U3262) );
  NAND2_X1 U13393 ( .A1(n10810), .A2(n14708), .ZN(n10812) );
  AND3_X1 U13394 ( .A1(n10813), .A2(n10812), .A3(n10811), .ZN(n10816) );
  INV_X1 U13395 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10814) );
  MUX2_X1 U13396 ( .A(n10816), .B(n10814), .S(n14713), .Z(n10815) );
  OAI21_X1 U13397 ( .B1(n10819), .B2(n14209), .A(n10815), .ZN(P1_U3495) );
  MUX2_X1 U13398 ( .A(n10817), .B(n10816), .S(n14730), .Z(n10818) );
  OAI21_X1 U13399 ( .B1(n10819), .B2(n14155), .A(n10818), .ZN(P1_U3540) );
  INV_X1 U13400 ( .A(n13550), .ZN(n10831) );
  NAND2_X1 U13401 ( .A1(n10821), .A2(n10820), .ZN(n10822) );
  AOI21_X1 U13402 ( .B1(n10823), .B2(n14708), .A(n10822), .ZN(n10824) );
  AND2_X1 U13403 ( .A1(n10825), .A2(n10824), .ZN(n10828) );
  INV_X1 U13404 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10826) );
  MUX2_X1 U13405 ( .A(n10828), .B(n10826), .S(n14713), .Z(n10827) );
  OAI21_X1 U13406 ( .B1(n10831), .B2(n14209), .A(n10827), .ZN(P1_U3498) );
  MUX2_X1 U13407 ( .A(n10829), .B(n10828), .S(n14730), .Z(n10830) );
  OAI21_X1 U13408 ( .B1(n10831), .B2(n14155), .A(n10830), .ZN(P1_U3541) );
  AOI22_X1 U13409 ( .A1(n11507), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n11506), 
        .B2(n14764), .ZN(n10833) );
  XNOR2_X1 U13410 ( .A(n13331), .B(n12883), .ZN(n12022) );
  XNOR2_X1 U13411 ( .A(n10876), .B(n12022), .ZN(n13336) );
  OAI22_X1 U13412 ( .A1(n13228), .A2(n10835), .B1(n11655), .B2(n13232), .ZN(
        n10850) );
  NAND2_X1 U13413 ( .A1(n10839), .A2(n10838), .ZN(n10880) );
  INV_X1 U13414 ( .A(n12022), .ZN(n10875) );
  XNOR2_X1 U13415 ( .A(n10840), .B(n10875), .ZN(n10846) );
  NAND2_X1 U13416 ( .A1(n11958), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n10845) );
  INV_X1 U13417 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12942) );
  OR2_X1 U13418 ( .A1(n11962), .A2(n12942), .ZN(n10844) );
  INV_X1 U13419 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n12811) );
  XNOR2_X1 U13420 ( .A(n10887), .B(n12811), .ZN(n12812) );
  OR2_X1 U13421 ( .A1(n11741), .A2(n12812), .ZN(n10843) );
  INV_X1 U13422 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10841) );
  OR2_X1 U13423 ( .A1(n11743), .A2(n10841), .ZN(n10842) );
  NAND4_X1 U13424 ( .A1(n10845), .A2(n10844), .A3(n10843), .A4(n10842), .ZN(
        n12882) );
  INV_X1 U13425 ( .A(n12882), .ZN(n13023) );
  OAI22_X1 U13426 ( .A1(n11868), .A2(n12775), .B1(n13023), .B2(n12988), .ZN(
        n11653) );
  AOI21_X1 U13427 ( .B1(n10846), .B2(n13251), .A(n11653), .ZN(n13335) );
  AOI21_X1 U13428 ( .B1(n13331), .B2(n10847), .A(n6800), .ZN(n13333) );
  NAND2_X1 U13429 ( .A1(n13333), .A2(n11702), .ZN(n10848) );
  AOI21_X1 U13430 ( .B1(n13335), .B2(n10848), .A(n6466), .ZN(n10849) );
  AOI211_X1 U13431 ( .C1(n13248), .C2(n13331), .A(n10850), .B(n10849), .ZN(
        n10851) );
  OAI21_X1 U13432 ( .B1(n13239), .B2(n13336), .A(n10851), .ZN(P2_U3250) );
  OAI22_X1 U13433 ( .A1(n6480), .A2(n10853), .B1(n10852), .B2(n15131), .ZN(
        n10855) );
  NAND2_X1 U13434 ( .A1(n10855), .A2(n10854), .ZN(n10856) );
  NAND2_X1 U13435 ( .A1(n10856), .A2(n6477), .ZN(n10859) );
  AOI21_X1 U13436 ( .B1(n10859), .B2(n10858), .A(n10857), .ZN(n10866) );
  NAND2_X1 U13437 ( .A1(n10861), .A2(n10860), .ZN(n10862) );
  AND2_X1 U13438 ( .A1(n10863), .A2(n10862), .ZN(n10865) );
  AOI21_X1 U13439 ( .B1(n10868), .B2(n15160), .A(n10867), .ZN(n10871) );
  MUX2_X1 U13440 ( .A(n10869), .B(n10871), .S(n15181), .Z(n10870) );
  OAI21_X1 U13441 ( .B1(n12705), .B2(n10874), .A(n10870), .ZN(P3_U3470) );
  INV_X1 U13442 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n10872) );
  MUX2_X1 U13443 ( .A(n10872), .B(n10871), .S(n15164), .Z(n10873) );
  OAI21_X1 U13444 ( .B1(n12757), .B2(n10874), .A(n10873), .ZN(P3_U3423) );
  INV_X1 U13445 ( .A(n13331), .ZN(n10881) );
  AOI22_X1 U13446 ( .A1(n11507), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n11506), 
        .B2(n14773), .ZN(n10877) );
  XNOR2_X1 U13447 ( .A(n13328), .B(n13023), .ZN(n12020) );
  NAND2_X1 U13448 ( .A1(n10879), .A2(n12020), .ZN(n13024) );
  OAI21_X1 U13449 ( .B1(n10879), .B2(n12020), .A(n13024), .ZN(n13330) );
  INV_X1 U13450 ( .A(n12020), .ZN(n10883) );
  OAI211_X1 U13451 ( .C1(n10884), .C2(n10883), .A(n12999), .B(n13251), .ZN(
        n10895) );
  INV_X1 U13452 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10885) );
  OAI21_X1 U13453 ( .B1(n10887), .B2(n12811), .A(n10885), .ZN(n10888) );
  NAND2_X1 U13454 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n10886) );
  NAND2_X1 U13455 ( .A1(n10888), .A2(n11197), .ZN(n13233) );
  OR2_X1 U13456 ( .A1(n13233), .A2(n11741), .ZN(n10892) );
  NAND2_X1 U13457 ( .A1(n11959), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n10891) );
  INV_X1 U13458 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13234) );
  OR2_X1 U13459 ( .A1(n11962), .A2(n13234), .ZN(n10890) );
  INV_X1 U13460 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n12957) );
  OR2_X1 U13461 ( .A1(n6950), .A2(n12957), .ZN(n10889) );
  NAND4_X1 U13462 ( .A1(n10892), .A2(n10891), .A3(n10890), .A4(n10889), .ZN(
        n12998) );
  NAND2_X1 U13463 ( .A1(n12998), .A2(n12858), .ZN(n10894) );
  NAND2_X1 U13464 ( .A1(n12883), .A2(n13020), .ZN(n10893) );
  AND2_X1 U13465 ( .A1(n10894), .A2(n10893), .ZN(n12810) );
  NAND2_X1 U13466 ( .A1(n10895), .A2(n12810), .ZN(n13326) );
  NAND2_X1 U13467 ( .A1(n13326), .A2(n13228), .ZN(n10900) );
  AOI211_X1 U13468 ( .C1(n13328), .C2(n10896), .A(n13243), .B(n7151), .ZN(
        n13327) );
  NOR2_X1 U13469 ( .A1(n7498), .A2(n13231), .ZN(n10898) );
  OAI22_X1 U13470 ( .A1(n13155), .A2(n12942), .B1(n12812), .B2(n13232), .ZN(
        n10897) );
  AOI211_X1 U13471 ( .C1(n13327), .C2(n13245), .A(n10898), .B(n10897), .ZN(
        n10899) );
  OAI211_X1 U13472 ( .C1(n13330), .C2(n13239), .A(n10900), .B(n10899), .ZN(
        P2_U3249) );
  INV_X1 U13473 ( .A(n10901), .ZN(n10902) );
  NAND2_X1 U13474 ( .A1(n13474), .A2(n10902), .ZN(n10903) );
  NAND2_X1 U13475 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14514)
         );
  OAI211_X1 U13476 ( .C1(n10904), .C2(n13462), .A(n10903), .B(n14514), .ZN(
        n10922) );
  AND2_X1 U13477 ( .A1(n11367), .A2(n13722), .ZN(n10905) );
  AOI21_X1 U13478 ( .B1(n13538), .B2(n11436), .A(n10905), .ZN(n11238) );
  NAND2_X1 U13479 ( .A1(n13538), .A2(n11422), .ZN(n10907) );
  NAND2_X1 U13480 ( .A1(n13722), .A2(n11436), .ZN(n10906) );
  NAND2_X1 U13481 ( .A1(n10907), .A2(n10906), .ZN(n10908) );
  XNOR2_X1 U13482 ( .A(n10908), .B(n11477), .ZN(n11240) );
  XOR2_X1 U13483 ( .A(n11238), .B(n11240), .Z(n10920) );
  AND2_X1 U13484 ( .A1(n11367), .A2(n13723), .ZN(n10909) );
  AOI21_X1 U13485 ( .B1(n14416), .B2(n11234), .A(n10909), .ZN(n10913) );
  INV_X1 U13486 ( .A(n10913), .ZN(n10918) );
  NAND2_X1 U13487 ( .A1(n14416), .A2(n11422), .ZN(n10911) );
  NAND2_X1 U13488 ( .A1(n13723), .A2(n11234), .ZN(n10910) );
  NAND2_X1 U13489 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  XNOR2_X1 U13490 ( .A(n10912), .B(n11477), .ZN(n10917) );
  XNOR2_X1 U13491 ( .A(n10917), .B(n10913), .ZN(n14406) );
  INV_X1 U13492 ( .A(n10914), .ZN(n10915) );
  NAND2_X1 U13493 ( .A1(n10916), .A2(n10915), .ZN(n14407) );
  NAND3_X1 U13494 ( .A1(n14408), .A2(n14406), .A3(n14407), .ZN(n14411) );
  OAI21_X1 U13495 ( .B1(n10918), .B2(n10917), .A(n14411), .ZN(n10919) );
  AOI211_X1 U13496 ( .C1(n10920), .C2(n10919), .A(n14410), .B(n11239), .ZN(
        n10921) );
  AOI211_X1 U13497 ( .C1(n13538), .C2(n14415), .A(n10922), .B(n10921), .ZN(
        n10923) );
  INV_X1 U13498 ( .A(n10923), .ZN(P1_U3224) );
  OR2_X1 U13499 ( .A1(n14445), .A2(n14428), .ZN(n13548) );
  NAND2_X1 U13500 ( .A1(n14445), .A2(n14428), .ZN(n13549) );
  NAND2_X1 U13501 ( .A1(n10926), .A2(n6468), .ZN(n10929) );
  AOI22_X1 U13502 ( .A1(n11284), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11283), 
        .B2(n10927), .ZN(n10928) );
  INV_X1 U13503 ( .A(n14447), .ZN(n14374) );
  NAND2_X1 U13504 ( .A1(n14145), .A2(n14374), .ZN(n13563) );
  NAND2_X1 U13505 ( .A1(n13562), .A2(n13563), .ZN(n13688) );
  XNOR2_X1 U13506 ( .A(n11614), .B(n11597), .ZN(n14146) );
  INV_X1 U13507 ( .A(n14146), .ZN(n10944) );
  XNOR2_X1 U13508 ( .A(n11598), .B(n11597), .ZN(n14151) );
  NAND2_X1 U13509 ( .A1(n14145), .A2(n6616), .ZN(n10931) );
  NAND2_X1 U13510 ( .A1(n10931), .A2(n14604), .ZN(n10932) );
  OR2_X1 U13511 ( .A1(n10932), .A2(n14025), .ZN(n14149) );
  AND2_X1 U13512 ( .A1(n10934), .A2(n10933), .ZN(n10935) );
  OR2_X1 U13513 ( .A1(n10935), .A2(n11272), .ZN(n14393) );
  INV_X1 U13514 ( .A(n9589), .ZN(n11631) );
  AOI22_X1 U13515 ( .A1(n11483), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11631), 
        .B2(P1_REG1_REG_16__SCAN_IN), .ZN(n10937) );
  NAND2_X1 U13516 ( .A1(n11632), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n10936) );
  OAI211_X1 U13517 ( .C1(n14393), .C2(n9585), .A(n10937), .B(n10936), .ZN(
        n14437) );
  OAI22_X1 U13518 ( .A1(n6464), .A2(n10726), .B1(n14435), .B2(n14599), .ZN(
        n10939) );
  NOR2_X1 U13519 ( .A1(n14029), .A2(n14428), .ZN(n10938) );
  AOI211_X1 U13520 ( .C1(n14032), .C2(n14437), .A(n10939), .B(n10938), .ZN(
        n10941) );
  NAND2_X1 U13521 ( .A1(n14145), .A2(n14601), .ZN(n10940) );
  OAI211_X1 U13522 ( .C1(n14149), .C2(n14035), .A(n10941), .B(n10940), .ZN(
        n10942) );
  AOI21_X1 U13523 ( .B1(n14151), .B2(n14624), .A(n10942), .ZN(n10943) );
  OAI21_X1 U13524 ( .B1(n10944), .B2(n14038), .A(n10943), .ZN(P1_U3278) );
  INV_X1 U13525 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11374) );
  OAI222_X1 U13526 ( .A1(n14223), .A2(n11374), .B1(n14221), .B2(n10945), .C1(
        n9095), .C2(P1_U3086), .ZN(P1_U3331) );
  NAND2_X1 U13527 ( .A1(n10947), .A2(n10946), .ZN(n14627) );
  INV_X1 U13528 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10950) );
  NOR2_X1 U13529 ( .A1(n10949), .A2(n10948), .ZN(n11165) );
  AOI22_X1 U13530 ( .A1(n14627), .A2(n10950), .B1(n11165), .B2(n9095), .ZN(
        P1_U3445) );
  INV_X1 U13531 ( .A(n11071), .ZN(n11067) );
  INV_X1 U13532 ( .A(n10951), .ZN(n11028) );
  INV_X1 U13533 ( .A(n11015), .ZN(n10953) );
  INV_X1 U13534 ( .A(n10956), .ZN(n10952) );
  MUX2_X1 U13535 ( .A(n10953), .B(n10952), .S(n11093), .Z(n10954) );
  NOR2_X1 U13536 ( .A1(n14352), .A2(n10954), .ZN(n11019) );
  NAND2_X1 U13537 ( .A1(n10956), .A2(n10955), .ZN(n10958) );
  AOI21_X1 U13538 ( .B1(n11019), .B2(n10958), .A(n10957), .ZN(n11022) );
  INV_X1 U13539 ( .A(n10959), .ZN(n10961) );
  NAND2_X1 U13540 ( .A1(n10961), .A2(n11160), .ZN(n10964) );
  NAND2_X1 U13541 ( .A1(n10961), .A2(n10960), .ZN(n10962) );
  NAND3_X1 U13542 ( .A1(n10968), .A2(n6476), .A3(n10962), .ZN(n10963) );
  OAI21_X1 U13543 ( .B1(n15090), .B2(n10964), .A(n10963), .ZN(n10967) );
  NAND2_X1 U13544 ( .A1(n15088), .A2(n10965), .ZN(n10966) );
  NAND2_X1 U13545 ( .A1(n10967), .A2(n10966), .ZN(n10971) );
  MUX2_X1 U13546 ( .A(n10969), .B(n10968), .S(n11093), .Z(n10970) );
  NAND3_X1 U13547 ( .A1(n10971), .A2(n15074), .A3(n10970), .ZN(n10978) );
  NAND2_X1 U13548 ( .A1(n10979), .A2(n10972), .ZN(n10975) );
  NAND2_X1 U13549 ( .A1(n10980), .A2(n10973), .ZN(n10974) );
  MUX2_X1 U13550 ( .A(n10975), .B(n10974), .S(n11093), .Z(n10976) );
  INV_X1 U13551 ( .A(n10976), .ZN(n10977) );
  NAND2_X1 U13552 ( .A1(n10978), .A2(n10977), .ZN(n10982) );
  MUX2_X1 U13553 ( .A(n10980), .B(n10979), .S(n11093), .Z(n10981) );
  NAND3_X1 U13554 ( .A1(n10982), .A2(n11131), .A3(n10981), .ZN(n10986) );
  MUX2_X1 U13555 ( .A(n10984), .B(n10983), .S(n6477), .Z(n10985) );
  NAND3_X1 U13556 ( .A1(n10986), .A2(n11130), .A3(n10985), .ZN(n10993) );
  NAND2_X1 U13557 ( .A1(n10994), .A2(n10987), .ZN(n10990) );
  NAND2_X1 U13558 ( .A1(n10995), .A2(n10988), .ZN(n10989) );
  MUX2_X1 U13559 ( .A(n10990), .B(n10989), .S(n11093), .Z(n10991) );
  INV_X1 U13560 ( .A(n10991), .ZN(n10992) );
  NAND2_X1 U13561 ( .A1(n10993), .A2(n10992), .ZN(n10997) );
  MUX2_X1 U13562 ( .A(n10995), .B(n10994), .S(n11093), .Z(n10996) );
  MUX2_X1 U13563 ( .A(n10999), .B(n10998), .S(n11093), .Z(n11000) );
  NAND3_X1 U13564 ( .A1(n11001), .A2(n11129), .A3(n11000), .ZN(n11005) );
  INV_X1 U13565 ( .A(n15042), .ZN(n11138) );
  MUX2_X1 U13566 ( .A(n11003), .B(n11002), .S(n6476), .Z(n11004) );
  NAND3_X1 U13567 ( .A1(n11005), .A2(n11138), .A3(n11004), .ZN(n11009) );
  NAND2_X1 U13568 ( .A1(n15024), .A2(n15048), .ZN(n11007) );
  NAND2_X1 U13569 ( .A1(n8297), .A2(n15152), .ZN(n11006) );
  MUX2_X1 U13570 ( .A(n11007), .B(n11006), .S(n11093), .Z(n11008) );
  NAND2_X1 U13571 ( .A1(n11009), .A2(n11008), .ZN(n11010) );
  INV_X1 U13572 ( .A(n15022), .ZN(n15015) );
  NAND2_X1 U13573 ( .A1(n11010), .A2(n15015), .ZN(n11013) );
  AND3_X1 U13574 ( .A1(n11013), .A2(n11137), .A3(n11011), .ZN(n11018) );
  NAND3_X1 U13575 ( .A1(n11013), .A2(n11137), .A3(n11012), .ZN(n11016) );
  NAND3_X1 U13576 ( .A1(n11016), .A2(n11015), .A3(n11014), .ZN(n11017) );
  NAND2_X1 U13577 ( .A1(n11020), .A2(n11019), .ZN(n11021) );
  OAI211_X1 U13578 ( .C1(n11093), .C2(n11022), .A(n11021), .B(n12629), .ZN(
        n11029) );
  INV_X1 U13579 ( .A(n12611), .ZN(n12607) );
  AOI21_X1 U13580 ( .B1(n11029), .B2(n11023), .A(n12607), .ZN(n11026) );
  NAND2_X1 U13581 ( .A1(n11036), .A2(n11024), .ZN(n11025) );
  OAI21_X1 U13582 ( .B1(n11026), .B2(n11025), .A(n6476), .ZN(n11033) );
  OAI22_X1 U13583 ( .A1(n11029), .A2(n11028), .B1(n6477), .B2(n11027), .ZN(
        n11030) );
  NAND2_X1 U13584 ( .A1(n11030), .A2(n12611), .ZN(n11032) );
  INV_X1 U13585 ( .A(n11035), .ZN(n11031) );
  AOI21_X1 U13586 ( .B1(n11033), .B2(n11032), .A(n11031), .ZN(n11038) );
  AOI21_X1 U13587 ( .B1(n11035), .B2(n11034), .A(n6476), .ZN(n11037) );
  OAI22_X1 U13588 ( .A1(n11038), .A2(n11037), .B1(n6476), .B2(n11036), .ZN(
        n11039) );
  NAND3_X1 U13589 ( .A1(n11039), .A2(n12565), .A3(n12587), .ZN(n11050) );
  INV_X1 U13590 ( .A(n11044), .ZN(n11042) );
  OAI211_X1 U13591 ( .C1(n11042), .C2(n11041), .A(n11052), .B(n11040), .ZN(
        n11047) );
  NAND2_X1 U13592 ( .A1(n12565), .A2(n11043), .ZN(n11045) );
  NAND3_X1 U13593 ( .A1(n11045), .A2(n12537), .A3(n11044), .ZN(n11046) );
  MUX2_X1 U13594 ( .A(n11047), .B(n11046), .S(n6477), .Z(n11048) );
  INV_X1 U13595 ( .A(n11048), .ZN(n11049) );
  NAND2_X1 U13596 ( .A1(n11050), .A2(n11049), .ZN(n11055) );
  INV_X1 U13597 ( .A(n12538), .ZN(n11054) );
  MUX2_X1 U13598 ( .A(n12537), .B(n11052), .S(n6477), .Z(n11053) );
  NAND3_X1 U13599 ( .A1(n11055), .A2(n11054), .A3(n11053), .ZN(n11059) );
  MUX2_X1 U13600 ( .A(n11057), .B(n11056), .S(n11093), .Z(n11058) );
  MUX2_X1 U13601 ( .A(n11061), .B(n11060), .S(n11093), .Z(n11062) );
  NAND3_X1 U13602 ( .A1(n11063), .A2(n12511), .A3(n11062), .ZN(n11070) );
  NAND4_X1 U13603 ( .A1(n11065), .A2(n11064), .A3(n12499), .A4(n11070), .ZN(
        n11066) );
  OAI21_X1 U13604 ( .B1(n12486), .B2(n11072), .A(n11071), .ZN(n11073) );
  INV_X1 U13605 ( .A(n11075), .ZN(n11076) );
  NOR2_X1 U13606 ( .A1(n12451), .A2(n11076), .ZN(n11079) );
  INV_X1 U13607 ( .A(n11077), .ZN(n11078) );
  AOI21_X1 U13608 ( .B1(n11085), .B2(n11079), .A(n11078), .ZN(n11087) );
  INV_X1 U13609 ( .A(n11080), .ZN(n11081) );
  NOR2_X1 U13610 ( .A1(n12451), .A2(n11081), .ZN(n11084) );
  INV_X1 U13611 ( .A(n11082), .ZN(n11083) );
  AOI21_X1 U13612 ( .B1(n11085), .B2(n11084), .A(n11083), .ZN(n11086) );
  MUX2_X1 U13613 ( .A(n11087), .B(n11086), .S(n11093), .Z(n11088) );
  INV_X1 U13614 ( .A(n12433), .ZN(n12439) );
  AOI21_X1 U13615 ( .B1(n12719), .B2(n12425), .A(n11094), .ZN(n11092) );
  NAND2_X1 U13616 ( .A1(n11089), .A2(n11093), .ZN(n11090) );
  OAI211_X1 U13617 ( .C1(n11092), .C2(n8189), .A(n11091), .B(n11090), .ZN(
        n11096) );
  NAND3_X1 U13618 ( .A1(n11094), .A2(n11093), .A3(n12421), .ZN(n11095) );
  NAND3_X1 U13619 ( .A1(n11096), .A2(n11123), .A3(n11095), .ZN(n11104) );
  INV_X1 U13620 ( .A(n11097), .ZN(n11098) );
  INV_X1 U13621 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12049) );
  INV_X1 U13622 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11952) );
  XNOR2_X1 U13623 ( .A(n11952), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11105) );
  XNOR2_X1 U13624 ( .A(n11106), .B(n11105), .ZN(n12045) );
  NAND2_X1 U13625 ( .A1(n12045), .A2(n11108), .ZN(n11102) );
  INV_X1 U13626 ( .A(SI_30_), .ZN(n12047) );
  OR2_X1 U13627 ( .A1(n11100), .A2(n12047), .ZN(n11101) );
  NAND2_X1 U13628 ( .A1(n11102), .A2(n11101), .ZN(n12637) );
  AND2_X1 U13629 ( .A1(n12713), .A2(n12221), .ZN(n11149) );
  INV_X1 U13630 ( .A(n11149), .ZN(n11103) );
  NAND3_X1 U13631 ( .A1(n11104), .A2(n11125), .A3(n11103), .ZN(n11120) );
  INV_X1 U13632 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14219) );
  XNOR2_X1 U13633 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11107) );
  OR2_X1 U13634 ( .A1(n7010), .A2(n15357), .ZN(n11109) );
  NAND2_X1 U13635 ( .A1(n6481), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U13636 ( .A1(n6479), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11112) );
  NAND2_X1 U13637 ( .A1(n7806), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n11111) );
  AND3_X1 U13638 ( .A1(n11113), .A2(n11112), .A3(n11111), .ZN(n11114) );
  OR2_X1 U13639 ( .A1(n12633), .A2(n11119), .ZN(n11118) );
  INV_X1 U13640 ( .A(n12221), .ZN(n11116) );
  NAND2_X1 U13641 ( .A1(n12637), .A2(n11116), .ZN(n11117) );
  NAND2_X1 U13642 ( .A1(n11118), .A2(n11117), .ZN(n11150) );
  INV_X1 U13643 ( .A(n11121), .ZN(n15103) );
  INV_X1 U13644 ( .A(n11122), .ZN(n11126) );
  OAI21_X1 U13645 ( .B1(n12713), .B2(n12407), .A(n11123), .ZN(n11124) );
  NAND4_X1 U13646 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11136) );
  NAND3_X1 U13647 ( .A1(n15074), .A2(n11132), .A3(n11131), .ZN(n11135) );
  NOR4_X1 U13648 ( .A1(n11136), .A2(n11135), .A3(n7833), .A4(n11134), .ZN(
        n11139) );
  NAND4_X1 U13649 ( .A1(n11139), .A2(n15015), .A3(n11138), .A4(n11137), .ZN(
        n11141) );
  NOR4_X1 U13650 ( .A1(n12607), .A2(n11141), .A3(n14352), .A4(n11140), .ZN(
        n11142) );
  NAND4_X1 U13651 ( .A1(n12587), .A2(n12629), .A3(n11142), .A4(n12600), .ZN(
        n11143) );
  NOR4_X1 U13652 ( .A1(n12538), .A2(n12561), .A3(n12552), .A4(n11143), .ZN(
        n11144) );
  NAND4_X1 U13653 ( .A1(n12499), .A2(n12511), .A3(n12524), .A4(n11144), .ZN(
        n11145) );
  NOR4_X1 U13654 ( .A1(n12451), .A2(n12467), .A3(n12486), .A4(n11145), .ZN(
        n11146) );
  NAND4_X1 U13655 ( .A1(n11147), .A2(n12421), .A3(n11146), .A4(n12433), .ZN(
        n11148) );
  NAND3_X1 U13656 ( .A1(n11158), .A2(n11157), .A3(n12369), .ZN(n11159) );
  OAI211_X1 U13657 ( .C1(n11160), .C2(n11162), .A(n11159), .B(P3_B_REG_SCAN_IN), .ZN(n11161) );
  OAI21_X1 U13658 ( .B1(n11163), .B2(n11162), .A(n11161), .ZN(P3_U3296) );
  OAI222_X1 U13659 ( .A1(n14223), .A2(n11395), .B1(n14221), .B2(n11164), .C1(
        n9097), .C2(P1_U3086), .ZN(P1_U3330) );
  INV_X1 U13660 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U13661 ( .A1(n14627), .A2(n11166), .B1(n11165), .B2(n9097), .ZN(
        P1_U3446) );
  INV_X1 U13662 ( .A(n11167), .ZN(n11168) );
  INV_X1 U13663 ( .A(n11170), .ZN(n11171) );
  NAND2_X1 U13664 ( .A1(n11171), .A2(SI_26_), .ZN(n11172) );
  MUX2_X1 U13665 ( .A(n14222), .B(n13367), .S(n11332), .Z(n11173) );
  XNOR2_X1 U13666 ( .A(n11173), .B(SI_27_), .ZN(n11443) );
  INV_X1 U13667 ( .A(n11173), .ZN(n11174) );
  NAND2_X1 U13668 ( .A1(n11174), .A2(SI_27_), .ZN(n11175) );
  MUX2_X1 U13669 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n11332), .Z(n11177) );
  XNOR2_X1 U13670 ( .A(n11177), .B(SI_28_), .ZN(n11465) );
  INV_X1 U13671 ( .A(n11177), .ZN(n11178) );
  NAND2_X1 U13672 ( .A1(n11178), .A2(n15243), .ZN(n11179) );
  INV_X1 U13673 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11649) );
  MUX2_X1 U13674 ( .A(n11649), .B(n12049), .S(n11332), .Z(n11180) );
  XNOR2_X1 U13675 ( .A(n11180), .B(SI_29_), .ZN(n11610) );
  MUX2_X1 U13676 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n11332), .Z(n11919) );
  XNOR2_X1 U13677 ( .A(n11919), .B(SI_30_), .ZN(n11921) );
  INV_X1 U13678 ( .A(n11921), .ZN(n11181) );
  INV_X1 U13679 ( .A(n13635), .ZN(n14218) );
  OAI222_X1 U13680 ( .A1(n13366), .A2(n14218), .B1(P2_U3088), .B2(n7022), .C1(
        n11952), .C2(n13368), .ZN(P2_U3297) );
  INV_X1 U13681 ( .A(n11182), .ZN(n11183) );
  OAI222_X1 U13682 ( .A1(n12770), .A2(n11183), .B1(n8212), .B2(P3_U3151), .C1(
        n15243), .C2(n12771), .ZN(P3_U3267) );
  XNOR2_X1 U13683 ( .A(n13331), .B(n11736), .ZN(n11189) );
  OR2_X1 U13684 ( .A1(n11187), .A2(n11702), .ZN(n11188) );
  AND2_X1 U13685 ( .A1(n11190), .A2(n11189), .ZN(n11191) );
  XNOR2_X1 U13686 ( .A(n13328), .B(n11736), .ZN(n11208) );
  NAND2_X1 U13687 ( .A1(n12882), .A2(n9668), .ZN(n11192) );
  XNOR2_X1 U13688 ( .A(n11208), .B(n11192), .ZN(n12806) );
  INV_X1 U13689 ( .A(n11192), .ZN(n11193) );
  AOI22_X1 U13690 ( .A1(n11507), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n11506), 
        .B2(n14789), .ZN(n11195) );
  XNOR2_X1 U13691 ( .A(n13323), .B(n11736), .ZN(n11500) );
  NAND2_X1 U13692 ( .A1(n12998), .A2(n9668), .ZN(n11498) );
  XNOR2_X1 U13693 ( .A(n11500), .B(n11498), .ZN(n11209) );
  AND2_X1 U13694 ( .A1(n11197), .A2(n12960), .ZN(n11198) );
  OR2_X1 U13695 ( .A1(n11198), .A2(n11510), .ZN(n13214) );
  INV_X1 U13696 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n11199) );
  OR2_X1 U13697 ( .A1(n6950), .A2(n11199), .ZN(n11202) );
  INV_X1 U13698 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n11200) );
  OR2_X1 U13699 ( .A1(n11743), .A2(n11200), .ZN(n11201) );
  AND2_X1 U13700 ( .A1(n11202), .A2(n11201), .ZN(n11204) );
  INV_X1 U13701 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13215) );
  OR2_X1 U13702 ( .A1(n11962), .A2(n13215), .ZN(n11203) );
  OAI211_X1 U13703 ( .C1(n13214), .C2(n11741), .A(n11204), .B(n11203), .ZN(
        n13000) );
  AOI22_X1 U13704 ( .A1(n13000), .A2(n12858), .B1(n12882), .B2(n13020), .ZN(
        n13225) );
  INV_X1 U13705 ( .A(n13225), .ZN(n11205) );
  AOI22_X1 U13706 ( .A1(n12871), .A2(n11205), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11206) );
  OAI21_X1 U13707 ( .B1(n13233), .B2(n12873), .A(n11206), .ZN(n11213) );
  INV_X1 U13708 ( .A(n11207), .ZN(n11211) );
  AOI22_X1 U13709 ( .A1(n11208), .A2(n12808), .B1(n11651), .B2(n12882), .ZN(
        n11210) );
  NOR3_X1 U13710 ( .A1(n11211), .A2(n11210), .A3(n11209), .ZN(n11212) );
  AOI211_X1 U13711 ( .C1(n13323), .C2(n12875), .A(n11213), .B(n11212), .ZN(
        n11214) );
  OAI21_X1 U13712 ( .B1(n11502), .B2(n12877), .A(n11214), .ZN(P2_U3200) );
  AOI21_X1 U13713 ( .B1(n11217), .B2(n11216), .A(n7435), .ZN(n11223) );
  INV_X1 U13714 ( .A(n12756), .ZN(n12628) );
  INV_X1 U13715 ( .A(n11218), .ZN(n12624) );
  INV_X1 U13716 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15244) );
  NOR2_X1 U13717 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15244), .ZN(n12278) );
  NOR2_X1 U13718 ( .A1(n12619), .A2(n12213), .ZN(n11219) );
  AOI211_X1 U13719 ( .C1(n12211), .C2(n8315), .A(n12278), .B(n11219), .ZN(
        n11220) );
  OAI21_X1 U13720 ( .B1(n12624), .B2(n12191), .A(n11220), .ZN(n11221) );
  AOI21_X1 U13721 ( .B1(n12628), .B2(n12193), .A(n11221), .ZN(n11222) );
  OAI21_X1 U13722 ( .B1(n11223), .B2(n12219), .A(n11222), .ZN(P3_U3155) );
  NAND2_X1 U13723 ( .A1(n11505), .A2(n6468), .ZN(n11225) );
  AOI22_X1 U13724 ( .A1(n11284), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11283), 
        .B2(n13489), .ZN(n11224) );
  OR2_X1 U13725 ( .A1(n11289), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11226) );
  NAND2_X1 U13726 ( .A1(n11305), .A2(n11226), .ZN(n13983) );
  INV_X1 U13727 ( .A(n13983), .ZN(n13403) );
  NAND2_X1 U13728 ( .A1(n13403), .A2(n11227), .ZN(n11233) );
  NAND2_X1 U13729 ( .A1(n11632), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U13730 ( .A1(n11483), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11228) );
  OAI211_X1 U13731 ( .C1(n9589), .C2(n11230), .A(n11229), .B(n11228), .ZN(
        n11231) );
  INV_X1 U13732 ( .A(n11231), .ZN(n11232) );
  AOI22_X1 U13733 ( .A1(n13981), .A2(n11436), .B1(n11367), .B2(n13994), .ZN(
        n11301) );
  NAND2_X1 U13734 ( .A1(n13981), .A2(n11422), .ZN(n11236) );
  OR2_X1 U13735 ( .A1(n14124), .A2(n11276), .ZN(n11235) );
  NAND2_X1 U13736 ( .A1(n11236), .A2(n11235), .ZN(n11237) );
  XNOR2_X1 U13737 ( .A(n11237), .B(n11477), .ZN(n11295) );
  INV_X1 U13738 ( .A(n11295), .ZN(n11300) );
  INV_X1 U13739 ( .A(n11238), .ZN(n11241) );
  AOI22_X1 U13740 ( .A1(n13550), .A2(n11422), .B1(n11234), .B2(n14446), .ZN(
        n11242) );
  XNOR2_X1 U13741 ( .A(n11242), .B(n11477), .ZN(n11249) );
  AND2_X1 U13742 ( .A1(n11367), .A2(n14446), .ZN(n11243) );
  AOI21_X1 U13743 ( .B1(n13550), .B2(n11436), .A(n11243), .ZN(n11248) );
  XNOR2_X1 U13744 ( .A(n11249), .B(n11248), .ZN(n13449) );
  NAND2_X1 U13745 ( .A1(n14445), .A2(n11422), .ZN(n11245) );
  OR2_X1 U13746 ( .A1(n14428), .A2(n11276), .ZN(n11244) );
  NAND2_X1 U13747 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  XNOR2_X1 U13748 ( .A(n11246), .B(n11410), .ZN(n11251) );
  NOR2_X1 U13749 ( .A1(n14428), .A2(n9289), .ZN(n11247) );
  AOI21_X1 U13750 ( .B1(n14445), .B2(n11436), .A(n11247), .ZN(n11250) );
  XNOR2_X1 U13751 ( .A(n11251), .B(n11250), .ZN(n14376) );
  NOR2_X1 U13752 ( .A1(n11249), .A2(n11248), .ZN(n14377) );
  NAND2_X1 U13753 ( .A1(n14145), .A2(n9068), .ZN(n11253) );
  NAND2_X1 U13754 ( .A1(n14447), .A2(n11459), .ZN(n11252) );
  NAND2_X1 U13755 ( .A1(n11253), .A2(n11252), .ZN(n11254) );
  XNOR2_X1 U13756 ( .A(n11254), .B(n11477), .ZN(n11256) );
  AOI22_X1 U13757 ( .A1(n14145), .A2(n11436), .B1(n11367), .B2(n14447), .ZN(
        n14421) );
  AOI22_X1 U13758 ( .A1(n11284), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11283), 
        .B2(n13796), .ZN(n11259) );
  INV_X1 U13759 ( .A(n14437), .ZN(n14425) );
  OAI22_X1 U13760 ( .A1(n14205), .A2(n11276), .B1(n14425), .B2(n9289), .ZN(
        n11265) );
  NAND2_X1 U13761 ( .A1(n14390), .A2(n11422), .ZN(n11262) );
  NAND2_X1 U13762 ( .A1(n14437), .A2(n11459), .ZN(n11261) );
  NAND2_X1 U13763 ( .A1(n11262), .A2(n11261), .ZN(n11263) );
  XNOR2_X1 U13764 ( .A(n11263), .B(n11477), .ZN(n11264) );
  XOR2_X1 U13765 ( .A(n11265), .B(n11264), .Z(n14386) );
  INV_X1 U13766 ( .A(n11264), .ZN(n11267) );
  INV_X1 U13767 ( .A(n11265), .ZN(n11266) );
  NAND2_X1 U13768 ( .A1(n11268), .A2(n6468), .ZN(n11271) );
  AOI22_X1 U13769 ( .A1(n11284), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11283), 
        .B2(n11269), .ZN(n11270) );
  NOR2_X1 U13770 ( .A1(n11272), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11273) );
  OR2_X1 U13771 ( .A1(n11287), .A2(n11273), .ZN(n14403) );
  AOI22_X1 U13772 ( .A1(n11632), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n11631), 
        .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n11275) );
  OR2_X1 U13773 ( .A1(n13638), .A2(n10410), .ZN(n11274) );
  OAI211_X1 U13774 ( .C1(n14403), .C2(n9585), .A(n11275), .B(n11274), .ZN(
        n14134) );
  INV_X1 U13775 ( .A(n14134), .ZN(n14123) );
  OAI22_X1 U13776 ( .A1(n14440), .A2(n11476), .B1(n14123), .B2(n11276), .ZN(
        n11277) );
  XNOR2_X1 U13777 ( .A(n11277), .B(n11410), .ZN(n11281) );
  OR2_X1 U13778 ( .A1(n14440), .A2(n11276), .ZN(n11279) );
  NAND2_X1 U13779 ( .A1(n14134), .A2(n11367), .ZN(n11278) );
  AND2_X1 U13780 ( .A1(n11279), .A2(n11278), .ZN(n11280) );
  NAND2_X1 U13781 ( .A1(n11281), .A2(n11280), .ZN(n14394) );
  NAND2_X1 U13782 ( .A1(n11495), .A2(n6468), .ZN(n11286) );
  AOI22_X1 U13783 ( .A1(n11284), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11283), 
        .B2(n11282), .ZN(n11285) );
  OR2_X1 U13784 ( .A1(n14201), .A2(n11276), .ZN(n11293) );
  NOR2_X1 U13785 ( .A1(n11287), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11288) );
  OR2_X1 U13786 ( .A1(n11289), .A2(n11288), .ZN(n13471) );
  AOI22_X1 U13787 ( .A1(n11632), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n11631), 
        .B2(P1_REG1_REG_18__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U13788 ( .A1(n11483), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11290) );
  OAI211_X1 U13789 ( .C1(n13471), .C2(n9585), .A(n11291), .B(n11290), .ZN(
        n13720) );
  NAND2_X1 U13790 ( .A1(n13720), .A2(n11367), .ZN(n11292) );
  NAND2_X1 U13791 ( .A1(n11293), .A2(n11292), .ZN(n11297) );
  INV_X1 U13792 ( .A(n13720), .ZN(n14397) );
  OAI22_X1 U13793 ( .A1(n14201), .A2(n11476), .B1(n14397), .B2(n11276), .ZN(
        n11294) );
  XNOR2_X1 U13794 ( .A(n11294), .B(n11477), .ZN(n11296) );
  XOR2_X1 U13795 ( .A(n11297), .B(n11296), .Z(n13469) );
  XNOR2_X1 U13796 ( .A(n11295), .B(n11301), .ZN(n13399) );
  INV_X1 U13797 ( .A(n11296), .ZN(n11299) );
  INV_X1 U13798 ( .A(n11297), .ZN(n11298) );
  NAND2_X1 U13799 ( .A1(n11299), .A2(n11298), .ZN(n13397) );
  NAND2_X1 U13800 ( .A1(n11518), .A2(n6468), .ZN(n11304) );
  OR2_X1 U13801 ( .A1(n13653), .A2(n11302), .ZN(n11303) );
  INV_X1 U13802 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13439) );
  NAND2_X1 U13803 ( .A1(n11305), .A2(n13439), .ZN(n11307) );
  INV_X1 U13804 ( .A(n11319), .ZN(n11306) );
  NAND2_X1 U13805 ( .A1(n11307), .A2(n11306), .ZN(n13969) );
  OR2_X1 U13806 ( .A1(n13969), .A2(n9585), .ZN(n11312) );
  INV_X1 U13807 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n13970) );
  NAND2_X1 U13808 ( .A1(n11632), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11309) );
  NAND2_X1 U13809 ( .A1(n11631), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11308) );
  OAI211_X1 U13810 ( .C1(n13638), .C2(n13970), .A(n11309), .B(n11308), .ZN(
        n11310) );
  INV_X1 U13811 ( .A(n11310), .ZN(n11311) );
  OAI22_X1 U13812 ( .A1(n14196), .A2(n11276), .B1(n13592), .B2(n9289), .ZN(
        n11315) );
  OAI22_X1 U13813 ( .A1(n14196), .A2(n11476), .B1(n13592), .B2(n11276), .ZN(
        n11313) );
  XNOR2_X1 U13814 ( .A(n11313), .B(n11477), .ZN(n11314) );
  XOR2_X1 U13815 ( .A(n11315), .B(n11314), .Z(n13437) );
  NAND2_X1 U13816 ( .A1(n11529), .A2(n6468), .ZN(n11318) );
  OR2_X1 U13817 ( .A1(n13653), .A2(n11316), .ZN(n11317) );
  NAND2_X1 U13818 ( .A1(n13950), .A2(n11422), .ZN(n11325) );
  NAND2_X1 U13819 ( .A1(n11483), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11323) );
  INV_X1 U13820 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14189) );
  OR2_X1 U13821 ( .A1(n13639), .A2(n14189), .ZN(n11322) );
  NAND2_X1 U13822 ( .A1(n11319), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11336) );
  OAI21_X1 U13823 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n11319), .A(n11336), 
        .ZN(n13409) );
  OR2_X1 U13824 ( .A1(n9585), .A2(n13409), .ZN(n11321) );
  INV_X1 U13825 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n14108) );
  OR2_X1 U13826 ( .A1(n9589), .A2(n14108), .ZN(n11320) );
  NAND4_X1 U13827 ( .A1(n11323), .A2(n11322), .A3(n11321), .A4(n11320), .ZN(
        n13718) );
  NAND2_X1 U13828 ( .A1(n13718), .A2(n11459), .ZN(n11324) );
  NAND2_X1 U13829 ( .A1(n11325), .A2(n11324), .ZN(n11326) );
  XNOR2_X1 U13830 ( .A(n11326), .B(n11477), .ZN(n11330) );
  NAND2_X1 U13831 ( .A1(n13950), .A2(n11459), .ZN(n11328) );
  NAND2_X1 U13832 ( .A1(n11367), .A2(n13718), .ZN(n11327) );
  NAND2_X1 U13833 ( .A1(n11328), .A2(n11327), .ZN(n11329) );
  NOR2_X1 U13834 ( .A1(n11330), .A2(n11329), .ZN(n11331) );
  AOI21_X1 U13835 ( .B1(n11330), .B2(n11329), .A(n11331), .ZN(n13406) );
  INV_X1 U13836 ( .A(n11331), .ZN(n13455) );
  NAND2_X1 U13837 ( .A1(n13601), .A2(n11422), .ZN(n11343) );
  NAND2_X1 U13838 ( .A1(n11483), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11341) );
  INV_X1 U13839 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n14186) );
  OR2_X1 U13840 ( .A1(n13639), .A2(n14186), .ZN(n11340) );
  OAI21_X1 U13841 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11337), .A(n11357), 
        .ZN(n13937) );
  OR2_X1 U13842 ( .A1(n9585), .A2(n13937), .ZN(n11339) );
  INV_X1 U13843 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n14100) );
  OR2_X1 U13844 ( .A1(n6463), .A2(n14100), .ZN(n11338) );
  NAND4_X1 U13845 ( .A1(n11341), .A2(n11340), .A3(n11339), .A4(n11338), .ZN(
        n13717) );
  NAND2_X1 U13846 ( .A1(n13717), .A2(n11459), .ZN(n11342) );
  NAND2_X1 U13847 ( .A1(n11343), .A2(n11342), .ZN(n11344) );
  XNOR2_X1 U13848 ( .A(n11344), .B(n11410), .ZN(n11346) );
  AND2_X1 U13849 ( .A1(n11367), .A2(n13717), .ZN(n11345) );
  AOI21_X1 U13850 ( .B1(n13601), .B2(n11234), .A(n11345), .ZN(n11347) );
  NAND2_X1 U13851 ( .A1(n11346), .A2(n11347), .ZN(n11351) );
  INV_X1 U13852 ( .A(n11346), .ZN(n11349) );
  INV_X1 U13853 ( .A(n11347), .ZN(n11348) );
  NAND2_X1 U13854 ( .A1(n11349), .A2(n11348), .ZN(n11350) );
  NAND2_X1 U13855 ( .A1(n11351), .A2(n11350), .ZN(n13454) );
  INV_X1 U13856 ( .A(n11351), .ZN(n13378) );
  NAND2_X1 U13857 ( .A1(n11575), .A2(n6468), .ZN(n11354) );
  OR2_X1 U13858 ( .A1(n13653), .A2(n11352), .ZN(n11353) );
  NAND2_X1 U13859 ( .A1(n13918), .A2(n11422), .ZN(n11365) );
  NAND2_X1 U13860 ( .A1(n11631), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11360) );
  INV_X1 U13861 ( .A(n11357), .ZN(n11355) );
  NAND2_X1 U13862 ( .A1(n11355), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11379) );
  INV_X1 U13863 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n11356) );
  NAND2_X1 U13864 ( .A1(n11357), .A2(n11356), .ZN(n11358) );
  NAND2_X1 U13865 ( .A1(n11379), .A2(n11358), .ZN(n13919) );
  OR2_X1 U13866 ( .A1(n9585), .A2(n13919), .ZN(n11359) );
  NAND2_X1 U13867 ( .A1(n11360), .A2(n11359), .ZN(n11363) );
  INV_X1 U13868 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13920) );
  NOR2_X1 U13869 ( .A1(n13638), .A2(n13920), .ZN(n11362) );
  INV_X1 U13870 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14183) );
  NOR2_X1 U13871 ( .A1(n13639), .A2(n14183), .ZN(n11361) );
  NAND2_X1 U13872 ( .A1(n13894), .A2(n11459), .ZN(n11364) );
  NAND2_X1 U13873 ( .A1(n11365), .A2(n11364), .ZN(n11366) );
  XNOR2_X1 U13874 ( .A(n11366), .B(n11410), .ZN(n11369) );
  AND2_X1 U13875 ( .A1(n13894), .A2(n11367), .ZN(n11368) );
  AOI21_X1 U13876 ( .B1(n13918), .B2(n11234), .A(n11368), .ZN(n11370) );
  NAND2_X1 U13877 ( .A1(n11369), .A2(n11370), .ZN(n13427) );
  INV_X1 U13878 ( .A(n11369), .ZN(n11372) );
  INV_X1 U13879 ( .A(n11370), .ZN(n11371) );
  NAND2_X1 U13880 ( .A1(n11372), .A2(n11371), .ZN(n11373) );
  AND2_X1 U13881 ( .A1(n13427), .A2(n11373), .ZN(n13377) );
  NAND2_X1 U13882 ( .A1(n11663), .A2(n6468), .ZN(n11376) );
  OR2_X1 U13883 ( .A1(n13653), .A2(n11374), .ZN(n11375) );
  NAND2_X1 U13884 ( .A1(n13903), .A2(n9068), .ZN(n11386) );
  NAND2_X1 U13885 ( .A1(n11632), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11384) );
  INV_X1 U13886 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14086) );
  OR2_X1 U13887 ( .A1(n9589), .A2(n14086), .ZN(n11383) );
  INV_X1 U13888 ( .A(n11379), .ZN(n11377) );
  NAND2_X1 U13889 ( .A1(n11377), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11401) );
  INV_X1 U13890 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U13891 ( .A1(n11379), .A2(n11378), .ZN(n11380) );
  NAND2_X1 U13892 ( .A1(n11401), .A2(n11380), .ZN(n13904) );
  OR2_X1 U13893 ( .A1(n9585), .A2(n13904), .ZN(n11382) );
  INV_X1 U13894 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n13905) );
  OR2_X1 U13895 ( .A1(n13638), .A2(n13905), .ZN(n11381) );
  NAND4_X1 U13896 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n13924) );
  NAND2_X1 U13897 ( .A1(n13924), .A2(n11459), .ZN(n11385) );
  NAND2_X1 U13898 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  XNOR2_X1 U13899 ( .A(n11387), .B(n11410), .ZN(n11389) );
  AND2_X1 U13900 ( .A1(n11367), .A2(n13924), .ZN(n11388) );
  AOI21_X1 U13901 ( .B1(n13903), .B2(n11234), .A(n11388), .ZN(n11390) );
  NAND2_X1 U13902 ( .A1(n11389), .A2(n11390), .ZN(n11394) );
  INV_X1 U13903 ( .A(n11389), .ZN(n11392) );
  INV_X1 U13904 ( .A(n11390), .ZN(n11391) );
  NAND2_X1 U13905 ( .A1(n11392), .A2(n11391), .ZN(n11393) );
  NAND2_X1 U13906 ( .A1(n11394), .A2(n11393), .ZN(n13426) );
  INV_X1 U13907 ( .A(n11394), .ZN(n13417) );
  NAND2_X1 U13908 ( .A1(n11671), .A2(n6468), .ZN(n11397) );
  OR2_X1 U13909 ( .A1(n13653), .A2(n11395), .ZN(n11396) );
  NAND2_X1 U13910 ( .A1(n14078), .A2(n9068), .ZN(n11409) );
  NAND2_X1 U13911 ( .A1(n11632), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11407) );
  INV_X1 U13912 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11398) );
  OR2_X1 U13913 ( .A1(n6463), .A2(n11398), .ZN(n11406) );
  INV_X1 U13914 ( .A(n11401), .ZN(n11399) );
  NAND2_X1 U13915 ( .A1(n11399), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11426) );
  INV_X1 U13916 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11400) );
  NAND2_X1 U13917 ( .A1(n11401), .A2(n11400), .ZN(n11402) );
  NAND2_X1 U13918 ( .A1(n11426), .A2(n11402), .ZN(n13883) );
  OR2_X1 U13919 ( .A1(n9585), .A2(n13883), .ZN(n11405) );
  INV_X1 U13920 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n11403) );
  OR2_X1 U13921 ( .A1(n13638), .A2(n11403), .ZN(n11404) );
  NAND4_X1 U13922 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n13895) );
  NAND2_X1 U13923 ( .A1(n13895), .A2(n11459), .ZN(n11408) );
  NAND2_X1 U13924 ( .A1(n11409), .A2(n11408), .ZN(n11411) );
  XNOR2_X1 U13925 ( .A(n11411), .B(n11410), .ZN(n11413) );
  AND2_X1 U13926 ( .A1(n11367), .A2(n13895), .ZN(n11412) );
  AOI21_X1 U13927 ( .B1(n14078), .B2(n11234), .A(n11412), .ZN(n11414) );
  NAND2_X1 U13928 ( .A1(n11413), .A2(n11414), .ZN(n11418) );
  INV_X1 U13929 ( .A(n11413), .ZN(n11416) );
  INV_X1 U13930 ( .A(n11414), .ZN(n11415) );
  NAND2_X1 U13931 ( .A1(n11416), .A2(n11415), .ZN(n11417) );
  NAND2_X1 U13932 ( .A1(n11688), .A2(n6468), .ZN(n11421) );
  OR2_X1 U13933 ( .A1(n13653), .A2(n11419), .ZN(n11420) );
  NAND2_X1 U13934 ( .A1(n14174), .A2(n11422), .ZN(n11434) );
  NAND2_X1 U13935 ( .A1(n11483), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11432) );
  INV_X1 U13936 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11423) );
  OR2_X1 U13937 ( .A1(n13639), .A2(n11423), .ZN(n11431) );
  INV_X1 U13938 ( .A(n11426), .ZN(n11424) );
  NAND2_X1 U13939 ( .A1(n11424), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11450) );
  INV_X1 U13940 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11425) );
  NAND2_X1 U13941 ( .A1(n11426), .A2(n11425), .ZN(n11427) );
  NAND2_X1 U13942 ( .A1(n11450), .A2(n11427), .ZN(n13868) );
  OR2_X1 U13943 ( .A1(n9585), .A2(n13868), .ZN(n11430) );
  INV_X1 U13944 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11428) );
  OR2_X1 U13945 ( .A1(n6463), .A2(n11428), .ZN(n11429) );
  NAND4_X1 U13946 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n13879) );
  NAND2_X1 U13947 ( .A1(n13879), .A2(n11459), .ZN(n11433) );
  NAND2_X1 U13948 ( .A1(n11434), .A2(n11433), .ZN(n11435) );
  XNOR2_X1 U13949 ( .A(n11435), .B(n11477), .ZN(n11440) );
  NAND2_X1 U13950 ( .A1(n14174), .A2(n11436), .ZN(n11438) );
  NAND2_X1 U13951 ( .A1(n11367), .A2(n13879), .ZN(n11437) );
  NAND2_X1 U13952 ( .A1(n11438), .A2(n11437), .ZN(n11439) );
  NOR2_X1 U13953 ( .A1(n11440), .A2(n11439), .ZN(n11441) );
  AOI21_X1 U13954 ( .B1(n11440), .B2(n11439), .A(n11441), .ZN(n13479) );
  INV_X1 U13955 ( .A(n11441), .ZN(n11442) );
  INV_X1 U13956 ( .A(n11443), .ZN(n11444) );
  NAND2_X1 U13957 ( .A1(n13364), .A2(n6468), .ZN(n11447) );
  OR2_X1 U13958 ( .A1(n13653), .A2(n14222), .ZN(n11446) );
  NAND2_X1 U13959 ( .A1(n13618), .A2(n9068), .ZN(n11457) );
  NAND2_X1 U13960 ( .A1(n11483), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11455) );
  INV_X1 U13961 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14170) );
  OR2_X1 U13962 ( .A1(n13639), .A2(n14170), .ZN(n11454) );
  INV_X1 U13963 ( .A(n11450), .ZN(n11448) );
  NAND2_X1 U13964 ( .A1(n11448), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11470) );
  INV_X1 U13965 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11449) );
  NAND2_X1 U13966 ( .A1(n11450), .A2(n11449), .ZN(n11451) );
  NAND2_X1 U13967 ( .A1(n11470), .A2(n11451), .ZN(n13851) );
  OR2_X1 U13968 ( .A1(n9585), .A2(n13851), .ZN(n11453) );
  INV_X1 U13969 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14069) );
  OR2_X1 U13970 ( .A1(n9589), .A2(n14069), .ZN(n11452) );
  NAND4_X1 U13971 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n13820) );
  NAND2_X1 U13972 ( .A1(n13820), .A2(n11459), .ZN(n11456) );
  NAND2_X1 U13973 ( .A1(n11457), .A2(n11456), .ZN(n11458) );
  XNOR2_X1 U13974 ( .A(n11458), .B(n11477), .ZN(n11463) );
  NAND2_X1 U13975 ( .A1(n13618), .A2(n11459), .ZN(n11461) );
  NAND2_X1 U13976 ( .A1(n11367), .A2(n13820), .ZN(n11460) );
  NAND2_X1 U13977 ( .A1(n11461), .A2(n11460), .ZN(n11462) );
  NOR2_X1 U13978 ( .A1(n11463), .A2(n11462), .ZN(n11464) );
  AOI21_X1 U13979 ( .B1(n11463), .B2(n11462), .A(n11464), .ZN(n13370) );
  NAND2_X1 U13980 ( .A1(n11721), .A2(n6468), .ZN(n11468) );
  INV_X1 U13981 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11595) );
  OR2_X1 U13982 ( .A1(n13653), .A2(n11595), .ZN(n11467) );
  NAND2_X1 U13983 ( .A1(n11483), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n11475) );
  INV_X1 U13984 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n14165) );
  OR2_X1 U13985 ( .A1(n13639), .A2(n14165), .ZN(n11474) );
  INV_X1 U13986 ( .A(n11470), .ZN(n11469) );
  NAND2_X1 U13987 ( .A1(n11469), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n11640) );
  INV_X1 U13988 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U13989 ( .A1(n11470), .A2(n11482), .ZN(n11471) );
  NAND2_X1 U13990 ( .A1(n11640), .A2(n11471), .ZN(n13833) );
  OR2_X1 U13991 ( .A1(n9585), .A2(n13833), .ZN(n11473) );
  INV_X1 U13992 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n14062) );
  OR2_X1 U13993 ( .A1(n9589), .A2(n14062), .ZN(n11472) );
  NAND4_X1 U13994 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n14050) );
  OAI22_X1 U13995 ( .A1(n14168), .A2(n11476), .B1(n13372), .B2(n11276), .ZN(
        n11478) );
  XNOR2_X1 U13996 ( .A(n11478), .B(n11477), .ZN(n11480) );
  OAI22_X1 U13997 ( .A1(n14168), .A2(n11276), .B1(n13372), .B2(n9289), .ZN(
        n11479) );
  XNOR2_X1 U13998 ( .A(n11480), .B(n11479), .ZN(n11481) );
  OAI22_X1 U13999 ( .A1(n14436), .A2(n13833), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11482), .ZN(n11492) );
  NAND2_X1 U14000 ( .A1(n11483), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11489) );
  INV_X1 U14001 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n11484) );
  OR2_X1 U14002 ( .A1(n13639), .A2(n11484), .ZN(n11488) );
  OR2_X1 U14003 ( .A1(n9585), .A2(n11640), .ZN(n11487) );
  INV_X1 U14004 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n11485) );
  OR2_X1 U14005 ( .A1(n6463), .A2(n11485), .ZN(n11486) );
  NAND4_X1 U14006 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n13821) );
  INV_X1 U14007 ( .A(n13821), .ZN(n11490) );
  INV_X1 U14008 ( .A(n13820), .ZN(n11627) );
  OAI22_X1 U14009 ( .A1(n11490), .A2(n14426), .B1(n14427), .B2(n11627), .ZN(
        n11491) );
  AOI211_X1 U14010 ( .C1(n13830), .C2(n14415), .A(n11492), .B(n11491), .ZN(
        n11493) );
  OAI21_X1 U14011 ( .B1(n11494), .B2(n14410), .A(n11493), .ZN(P1_U3220) );
  AOI22_X1 U14012 ( .A1(n11507), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n11506), 
        .B2(n12972), .ZN(n11496) );
  XNOR2_X1 U14013 ( .A(n13318), .B(n11736), .ZN(n11503) );
  NAND2_X1 U14014 ( .A1(n13000), .A2(n9668), .ZN(n11504) );
  INV_X1 U14015 ( .A(n11498), .ZN(n11499) );
  XOR2_X1 U14016 ( .A(n11504), .B(n11503), .Z(n12854) );
  AOI22_X1 U14017 ( .A1(n11507), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11506), 
        .B2(n8916), .ZN(n11508) );
  XNOR2_X1 U14018 ( .A(n13202), .B(n11736), .ZN(n11514) );
  NOR2_X1 U14019 ( .A1(n11510), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n11511) );
  OR2_X1 U14020 ( .A1(n11522), .A2(n11511), .ZN(n13198) );
  AOI22_X1 U14021 ( .A1(n8982), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n11958), 
        .B2(P2_REG1_REG_19__SCAN_IN), .ZN(n11513) );
  NAND2_X1 U14022 ( .A1(n11959), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n11512) );
  OAI211_X1 U14023 ( .C1(n13198), .C2(n11741), .A(n11513), .B(n11512), .ZN(
        n13003) );
  NAND2_X1 U14024 ( .A1(n13003), .A2(n9668), .ZN(n11515) );
  NAND2_X1 U14025 ( .A1(n11514), .A2(n11515), .ZN(n12782) );
  INV_X1 U14026 ( .A(n11514), .ZN(n11517) );
  INV_X1 U14027 ( .A(n11515), .ZN(n11516) );
  NAND2_X1 U14028 ( .A1(n11517), .A2(n11516), .ZN(n12781) );
  NAND2_X1 U14029 ( .A1(n11518), .A2(n11951), .ZN(n11521) );
  OR2_X1 U14030 ( .A1(n11953), .A2(n11519), .ZN(n11520) );
  XNOR2_X1 U14031 ( .A(n13309), .B(n11579), .ZN(n11527) );
  NOR2_X1 U14032 ( .A1(n11522), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n11523) );
  OR2_X1 U14033 ( .A1(n11533), .A2(n11523), .ZN(n13183) );
  AOI22_X1 U14034 ( .A1(n8982), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n11958), 
        .B2(P2_REG1_REG_20__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U14035 ( .A1(n11959), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n11524) );
  OAI211_X1 U14036 ( .C1(n13183), .C2(n11741), .A(n11525), .B(n11524), .ZN(
        n13029) );
  NAND2_X1 U14037 ( .A1(n13029), .A2(n9668), .ZN(n11526) );
  NAND2_X1 U14038 ( .A1(n11527), .A2(n11526), .ZN(n11528) );
  OAI21_X1 U14039 ( .B1(n11527), .B2(n11526), .A(n11528), .ZN(n12847) );
  NAND2_X1 U14040 ( .A1(n11529), .A2(n11951), .ZN(n11532) );
  OR2_X1 U14041 ( .A1(n11953), .A2(n11530), .ZN(n11531) );
  XNOR2_X1 U14042 ( .A(n13304), .B(n11736), .ZN(n11540) );
  OR2_X1 U14043 ( .A1(n11533), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n11534) );
  NAND2_X1 U14044 ( .A1(n11533), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n11547) );
  AND2_X1 U14045 ( .A1(n11534), .A2(n11547), .ZN(n13170) );
  INV_X1 U14046 ( .A(n11741), .ZN(n11535) );
  NAND2_X1 U14047 ( .A1(n13170), .A2(n11535), .ZN(n11538) );
  AOI22_X1 U14048 ( .A1(n8982), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n11958), 
        .B2(P2_REG1_REG_21__SCAN_IN), .ZN(n11537) );
  NAND2_X1 U14049 ( .A1(n11959), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n11536) );
  NOR2_X1 U14050 ( .A1(n12848), .A2(n11702), .ZN(n11539) );
  XNOR2_X1 U14051 ( .A(n11540), .B(n11539), .ZN(n12790) );
  NAND2_X1 U14052 ( .A1(n11540), .A2(n11539), .ZN(n11541) );
  NAND2_X1 U14053 ( .A1(n11542), .A2(n11951), .ZN(n11545) );
  OR2_X1 U14054 ( .A1(n11953), .A2(n11543), .ZN(n11544) );
  XNOR2_X1 U14055 ( .A(n13157), .B(n11579), .ZN(n11571) );
  NAND2_X1 U14056 ( .A1(n8982), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n11553) );
  INV_X1 U14057 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n11546) );
  OR2_X1 U14058 ( .A1(n6950), .A2(n11546), .ZN(n11552) );
  OAI21_X1 U14059 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n11548), .A(n11558), 
        .ZN(n13153) );
  OR2_X1 U14060 ( .A1(n11741), .A2(n13153), .ZN(n11551) );
  INV_X1 U14061 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n11549) );
  OR2_X1 U14062 ( .A1(n11743), .A2(n11549), .ZN(n11550) );
  NAND4_X1 U14063 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n13034) );
  NAND2_X1 U14064 ( .A1(n13034), .A2(n9668), .ZN(n11554) );
  NAND2_X1 U14065 ( .A1(n11566), .A2(n11554), .ZN(n11574) );
  NAND2_X1 U14066 ( .A1(n8982), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n11564) );
  INV_X1 U14067 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n11555) );
  OR2_X1 U14068 ( .A1(n6950), .A2(n11555), .ZN(n11563) );
  INV_X1 U14069 ( .A(n11558), .ZN(n11556) );
  NAND2_X1 U14070 ( .A1(n11556), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n11583) );
  INV_X1 U14071 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U14072 ( .A1(n11558), .A2(n11557), .ZN(n11559) );
  NAND2_X1 U14073 ( .A1(n11583), .A2(n11559), .ZN(n13137) );
  OR2_X1 U14074 ( .A1(n11741), .A2(n13137), .ZN(n11562) );
  INV_X1 U14075 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n11560) );
  OR2_X1 U14076 ( .A1(n11743), .A2(n11560), .ZN(n11561) );
  OAI22_X1 U14077 ( .A1(n12848), .A2(n12775), .B1(n13006), .B2(n12988), .ZN(
        n13147) );
  AOI22_X1 U14078 ( .A1(n13147), .A2(n12871), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11565) );
  OAI21_X1 U14079 ( .B1(n13153), .B2(n12873), .A(n11565), .ZN(n11568) );
  INV_X1 U14080 ( .A(n13034), .ZN(n12002) );
  NOR3_X1 U14081 ( .A1(n11566), .A2(n12002), .A3(n12828), .ZN(n11567) );
  AOI211_X1 U14082 ( .C1(n13157), .C2(n12875), .A(n11568), .B(n11567), .ZN(
        n11569) );
  OAI21_X1 U14083 ( .B1(n11574), .B2(n12877), .A(n11569), .ZN(P2_U3207) );
  INV_X1 U14084 ( .A(n11570), .ZN(n11572) );
  NAND2_X1 U14085 ( .A1(n11572), .A2(n11571), .ZN(n11573) );
  NAND2_X1 U14086 ( .A1(n11575), .A2(n11951), .ZN(n11578) );
  OR2_X1 U14087 ( .A1(n11953), .A2(n11576), .ZN(n11577) );
  XNOR2_X1 U14088 ( .A(n12983), .B(n11579), .ZN(n11660) );
  NAND2_X1 U14089 ( .A1(n13035), .A2(n9668), .ZN(n11580) );
  NAND2_X1 U14090 ( .A1(n11958), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n11588) );
  INV_X1 U14091 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n11581) );
  OR2_X1 U14092 ( .A1(n11743), .A2(n11581), .ZN(n11587) );
  INV_X1 U14093 ( .A(n11583), .ZN(n11582) );
  NAND2_X1 U14094 ( .A1(n11582), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n11677) );
  INV_X1 U14095 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12841) );
  NAND2_X1 U14096 ( .A1(n11583), .A2(n12841), .ZN(n11584) );
  NAND2_X1 U14097 ( .A1(n11677), .A2(n11584), .ZN(n13119) );
  OR2_X1 U14098 ( .A1(n11741), .A2(n13119), .ZN(n11586) );
  INV_X1 U14099 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13120) );
  OR2_X1 U14100 ( .A1(n11962), .A2(n13120), .ZN(n11585) );
  NAND4_X1 U14101 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n12881) );
  INV_X1 U14102 ( .A(n12881), .ZN(n13036) );
  OAI22_X1 U14103 ( .A1(n12002), .A2(n12775), .B1(n13036), .B2(n12988), .ZN(
        n13135) );
  AOI22_X1 U14104 ( .A1(n12871), .A2(n13135), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11589) );
  OAI21_X1 U14105 ( .B1(n13137), .B2(n12873), .A(n11589), .ZN(n11592) );
  NOR3_X1 U14106 ( .A1(n11590), .A2(n13006), .A3(n12828), .ZN(n11591) );
  AOI211_X1 U14107 ( .C1(n13292), .C2(n12875), .A(n11592), .B(n11591), .ZN(
        n11593) );
  OAI21_X1 U14108 ( .B1(n11662), .B2(n12877), .A(n11593), .ZN(P2_U3188) );
  INV_X1 U14109 ( .A(n11721), .ZN(n13363) );
  OAI222_X1 U14110 ( .A1(n14223), .A2(n11595), .B1(n14221), .B2(n13363), .C1(
        P1_U3086), .C2(n11594), .ZN(P1_U3327) );
  OR2_X1 U14111 ( .A1(n14145), .A2(n14447), .ZN(n11596) );
  XNOR2_X1 U14112 ( .A(n14390), .B(n14437), .ZN(n13686) );
  NAND2_X1 U14113 ( .A1(n14022), .A2(n14021), .ZN(n14024) );
  OR2_X1 U14114 ( .A1(n14390), .A2(n14437), .ZN(n11599) );
  OR2_X1 U14115 ( .A1(n7206), .A2(n14134), .ZN(n13670) );
  INV_X1 U14116 ( .A(n13670), .ZN(n11600) );
  NAND2_X1 U14117 ( .A1(n7206), .A2(n14134), .ZN(n13669) );
  AND2_X1 U14118 ( .A1(n14001), .A2(n13720), .ZN(n13587) );
  OR2_X1 U14119 ( .A1(n14001), .A2(n13720), .ZN(n13586) );
  XNOR2_X1 U14120 ( .A(n13981), .B(n14124), .ZN(n13987) );
  OR2_X1 U14121 ( .A1(n13981), .A2(n13994), .ZN(n11601) );
  NAND2_X1 U14122 ( .A1(n11602), .A2(n11601), .ZN(n13966) );
  XNOR2_X1 U14123 ( .A(n13973), .B(n13719), .ZN(n13967) );
  OR2_X1 U14124 ( .A1(n14196), .A2(n13592), .ZN(n11603) );
  INV_X1 U14125 ( .A(n13718), .ZN(n11621) );
  XNOR2_X1 U14126 ( .A(n13950), .B(n11621), .ZN(n13953) );
  OR2_X1 U14127 ( .A1(n13601), .A2(n13717), .ZN(n11604) );
  INV_X1 U14128 ( .A(n13894), .ZN(n13431) );
  XNOR2_X1 U14129 ( .A(n13918), .B(n13431), .ZN(n13912) );
  NAND2_X1 U14130 ( .A1(n13918), .A2(n13894), .ZN(n11605) );
  NAND2_X1 U14131 ( .A1(n13911), .A2(n11605), .ZN(n13893) );
  NAND2_X1 U14132 ( .A1(n14078), .A2(n13895), .ZN(n11607) );
  OR2_X1 U14133 ( .A1(n14078), .A2(n13895), .ZN(n11606) );
  XNOR2_X1 U14134 ( .A(n14174), .B(n13879), .ZN(n13861) );
  INV_X1 U14135 ( .A(n13861), .ZN(n13858) );
  NAND2_X1 U14136 ( .A1(n13859), .A2(n13858), .ZN(n11609) );
  NAND2_X1 U14137 ( .A1(n14174), .A2(n13879), .ZN(n11608) );
  NAND2_X1 U14138 ( .A1(n11609), .A2(n11608), .ZN(n13844) );
  XNOR2_X1 U14139 ( .A(n13618), .B(n11627), .ZN(n13695) );
  XNOR2_X1 U14140 ( .A(n13830), .B(n13372), .ZN(n13818) );
  NAND2_X1 U14141 ( .A1(n11931), .A2(n6468), .ZN(n11613) );
  OR2_X1 U14142 ( .A1(n13653), .A2(n11649), .ZN(n11612) );
  XNOR2_X1 U14143 ( .A(n13629), .B(n13821), .ZN(n13696) );
  NOR2_X1 U14144 ( .A1(n14440), .A2(n14134), .ZN(n11615) );
  XNOR2_X1 U14145 ( .A(n14001), .B(n13720), .ZN(n13993) );
  NAND2_X1 U14146 ( .A1(n13992), .A2(n13993), .ZN(n11617) );
  NAND2_X1 U14147 ( .A1(n14201), .A2(n13720), .ZN(n11616) );
  NAND2_X1 U14148 ( .A1(n13981), .A2(n14124), .ZN(n11618) );
  INV_X1 U14149 ( .A(n13967), .ZN(n11619) );
  OR2_X2 U14150 ( .A1(n13959), .A2(n11619), .ZN(n13960) );
  NAND2_X1 U14151 ( .A1(n14196), .A2(n13719), .ZN(n11620) );
  NOR2_X1 U14152 ( .A1(n13950), .A2(n11621), .ZN(n11622) );
  INV_X1 U14153 ( .A(n13930), .ZN(n13933) );
  INV_X1 U14154 ( .A(n13717), .ZN(n13921) );
  NAND2_X1 U14155 ( .A1(n13915), .A2(n13914), .ZN(n13913) );
  NAND2_X1 U14156 ( .A1(n13918), .A2(n13431), .ZN(n11623) );
  INV_X1 U14157 ( .A(n13924), .ZN(n13420) );
  OR2_X1 U14158 ( .A1(n13903), .A2(n13420), .ZN(n13875) );
  AND2_X1 U14159 ( .A1(n13877), .A2(n13875), .ZN(n11624) );
  NAND2_X1 U14160 ( .A1(n13896), .A2(n11624), .ZN(n13876) );
  INV_X1 U14161 ( .A(n13895), .ZN(n13432) );
  NAND2_X1 U14162 ( .A1(n14078), .A2(n13432), .ZN(n11625) );
  NAND2_X1 U14163 ( .A1(n13876), .A2(n11625), .ZN(n13862) );
  NAND2_X1 U14164 ( .A1(n13862), .A2(n13861), .ZN(n13860) );
  INV_X1 U14165 ( .A(n13879), .ZN(n13421) );
  NAND2_X1 U14166 ( .A1(n14174), .A2(n13421), .ZN(n11626) );
  NAND2_X1 U14167 ( .A1(n13860), .A2(n11626), .ZN(n13840) );
  NAND2_X1 U14168 ( .A1(n13840), .A2(n13843), .ZN(n13839) );
  NAND2_X1 U14169 ( .A1(n13618), .A2(n11627), .ZN(n11628) );
  XNOR2_X1 U14170 ( .A(n11629), .B(n13696), .ZN(n14054) );
  NAND2_X1 U14171 ( .A1(n13979), .A2(n14196), .ZN(n13946) );
  NOR2_X1 U14172 ( .A1(n14174), .A2(n13881), .ZN(n13867) );
  NAND2_X1 U14173 ( .A1(n14066), .A2(n13867), .ZN(n13850) );
  AOI21_X1 U14174 ( .B1(n13629), .B2(n13831), .A(n13980), .ZN(n11630) );
  NAND2_X1 U14175 ( .A1(n11630), .A2(n13811), .ZN(n14052) );
  NOR2_X1 U14176 ( .A1(n14052), .A2(n14035), .ZN(n11647) );
  INV_X1 U14177 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13813) );
  NAND2_X1 U14178 ( .A1(n11631), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U14179 ( .A1(n11632), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11633) );
  OAI211_X1 U14180 ( .C1(n13638), .C2(n13813), .A(n11634), .B(n11633), .ZN(
        n13716) );
  INV_X1 U14181 ( .A(n13716), .ZN(n11637) );
  INV_X1 U14182 ( .A(P1_B_REG_SCAN_IN), .ZN(n11635) );
  OR2_X1 U14183 ( .A1(n14496), .A2(n11635), .ZN(n11636) );
  NAND2_X1 U14184 ( .A1(n14635), .A2(n11636), .ZN(n13805) );
  NOR2_X1 U14185 ( .A1(n11637), .A2(n13805), .ZN(n14049) );
  INV_X1 U14186 ( .A(n11638), .ZN(n11639) );
  NAND2_X1 U14187 ( .A1(n14049), .A2(n11639), .ZN(n11642) );
  OAI22_X1 U14188 ( .A1(n11642), .A2(n11641), .B1(n11640), .B2(n14599), .ZN(
        n11644) );
  NOR2_X1 U14189 ( .A1(n14029), .A2(n13372), .ZN(n11643) );
  AOI211_X1 U14190 ( .C1(n14016), .C2(P1_REG2_REG_29__SCAN_IN), .A(n11644), 
        .B(n11643), .ZN(n11645) );
  OAI21_X1 U14191 ( .B1(n7198), .B2(n13982), .A(n11645), .ZN(n11646) );
  AOI211_X1 U14192 ( .C1(n14054), .C2(n14623), .A(n11647), .B(n11646), .ZN(
        n11648) );
  OAI21_X1 U14193 ( .B1(n14056), .B2(n14004), .A(n11648), .ZN(P1_U3356) );
  INV_X1 U14194 ( .A(n11931), .ZN(n12050) );
  OAI222_X1 U14195 ( .A1(n14223), .A2(n11649), .B1(n14221), .B2(n12050), .C1(
        n9050), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U14196 ( .A(n11650), .ZN(n11652) );
  AOI22_X1 U14197 ( .A1(n11652), .A2(n12808), .B1(n11651), .B2(n12883), .ZN(
        n11658) );
  AOI22_X1 U14198 ( .A1(n12871), .A2(n11653), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11654) );
  OAI21_X1 U14199 ( .B1(n11655), .B2(n12873), .A(n11654), .ZN(n11656) );
  AOI21_X1 U14200 ( .B1(n13331), .B2(n12875), .A(n11656), .ZN(n11657) );
  OAI21_X1 U14201 ( .B1(n11659), .B2(n11658), .A(n11657), .ZN(P2_U3213) );
  NAND2_X1 U14202 ( .A1(n12881), .A2(n9668), .ZN(n11667) );
  NAND2_X1 U14203 ( .A1(n11663), .A2(n11951), .ZN(n11666) );
  OR2_X1 U14204 ( .A1(n11953), .A2(n11664), .ZN(n11665) );
  XNOR2_X1 U14205 ( .A(n13287), .B(n11736), .ZN(n11669) );
  XOR2_X1 U14206 ( .A(n11667), .B(n11669), .Z(n12838) );
  INV_X1 U14207 ( .A(n11667), .ZN(n11668) );
  NAND2_X1 U14208 ( .A1(n11669), .A2(n11668), .ZN(n11670) );
  NAND2_X1 U14209 ( .A1(n11671), .A2(n11951), .ZN(n11674) );
  OR2_X1 U14210 ( .A1(n11953), .A2(n11672), .ZN(n11673) );
  XNOR2_X1 U14211 ( .A(n13282), .B(n11736), .ZN(n11686) );
  NAND2_X1 U14212 ( .A1(n11958), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n11683) );
  INV_X1 U14213 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13104) );
  OR2_X1 U14214 ( .A1(n11962), .A2(n13104), .ZN(n11682) );
  INV_X1 U14215 ( .A(n11677), .ZN(n11675) );
  NAND2_X1 U14216 ( .A1(n11675), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n11695) );
  INV_X1 U14217 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n11676) );
  NAND2_X1 U14218 ( .A1(n11677), .A2(n11676), .ZN(n11678) );
  NAND2_X1 U14219 ( .A1(n11695), .A2(n11678), .ZN(n13103) );
  OR2_X1 U14220 ( .A1(n11741), .A2(n13103), .ZN(n11681) );
  INV_X1 U14221 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n11679) );
  OR2_X1 U14222 ( .A1(n11743), .A2(n11679), .ZN(n11680) );
  NAND4_X1 U14223 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n13038) );
  NAND2_X1 U14224 ( .A1(n13038), .A2(n9668), .ZN(n11684) );
  XNOR2_X1 U14225 ( .A(n11686), .B(n11684), .ZN(n12797) );
  INV_X1 U14226 ( .A(n11684), .ZN(n11685) );
  NAND2_X1 U14227 ( .A1(n11686), .A2(n11685), .ZN(n11687) );
  NAND2_X1 U14228 ( .A1(n11688), .A2(n11951), .ZN(n11691) );
  OR2_X1 U14229 ( .A1(n11953), .A2(n11689), .ZN(n11690) );
  XNOR2_X1 U14230 ( .A(n13090), .B(n11736), .ZN(n11704) );
  NAND2_X1 U14231 ( .A1(n8982), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n11701) );
  INV_X1 U14232 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n11692) );
  OR2_X1 U14233 ( .A1(n6950), .A2(n11692), .ZN(n11700) );
  INV_X1 U14234 ( .A(n11695), .ZN(n11693) );
  NAND2_X1 U14235 ( .A1(n11693), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n11712) );
  INV_X1 U14236 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U14237 ( .A1(n11695), .A2(n11694), .ZN(n11696) );
  NAND2_X1 U14238 ( .A1(n11712), .A2(n11696), .ZN(n13087) );
  OR2_X1 U14239 ( .A1(n11741), .A2(n13087), .ZN(n11699) );
  INV_X1 U14240 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n11697) );
  OR2_X1 U14241 ( .A1(n11743), .A2(n11697), .ZN(n11698) );
  OR2_X1 U14242 ( .A1(n12799), .A2(n11702), .ZN(n11703) );
  NAND2_X1 U14243 ( .A1(n11704), .A2(n11703), .ZN(n11706) );
  OAI21_X1 U14244 ( .B1(n11704), .B2(n11703), .A(n11706), .ZN(n12868) );
  NAND2_X1 U14245 ( .A1(n13364), .A2(n11951), .ZN(n11708) );
  OR2_X1 U14246 ( .A1(n11953), .A2(n13367), .ZN(n11707) );
  XNOR2_X1 U14247 ( .A(n13076), .B(n11736), .ZN(n11720) );
  NAND2_X1 U14248 ( .A1(n8982), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n11718) );
  INV_X1 U14249 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n11709) );
  OR2_X1 U14250 ( .A1(n6950), .A2(n11709), .ZN(n11717) );
  INV_X1 U14251 ( .A(n11712), .ZN(n11710) );
  INV_X1 U14252 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n11711) );
  NAND2_X1 U14253 ( .A1(n11712), .A2(n11711), .ZN(n11713) );
  NAND2_X1 U14254 ( .A1(n11729), .A2(n11713), .ZN(n13073) );
  OR2_X1 U14255 ( .A1(n11741), .A2(n13073), .ZN(n11716) );
  INV_X1 U14256 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n11714) );
  OR2_X1 U14257 ( .A1(n11743), .A2(n11714), .ZN(n11715) );
  INV_X1 U14258 ( .A(n13042), .ZN(n12880) );
  NAND2_X1 U14259 ( .A1(n12880), .A2(n9668), .ZN(n11719) );
  XNOR2_X1 U14260 ( .A(n11720), .B(n11719), .ZN(n12774) );
  NAND2_X1 U14261 ( .A1(n11721), .A2(n11951), .ZN(n11724) );
  OR2_X1 U14262 ( .A1(n11953), .A2(n11722), .ZN(n11723) );
  NAND2_X1 U14263 ( .A1(n8982), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n11735) );
  INV_X1 U14264 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n11725) );
  OR2_X1 U14265 ( .A1(n6950), .A2(n11725), .ZN(n11734) );
  NAND2_X1 U14266 ( .A1(n11727), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13048) );
  INV_X1 U14267 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11728) );
  NAND2_X1 U14268 ( .A1(n11729), .A2(n11728), .ZN(n11730) );
  NAND2_X1 U14269 ( .A1(n13048), .A2(n11730), .ZN(n13059) );
  OR2_X1 U14270 ( .A1(n11741), .A2(n13059), .ZN(n11733) );
  INV_X1 U14271 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n11731) );
  OR2_X1 U14272 ( .A1(n11743), .A2(n11731), .ZN(n11732) );
  NAND4_X1 U14273 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n13043) );
  NAND2_X1 U14274 ( .A1(n13043), .A2(n9668), .ZN(n11737) );
  XNOR2_X1 U14275 ( .A(n11737), .B(n11736), .ZN(n11738) );
  XNOR2_X1 U14276 ( .A(n13267), .B(n11738), .ZN(n11739) );
  XNOR2_X1 U14277 ( .A(n11740), .B(n11739), .ZN(n11752) );
  NAND2_X1 U14278 ( .A1(n8982), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U14279 ( .A1(n11958), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11746) );
  OR2_X1 U14280 ( .A1(n11741), .A2(n13048), .ZN(n11745) );
  INV_X1 U14281 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n11742) );
  OR2_X1 U14282 ( .A1(n11743), .A2(n11742), .ZN(n11744) );
  NAND4_X1 U14283 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n12879) );
  INV_X1 U14284 ( .A(n12879), .ZN(n11748) );
  OAI22_X1 U14285 ( .A1(n11748), .A2(n12988), .B1(n13042), .B2(n12775), .ZN(
        n13058) );
  AOI22_X1 U14286 ( .A1(n12871), .A2(n13058), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11749) );
  OAI21_X1 U14287 ( .B1(n13059), .B2(n12873), .A(n11749), .ZN(n11750) );
  AOI21_X1 U14288 ( .B1(n13267), .B2(n12875), .A(n11750), .ZN(n11751) );
  OAI21_X1 U14289 ( .B1(n11752), .B2(n12877), .A(n11751), .ZN(P2_U3192) );
  INV_X1 U14290 ( .A(n11753), .ZN(n11754) );
  OAI222_X1 U14291 ( .A1(n12369), .A2(P3_U3151), .B1(n12770), .B2(n11754), 
        .C1(n15347), .C2(n12771), .ZN(P3_U3268) );
  INV_X1 U14292 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n11756) );
  OR2_X4 U14293 ( .A1(n14881), .A2(n12031), .ZN(n11782) );
  NAND2_X1 U14294 ( .A1(n11837), .A2(n11782), .ZN(n11759) );
  NAND2_X1 U14295 ( .A1(n12888), .A2(n11965), .ZN(n11758) );
  NAND2_X1 U14296 ( .A1(n11759), .A2(n11758), .ZN(n11841) );
  NAND2_X1 U14297 ( .A1(n13244), .A2(n11762), .ZN(n11760) );
  INV_X1 U14298 ( .A(n11764), .ZN(n11761) );
  NAND2_X1 U14299 ( .A1(n11761), .A2(n11782), .ZN(n11766) );
  NAND2_X1 U14300 ( .A1(n11762), .A2(n11956), .ZN(n11992) );
  OAI22_X1 U14301 ( .A1(n13244), .A2(n11762), .B1(n11992), .B2(n8963), .ZN(
        n11763) );
  NAND2_X1 U14302 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  NAND2_X1 U14303 ( .A1(n11766), .A2(n11765), .ZN(n11772) );
  NAND2_X1 U14304 ( .A1(n11902), .A2(n14814), .ZN(n11773) );
  NAND2_X1 U14305 ( .A1(n11774), .A2(n11773), .ZN(n11767) );
  NAND2_X1 U14306 ( .A1(n12897), .A2(n6470), .ZN(n11770) );
  NAND2_X1 U14307 ( .A1(n11782), .A2(n14814), .ZN(n11769) );
  NAND2_X1 U14308 ( .A1(n11770), .A2(n11769), .ZN(n11771) );
  INV_X1 U14309 ( .A(n11772), .ZN(n11776) );
  AND2_X1 U14310 ( .A1(n11774), .A2(n11773), .ZN(n11775) );
  NAND2_X1 U14311 ( .A1(n11776), .A2(n11775), .ZN(n11777) );
  NAND2_X1 U14312 ( .A1(n11778), .A2(n11777), .ZN(n11785) );
  NAND2_X1 U14313 ( .A1(n12896), .A2(n6471), .ZN(n11780) );
  NAND2_X1 U14314 ( .A1(n11781), .A2(n11782), .ZN(n11779) );
  NAND2_X1 U14315 ( .A1(n11780), .A2(n11779), .ZN(n11784) );
  INV_X1 U14316 ( .A(n6510), .ZN(n11902) );
  AOI22_X1 U14317 ( .A1(n12896), .A2(n11782), .B1(n11902), .B2(n11781), .ZN(
        n11783) );
  NAND2_X1 U14318 ( .A1(n12895), .A2(n11782), .ZN(n11788) );
  NAND2_X1 U14319 ( .A1(n11786), .A2(n6472), .ZN(n11787) );
  NAND2_X1 U14320 ( .A1(n11788), .A2(n11787), .ZN(n11794) );
  NAND2_X1 U14321 ( .A1(n11793), .A2(n11794), .ZN(n11792) );
  NAND2_X1 U14322 ( .A1(n12895), .A2(n6472), .ZN(n11789) );
  OAI21_X1 U14323 ( .B1(n11790), .B2(n11984), .A(n11789), .ZN(n11791) );
  NAND2_X1 U14324 ( .A1(n11792), .A2(n11791), .ZN(n11798) );
  INV_X1 U14325 ( .A(n11793), .ZN(n11796) );
  INV_X1 U14326 ( .A(n11794), .ZN(n11795) );
  NAND2_X1 U14327 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  NAND2_X1 U14328 ( .A1(n12894), .A2(n6471), .ZN(n11800) );
  NAND2_X1 U14329 ( .A1(n11801), .A2(n11782), .ZN(n11799) );
  NAND2_X1 U14330 ( .A1(n11800), .A2(n11799), .ZN(n11803) );
  NAND2_X1 U14331 ( .A1(n12893), .A2(n11782), .ZN(n11806) );
  NAND2_X1 U14332 ( .A1(n12824), .A2(n6472), .ZN(n11805) );
  NAND2_X1 U14333 ( .A1(n11806), .A2(n11805), .ZN(n11809) );
  NAND2_X1 U14334 ( .A1(n12893), .A2(n6471), .ZN(n11807) );
  OAI21_X1 U14335 ( .B1(n14836), .B2(n11984), .A(n11807), .ZN(n11808) );
  NAND2_X1 U14336 ( .A1(n11812), .A2(n11782), .ZN(n11811) );
  NAND2_X1 U14337 ( .A1(n12892), .A2(n6472), .ZN(n11810) );
  NAND2_X1 U14338 ( .A1(n11811), .A2(n11810), .ZN(n11814) );
  AOI22_X1 U14339 ( .A1(n6471), .A2(n11812), .B1(n12892), .B2(n11782), .ZN(
        n11813) );
  NAND2_X1 U14340 ( .A1(n11820), .A2(n6472), .ZN(n11817) );
  NAND2_X1 U14341 ( .A1(n12891), .A2(n11782), .ZN(n11816) );
  NAND2_X1 U14342 ( .A1(n11817), .A2(n11816), .ZN(n11819) );
  INV_X1 U14343 ( .A(n11819), .ZN(n11818) );
  INV_X1 U14344 ( .A(n11902), .ZN(n11949) );
  NAND2_X1 U14345 ( .A1(n11820), .A2(n11782), .ZN(n11821) );
  OAI21_X1 U14346 ( .B1(n11822), .B2(n11949), .A(n11821), .ZN(n11823) );
  NAND2_X1 U14347 ( .A1(n11826), .A2(n11782), .ZN(n11825) );
  NAND2_X1 U14348 ( .A1(n12890), .A2(n11965), .ZN(n11824) );
  NAND2_X1 U14349 ( .A1(n11825), .A2(n11824), .ZN(n11828) );
  AOI22_X1 U14350 ( .A1(n11826), .A2(n11965), .B1(n12890), .B2(n11782), .ZN(
        n11827) );
  NOR2_X1 U14351 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  NAND2_X1 U14352 ( .A1(n14860), .A2(n11965), .ZN(n11833) );
  NAND2_X1 U14353 ( .A1(n12889), .A2(n11782), .ZN(n11832) );
  NAND2_X1 U14354 ( .A1(n11833), .A2(n11832), .ZN(n11835) );
  AOI22_X1 U14355 ( .A1(n14860), .A2(n11782), .B1(n11965), .B2(n12889), .ZN(
        n11834) );
  NAND2_X1 U14356 ( .A1(n11837), .A2(n6472), .ZN(n11838) );
  OAI21_X1 U14357 ( .B1(n11839), .B2(n11984), .A(n11838), .ZN(n11840) );
  NAND2_X1 U14358 ( .A1(n14878), .A2(n6471), .ZN(n11843) );
  NAND2_X1 U14359 ( .A1(n12887), .A2(n11782), .ZN(n11842) );
  NAND2_X1 U14360 ( .A1(n11843), .A2(n11842), .ZN(n11846) );
  INV_X1 U14361 ( .A(n6510), .ZN(n11965) );
  AOI22_X1 U14362 ( .A1(n14878), .A2(n11782), .B1(n11965), .B2(n12887), .ZN(
        n11844) );
  INV_X1 U14363 ( .A(n11845), .ZN(n11848) );
  NAND2_X1 U14364 ( .A1(n11848), .A2(n7687), .ZN(n11856) );
  NAND2_X1 U14365 ( .A1(n11851), .A2(n11782), .ZN(n11850) );
  NAND2_X1 U14366 ( .A1(n12886), .A2(n11965), .ZN(n11849) );
  NAND2_X1 U14367 ( .A1(n11850), .A2(n11849), .ZN(n11857) );
  NAND2_X1 U14368 ( .A1(n11851), .A2(n11965), .ZN(n11852) );
  OAI21_X1 U14369 ( .B1(n11853), .B2(n11984), .A(n11852), .ZN(n11854) );
  NAND2_X1 U14370 ( .A1(n11860), .A2(n11965), .ZN(n11859) );
  NAND2_X1 U14371 ( .A1(n12885), .A2(n11782), .ZN(n11858) );
  NAND2_X1 U14372 ( .A1(n11859), .A2(n11858), .ZN(n11862) );
  AOI22_X1 U14373 ( .A1(n11860), .A2(n11782), .B1(n11965), .B2(n12885), .ZN(
        n11861) );
  NAND2_X1 U14374 ( .A1(n11866), .A2(n11782), .ZN(n11865) );
  NAND2_X1 U14375 ( .A1(n12884), .A2(n6472), .ZN(n11864) );
  NAND2_X1 U14376 ( .A1(n11865), .A2(n11864), .ZN(n11872) );
  NAND2_X1 U14377 ( .A1(n11866), .A2(n6471), .ZN(n11867) );
  OAI21_X1 U14378 ( .B1(n11868), .B2(n11984), .A(n11867), .ZN(n11869) );
  NAND2_X1 U14379 ( .A1(n11870), .A2(n11869), .ZN(n11874) );
  NAND2_X1 U14380 ( .A1(n13331), .A2(n6472), .ZN(n11876) );
  NAND2_X1 U14381 ( .A1(n12883), .A2(n11782), .ZN(n11875) );
  NAND2_X1 U14382 ( .A1(n11876), .A2(n11875), .ZN(n11881) );
  AND2_X1 U14383 ( .A1(n12882), .A2(n11965), .ZN(n11877) );
  AOI21_X1 U14384 ( .B1(n13328), .B2(n11782), .A(n11877), .ZN(n11885) );
  NAND2_X1 U14385 ( .A1(n13328), .A2(n11965), .ZN(n11879) );
  NAND2_X1 U14386 ( .A1(n12882), .A2(n11782), .ZN(n11878) );
  NAND2_X1 U14387 ( .A1(n11879), .A2(n11878), .ZN(n11884) );
  AOI22_X1 U14388 ( .A1(n13331), .A2(n11782), .B1(n6471), .B2(n12883), .ZN(
        n11880) );
  AOI22_X1 U14389 ( .A1(n13323), .A2(n11782), .B1(n11965), .B2(n12998), .ZN(
        n11886) );
  NAND2_X1 U14390 ( .A1(n13323), .A2(n11965), .ZN(n11883) );
  NAND2_X1 U14391 ( .A1(n12998), .A2(n11782), .ZN(n11882) );
  NAND2_X1 U14392 ( .A1(n11883), .A2(n11882), .ZN(n11889) );
  AOI22_X1 U14393 ( .A1(n11886), .A2(n11889), .B1(n11885), .B2(n11884), .ZN(
        n11887) );
  NOR2_X1 U14394 ( .A1(n13323), .A2(n12998), .ZN(n11888) );
  AND2_X1 U14395 ( .A1(n13000), .A2(n11965), .ZN(n11890) );
  AOI21_X1 U14396 ( .B1(n13318), .B2(n11782), .A(n11890), .ZN(n11893) );
  NAND2_X1 U14397 ( .A1(n11894), .A2(n11893), .ZN(n11896) );
  AOI22_X1 U14398 ( .A1(n13318), .A2(n11965), .B1(n13000), .B2(n11782), .ZN(
        n11891) );
  NAND2_X1 U14399 ( .A1(n11896), .A2(n11895), .ZN(n11899) );
  INV_X1 U14400 ( .A(n11899), .ZN(n11901) );
  INV_X1 U14401 ( .A(n13003), .ZN(n13002) );
  OAI22_X1 U14402 ( .A1(n13202), .A2(n11949), .B1(n13002), .B2(n11984), .ZN(
        n11898) );
  INV_X1 U14403 ( .A(n11898), .ZN(n11900) );
  AOI22_X1 U14404 ( .A1(n7148), .A2(n11782), .B1(n11965), .B2(n13003), .ZN(
        n11897) );
  AOI22_X1 U14405 ( .A1(n13309), .A2(n11782), .B1(n11902), .B2(n13029), .ZN(
        n11903) );
  AOI22_X1 U14406 ( .A1(n13309), .A2(n6472), .B1(n13029), .B2(n11782), .ZN(
        n11904) );
  OAI22_X1 U14407 ( .A1(n13173), .A2(n11949), .B1(n12848), .B2(n11984), .ZN(
        n11905) );
  OAI22_X1 U14408 ( .A1(n13173), .A2(n11984), .B1(n12848), .B2(n11949), .ZN(
        n11906) );
  AOI22_X1 U14409 ( .A1(n13157), .A2(n11782), .B1(n6472), .B2(n13034), .ZN(
        n11908) );
  INV_X1 U14410 ( .A(n13157), .ZN(n13298) );
  OAI22_X1 U14411 ( .A1(n13298), .A2(n11949), .B1(n12002), .B2(n11984), .ZN(
        n11907) );
  OAI21_X1 U14412 ( .B1(n11909), .B2(n11908), .A(n11907), .ZN(n11911) );
  NAND2_X1 U14413 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  OAI22_X1 U14414 ( .A1(n12983), .A2(n11949), .B1(n13006), .B2(n11984), .ZN(
        n11912) );
  OAI22_X1 U14415 ( .A1(n12983), .A2(n11984), .B1(n13006), .B2(n11949), .ZN(
        n11913) );
  AOI22_X1 U14416 ( .A1(n13287), .A2(n11782), .B1(n11965), .B2(n12881), .ZN(
        n11915) );
  INV_X1 U14417 ( .A(n13287), .ZN(n13037) );
  OAI22_X1 U14418 ( .A1(n13037), .A2(n11949), .B1(n13036), .B2(n11984), .ZN(
        n11914) );
  AOI22_X1 U14419 ( .A1(n13282), .A2(n11965), .B1(n13038), .B2(n11782), .ZN(
        n11918) );
  INV_X1 U14420 ( .A(n11918), .ZN(n11917) );
  AOI22_X1 U14421 ( .A1(n13282), .A2(n11782), .B1(n11965), .B2(n13038), .ZN(
        n11916) );
  INV_X1 U14422 ( .A(n12799), .ZN(n13039) );
  AOI22_X1 U14423 ( .A1(n13276), .A2(n11965), .B1(n13039), .B2(n11782), .ZN(
        n11944) );
  OAI22_X1 U14424 ( .A1(n13090), .A2(n11984), .B1(n12799), .B2(n11949), .ZN(
        n11943) );
  NAND2_X1 U14425 ( .A1(n11919), .A2(SI_30_), .ZN(n11920) );
  MUX2_X1 U14426 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8494), .Z(n11923) );
  XNOR2_X1 U14427 ( .A(n11923), .B(SI_31_), .ZN(n11924) );
  NAND2_X1 U14428 ( .A1(n14216), .A2(n11951), .ZN(n11928) );
  INV_X1 U14429 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n11926) );
  OR2_X1 U14430 ( .A1(n11953), .A2(n11926), .ZN(n11927) );
  INV_X1 U14431 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n12985) );
  NAND2_X1 U14432 ( .A1(n11958), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U14433 ( .A1(n11959), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n11929) );
  OAI211_X1 U14434 ( .C1(n11962), .C2(n12985), .A(n11930), .B(n11929), .ZN(
        n12989) );
  XNOR2_X1 U14435 ( .A(n13256), .B(n12989), .ZN(n12029) );
  NAND2_X1 U14436 ( .A1(n11931), .A2(n11951), .ZN(n11933) );
  OR2_X1 U14437 ( .A1(n11953), .A2(n12049), .ZN(n11932) );
  AND2_X1 U14438 ( .A1(n12879), .A2(n11782), .ZN(n11934) );
  AOI21_X1 U14439 ( .B1(n13263), .B2(n11965), .A(n11934), .ZN(n11969) );
  NAND2_X1 U14440 ( .A1(n13263), .A2(n11782), .ZN(n11936) );
  NAND2_X1 U14441 ( .A1(n12879), .A2(n6471), .ZN(n11935) );
  NAND2_X1 U14442 ( .A1(n11936), .A2(n11935), .ZN(n11968) );
  NAND2_X1 U14443 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  AND2_X1 U14444 ( .A1(n13043), .A2(n11782), .ZN(n11937) );
  AOI21_X1 U14445 ( .B1(n13267), .B2(n6471), .A(n11937), .ZN(n11972) );
  NAND2_X1 U14446 ( .A1(n13267), .A2(n11782), .ZN(n11940) );
  NAND2_X1 U14447 ( .A1(n13043), .A2(n6472), .ZN(n11939) );
  NAND2_X1 U14448 ( .A1(n11940), .A2(n11939), .ZN(n11971) );
  NAND2_X1 U14449 ( .A1(n11972), .A2(n11971), .ZN(n11941) );
  AND2_X1 U14450 ( .A1(n11970), .A2(n11941), .ZN(n11942) );
  OAI22_X1 U14451 ( .A1(n13076), .A2(n11984), .B1(n13042), .B2(n11949), .ZN(
        n11976) );
  AOI22_X1 U14452 ( .A1(n13271), .A2(n11965), .B1(n12880), .B2(n11782), .ZN(
        n11977) );
  AOI22_X1 U14453 ( .A1(n11976), .A2(n11977), .B1(n11944), .B2(n11943), .ZN(
        n11945) );
  INV_X1 U14454 ( .A(n12989), .ZN(n11950) );
  MUX2_X1 U14455 ( .A(n12989), .B(n11984), .S(n13256), .Z(n11948) );
  OAI21_X1 U14456 ( .B1(n11950), .B2(n11949), .A(n11948), .ZN(n11979) );
  NAND2_X1 U14457 ( .A1(n13635), .A2(n11951), .ZN(n11955) );
  OR2_X1 U14458 ( .A1(n11953), .A2(n11952), .ZN(n11954) );
  NAND2_X1 U14459 ( .A1(n12989), .A2(n11782), .ZN(n11985) );
  OR2_X1 U14460 ( .A1(n9459), .A2(n11956), .ZN(n11996) );
  NAND4_X1 U14461 ( .A1(n11985), .A2(n11957), .A3(n11996), .A4(n11993), .ZN(
        n11963) );
  INV_X1 U14462 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12993) );
  NAND2_X1 U14463 ( .A1(n11958), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U14464 ( .A1(n11959), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11960) );
  OAI211_X1 U14465 ( .C1(n11962), .C2(n12993), .A(n11961), .B(n11960), .ZN(
        n13019) );
  AND2_X1 U14466 ( .A1(n11963), .A2(n13019), .ZN(n11964) );
  AOI21_X1 U14467 ( .B1(n12996), .B2(n11965), .A(n11964), .ZN(n11981) );
  NAND2_X1 U14468 ( .A1(n12996), .A2(n11782), .ZN(n11967) );
  NAND2_X1 U14469 ( .A1(n13019), .A2(n11965), .ZN(n11966) );
  NAND2_X1 U14470 ( .A1(n11967), .A2(n11966), .ZN(n11980) );
  OAI22_X1 U14471 ( .A1(n11981), .A2(n11980), .B1(n11969), .B2(n11968), .ZN(
        n11978) );
  INV_X1 U14472 ( .A(n12029), .ZN(n11974) );
  INV_X1 U14473 ( .A(n11970), .ZN(n11973) );
  INV_X1 U14474 ( .A(n11980), .ZN(n11983) );
  INV_X1 U14475 ( .A(n11981), .ZN(n11982) );
  AND2_X1 U14476 ( .A1(n11984), .A2(n12989), .ZN(n11988) );
  INV_X1 U14477 ( .A(n11985), .ZN(n11986) );
  NOR2_X1 U14478 ( .A1(n11986), .A2(n6471), .ZN(n11987) );
  MUX2_X1 U14479 ( .A(n11988), .B(n11987), .S(n13256), .Z(n11989) );
  OAI211_X1 U14480 ( .C1(n8916), .C2(n12031), .A(n11993), .B(n11992), .ZN(
        n11994) );
  INV_X1 U14481 ( .A(n11994), .ZN(n11995) );
  OAI21_X1 U14482 ( .B1(n11997), .B2(n8963), .A(n11996), .ZN(n11998) );
  NAND2_X1 U14483 ( .A1(n12000), .A2(n11998), .ZN(n11999) );
  INV_X1 U14484 ( .A(n12000), .ZN(n12034) );
  INV_X1 U14485 ( .A(n13043), .ZN(n12776) );
  NAND2_X1 U14486 ( .A1(n13267), .A2(n12776), .ZN(n12001) );
  NAND2_X1 U14487 ( .A1(n13276), .A2(n12799), .ZN(n13013) );
  XNOR2_X1 U14488 ( .A(n13157), .B(n12002), .ZN(n13145) );
  XNOR2_X1 U14489 ( .A(n13304), .B(n12848), .ZN(n13163) );
  INV_X1 U14490 ( .A(n13029), .ZN(n13030) );
  XNOR2_X1 U14491 ( .A(n13309), .B(n13030), .ZN(n13178) );
  OR2_X1 U14492 ( .A1(n7148), .A2(n13003), .ZN(n13028) );
  NAND2_X1 U14493 ( .A1(n7148), .A2(n13003), .ZN(n13027) );
  NAND2_X1 U14494 ( .A1(n13028), .A2(n13027), .ZN(n13192) );
  XOR2_X1 U14495 ( .A(n12998), .B(n13323), .Z(n13224) );
  NAND3_X1 U14496 ( .A1(n14806), .A2(n12003), .A3(n6953), .ZN(n12004) );
  NOR4_X1 U14497 ( .A1(n12006), .A2(n12005), .A3(n12004), .A4(n7021), .ZN(
        n12010) );
  NAND4_X1 U14498 ( .A1(n12010), .A2(n12009), .A3(n12008), .A4(n12007), .ZN(
        n12011) );
  NOR4_X1 U14499 ( .A1(n12014), .A2(n12013), .A3(n12012), .A4(n12011), .ZN(
        n12017) );
  NAND4_X1 U14500 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12019) );
  NOR4_X1 U14501 ( .A1(n12021), .A2(n12020), .A3(n13224), .A4(n12019), .ZN(
        n12023) );
  XNOR2_X1 U14502 ( .A(n13318), .B(n13000), .ZN(n13207) );
  NAND4_X1 U14503 ( .A1(n13192), .A2(n12023), .A3(n13207), .A4(n12022), .ZN(
        n12024) );
  NOR4_X1 U14504 ( .A1(n13145), .A2(n13163), .A3(n13178), .A4(n12024), .ZN(
        n12025) );
  XNOR2_X1 U14505 ( .A(n13292), .B(n13035), .ZN(n13133) );
  XNOR2_X1 U14506 ( .A(n13287), .B(n12881), .ZN(n13115) );
  NAND4_X1 U14507 ( .A1(n13091), .A2(n12025), .A3(n13133), .A4(n13115), .ZN(
        n12026) );
  INV_X1 U14508 ( .A(n13038), .ZN(n13009) );
  XNOR2_X1 U14509 ( .A(n13282), .B(n13009), .ZN(n13008) );
  NOR4_X1 U14510 ( .A1(n13056), .A2(n13077), .A3(n12026), .A4(n13008), .ZN(
        n12028) );
  XNOR2_X1 U14511 ( .A(n12996), .B(n13019), .ZN(n12027) );
  XNOR2_X1 U14512 ( .A(n13263), .B(n12879), .ZN(n13044) );
  NAND4_X1 U14513 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n13044), .ZN(
        n12030) );
  XNOR2_X1 U14514 ( .A(n12030), .B(n8916), .ZN(n12032) );
  NAND2_X1 U14515 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  INV_X1 U14516 ( .A(n12041), .ZN(n12035) );
  OAI21_X1 U14517 ( .B1(n12037), .B2(n12036), .A(n12035), .ZN(n12044) );
  NAND4_X1 U14518 ( .A1(n14805), .A2(n12039), .A3(n12038), .A4(n13020), .ZN(
        n12040) );
  OAI211_X1 U14519 ( .C1(n12042), .C2(n12041), .A(n12040), .B(P2_B_REG_SCAN_IN), .ZN(n12043) );
  NAND2_X1 U14520 ( .A1(n12044), .A2(n12043), .ZN(P2_U3328) );
  INV_X1 U14521 ( .A(n12045), .ZN(n12046) );
  OAI222_X1 U14522 ( .A1(P3_U3151), .A2(n12048), .B1(n12771), .B2(n12047), 
        .C1(n12770), .C2(n12046), .ZN(P3_U3265) );
  OAI222_X1 U14523 ( .A1(n13366), .A2(n12050), .B1(P2_U3088), .B2(n8902), .C1(
        n12049), .C2(n13368), .ZN(P2_U3298) );
  XNOR2_X1 U14524 ( .A(n12421), .B(n12051), .ZN(n12058) );
  INV_X1 U14525 ( .A(n12058), .ZN(n12052) );
  NAND2_X1 U14526 ( .A1(n12052), .A2(n12203), .ZN(n12065) );
  INV_X1 U14527 ( .A(n12053), .ZN(n12054) );
  NAND4_X1 U14528 ( .A1(n12064), .A2(n12054), .A3(n12203), .A4(n12058), .ZN(
        n12063) );
  AOI22_X1 U14529 ( .A1(n12428), .A2(n12217), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12056) );
  NAND2_X1 U14530 ( .A1(n12425), .A2(n12189), .ZN(n12055) );
  OAI211_X1 U14531 ( .C1(n12427), .C2(n12187), .A(n12056), .B(n12055), .ZN(
        n12060) );
  NOR4_X1 U14532 ( .A1(n12058), .A2(n12219), .A3(n12057), .A4(n12425), .ZN(
        n12059) );
  AOI211_X1 U14533 ( .C1(n12193), .C2(n12061), .A(n12060), .B(n12059), .ZN(
        n12062) );
  OAI211_X1 U14534 ( .C1(n12065), .C2(n12064), .A(n12063), .B(n12062), .ZN(
        P3_U3160) );
  OAI211_X1 U14535 ( .C1(n12068), .C2(n12067), .A(n12066), .B(n12203), .ZN(
        n12074) );
  INV_X1 U14536 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15338) );
  NOR2_X1 U14537 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15338), .ZN(n14951) );
  AOI21_X1 U14538 ( .B1(n12193), .B2(n12069), .A(n14951), .ZN(n12073) );
  AOI22_X1 U14539 ( .A1(n12229), .A2(n12189), .B1(n12211), .B2(n15044), .ZN(
        n12072) );
  NAND2_X1 U14540 ( .A1(n12217), .A2(n12070), .ZN(n12071) );
  NAND4_X1 U14541 ( .A1(n12074), .A2(n12073), .A3(n12072), .A4(n12071), .ZN(
        P3_U3153) );
  AOI21_X1 U14542 ( .B1(n12509), .B2(n12075), .A(n6517), .ZN(n12080) );
  AOI22_X1 U14543 ( .A1(n12496), .A2(n12189), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12077) );
  NAND2_X1 U14544 ( .A1(n12502), .A2(n12217), .ZN(n12076) );
  OAI211_X1 U14545 ( .C1(n7366), .C2(n12187), .A(n12077), .B(n12076), .ZN(
        n12078) );
  AOI21_X1 U14546 ( .B1(n12501), .B2(n12193), .A(n12078), .ZN(n12079) );
  OAI21_X1 U14547 ( .B1(n12080), .B2(n12219), .A(n12079), .ZN(P3_U3156) );
  XNOR2_X1 U14548 ( .A(n12081), .B(n12082), .ZN(n12087) );
  NAND2_X1 U14549 ( .A1(n12584), .A2(n12189), .ZN(n12083) );
  NAND2_X1 U14550 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12392)
         );
  OAI211_X1 U14551 ( .C1(n12522), .C2(n12187), .A(n12083), .B(n12392), .ZN(
        n12085) );
  NOR2_X1 U14552 ( .A1(n12556), .A2(n12214), .ZN(n12084) );
  AOI211_X1 U14553 ( .C1(n12554), .C2(n12217), .A(n12085), .B(n12084), .ZN(
        n12086) );
  OAI21_X1 U14554 ( .B1(n12087), .B2(n12219), .A(n12086), .ZN(P3_U3159) );
  OAI211_X1 U14555 ( .C1(n12090), .C2(n12089), .A(n12088), .B(n12203), .ZN(
        n12097) );
  AOI21_X1 U14556 ( .B1(n12193), .B2(n12092), .A(n12091), .ZN(n12096) );
  AOI22_X1 U14557 ( .A1(n12228), .A2(n12189), .B1(n12211), .B2(n15024), .ZN(
        n12095) );
  NAND2_X1 U14558 ( .A1(n12217), .A2(n12093), .ZN(n12094) );
  NAND4_X1 U14559 ( .A1(n12097), .A2(n12096), .A3(n12095), .A4(n12094), .ZN(
        P3_U3161) );
  AOI21_X1 U14560 ( .B1(n12099), .B2(n12098), .A(n6562), .ZN(n12104) );
  AOI22_X1 U14561 ( .A1(n12548), .A2(n12189), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12101) );
  NAND2_X1 U14562 ( .A1(n12217), .A2(n12527), .ZN(n12100) );
  OAI211_X1 U14563 ( .C1(n12523), .C2(n12187), .A(n12101), .B(n12100), .ZN(
        n12102) );
  AOI21_X1 U14564 ( .B1(n12526), .B2(n12193), .A(n12102), .ZN(n12103) );
  OAI21_X1 U14565 ( .B1(n12104), .B2(n12219), .A(n12103), .ZN(P3_U3163) );
  XNOR2_X1 U14566 ( .A(n12105), .B(n12106), .ZN(n12174) );
  OAI22_X1 U14567 ( .A1(n12174), .A2(n15025), .B1(n12105), .B2(n12106), .ZN(
        n12109) );
  XNOR2_X1 U14568 ( .A(n12107), .B(n14356), .ZN(n12108) );
  XNOR2_X1 U14569 ( .A(n12109), .B(n12108), .ZN(n12117) );
  NOR2_X1 U14570 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12110), .ZN(n14995) );
  AOI21_X1 U14571 ( .B1(n15025), .B2(n12189), .A(n14995), .ZN(n12115) );
  OR2_X1 U14572 ( .A1(n14366), .A2(n12214), .ZN(n12114) );
  NAND2_X1 U14573 ( .A1(n12217), .A2(n12111), .ZN(n12113) );
  NAND2_X1 U14574 ( .A1(n12226), .A2(n12211), .ZN(n12112) );
  NAND4_X1 U14575 ( .A1(n12115), .A2(n12114), .A3(n12113), .A4(n12112), .ZN(
        n12116) );
  AOI21_X1 U14576 ( .B1(n12117), .B2(n12203), .A(n12116), .ZN(n12118) );
  INV_X1 U14577 ( .A(n12118), .ZN(P3_U3164) );
  XNOR2_X1 U14578 ( .A(n12119), .B(n8315), .ZN(n12210) );
  AOI22_X1 U14579 ( .A1(n12210), .A2(n12120), .B1(n12620), .B2(n12119), .ZN(
        n12125) );
  INV_X1 U14580 ( .A(n12121), .ZN(n12122) );
  NOR2_X1 U14581 ( .A1(n12123), .A2(n12122), .ZN(n12124) );
  XNOR2_X1 U14582 ( .A(n12125), .B(n12124), .ZN(n12131) );
  NAND2_X1 U14583 ( .A1(n12211), .A2(n12570), .ZN(n12126) );
  NAND2_X1 U14584 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12328)
         );
  OAI211_X1 U14585 ( .C1(n12620), .C2(n12213), .A(n12126), .B(n12328), .ZN(
        n12129) );
  INV_X1 U14586 ( .A(n12127), .ZN(n12748) );
  NOR2_X1 U14587 ( .A1(n12748), .A2(n12214), .ZN(n12128) );
  AOI211_X1 U14588 ( .C1(n12602), .C2(n12217), .A(n12129), .B(n12128), .ZN(
        n12130) );
  OAI21_X1 U14589 ( .B1(n12131), .B2(n12219), .A(n12130), .ZN(P3_U3166) );
  XNOR2_X1 U14590 ( .A(n12133), .B(n12132), .ZN(n12138) );
  NOR2_X1 U14591 ( .A1(n15255), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12352) );
  AOI21_X1 U14592 ( .B1(n12584), .B2(n12211), .A(n12352), .ZN(n12134) );
  OAI21_X1 U14593 ( .B1(n12610), .B2(n12213), .A(n12134), .ZN(n12136) );
  NOR2_X1 U14594 ( .A1(n12689), .A2(n12214), .ZN(n12135) );
  AOI211_X1 U14595 ( .C1(n12591), .C2(n12217), .A(n12136), .B(n12135), .ZN(
        n12137) );
  OAI21_X1 U14596 ( .B1(n12138), .B2(n12219), .A(n12137), .ZN(P3_U3168) );
  INV_X1 U14597 ( .A(n12139), .ZN(n12141) );
  NOR3_X1 U14598 ( .A1(n6517), .A2(n12141), .A3(n12140), .ZN(n12144) );
  INV_X1 U14599 ( .A(n12142), .ZN(n12143) );
  INV_X1 U14600 ( .A(n12490), .ZN(n12146) );
  AOI22_X1 U14601 ( .A1(n12509), .A2(n12189), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12145) );
  OAI21_X1 U14602 ( .B1(n12146), .B2(n12191), .A(n12145), .ZN(n12147) );
  AOI21_X1 U14603 ( .B1(n12224), .B2(n12211), .A(n12147), .ZN(n12148) );
  OAI211_X1 U14604 ( .C1(n12214), .C2(n12725), .A(n12149), .B(n12148), .ZN(
        P3_U3169) );
  XNOR2_X1 U14605 ( .A(n12151), .B(n12150), .ZN(n12156) );
  AOI22_X1 U14606 ( .A1(n12508), .A2(n12211), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12153) );
  NAND2_X1 U14607 ( .A1(n12217), .A2(n12542), .ZN(n12152) );
  OAI211_X1 U14608 ( .C1(n12534), .C2(n12213), .A(n12153), .B(n12152), .ZN(
        n12154) );
  AOI21_X1 U14609 ( .B1(n12536), .B2(n12193), .A(n12154), .ZN(n12155) );
  OAI21_X1 U14610 ( .B1(n12156), .B2(n12219), .A(n12155), .ZN(P3_U3173) );
  XNOR2_X1 U14611 ( .A(n12157), .B(n12226), .ZN(n12158) );
  XNOR2_X1 U14612 ( .A(n12159), .B(n12158), .ZN(n12164) );
  NOR2_X1 U14613 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7689), .ZN(n12259) );
  AOI21_X1 U14614 ( .B1(n12211), .B2(n12225), .A(n12259), .ZN(n12160) );
  OAI21_X1 U14615 ( .B1(n14356), .B2(n12213), .A(n12160), .ZN(n12162) );
  NOR2_X1 U14616 ( .A1(n14357), .A2(n12214), .ZN(n12161) );
  AOI211_X1 U14617 ( .C1(n14358), .C2(n12217), .A(n12162), .B(n12161), .ZN(
        n12163) );
  OAI21_X1 U14618 ( .B1(n12164), .B2(n12219), .A(n12163), .ZN(P3_U3174) );
  INV_X1 U14619 ( .A(n12165), .ZN(n12166) );
  AOI21_X1 U14620 ( .B1(n12496), .B2(n12167), .A(n12166), .ZN(n12172) );
  AOI22_X1 U14621 ( .A1(n12508), .A2(n12189), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12169) );
  NAND2_X1 U14622 ( .A1(n12513), .A2(n12217), .ZN(n12168) );
  OAI211_X1 U14623 ( .C1(n12479), .C2(n12187), .A(n12169), .B(n12168), .ZN(
        n12170) );
  AOI21_X1 U14624 ( .B1(n12665), .B2(n12193), .A(n12170), .ZN(n12171) );
  OAI21_X1 U14625 ( .B1(n12172), .B2(n12219), .A(n12171), .ZN(P3_U3175) );
  XNOR2_X1 U14626 ( .A(n12174), .B(n12173), .ZN(n12183) );
  NAND2_X1 U14627 ( .A1(n12217), .A2(n12175), .ZN(n12178) );
  AOI21_X1 U14628 ( .B1(n12211), .B2(n12227), .A(n12176), .ZN(n12177) );
  OAI211_X1 U14629 ( .C1(n12179), .C2(n12213), .A(n12178), .B(n12177), .ZN(
        n12180) );
  AOI21_X1 U14630 ( .B1(n12181), .B2(n12193), .A(n12180), .ZN(n12182) );
  OAI21_X1 U14631 ( .B1(n12183), .B2(n12219), .A(n12182), .ZN(P3_U3176) );
  XNOR2_X1 U14632 ( .A(n12185), .B(n12184), .ZN(n12195) );
  INV_X1 U14633 ( .A(n12186), .ZN(n12574) );
  NAND2_X1 U14634 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12368)
         );
  OAI21_X1 U14635 ( .B1(n12187), .B2(n12534), .A(n12368), .ZN(n12188) );
  AOI21_X1 U14636 ( .B1(n12189), .B2(n12570), .A(n12188), .ZN(n12190) );
  OAI21_X1 U14637 ( .B1(n12574), .B2(n12191), .A(n12190), .ZN(n12192) );
  AOI21_X1 U14638 ( .B1(n12681), .B2(n12193), .A(n12192), .ZN(n12194) );
  OAI21_X1 U14639 ( .B1(n12195), .B2(n12219), .A(n12194), .ZN(P3_U3178) );
  INV_X1 U14640 ( .A(n12648), .ZN(n12461) );
  NAND2_X1 U14641 ( .A1(n12197), .A2(n12196), .ZN(n12201) );
  AND2_X1 U14642 ( .A1(n12199), .A2(n12198), .ZN(n12200) );
  OAI21_X1 U14643 ( .B1(n12202), .B2(n12201), .A(n12200), .ZN(n12204) );
  NAND2_X1 U14644 ( .A1(n12204), .A2(n12203), .ZN(n12208) );
  AOI22_X1 U14645 ( .A1(n12459), .A2(n12217), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12205) );
  OAI21_X1 U14646 ( .B1(n12480), .B2(n12213), .A(n12205), .ZN(n12206) );
  AOI21_X1 U14647 ( .B1(n12425), .B2(n12211), .A(n12206), .ZN(n12207) );
  OAI211_X1 U14648 ( .C1(n12461), .C2(n12214), .A(n12208), .B(n12207), .ZN(
        P3_U3180) );
  XNOR2_X1 U14649 ( .A(n12210), .B(n12209), .ZN(n12220) );
  NAND2_X1 U14650 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12299)
         );
  NAND2_X1 U14651 ( .A1(n12211), .A2(n12583), .ZN(n12212) );
  OAI211_X1 U14652 ( .C1(n14355), .C2(n12213), .A(n12299), .B(n12212), .ZN(
        n12216) );
  NOR2_X1 U14653 ( .A1(n12752), .A2(n12214), .ZN(n12215) );
  AOI211_X1 U14654 ( .C1(n12613), .C2(n12217), .A(n12216), .B(n12215), .ZN(
        n12218) );
  OAI21_X1 U14655 ( .B1(n12220), .B2(n12219), .A(n12218), .ZN(P3_U3181) );
  MUX2_X1 U14656 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12407), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14657 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12221), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14658 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12222), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14659 ( .A(n12425), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12235), .Z(
        P3_U3518) );
  MUX2_X1 U14660 ( .A(n12223), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12235), .Z(
        P3_U3517) );
  MUX2_X1 U14661 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12224), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14662 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12469), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14663 ( .A(n12509), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12235), .Z(
        P3_U3514) );
  MUX2_X1 U14664 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12496), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14665 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12508), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14666 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12548), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14667 ( .A(n12571), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12235), .Z(
        P3_U3510) );
  MUX2_X1 U14668 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12584), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14669 ( .A(n12570), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12235), .Z(
        P3_U3508) );
  MUX2_X1 U14670 ( .A(n12583), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12235), .Z(
        P3_U3507) );
  MUX2_X1 U14671 ( .A(n8315), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12235), .Z(
        P3_U3506) );
  MUX2_X1 U14672 ( .A(n12225), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12235), .Z(
        P3_U3505) );
  MUX2_X1 U14673 ( .A(n12226), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12235), .Z(
        P3_U3504) );
  MUX2_X1 U14674 ( .A(n12227), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12235), .Z(
        P3_U3503) );
  MUX2_X1 U14675 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n15025), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14676 ( .A(n8302), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12235), .Z(
        P3_U3501) );
  MUX2_X1 U14677 ( .A(n15024), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12235), .Z(
        P3_U3500) );
  MUX2_X1 U14678 ( .A(n15044), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12235), .Z(
        P3_U3499) );
  MUX2_X1 U14679 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12228), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14680 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12229), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14681 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12230), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14682 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12231), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14683 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12232), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14684 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12233), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14685 ( .A(n12234), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12235), .Z(
        P3_U3492) );
  MUX2_X1 U14686 ( .A(n15094), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12235), .Z(
        P3_U3491) );
  INV_X1 U14687 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14360) );
  NAND2_X1 U14688 ( .A1(n12253), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12239) );
  INV_X1 U14689 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U14690 ( .A1(n14992), .A2(n12237), .ZN(n12238) );
  AND2_X1 U14691 ( .A1(n12239), .A2(n12238), .ZN(n14998) );
  AOI21_X1 U14692 ( .B1(n14360), .B2(n12240), .A(n12274), .ZN(n12266) );
  INV_X1 U14693 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14365) );
  INV_X1 U14694 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U14695 ( .A1(n14992), .A2(n12244), .ZN(n12243) );
  OAI21_X1 U14696 ( .B1(n14992), .B2(n12244), .A(n12243), .ZN(n15003) );
  INV_X1 U14697 ( .A(n15003), .ZN(n12245) );
  NAND2_X1 U14698 ( .A1(n14992), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12246) );
  AOI21_X1 U14699 ( .B1(n14365), .B2(n12247), .A(n12268), .ZN(n12248) );
  NOR2_X1 U14700 ( .A1(n12248), .A2(n14977), .ZN(n12264) );
  MUX2_X1 U14701 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12369), .Z(n12281) );
  XNOR2_X1 U14702 ( .A(n12281), .B(n12280), .ZN(n12257) );
  MUX2_X1 U14703 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12369), .Z(n12254) );
  NAND2_X1 U14704 ( .A1(n12254), .A2(n14992), .ZN(n12255) );
  INV_X1 U14705 ( .A(n12249), .ZN(n12252) );
  XNOR2_X1 U14706 ( .A(n12254), .B(n12253), .ZN(n15009) );
  NAND2_X1 U14707 ( .A1(n12257), .A2(n12256), .ZN(n12258) );
  AOI21_X1 U14708 ( .B1(n12258), .B2(n7133), .A(n14911), .ZN(n12263) );
  INV_X1 U14709 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U14710 ( .A1(n14983), .A2(n7163), .ZN(n12261) );
  INV_X1 U14711 ( .A(n12259), .ZN(n12260) );
  OAI211_X1 U14712 ( .C1(n14258), .C2(n14974), .A(n12261), .B(n12260), .ZN(
        n12262) );
  NOR3_X1 U14713 ( .A1(n12264), .A2(n12263), .A3(n12262), .ZN(n12265) );
  OAI21_X1 U14714 ( .B1(n12266), .B2(n14990), .A(n12265), .ZN(P3_U3195) );
  NOR2_X1 U14715 ( .A1(n7163), .A2(n12267), .ZN(n12269) );
  NAND2_X1 U14716 ( .A1(n12289), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12300) );
  OR2_X1 U14717 ( .A1(n12289), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U14718 ( .A1(n12300), .A2(n12270), .ZN(n12282) );
  NAND2_X1 U14719 ( .A1(n12271), .A2(n12282), .ZN(n12272) );
  AOI21_X1 U14720 ( .B1(n12292), .B2(n12272), .A(n14977), .ZN(n12291) );
  NOR2_X1 U14721 ( .A1(n7163), .A2(n12273), .ZN(n12275) );
  NAND2_X1 U14722 ( .A1(n12289), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12301) );
  OR2_X1 U14723 ( .A1(n12289), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12276) );
  NAND2_X1 U14724 ( .A1(n12301), .A2(n12276), .ZN(n12294) );
  XNOR2_X1 U14725 ( .A(n12295), .B(n12294), .ZN(n12279) );
  INV_X1 U14726 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14261) );
  NOR2_X1 U14727 ( .A1(n14974), .A2(n14261), .ZN(n12277) );
  AOI211_X1 U14728 ( .C1(n12279), .C2(n14997), .A(n12278), .B(n12277), .ZN(
        n12288) );
  NOR2_X1 U14729 ( .A1(n12281), .A2(n12280), .ZN(n12285) );
  MUX2_X1 U14730 ( .A(n12294), .B(n12282), .S(n12369), .Z(n12284) );
  OAI21_X1 U14731 ( .B1(n12285), .B2(n12283), .A(n12284), .ZN(n12286) );
  NAND3_X1 U14732 ( .A1(n12286), .A2(n15007), .A3(n12303), .ZN(n12287) );
  OAI211_X1 U14733 ( .C1(n14993), .C2(n12289), .A(n12288), .B(n12287), .ZN(
        n12290) );
  OR2_X1 U14734 ( .A1(n12291), .A2(n12290), .ZN(P3_U3196) );
  INV_X1 U14735 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12698) );
  AOI21_X1 U14736 ( .B1(n12698), .B2(n12293), .A(n12332), .ZN(n12314) );
  INV_X1 U14737 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12297) );
  AOI21_X1 U14738 ( .B1(n12297), .B2(n12296), .A(n12318), .ZN(n12298) );
  OR2_X1 U14739 ( .A1(n12298), .A2(n14990), .ZN(n12313) );
  INV_X1 U14740 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14324) );
  OAI21_X1 U14741 ( .B1(n14974), .B2(n14324), .A(n12299), .ZN(n12311) );
  MUX2_X1 U14742 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12369), .Z(n12308) );
  MUX2_X1 U14743 ( .A(n12301), .B(n12300), .S(n12369), .Z(n12302) );
  AOI21_X1 U14744 ( .B1(n12305), .B2(n12304), .A(n12323), .ZN(n12306) );
  AOI21_X1 U14745 ( .B1(n12308), .B2(n12307), .A(n12322), .ZN(n12309) );
  NOR2_X1 U14746 ( .A1(n12309), .A2(n14911), .ZN(n12310) );
  AOI211_X1 U14747 ( .C1(n14983), .C2(n12331), .A(n12311), .B(n12310), .ZN(
        n12312) );
  OAI211_X1 U14748 ( .C1(n12314), .C2(n14977), .A(n12313), .B(n12312), .ZN(
        P3_U3197) );
  NAND2_X1 U14749 ( .A1(n12333), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12315) );
  OAI21_X1 U14750 ( .B1(n12333), .B2(P3_REG2_REG_16__SCAN_IN), .A(n12315), 
        .ZN(n12316) );
  INV_X1 U14751 ( .A(n12316), .ZN(n12321) );
  INV_X1 U14752 ( .A(n12349), .ZN(n12319) );
  AOI21_X1 U14753 ( .B1(n12321), .B2(n12320), .A(n12319), .ZN(n12342) );
  INV_X1 U14754 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12324) );
  INV_X1 U14755 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12694) );
  MUX2_X1 U14756 ( .A(n12324), .B(n12694), .S(n12369), .Z(n12325) );
  NAND2_X1 U14757 ( .A1(n12325), .A2(n12333), .ZN(n12355) );
  MUX2_X1 U14758 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12369), .Z(n12326) );
  NAND2_X1 U14759 ( .A1(n12355), .A2(n6640), .ZN(n12327) );
  XNOR2_X1 U14760 ( .A(n12356), .B(n12327), .ZN(n12340) );
  INV_X1 U14761 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14228) );
  NAND2_X1 U14762 ( .A1(n14983), .A2(n12333), .ZN(n12329) );
  OAI211_X1 U14763 ( .C1(n14228), .C2(n14974), .A(n12329), .B(n12328), .ZN(
        n12339) );
  NAND2_X1 U14764 ( .A1(n12347), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12343) );
  NAND2_X1 U14765 ( .A1(n12333), .A2(n12694), .ZN(n12334) );
  NAND2_X1 U14766 ( .A1(n12343), .A2(n12334), .ZN(n12335) );
  NAND2_X1 U14767 ( .A1(n12336), .A2(n12335), .ZN(n12337) );
  AOI21_X1 U14768 ( .B1(n12344), .B2(n12337), .A(n14977), .ZN(n12338) );
  AOI211_X1 U14769 ( .C1(n15007), .C2(n12340), .A(n12339), .B(n12338), .ZN(
        n12341) );
  OAI21_X1 U14770 ( .B1(n12342), .B2(n14990), .A(n12341), .ZN(P3_U3198) );
  INV_X1 U14771 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12346) );
  AOI21_X1 U14772 ( .B1(n12346), .B2(n12345), .A(n12377), .ZN(n12362) );
  NAND2_X1 U14773 ( .A1(n12347), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12348) );
  INV_X1 U14774 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12350) );
  AOI21_X1 U14775 ( .B1(n12351), .B2(n12350), .A(n12364), .ZN(n12354) );
  AOI21_X1 U14776 ( .B1(n14996), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12352), 
        .ZN(n12353) );
  OAI21_X1 U14777 ( .B1(n14990), .B2(n12354), .A(n12353), .ZN(n12360) );
  MUX2_X1 U14778 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12369), .Z(n12372) );
  XNOR2_X1 U14779 ( .A(n12372), .B(n12371), .ZN(n12357) );
  NOR2_X1 U14780 ( .A1(n12358), .A2(n12357), .ZN(n12370) );
  AOI211_X1 U14781 ( .C1(n12358), .C2(n12357), .A(n12370), .B(n14911), .ZN(
        n12359) );
  AOI211_X1 U14782 ( .C1(n14983), .C2(n7035), .A(n12360), .B(n12359), .ZN(
        n12361) );
  OAI21_X1 U14783 ( .B1(n12362), .B2(n14977), .A(n12361), .ZN(P3_U3199) );
  NOR2_X1 U14784 ( .A1(n7035), .A2(n12363), .ZN(n12365) );
  NOR2_X1 U14785 ( .A1(n12365), .A2(n12364), .ZN(n12367) );
  NAND2_X1 U14786 ( .A1(n12378), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12387) );
  OAI21_X1 U14787 ( .B1(n12378), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12387), 
        .ZN(n12366) );
  NOR2_X1 U14788 ( .A1(n12367), .A2(n12366), .ZN(n12389) );
  AOI21_X1 U14789 ( .B1(n12367), .B2(n12366), .A(n12389), .ZN(n12381) );
  INV_X1 U14790 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15187) );
  OAI21_X1 U14791 ( .B1(n14974), .B2(n15187), .A(n12368), .ZN(n12375) );
  MUX2_X1 U14792 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12369), .Z(n12374) );
  XNOR2_X1 U14793 ( .A(n12396), .B(n12395), .ZN(n12373) );
  NOR2_X1 U14794 ( .A1(n12373), .A2(n12374), .ZN(n12394) );
  NAND2_X1 U14795 ( .A1(n12378), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12382) );
  OAI21_X1 U14796 ( .B1(n12378), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12382), 
        .ZN(n12379) );
  INV_X1 U14797 ( .A(n12382), .ZN(n12383) );
  NOR2_X1 U14798 ( .A1(n12384), .A2(n12383), .ZN(n12385) );
  XNOR2_X1 U14799 ( .A(n6480), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12399) );
  XNOR2_X1 U14800 ( .A(n12385), .B(n12399), .ZN(n12405) );
  INV_X1 U14801 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12386) );
  MUX2_X1 U14802 ( .A(n12386), .B(P3_REG2_REG_19__SCAN_IN), .S(n6480), .Z(
        n12398) );
  INV_X1 U14803 ( .A(n12387), .ZN(n12388) );
  NOR2_X1 U14804 ( .A1(n12389), .A2(n12388), .ZN(n12390) );
  XOR2_X1 U14805 ( .A(n12398), .B(n12390), .Z(n12391) );
  NAND2_X1 U14806 ( .A1(n12391), .A2(n14997), .ZN(n12404) );
  INV_X1 U14807 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n12393) );
  OAI21_X1 U14808 ( .B1(n14974), .B2(n12393), .A(n12392), .ZN(n12401) );
  MUX2_X1 U14809 ( .A(n12399), .B(n12398), .S(n6812), .Z(n12400) );
  OAI211_X1 U14810 ( .C1(n12405), .C2(n14977), .A(n12404), .B(n12403), .ZN(
        P3_U3201) );
  NAND2_X1 U14811 ( .A1(n12407), .A2(n12406), .ZN(n12708) );
  NAND2_X1 U14812 ( .A1(n12408), .A2(n15102), .ZN(n12414) );
  OAI21_X1 U14813 ( .B1(n12708), .B2(n15068), .A(n12414), .ZN(n12410) );
  AOI21_X1 U14814 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15068), .A(n12410), 
        .ZN(n12409) );
  OAI21_X1 U14815 ( .B1(n12710), .B2(n15049), .A(n12409), .ZN(P3_U3202) );
  AOI21_X1 U14816 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15068), .A(n12410), 
        .ZN(n12411) );
  OAI21_X1 U14817 ( .B1(n12713), .B2(n15049), .A(n12411), .ZN(P3_U3203) );
  INV_X1 U14818 ( .A(n12412), .ZN(n12419) );
  OAI21_X1 U14819 ( .B1(n15107), .B2(n12415), .A(n12414), .ZN(n12416) );
  AOI21_X1 U14820 ( .B1(n12417), .B2(n12627), .A(n12416), .ZN(n12418) );
  NAND2_X1 U14821 ( .A1(n12436), .A2(n12420), .ZN(n12422) );
  XNOR2_X1 U14822 ( .A(n12422), .B(n12421), .ZN(n12642) );
  INV_X1 U14823 ( .A(n12642), .ZN(n12432) );
  AOI22_X1 U14824 ( .A1(n12428), .A2(n15102), .B1(n15068), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12429) );
  OAI21_X1 U14825 ( .B1(n12716), .B2(n15049), .A(n12429), .ZN(n12430) );
  AOI21_X1 U14826 ( .B1(n12641), .B2(n15107), .A(n12430), .ZN(n12431) );
  OAI21_X1 U14827 ( .B1(n12432), .B2(n12579), .A(n12431), .ZN(P3_U3205) );
  OR2_X1 U14828 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  OAI22_X1 U14829 ( .A1(n12440), .A2(n15096), .B1(n12472), .B2(n15072), .ZN(
        n12441) );
  AOI22_X1 U14830 ( .A1(n12443), .A2(n15102), .B1(n15068), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12446) );
  NAND2_X1 U14831 ( .A1(n12444), .A2(n12627), .ZN(n12445) );
  OAI211_X1 U14832 ( .C1(n12644), .C2(n12447), .A(n12446), .B(n12445), .ZN(
        n12448) );
  AOI21_X1 U14833 ( .B1(n12645), .B2(n15107), .A(n12448), .ZN(n12449) );
  INV_X1 U14834 ( .A(n12449), .ZN(P3_U3206) );
  XOR2_X1 U14835 ( .A(n12450), .B(n12451), .Z(n12457) );
  XNOR2_X1 U14836 ( .A(n12452), .B(n12451), .ZN(n12458) );
  NOR2_X1 U14837 ( .A1(n12458), .A2(n12453), .ZN(n12456) );
  OAI22_X1 U14838 ( .A1(n12454), .A2(n15096), .B1(n12480), .B2(n15072), .ZN(
        n12455) );
  INV_X1 U14839 ( .A(n12458), .ZN(n12649) );
  AOI22_X1 U14840 ( .A1(n12459), .A2(n15102), .B1(n15068), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12460) );
  OAI21_X1 U14841 ( .B1(n12461), .B2(n15049), .A(n12460), .ZN(n12462) );
  AOI21_X1 U14842 ( .B1(n12649), .B2(n15030), .A(n12462), .ZN(n12463) );
  OAI21_X1 U14843 ( .B1(n12651), .B2(n15068), .A(n12463), .ZN(P3_U3207) );
  XNOR2_X1 U14844 ( .A(n12464), .B(n12467), .ZN(n12655) );
  NAND2_X1 U14845 ( .A1(n12478), .A2(n12486), .ZN(n12477) );
  NAND2_X1 U14846 ( .A1(n12477), .A2(n12465), .ZN(n12468) );
  OAI211_X1 U14847 ( .C1(n12468), .C2(n12467), .A(n12466), .B(n15099), .ZN(
        n12471) );
  NAND2_X1 U14848 ( .A1(n12469), .A2(n15093), .ZN(n12470) );
  OAI211_X1 U14849 ( .C1(n12472), .C2(n15096), .A(n12471), .B(n12470), .ZN(
        n12652) );
  AOI22_X1 U14850 ( .A1(n12473), .A2(n15102), .B1(n15068), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12474) );
  OAI21_X1 U14851 ( .B1(n8397), .B2(n15049), .A(n12474), .ZN(n12475) );
  AOI21_X1 U14852 ( .B1(n12652), .B2(n15107), .A(n12475), .ZN(n12476) );
  OAI21_X1 U14853 ( .B1(n12579), .B2(n12655), .A(n12476), .ZN(P3_U3208) );
  OAI211_X1 U14854 ( .C1(n12486), .C2(n12478), .A(n12477), .B(n15099), .ZN(
        n12483) );
  OAI22_X1 U14855 ( .A1(n12480), .A2(n15096), .B1(n12479), .B2(n15072), .ZN(
        n12481) );
  INV_X1 U14856 ( .A(n12481), .ZN(n12482) );
  AND2_X1 U14857 ( .A1(n12483), .A2(n12482), .ZN(n12658) );
  NAND2_X1 U14858 ( .A1(n12485), .A2(n12484), .ZN(n12487) );
  NAND2_X1 U14859 ( .A1(n12487), .A2(n12486), .ZN(n12489) );
  NAND2_X1 U14860 ( .A1(n12489), .A2(n12488), .ZN(n12656) );
  AOI22_X1 U14861 ( .A1(n12490), .A2(n15102), .B1(n15068), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12491) );
  OAI21_X1 U14862 ( .B1(n12725), .B2(n15049), .A(n12491), .ZN(n12492) );
  AOI21_X1 U14863 ( .B1(n12656), .B2(n15065), .A(n12492), .ZN(n12493) );
  OAI21_X1 U14864 ( .B1(n12658), .B2(n15068), .A(n12493), .ZN(P3_U3209) );
  OAI211_X1 U14865 ( .C1(n12495), .C2(n8130), .A(n12494), .B(n15099), .ZN(
        n12498) );
  NAND2_X1 U14866 ( .A1(n12496), .A2(n15093), .ZN(n12497) );
  OAI211_X1 U14867 ( .C1(n7366), .C2(n15096), .A(n12498), .B(n12497), .ZN(
        n12661) );
  INV_X1 U14868 ( .A(n12661), .ZN(n12506) );
  XOR2_X1 U14869 ( .A(n12500), .B(n12499), .Z(n12662) );
  INV_X1 U14870 ( .A(n12501), .ZN(n12729) );
  AOI22_X1 U14871 ( .A1(n12502), .A2(n15102), .B1(n15068), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12503) );
  OAI21_X1 U14872 ( .B1(n12729), .B2(n15049), .A(n12503), .ZN(n12504) );
  AOI21_X1 U14873 ( .B1(n12662), .B2(n15065), .A(n12504), .ZN(n12505) );
  OAI21_X1 U14874 ( .B1(n12506), .B2(n15068), .A(n12505), .ZN(P3_U3210) );
  XOR2_X1 U14875 ( .A(n12507), .B(n12511), .Z(n12510) );
  AOI222_X1 U14876 ( .A1(n15099), .A2(n12510), .B1(n12509), .B2(n15045), .C1(
        n12508), .C2(n15093), .ZN(n12667) );
  XNOR2_X1 U14877 ( .A(n12512), .B(n12511), .ZN(n12668) );
  AOI22_X1 U14878 ( .A1(n12513), .A2(n15102), .B1(n15068), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n12515) );
  NAND2_X1 U14879 ( .A1(n12665), .A2(n12627), .ZN(n12514) );
  OAI211_X1 U14880 ( .C1(n12668), .C2(n12579), .A(n12515), .B(n12514), .ZN(
        n12516) );
  INV_X1 U14881 ( .A(n12516), .ZN(n12517) );
  OAI21_X1 U14882 ( .B1(n12667), .B2(n15068), .A(n12517), .ZN(P3_U3211) );
  INV_X1 U14883 ( .A(n12518), .ZN(n12519) );
  AOI21_X1 U14884 ( .B1(n12524), .B2(n12520), .A(n12519), .ZN(n12521) );
  OAI222_X1 U14885 ( .A1(n15096), .A2(n12523), .B1(n15072), .B2(n12522), .C1(
        n15075), .C2(n12521), .ZN(n12669) );
  INV_X1 U14886 ( .A(n12669), .ZN(n12531) );
  XOR2_X1 U14887 ( .A(n12525), .B(n12524), .Z(n12670) );
  INV_X1 U14888 ( .A(n12526), .ZN(n12734) );
  AOI22_X1 U14889 ( .A1(n15068), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12527), 
        .B2(n15102), .ZN(n12528) );
  OAI21_X1 U14890 ( .B1(n12734), .B2(n15049), .A(n12528), .ZN(n12529) );
  AOI21_X1 U14891 ( .B1(n12670), .B2(n15065), .A(n12529), .ZN(n12530) );
  OAI21_X1 U14892 ( .B1(n12531), .B2(n15068), .A(n12530), .ZN(P3_U3212) );
  XNOR2_X1 U14893 ( .A(n12532), .B(n12538), .ZN(n12533) );
  OAI222_X1 U14894 ( .A1(n15096), .A2(n12535), .B1(n15072), .B2(n12534), .C1(
        n12533), .C2(n15075), .ZN(n12673) );
  INV_X1 U14895 ( .A(n12536), .ZN(n12738) );
  NAND2_X1 U14896 ( .A1(n12550), .A2(n12537), .ZN(n12539) );
  NAND2_X1 U14897 ( .A1(n12539), .A2(n12538), .ZN(n12541) );
  AND2_X1 U14898 ( .A1(n12541), .A2(n12540), .ZN(n12674) );
  NAND2_X1 U14899 ( .A1(n12674), .A2(n15065), .ZN(n12544) );
  AOI22_X1 U14900 ( .A1(n15068), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15102), 
        .B2(n12542), .ZN(n12543) );
  OAI211_X1 U14901 ( .C1(n12738), .C2(n15049), .A(n12544), .B(n12543), .ZN(
        n12545) );
  AOI21_X1 U14902 ( .B1(n12673), .B2(n15107), .A(n12545), .ZN(n12546) );
  INV_X1 U14903 ( .A(n12546), .ZN(P3_U3213) );
  XNOR2_X1 U14904 ( .A(n12547), .B(n12552), .ZN(n12549) );
  AOI222_X1 U14905 ( .A1(n15099), .A2(n12549), .B1(n12548), .B2(n15045), .C1(
        n12584), .C2(n15093), .ZN(n12679) );
  INV_X1 U14906 ( .A(n12550), .ZN(n12551) );
  AOI21_X1 U14907 ( .B1(n12553), .B2(n12552), .A(n12551), .ZN(n12680) );
  INV_X1 U14908 ( .A(n12680), .ZN(n12558) );
  AOI22_X1 U14909 ( .A1(n15068), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15102), 
        .B2(n12554), .ZN(n12555) );
  OAI21_X1 U14910 ( .B1(n12556), .B2(n15049), .A(n12555), .ZN(n12557) );
  AOI21_X1 U14911 ( .B1(n12558), .B2(n15065), .A(n12557), .ZN(n12559) );
  OAI21_X1 U14912 ( .B1(n12679), .B2(n15068), .A(n12559), .ZN(P3_U3214) );
  NAND2_X1 U14913 ( .A1(n12590), .A2(n12560), .ZN(n12562) );
  NAND2_X1 U14914 ( .A1(n12562), .A2(n12561), .ZN(n12564) );
  NAND2_X1 U14915 ( .A1(n12564), .A2(n12563), .ZN(n12682) );
  NAND2_X1 U14916 ( .A1(n12566), .A2(n12565), .ZN(n12567) );
  NAND2_X1 U14917 ( .A1(n12568), .A2(n12567), .ZN(n12569) );
  NAND2_X1 U14918 ( .A1(n12569), .A2(n15099), .ZN(n12573) );
  AOI22_X1 U14919 ( .A1(n12571), .A2(n15045), .B1(n12570), .B2(n15093), .ZN(
        n12572) );
  NAND2_X1 U14920 ( .A1(n12573), .A2(n12572), .ZN(n12684) );
  NAND2_X1 U14921 ( .A1(n12684), .A2(n15107), .ZN(n12578) );
  INV_X1 U14922 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12575) );
  OAI22_X1 U14923 ( .A1(n15107), .A2(n12575), .B1(n12574), .B2(n15053), .ZN(
        n12576) );
  AOI21_X1 U14924 ( .B1(n12681), .B2(n12627), .A(n12576), .ZN(n12577) );
  OAI211_X1 U14925 ( .C1(n12682), .C2(n12579), .A(n12578), .B(n12577), .ZN(
        P3_U3215) );
  NAND2_X1 U14926 ( .A1(n12580), .A2(n12587), .ZN(n12581) );
  NAND3_X1 U14927 ( .A1(n12582), .A2(n15099), .A3(n12581), .ZN(n12586) );
  AOI22_X1 U14928 ( .A1(n12584), .A2(n15045), .B1(n15093), .B2(n12583), .ZN(
        n12585) );
  NAND2_X1 U14929 ( .A1(n12586), .A2(n12585), .ZN(n12691) );
  INV_X1 U14930 ( .A(n12691), .ZN(n12595) );
  OR2_X1 U14931 ( .A1(n12588), .A2(n12587), .ZN(n12589) );
  NAND2_X1 U14932 ( .A1(n12590), .A2(n12589), .ZN(n12687) );
  AOI22_X1 U14933 ( .A1(n15068), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15102), 
        .B2(n12591), .ZN(n12592) );
  OAI21_X1 U14934 ( .B1(n12689), .B2(n15049), .A(n12592), .ZN(n12593) );
  AOI21_X1 U14935 ( .B1(n12687), .B2(n15065), .A(n12593), .ZN(n12594) );
  OAI21_X1 U14936 ( .B1(n12595), .B2(n15068), .A(n12594), .ZN(P3_U3216) );
  XOR2_X1 U14937 ( .A(n12596), .B(n12600), .Z(n12597) );
  OAI222_X1 U14938 ( .A1(n15096), .A2(n12598), .B1(n15072), .B2(n12620), .C1(
        n12597), .C2(n15075), .ZN(n12692) );
  INV_X1 U14939 ( .A(n12692), .ZN(n12606) );
  OAI21_X1 U14940 ( .B1(n12601), .B2(n12600), .A(n12599), .ZN(n12693) );
  AOI22_X1 U14941 ( .A1(n15068), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15102), 
        .B2(n12602), .ZN(n12603) );
  OAI21_X1 U14942 ( .B1(n12748), .B2(n15049), .A(n12603), .ZN(n12604) );
  AOI21_X1 U14943 ( .B1(n12693), .B2(n15065), .A(n12604), .ZN(n12605) );
  OAI21_X1 U14944 ( .B1(n12606), .B2(n15068), .A(n12605), .ZN(P3_U3217) );
  XNOR2_X1 U14945 ( .A(n12608), .B(n12607), .ZN(n12609) );
  OAI222_X1 U14946 ( .A1(n15096), .A2(n12610), .B1(n15072), .B2(n14355), .C1(
        n12609), .C2(n15075), .ZN(n12696) );
  INV_X1 U14947 ( .A(n12696), .ZN(n12617) );
  XNOR2_X1 U14948 ( .A(n12612), .B(n12611), .ZN(n12697) );
  AOI22_X1 U14949 ( .A1(n15068), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15102), 
        .B2(n12613), .ZN(n12614) );
  OAI21_X1 U14950 ( .B1(n12752), .B2(n15049), .A(n12614), .ZN(n12615) );
  AOI21_X1 U14951 ( .B1(n12697), .B2(n15065), .A(n12615), .ZN(n12616) );
  OAI21_X1 U14952 ( .B1(n12617), .B2(n15068), .A(n12616), .ZN(P3_U3218) );
  AOI21_X1 U14953 ( .B1(n12618), .B2(n12629), .A(n15075), .ZN(n12623) );
  OAI22_X1 U14954 ( .A1(n12620), .A2(n15096), .B1(n12619), .B2(n15072), .ZN(
        n12621) );
  AOI21_X1 U14955 ( .B1(n12623), .B2(n12622), .A(n12621), .ZN(n12702) );
  INV_X1 U14956 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12625) );
  OAI22_X1 U14957 ( .A1(n15107), .A2(n12625), .B1(n12624), .B2(n15053), .ZN(
        n12626) );
  AOI21_X1 U14958 ( .B1(n12628), .B2(n12627), .A(n12626), .ZN(n12632) );
  XNOR2_X1 U14959 ( .A(n12630), .B(n7564), .ZN(n12700) );
  NAND2_X1 U14960 ( .A1(n12700), .A2(n15065), .ZN(n12631) );
  OAI211_X1 U14961 ( .C1(n12702), .C2(n15068), .A(n12632), .B(n12631), .ZN(
        P3_U3219) );
  INV_X1 U14962 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12636) );
  NAND2_X1 U14963 ( .A1(n12633), .A2(n7570), .ZN(n12635) );
  INV_X1 U14964 ( .A(n12708), .ZN(n12634) );
  NAND2_X1 U14965 ( .A1(n12634), .A2(n15181), .ZN(n12638) );
  OAI211_X1 U14966 ( .C1(n15181), .C2(n12636), .A(n12635), .B(n12638), .ZN(
        P3_U3490) );
  INV_X1 U14967 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U14968 ( .A1(n12637), .A2(n7570), .ZN(n12639) );
  OAI211_X1 U14969 ( .C1(n15181), .C2(n12640), .A(n12639), .B(n12638), .ZN(
        P3_U3489) );
  INV_X1 U14970 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12643) );
  INV_X1 U14971 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12647) );
  INV_X1 U14972 ( .A(n12644), .ZN(n12646) );
  AOI22_X1 U14973 ( .A1(n12649), .A2(n15148), .B1(n15151), .B2(n12648), .ZN(
        n12650) );
  NAND2_X1 U14974 ( .A1(n12651), .A2(n12650), .ZN(n12720) );
  MUX2_X1 U14975 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n12720), .S(n15181), .Z(
        P3_U3485) );
  AOI21_X1 U14976 ( .B1(n15151), .B2(n12653), .A(n12652), .ZN(n12654) );
  OAI21_X1 U14977 ( .B1(n15156), .B2(n12655), .A(n12654), .ZN(n12721) );
  MUX2_X1 U14978 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12721), .S(n15181), .Z(
        P3_U3484) );
  NAND2_X1 U14979 ( .A1(n12656), .A2(n15160), .ZN(n12657) );
  INV_X1 U14980 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12659) );
  MUX2_X1 U14981 ( .A(n12723), .B(n12659), .S(n6961), .Z(n12660) );
  OAI21_X1 U14982 ( .B1(n12705), .B2(n12725), .A(n12660), .ZN(P3_U3483) );
  INV_X1 U14983 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12663) );
  AOI21_X1 U14984 ( .B1(n12662), .B2(n15160), .A(n12661), .ZN(n12726) );
  MUX2_X1 U14985 ( .A(n12663), .B(n12726), .S(n15181), .Z(n12664) );
  OAI21_X1 U14986 ( .B1(n12729), .B2(n12705), .A(n12664), .ZN(P3_U3482) );
  NAND2_X1 U14987 ( .A1(n12665), .A2(n15151), .ZN(n12666) );
  OAI211_X1 U14988 ( .C1(n15156), .C2(n12668), .A(n12667), .B(n12666), .ZN(
        n12730) );
  MUX2_X1 U14989 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n12730), .S(n15181), .Z(
        P3_U3481) );
  INV_X1 U14990 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12671) );
  AOI21_X1 U14991 ( .B1(n15160), .B2(n12670), .A(n12669), .ZN(n12731) );
  MUX2_X1 U14992 ( .A(n12671), .B(n12731), .S(n15181), .Z(n12672) );
  OAI21_X1 U14993 ( .B1(n12734), .B2(n12705), .A(n12672), .ZN(P3_U3480) );
  INV_X1 U14994 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12675) );
  AOI21_X1 U14995 ( .B1(n12674), .B2(n15160), .A(n12673), .ZN(n12735) );
  MUX2_X1 U14996 ( .A(n12675), .B(n12735), .S(n15181), .Z(n12676) );
  OAI21_X1 U14997 ( .B1(n12738), .B2(n12705), .A(n12676), .ZN(P3_U3479) );
  NAND2_X1 U14998 ( .A1(n12677), .A2(n15151), .ZN(n12678) );
  OAI211_X1 U14999 ( .C1(n15156), .C2(n12680), .A(n12679), .B(n12678), .ZN(
        n12739) );
  MUX2_X1 U15000 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12739), .S(n15181), .Z(
        P3_U3478) );
  INV_X1 U15001 ( .A(n12681), .ZN(n12743) );
  INV_X1 U15002 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12685) );
  NOR2_X1 U15003 ( .A1(n12682), .A2(n15156), .ZN(n12683) );
  NOR2_X1 U15004 ( .A1(n12684), .A2(n12683), .ZN(n12740) );
  MUX2_X1 U15005 ( .A(n12685), .B(n12740), .S(n15181), .Z(n12686) );
  OAI21_X1 U15006 ( .B1(n12743), .B2(n12705), .A(n12686), .ZN(P3_U3477) );
  NAND2_X1 U15007 ( .A1(n12687), .A2(n15160), .ZN(n12688) );
  OAI21_X1 U15008 ( .B1(n15131), .B2(n12689), .A(n12688), .ZN(n12690) );
  MUX2_X1 U15009 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12744), .S(n15181), .Z(
        P3_U3476) );
  AOI21_X1 U15010 ( .B1(n15160), .B2(n12693), .A(n12692), .ZN(n12745) );
  MUX2_X1 U15011 ( .A(n12694), .B(n12745), .S(n15181), .Z(n12695) );
  OAI21_X1 U15012 ( .B1(n12748), .B2(n12705), .A(n12695), .ZN(P3_U3475) );
  AOI21_X1 U15013 ( .B1(n12697), .B2(n15160), .A(n12696), .ZN(n12749) );
  MUX2_X1 U15014 ( .A(n12698), .B(n12749), .S(n15181), .Z(n12699) );
  OAI21_X1 U15015 ( .B1(n12705), .B2(n12752), .A(n12699), .ZN(P3_U3474) );
  INV_X1 U15016 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12703) );
  NAND2_X1 U15017 ( .A1(n12700), .A2(n15160), .ZN(n12701) );
  AND2_X1 U15018 ( .A1(n12702), .A2(n12701), .ZN(n12753) );
  MUX2_X1 U15019 ( .A(n12703), .B(n12753), .S(n15181), .Z(n12704) );
  OAI21_X1 U15020 ( .B1(n12705), .B2(n12756), .A(n12704), .ZN(P3_U3473) );
  OAI21_X1 U15021 ( .B1(n12707), .B2(n15131), .A(n12706), .ZN(n12758) );
  MUX2_X1 U15022 ( .A(P3_REG1_REG_0__SCAN_IN), .B(n12758), .S(n15181), .Z(
        P3_U3459) );
  NOR2_X1 U15023 ( .A1(n12708), .A2(n15162), .ZN(n12711) );
  AOI21_X1 U15024 ( .B1(n15162), .B2(P3_REG0_REG_31__SCAN_IN), .A(n12711), 
        .ZN(n12709) );
  OAI21_X1 U15025 ( .B1(n12710), .B2(n12757), .A(n12709), .ZN(P3_U3458) );
  AOI21_X1 U15026 ( .B1(n15162), .B2(P3_REG0_REG_30__SCAN_IN), .A(n12711), 
        .ZN(n12712) );
  OAI21_X1 U15027 ( .B1(n12713), .B2(n12757), .A(n12712), .ZN(P3_U3457) );
  INV_X1 U15028 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12715) );
  INV_X1 U15029 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12718) );
  MUX2_X1 U15030 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n12720), .S(n15164), .Z(
        P3_U3453) );
  MUX2_X1 U15031 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12721), .S(n15164), .Z(
        P3_U3452) );
  INV_X1 U15032 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12722) );
  MUX2_X1 U15033 ( .A(n12723), .B(n12722), .S(n15162), .Z(n12724) );
  OAI21_X1 U15034 ( .B1(n12757), .B2(n12725), .A(n12724), .ZN(P3_U3451) );
  INV_X1 U15035 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12727) );
  MUX2_X1 U15036 ( .A(n12727), .B(n12726), .S(n15164), .Z(n12728) );
  OAI21_X1 U15037 ( .B1(n12729), .B2(n12757), .A(n12728), .ZN(P3_U3450) );
  MUX2_X1 U15038 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n12730), .S(n15164), .Z(
        P3_U3449) );
  INV_X1 U15039 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12732) );
  MUX2_X1 U15040 ( .A(n12732), .B(n12731), .S(n15164), .Z(n12733) );
  OAI21_X1 U15041 ( .B1(n12734), .B2(n12757), .A(n12733), .ZN(P3_U3448) );
  INV_X1 U15042 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12736) );
  MUX2_X1 U15043 ( .A(n12736), .B(n12735), .S(n15164), .Z(n12737) );
  OAI21_X1 U15044 ( .B1(n12738), .B2(n12757), .A(n12737), .ZN(P3_U3447) );
  MUX2_X1 U15045 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n12739), .S(n15164), .Z(
        P3_U3446) );
  INV_X1 U15046 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12741) );
  MUX2_X1 U15047 ( .A(n12741), .B(n12740), .S(n15164), .Z(n12742) );
  OAI21_X1 U15048 ( .B1(n12743), .B2(n12757), .A(n12742), .ZN(P3_U3444) );
  MUX2_X1 U15049 ( .A(n12744), .B(P3_REG0_REG_17__SCAN_IN), .S(n15162), .Z(
        P3_U3441) );
  INV_X1 U15050 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12746) );
  MUX2_X1 U15051 ( .A(n12746), .B(n12745), .S(n15164), .Z(n12747) );
  OAI21_X1 U15052 ( .B1(n12748), .B2(n12757), .A(n12747), .ZN(P3_U3438) );
  INV_X1 U15053 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12750) );
  MUX2_X1 U15054 ( .A(n12750), .B(n12749), .S(n15164), .Z(n12751) );
  OAI21_X1 U15055 ( .B1(n12757), .B2(n12752), .A(n12751), .ZN(P3_U3435) );
  INV_X1 U15056 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12754) );
  MUX2_X1 U15057 ( .A(n12754), .B(n12753), .S(n15164), .Z(n12755) );
  OAI21_X1 U15058 ( .B1(n12757), .B2(n12756), .A(n12755), .ZN(P3_U3432) );
  MUX2_X1 U15059 ( .A(P3_REG0_REG_0__SCAN_IN), .B(n12758), .S(n15164), .Z(
        P3_U3390) );
  MUX2_X1 U15060 ( .A(P3_D_REG_0__SCAN_IN), .B(n12760), .S(n12759), .Z(
        P3_U3376) );
  INV_X1 U15061 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12761) );
  NAND3_X1 U15062 ( .A1(n12761), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n12762) );
  OAI22_X1 U15063 ( .A1(n7721), .A2(n12762), .B1(n15357), .B2(n12771), .ZN(
        n12763) );
  AOI21_X1 U15064 ( .B1(n12765), .B2(n12764), .A(n12763), .ZN(n12766) );
  INV_X1 U15065 ( .A(n12766), .ZN(P3_U3264) );
  INV_X1 U15066 ( .A(n12767), .ZN(n12769) );
  OAI222_X1 U15067 ( .A1(n12771), .A2(n15364), .B1(n12770), .B2(n12769), .C1(
        P3_U3151), .C2(n12768), .ZN(P3_U3266) );
  XNOR2_X1 U15068 ( .A(n12773), .B(n12774), .ZN(n12780) );
  OAI22_X1 U15069 ( .A1(n12776), .A2(n12988), .B1(n12799), .B2(n12775), .ZN(
        n13070) );
  AOI22_X1 U15070 ( .A1(n12871), .A2(n13070), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12777) );
  OAI21_X1 U15071 ( .B1(n13073), .B2(n12873), .A(n12777), .ZN(n12778) );
  AOI21_X1 U15072 ( .B1(n13271), .B2(n12875), .A(n12778), .ZN(n12779) );
  OAI21_X1 U15073 ( .B1(n12780), .B2(n12877), .A(n12779), .ZN(P2_U3186) );
  NAND2_X1 U15074 ( .A1(n12782), .A2(n12781), .ZN(n12784) );
  XOR2_X1 U15075 ( .A(n12784), .B(n12783), .Z(n12789) );
  AOI22_X1 U15076 ( .A1(n13029), .A2(n12858), .B1(n13020), .B2(n13000), .ZN(
        n13193) );
  INV_X1 U15077 ( .A(n13193), .ZN(n12785) );
  AOI22_X1 U15078 ( .A1(n12785), .A2(n12871), .B1(P2_REG3_REG_19__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12786) );
  OAI21_X1 U15079 ( .B1(n13198), .B2(n12873), .A(n12786), .ZN(n12787) );
  AOI21_X1 U15080 ( .B1(n7148), .B2(n12875), .A(n12787), .ZN(n12788) );
  OAI21_X1 U15081 ( .B1(n12789), .B2(n12877), .A(n12788), .ZN(P2_U3191) );
  XNOR2_X1 U15082 ( .A(n12791), .B(n12790), .ZN(n12796) );
  AOI22_X1 U15083 ( .A1(n13029), .A2(n13020), .B1(n12858), .B2(n13034), .ZN(
        n13165) );
  INV_X1 U15084 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12792) );
  OAI22_X1 U15085 ( .A1(n12859), .A2(n13165), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12792), .ZN(n12794) );
  NOR2_X1 U15086 ( .A1(n13173), .A2(n12865), .ZN(n12793) );
  AOI211_X1 U15087 ( .C1(n12861), .C2(n13170), .A(n12794), .B(n12793), .ZN(
        n12795) );
  OAI21_X1 U15088 ( .B1(n12796), .B2(n12877), .A(n12795), .ZN(P2_U3195) );
  XNOR2_X1 U15089 ( .A(n12798), .B(n12797), .ZN(n12805) );
  OR2_X1 U15090 ( .A1(n12799), .A2(n12988), .ZN(n12801) );
  NAND2_X1 U15091 ( .A1(n12881), .A2(n13020), .ZN(n12800) );
  NAND2_X1 U15092 ( .A1(n12801), .A2(n12800), .ZN(n13097) );
  AOI22_X1 U15093 ( .A1(n12871), .A2(n13097), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12802) );
  OAI21_X1 U15094 ( .B1(n13103), .B2(n12873), .A(n12802), .ZN(n12803) );
  AOI21_X1 U15095 ( .B1(n13282), .B2(n12875), .A(n12803), .ZN(n12804) );
  OAI21_X1 U15096 ( .B1(n12805), .B2(n12877), .A(n12804), .ZN(P2_U3197) );
  OAI21_X1 U15097 ( .B1(n12807), .B2(n12806), .A(n11207), .ZN(n12809) );
  NAND2_X1 U15098 ( .A1(n12809), .A2(n12808), .ZN(n12817) );
  INV_X1 U15099 ( .A(n12810), .ZN(n12815) );
  NOR2_X1 U15100 ( .A1(n12811), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12814) );
  NOR2_X1 U15101 ( .A1(n12873), .A2(n12812), .ZN(n12813) );
  AOI211_X1 U15102 ( .C1(n12871), .C2(n12815), .A(n12814), .B(n12813), .ZN(
        n12816) );
  OAI211_X1 U15103 ( .C1(n7498), .C2(n12865), .A(n12817), .B(n12816), .ZN(
        P2_U3198) );
  OR2_X1 U15104 ( .A1(n12818), .A2(n12877), .ZN(n12836) );
  INV_X1 U15105 ( .A(n12819), .ZN(n12820) );
  AOI21_X1 U15106 ( .B1(n12871), .B2(n12821), .A(n12820), .ZN(n12835) );
  INV_X1 U15107 ( .A(n12822), .ZN(n12823) );
  AOI22_X1 U15108 ( .A1(n12824), .A2(n12875), .B1(n12861), .B2(n12823), .ZN(
        n12834) );
  INV_X1 U15109 ( .A(n12825), .ZN(n12826) );
  OAI22_X1 U15110 ( .A1(n12828), .A2(n12827), .B1(n12826), .B2(n12877), .ZN(
        n12831) );
  INV_X1 U15111 ( .A(n12829), .ZN(n12830) );
  NAND3_X1 U15112 ( .A1(n12832), .A2(n12831), .A3(n12830), .ZN(n12833) );
  NAND4_X1 U15113 ( .A1(n12836), .A2(n12835), .A3(n12834), .A4(n12833), .ZN(
        P2_U3199) );
  AOI21_X1 U15114 ( .B1(n12837), .B2(n12838), .A(n12877), .ZN(n12840) );
  NAND2_X1 U15115 ( .A1(n12840), .A2(n12839), .ZN(n12845) );
  INV_X1 U15116 ( .A(n13119), .ZN(n12843) );
  AOI22_X1 U15117 ( .A1(n13035), .A2(n13020), .B1(n12858), .B2(n13038), .ZN(
        n13111) );
  OAI22_X1 U15118 ( .A1(n12859), .A2(n13111), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12841), .ZN(n12842) );
  AOI21_X1 U15119 ( .B1(n12843), .B2(n12861), .A(n12842), .ZN(n12844) );
  OAI211_X1 U15120 ( .C1(n13037), .C2(n12865), .A(n12845), .B(n12844), .ZN(
        P2_U3201) );
  AOI21_X1 U15121 ( .B1(n12847), .B2(n12846), .A(n6618), .ZN(n12853) );
  INV_X1 U15122 ( .A(n12848), .ZN(n13032) );
  AOI22_X1 U15123 ( .A1(n13032), .A2(n12858), .B1(n13020), .B2(n13003), .ZN(
        n13180) );
  INV_X1 U15124 ( .A(n13180), .ZN(n12849) );
  AOI22_X1 U15125 ( .A1(n12849), .A2(n12871), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12850) );
  OAI21_X1 U15126 ( .B1(n13183), .B2(n12873), .A(n12850), .ZN(n12851) );
  AOI21_X1 U15127 ( .B1(n13309), .B2(n12875), .A(n12851), .ZN(n12852) );
  OAI21_X1 U15128 ( .B1(n12853), .B2(n12877), .A(n12852), .ZN(P2_U3205) );
  AOI21_X1 U15129 ( .B1(n12855), .B2(n12854), .A(n12877), .ZN(n12857) );
  NAND2_X1 U15130 ( .A1(n12857), .A2(n12856), .ZN(n12864) );
  INV_X1 U15131 ( .A(n13214), .ZN(n12862) );
  AOI22_X1 U15132 ( .A1(n13003), .A2(n12858), .B1(n13020), .B2(n12998), .ZN(
        n13209) );
  OAI22_X1 U15133 ( .A1(n12859), .A2(n13209), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12960), .ZN(n12860) );
  AOI21_X1 U15134 ( .B1(n12862), .B2(n12861), .A(n12860), .ZN(n12863) );
  OAI211_X1 U15135 ( .C1(n13213), .C2(n12865), .A(n12864), .B(n12863), .ZN(
        P2_U3210) );
  AOI21_X1 U15136 ( .B1(n12866), .B2(n12868), .A(n12867), .ZN(n12878) );
  OR2_X1 U15137 ( .A1(n13042), .A2(n12988), .ZN(n12870) );
  NAND2_X1 U15138 ( .A1(n13038), .A2(n13020), .ZN(n12869) );
  NAND2_X1 U15139 ( .A1(n12870), .A2(n12869), .ZN(n13083) );
  AOI22_X1 U15140 ( .A1(n12871), .A2(n13083), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12872) );
  OAI21_X1 U15141 ( .B1(n13087), .B2(n12873), .A(n12872), .ZN(n12874) );
  AOI21_X1 U15142 ( .B1(n13276), .B2(n12875), .A(n12874), .ZN(n12876) );
  OAI21_X1 U15143 ( .B1(n12878), .B2(n12877), .A(n12876), .ZN(P2_U3212) );
  MUX2_X1 U15144 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n12989), .S(n6467), .Z(
        P2_U3562) );
  MUX2_X1 U15145 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13019), .S(n6467), .Z(
        P2_U3561) );
  MUX2_X1 U15146 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n12879), .S(n6467), .Z(
        P2_U3560) );
  MUX2_X1 U15147 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13043), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15148 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n12880), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15149 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13039), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15150 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13038), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15151 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n12881), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15152 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13035), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15153 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13034), .S(n6467), .Z(
        P2_U3553) );
  MUX2_X1 U15154 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13032), .S(n6467), .Z(
        P2_U3552) );
  MUX2_X1 U15155 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13029), .S(n6467), .Z(
        P2_U3551) );
  MUX2_X1 U15156 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13003), .S(n6467), .Z(
        P2_U3550) );
  MUX2_X1 U15157 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13000), .S(n6467), .Z(
        P2_U3549) );
  MUX2_X1 U15158 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n12998), .S(n6467), .Z(
        P2_U3548) );
  MUX2_X1 U15159 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n12882), .S(n6467), .Z(
        P2_U3547) );
  MUX2_X1 U15160 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n12883), .S(n6467), .Z(
        P2_U3546) );
  MUX2_X1 U15161 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n12884), .S(n6467), .Z(
        P2_U3545) );
  MUX2_X1 U15162 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n12885), .S(n6467), .Z(
        P2_U3544) );
  MUX2_X1 U15163 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n12886), .S(n6467), .Z(
        P2_U3543) );
  MUX2_X1 U15164 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n12887), .S(n6467), .Z(
        P2_U3542) );
  MUX2_X1 U15165 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n12888), .S(n6467), .Z(
        P2_U3541) );
  MUX2_X1 U15166 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n12889), .S(n6467), .Z(
        P2_U3540) );
  MUX2_X1 U15167 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n12890), .S(n6467), .Z(
        P2_U3539) );
  MUX2_X1 U15168 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n12891), .S(n6467), .Z(
        P2_U3538) );
  MUX2_X1 U15169 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n12892), .S(n6467), .Z(
        P2_U3537) );
  MUX2_X1 U15170 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n12893), .S(n6467), .Z(
        P2_U3536) );
  MUX2_X1 U15171 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n12894), .S(n6467), .Z(
        P2_U3535) );
  MUX2_X1 U15172 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n12895), .S(n6467), .Z(
        P2_U3534) );
  MUX2_X1 U15173 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n12896), .S(n6467), .Z(
        P2_U3533) );
  MUX2_X1 U15174 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n12897), .S(n6467), .Z(
        P2_U3532) );
  MUX2_X1 U15175 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n12898), .S(n6467), .Z(
        P2_U3531) );
  AND3_X1 U15176 ( .A1(n12901), .A2(n12900), .A3(n12899), .ZN(n12902) );
  NOR3_X1 U15177 ( .A1(n14733), .A2(n12903), .A3(n12902), .ZN(n12904) );
  AOI21_X1 U15178 ( .B1(n14790), .B2(n12905), .A(n12904), .ZN(n12916) );
  MUX2_X1 U15179 ( .A(n12906), .B(P2_REG1_REG_3__SCAN_IN), .S(n12905), .Z(
        n12909) );
  INV_X1 U15180 ( .A(n12907), .ZN(n12908) );
  NAND2_X1 U15181 ( .A1(n12909), .A2(n12908), .ZN(n12911) );
  OAI211_X1 U15182 ( .C1(n12912), .C2(n12911), .A(n14785), .B(n12910), .ZN(
        n12914) );
  NAND2_X1 U15183 ( .A1(n14784), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n12913) );
  NAND4_X1 U15184 ( .A1(n12916), .A2(n12915), .A3(n12914), .A4(n12913), .ZN(
        P2_U3217) );
  OAI21_X1 U15185 ( .B1(n12919), .B2(n12918), .A(n12917), .ZN(n12920) );
  NAND2_X1 U15186 ( .A1(n12920), .A2(n14791), .ZN(n12930) );
  AND2_X1 U15187 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n12921) );
  AOI21_X1 U15188 ( .B1(n14784), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n12921), .ZN(
        n12929) );
  OAI21_X1 U15189 ( .B1(n12924), .B2(n12923), .A(n12922), .ZN(n12925) );
  NAND2_X1 U15190 ( .A1(n12925), .A2(n14785), .ZN(n12928) );
  NAND2_X1 U15191 ( .A1(n14790), .A2(n12926), .ZN(n12927) );
  NAND4_X1 U15192 ( .A1(n12930), .A2(n12929), .A3(n12928), .A4(n12927), .ZN(
        P2_U3223) );
  NAND2_X1 U15193 ( .A1(n14789), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U15194 ( .A1(n14746), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12936) );
  INV_X1 U15195 ( .A(n12936), .ZN(n12934) );
  AOI21_X1 U15196 ( .B1(n10527), .B2(n12935), .A(n12934), .ZN(n14739) );
  NAND2_X1 U15197 ( .A1(n14740), .A2(n14739), .ZN(n14738) );
  NAND2_X1 U15198 ( .A1(n12949), .A2(n12937), .ZN(n12938) );
  NAND2_X1 U15199 ( .A1(n14764), .A2(n12939), .ZN(n12941) );
  XNOR2_X1 U15200 ( .A(n12940), .B(n12939), .ZN(n14766) );
  NOR2_X1 U15201 ( .A1(n12953), .A2(n12942), .ZN(n12943) );
  AOI21_X1 U15202 ( .B1(n12942), .B2(n12953), .A(n12943), .ZN(n14775) );
  INV_X1 U15203 ( .A(n12945), .ZN(n12944) );
  AOI21_X1 U15204 ( .B1(n13234), .B2(n12956), .A(n12944), .ZN(n14793) );
  NAND2_X1 U15205 ( .A1(n14794), .A2(n14793), .ZN(n14792) );
  AOI21_X1 U15206 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n12946), .A(n12969), 
        .ZN(n12966) );
  OAI21_X1 U15207 ( .B1(n12948), .B2(P2_REG1_REG_12__SCAN_IN), .A(n12947), 
        .ZN(n14743) );
  MUX2_X1 U15208 ( .A(n10310), .B(P2_REG1_REG_13__SCAN_IN), .S(n14746), .Z(
        n14744) );
  NOR2_X1 U15209 ( .A1(n14743), .A2(n14744), .ZN(n14741) );
  AOI21_X1 U15210 ( .B1(n14746), .B2(P2_REG1_REG_13__SCAN_IN), .A(n14741), 
        .ZN(n14757) );
  XNOR2_X1 U15211 ( .A(n12949), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14758) );
  INV_X1 U15212 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12950) );
  OAI22_X1 U15213 ( .A1(n14757), .A2(n14758), .B1(n14752), .B2(n12950), .ZN(
        n12951) );
  NAND2_X1 U15214 ( .A1(n14764), .A2(n12951), .ZN(n12952) );
  XOR2_X1 U15215 ( .A(n14764), .B(n12951), .Z(n14768) );
  NAND2_X1 U15216 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14768), .ZN(n14767) );
  NAND2_X1 U15217 ( .A1(n12952), .A2(n14767), .ZN(n14778) );
  INV_X1 U15218 ( .A(n14778), .ZN(n12955) );
  XNOR2_X1 U15219 ( .A(n14773), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14777) );
  INV_X1 U15220 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12954) );
  OAI22_X1 U15221 ( .A1(n12955), .A2(n14777), .B1(n12954), .B2(n12953), .ZN(
        n14788) );
  XNOR2_X1 U15222 ( .A(n12956), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14787) );
  NAND2_X1 U15223 ( .A1(n14788), .A2(n14787), .ZN(n14786) );
  OAI21_X1 U15224 ( .B1(n12957), .B2(n12956), .A(n14786), .ZN(n12971) );
  XNOR2_X1 U15225 ( .A(n12958), .B(n12971), .ZN(n12959) );
  NAND2_X1 U15226 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n12959), .ZN(n12973) );
  OAI211_X1 U15227 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n12959), .A(n14785), 
        .B(n12973), .ZN(n12963) );
  NOR2_X1 U15228 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12960), .ZN(n12961) );
  AOI21_X1 U15229 ( .B1(n14784), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n12961), 
        .ZN(n12962) );
  NAND2_X1 U15230 ( .A1(n12963), .A2(n12962), .ZN(n12964) );
  AOI21_X1 U15231 ( .B1(n12972), .B2(n14790), .A(n12964), .ZN(n12965) );
  OAI21_X1 U15232 ( .B1(n12966), .B2(n14733), .A(n12965), .ZN(P2_U3232) );
  INV_X1 U15233 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n12982) );
  NOR2_X1 U15234 ( .A1(n12972), .A2(n12967), .ZN(n12968) );
  INV_X1 U15235 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n12976) );
  NAND2_X1 U15236 ( .A1(n12972), .A2(n12971), .ZN(n12974) );
  NAND2_X1 U15237 ( .A1(n12974), .A2(n12973), .ZN(n12975) );
  XNOR2_X1 U15238 ( .A(n12976), .B(n12975), .ZN(n12979) );
  NOR2_X1 U15239 ( .A1(n12979), .A2(n14742), .ZN(n12977) );
  AOI211_X1 U15240 ( .C1(n12978), .C2(n14791), .A(n14790), .B(n12977), .ZN(
        n12980) );
  NAND2_X1 U15241 ( .A1(n14784), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n12981) );
  NOR2_X1 U15242 ( .A1(n13195), .A2(n13309), .ZN(n13182) );
  NAND2_X1 U15243 ( .A1(n13182), .A2(n13173), .ZN(n13167) );
  INV_X1 U15244 ( .A(n13267), .ZN(n13064) );
  NAND2_X1 U15245 ( .A1(n12984), .A2(n13332), .ZN(n13257) );
  NOR2_X1 U15246 ( .A1(n13228), .A2(n12985), .ZN(n12990) );
  INV_X1 U15247 ( .A(P2_B_REG_SCAN_IN), .ZN(n12986) );
  NOR2_X1 U15248 ( .A1(n13365), .A2(n12986), .ZN(n12987) );
  NOR2_X1 U15249 ( .A1(n12988), .A2(n12987), .ZN(n13018) );
  NAND2_X1 U15250 ( .A1(n12989), .A2(n13018), .ZN(n13258) );
  NOR2_X1 U15251 ( .A1(n6466), .A2(n13258), .ZN(n12994) );
  AOI211_X1 U15252 ( .C1(n13256), .C2(n13248), .A(n12990), .B(n12994), .ZN(
        n12991) );
  OAI21_X1 U15253 ( .B1(n13257), .B2(n13159), .A(n12991), .ZN(P2_U3234) );
  OAI211_X1 U15254 ( .C1(n13047), .C2(n13260), .A(n13332), .B(n12992), .ZN(
        n13259) );
  NOR2_X1 U15255 ( .A1(n13228), .A2(n12993), .ZN(n12995) );
  AOI211_X1 U15256 ( .C1(n12996), .C2(n13248), .A(n12995), .B(n12994), .ZN(
        n12997) );
  OAI21_X1 U15257 ( .B1(n13259), .B2(n13159), .A(n12997), .ZN(P2_U3235) );
  INV_X1 U15258 ( .A(n12998), .ZN(n13025) );
  INV_X1 U15259 ( .A(n13000), .ZN(n13026) );
  NAND2_X1 U15260 ( .A1(n13318), .A2(n13026), .ZN(n13001) );
  INV_X1 U15261 ( .A(n13178), .ZN(n13176) );
  INV_X1 U15262 ( .A(n13309), .ZN(n13187) );
  INV_X1 U15263 ( .A(n13163), .ZN(n13033) );
  NOR2_X1 U15264 ( .A1(n13173), .A2(n13032), .ZN(n13005) );
  INV_X1 U15265 ( .A(n13145), .ZN(n13150) );
  NAND2_X1 U15266 ( .A1(n13292), .A2(n13006), .ZN(n13007) );
  NAND2_X1 U15267 ( .A1(n13096), .A2(n13100), .ZN(n13011) );
  NAND2_X1 U15268 ( .A1(n13282), .A2(n13009), .ZN(n13010) );
  NAND2_X1 U15269 ( .A1(n13082), .A2(n13012), .ZN(n13014) );
  NAND2_X1 U15270 ( .A1(n13271), .A2(n13042), .ZN(n13015) );
  AOI22_X1 U15271 ( .A1(n13020), .A2(n13043), .B1(n13019), .B2(n13018), .ZN(
        n13021) );
  NAND2_X1 U15272 ( .A1(n13309), .A2(n13029), .ZN(n13031) );
  OAI21_X1 U15273 ( .B1(n13035), .B2(n13292), .A(n13128), .ZN(n13114) );
  NOR2_X1 U15274 ( .A1(n13276), .A2(n13039), .ZN(n13041) );
  NAND2_X1 U15275 ( .A1(n13276), .A2(n13039), .ZN(n13040) );
  INV_X1 U15276 ( .A(n13044), .ZN(n13045) );
  INV_X1 U15277 ( .A(n13263), .ZN(n13052) );
  AOI211_X1 U15278 ( .C1(n13263), .C2(n13061), .A(n13243), .B(n13047), .ZN(
        n13262) );
  NAND2_X1 U15279 ( .A1(n13262), .A2(n13245), .ZN(n13051) );
  INV_X1 U15280 ( .A(n13048), .ZN(n13049) );
  AOI22_X1 U15281 ( .A1(n6466), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n13049), 
        .B2(n13247), .ZN(n13050) );
  OAI211_X1 U15282 ( .C1(n13052), .C2(n13231), .A(n13051), .B(n13050), .ZN(
        n13053) );
  AOI21_X1 U15283 ( .B1(n13261), .B2(n13246), .A(n13053), .ZN(n13054) );
  OAI21_X1 U15284 ( .B1(n13265), .B2(n6466), .A(n13054), .ZN(P2_U3236) );
  OAI21_X1 U15285 ( .B1(n13059), .B2(n13232), .A(n13268), .ZN(n13060) );
  NAND2_X1 U15286 ( .A1(n13060), .A2(n13228), .ZN(n13067) );
  AOI211_X1 U15287 ( .C1(n13267), .C2(n6796), .A(n13243), .B(n13062), .ZN(
        n13266) );
  INV_X1 U15288 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13063) );
  OAI22_X1 U15289 ( .A1(n13064), .A2(n13231), .B1(n13228), .B2(n13063), .ZN(
        n13065) );
  AOI21_X1 U15290 ( .B1(n13266), .B2(n13245), .A(n13065), .ZN(n13066) );
  OAI211_X1 U15291 ( .C1(n13239), .C2(n13269), .A(n13067), .B(n13066), .ZN(
        P2_U3237) );
  XNOR2_X1 U15292 ( .A(n13069), .B(n13068), .ZN(n13071) );
  AOI211_X1 U15293 ( .C1(n13271), .C2(n13086), .A(n13243), .B(n13072), .ZN(
        n13270) );
  INV_X1 U15294 ( .A(n13073), .ZN(n13074) );
  AOI22_X1 U15295 ( .A1(n6466), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n13074), 
        .B2(n13247), .ZN(n13075) );
  OAI21_X1 U15296 ( .B1(n13076), .B2(n13231), .A(n13075), .ZN(n13080) );
  XNOR2_X1 U15297 ( .A(n13078), .B(n13077), .ZN(n13274) );
  NOR2_X1 U15298 ( .A1(n13274), .A2(n13239), .ZN(n13079) );
  AOI211_X1 U15299 ( .C1(n13245), .C2(n13270), .A(n13080), .B(n13079), .ZN(
        n13081) );
  OAI21_X1 U15300 ( .B1(n13273), .B2(n6466), .A(n13081), .ZN(P2_U3238) );
  XNOR2_X1 U15301 ( .A(n13082), .B(n13091), .ZN(n13084) );
  AOI21_X1 U15302 ( .B1(n13084), .B2(n13251), .A(n13083), .ZN(n13278) );
  OR2_X1 U15303 ( .A1(n13090), .A2(n13102), .ZN(n13085) );
  AND3_X1 U15304 ( .A1(n13086), .A2(n13085), .A3(n13332), .ZN(n13275) );
  INV_X1 U15305 ( .A(n13087), .ZN(n13088) );
  AOI22_X1 U15306 ( .A1(n6466), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13088), 
        .B2(n13247), .ZN(n13089) );
  OAI21_X1 U15307 ( .B1(n13090), .B2(n13231), .A(n13089), .ZN(n13094) );
  XNOR2_X1 U15308 ( .A(n13092), .B(n13091), .ZN(n13279) );
  NOR2_X1 U15309 ( .A1(n13279), .A2(n13239), .ZN(n13093) );
  AOI211_X1 U15310 ( .C1(n13275), .C2(n13245), .A(n13094), .B(n13093), .ZN(
        n13095) );
  OAI21_X1 U15311 ( .B1(n6466), .B2(n13278), .A(n13095), .ZN(P2_U3239) );
  XNOR2_X1 U15312 ( .A(n13096), .B(n13100), .ZN(n13098) );
  AOI21_X1 U15313 ( .B1(n13098), .B2(n13251), .A(n13097), .ZN(n13284) );
  AOI21_X1 U15314 ( .B1(n13100), .B2(n13099), .A(n6560), .ZN(n13285) );
  INV_X1 U15315 ( .A(n13285), .ZN(n13108) );
  AND2_X1 U15316 ( .A1(n13282), .A2(n13122), .ZN(n13101) );
  OR3_X1 U15317 ( .A1(n13102), .A2(n13101), .A3(n13243), .ZN(n13280) );
  OAI22_X1 U15318 ( .A1(n13155), .A2(n13104), .B1(n13103), .B2(n13232), .ZN(
        n13105) );
  AOI21_X1 U15319 ( .B1(n13282), .B2(n13248), .A(n13105), .ZN(n13106) );
  OAI21_X1 U15320 ( .B1(n13280), .B2(n13159), .A(n13106), .ZN(n13107) );
  AOI21_X1 U15321 ( .B1(n13108), .B2(n13246), .A(n13107), .ZN(n13109) );
  OAI21_X1 U15322 ( .B1(n6466), .B2(n13284), .A(n13109), .ZN(P2_U3240) );
  XNOR2_X1 U15323 ( .A(n13110), .B(n13115), .ZN(n13113) );
  INV_X1 U15324 ( .A(n13111), .ZN(n13112) );
  AOI21_X1 U15325 ( .B1(n13113), .B2(n13251), .A(n13112), .ZN(n13289) );
  INV_X1 U15326 ( .A(n13114), .ZN(n13118) );
  INV_X1 U15327 ( .A(n13115), .ZN(n13117) );
  OAI21_X1 U15328 ( .B1(n13118), .B2(n13117), .A(n13116), .ZN(n13290) );
  OAI22_X1 U15329 ( .A1(n13155), .A2(n13120), .B1(n13119), .B2(n13232), .ZN(
        n13121) );
  AOI21_X1 U15330 ( .B1(n13287), .B2(n13248), .A(n13121), .ZN(n13125) );
  AOI21_X1 U15331 ( .B1(n13287), .B2(n13138), .A(n13243), .ZN(n13123) );
  AND2_X1 U15332 ( .A1(n13123), .A2(n13122), .ZN(n13286) );
  NAND2_X1 U15333 ( .A1(n13286), .A2(n13245), .ZN(n13124) );
  OAI211_X1 U15334 ( .C1(n13290), .C2(n13239), .A(n13125), .B(n13124), .ZN(
        n13126) );
  INV_X1 U15335 ( .A(n13126), .ZN(n13127) );
  OAI21_X1 U15336 ( .B1(n6466), .B2(n13289), .A(n13127), .ZN(P2_U3241) );
  OAI21_X1 U15337 ( .B1(n13130), .B2(n13129), .A(n13128), .ZN(n13131) );
  INV_X1 U15338 ( .A(n13131), .ZN(n13295) );
  OAI21_X1 U15339 ( .B1(n13134), .B2(n13133), .A(n13132), .ZN(n13136) );
  AOI21_X1 U15340 ( .B1(n13136), .B2(n13251), .A(n13135), .ZN(n13294) );
  OAI21_X1 U15341 ( .B1(n13137), .B2(n13232), .A(n13294), .ZN(n13143) );
  INV_X1 U15342 ( .A(n13152), .ZN(n13139) );
  AOI211_X1 U15343 ( .C1(n13292), .C2(n13139), .A(n13243), .B(n6799), .ZN(
        n13291) );
  INV_X1 U15344 ( .A(n13291), .ZN(n13141) );
  AOI22_X1 U15345 ( .A1(n13292), .A2(n13248), .B1(n6466), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13140) );
  OAI21_X1 U15346 ( .B1(n13141), .B2(n13159), .A(n13140), .ZN(n13142) );
  AOI21_X1 U15347 ( .B1(n13143), .B2(n13228), .A(n13142), .ZN(n13144) );
  OAI21_X1 U15348 ( .B1(n13295), .B2(n13239), .A(n13144), .ZN(P2_U3242) );
  XNOR2_X1 U15349 ( .A(n13146), .B(n13145), .ZN(n13148) );
  AOI21_X1 U15350 ( .B1(n13148), .B2(n13251), .A(n13147), .ZN(n13297) );
  AOI21_X1 U15351 ( .B1(n13150), .B2(n13149), .A(n6561), .ZN(n13300) );
  AND2_X1 U15352 ( .A1(n13167), .A2(n13157), .ZN(n13151) );
  OR3_X1 U15353 ( .A1(n13152), .A2(n13151), .A3(n13243), .ZN(n13296) );
  INV_X1 U15354 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13154) );
  OAI22_X1 U15355 ( .A1(n13155), .A2(n13154), .B1(n13153), .B2(n13232), .ZN(
        n13156) );
  AOI21_X1 U15356 ( .B1(n13157), .B2(n13248), .A(n13156), .ZN(n13158) );
  OAI21_X1 U15357 ( .B1(n13296), .B2(n13159), .A(n13158), .ZN(n13160) );
  AOI21_X1 U15358 ( .B1(n13300), .B2(n13246), .A(n13160), .ZN(n13161) );
  OAI21_X1 U15359 ( .B1(n13297), .B2(n6466), .A(n13161), .ZN(P2_U3243) );
  XNOR2_X1 U15360 ( .A(n13162), .B(n13163), .ZN(n13306) );
  XNOR2_X1 U15361 ( .A(n13164), .B(n13163), .ZN(n13166) );
  OAI21_X1 U15362 ( .B1(n13166), .B2(n13226), .A(n13165), .ZN(n13302) );
  INV_X1 U15363 ( .A(n13182), .ZN(n13169) );
  INV_X1 U15364 ( .A(n13167), .ZN(n13168) );
  AOI211_X1 U15365 ( .C1(n13304), .C2(n13169), .A(n13243), .B(n13168), .ZN(
        n13303) );
  NAND2_X1 U15366 ( .A1(n13303), .A2(n13245), .ZN(n13172) );
  AOI22_X1 U15367 ( .A1(n6466), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13170), 
        .B2(n13247), .ZN(n13171) );
  OAI211_X1 U15368 ( .C1(n13173), .C2(n13231), .A(n13172), .B(n13171), .ZN(
        n13174) );
  AOI21_X1 U15369 ( .B1(n13302), .B2(n13228), .A(n13174), .ZN(n13175) );
  OAI21_X1 U15370 ( .B1(n13239), .B2(n13306), .A(n13175), .ZN(P2_U3244) );
  XNOR2_X1 U15371 ( .A(n13177), .B(n13176), .ZN(n13311) );
  XNOR2_X1 U15372 ( .A(n13179), .B(n13178), .ZN(n13181) );
  OAI21_X1 U15373 ( .B1(n13181), .B2(n13226), .A(n13180), .ZN(n13307) );
  AOI211_X1 U15374 ( .C1(n13309), .C2(n13195), .A(n13243), .B(n13182), .ZN(
        n13308) );
  NAND2_X1 U15375 ( .A1(n13308), .A2(n13245), .ZN(n13186) );
  INV_X1 U15376 ( .A(n13183), .ZN(n13184) );
  AOI22_X1 U15377 ( .A1(n6466), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13184), 
        .B2(n13247), .ZN(n13185) );
  OAI211_X1 U15378 ( .C1(n13187), .C2(n13231), .A(n13186), .B(n13185), .ZN(
        n13188) );
  AOI21_X1 U15379 ( .B1(n13307), .B2(n13228), .A(n13188), .ZN(n13189) );
  OAI21_X1 U15380 ( .B1(n13239), .B2(n13311), .A(n13189), .ZN(P2_U3245) );
  XOR2_X1 U15381 ( .A(n13192), .B(n13190), .Z(n13315) );
  XOR2_X1 U15382 ( .A(n13192), .B(n13191), .Z(n13194) );
  OAI21_X1 U15383 ( .B1(n13194), .B2(n13226), .A(n13193), .ZN(n13312) );
  INV_X1 U15384 ( .A(n13211), .ZN(n13197) );
  INV_X1 U15385 ( .A(n13195), .ZN(n13196) );
  AOI211_X1 U15386 ( .C1(n7148), .C2(n13197), .A(n13243), .B(n13196), .ZN(
        n13313) );
  NAND2_X1 U15387 ( .A1(n13313), .A2(n13245), .ZN(n13201) );
  INV_X1 U15388 ( .A(n13198), .ZN(n13199) );
  AOI22_X1 U15389 ( .A1(n6466), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13199), 
        .B2(n13247), .ZN(n13200) );
  OAI211_X1 U15390 ( .C1(n13202), .C2(n13231), .A(n13201), .B(n13200), .ZN(
        n13203) );
  AOI21_X1 U15391 ( .B1(n13312), .B2(n13228), .A(n13203), .ZN(n13204) );
  OAI21_X1 U15392 ( .B1(n13239), .B2(n13315), .A(n13204), .ZN(P2_U3246) );
  AOI21_X1 U15393 ( .B1(n13207), .B2(n13206), .A(n13205), .ZN(n13320) );
  XNOR2_X1 U15394 ( .A(n13208), .B(n13207), .ZN(n13210) );
  OAI21_X1 U15395 ( .B1(n13210), .B2(n13226), .A(n13209), .ZN(n13316) );
  NAND2_X1 U15396 ( .A1(n13316), .A2(n13228), .ZN(n13219) );
  INV_X1 U15397 ( .A(n13229), .ZN(n13212) );
  AOI211_X1 U15398 ( .C1(n13318), .C2(n13212), .A(n13243), .B(n13211), .ZN(
        n13317) );
  NOR2_X1 U15399 ( .A1(n13213), .A2(n13231), .ZN(n13217) );
  OAI22_X1 U15400 ( .A1(n13155), .A2(n13215), .B1(n13214), .B2(n13232), .ZN(
        n13216) );
  AOI211_X1 U15401 ( .C1(n13317), .C2(n13245), .A(n13217), .B(n13216), .ZN(
        n13218) );
  OAI211_X1 U15402 ( .C1(n13320), .C2(n13239), .A(n13219), .B(n13218), .ZN(
        P2_U3247) );
  OAI21_X1 U15403 ( .B1(n13221), .B2(n13224), .A(n13220), .ZN(n13325) );
  AOI21_X1 U15404 ( .B1(n13224), .B2(n13223), .A(n13222), .ZN(n13227) );
  OAI21_X1 U15405 ( .B1(n13227), .B2(n13226), .A(n13225), .ZN(n13321) );
  NAND2_X1 U15406 ( .A1(n13321), .A2(n13228), .ZN(n13238) );
  AOI211_X1 U15407 ( .C1(n13323), .C2(n13230), .A(n13243), .B(n13229), .ZN(
        n13322) );
  NOR2_X1 U15408 ( .A1(n7150), .A2(n13231), .ZN(n13236) );
  OAI22_X1 U15409 ( .A1(n13155), .A2(n13234), .B1(n13233), .B2(n13232), .ZN(
        n13235) );
  AOI211_X1 U15410 ( .C1(n13322), .C2(n13245), .A(n13236), .B(n13235), .ZN(
        n13237) );
  OAI211_X1 U15411 ( .C1(n13325), .C2(n13239), .A(n13238), .B(n13237), .ZN(
        P2_U3248) );
  OAI21_X1 U15412 ( .B1(n6940), .B2(n13241), .A(n13240), .ZN(n14819) );
  AOI211_X1 U15413 ( .C1(n13244), .C2(n14814), .A(n13243), .B(n13242), .ZN(
        n14813) );
  AOI22_X1 U15414 ( .A1(n13246), .A2(n14819), .B1(n13245), .B2(n14813), .ZN(
        n13255) );
  AOI22_X1 U15415 ( .A1(n13248), .A2(n14814), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13247), .ZN(n13254) );
  XNOR2_X1 U15416 ( .A(n13249), .B(n6953), .ZN(n13252) );
  AOI21_X1 U15417 ( .B1(n13252), .B2(n13251), .A(n13250), .ZN(n14812) );
  MUX2_X1 U15418 ( .A(n8629), .B(n14812), .S(n13228), .Z(n13253) );
  NAND3_X1 U15419 ( .A1(n13255), .A2(n13254), .A3(n13253), .ZN(P2_U3264) );
  OAI211_X1 U15420 ( .C1(n7145), .C2(n14867), .A(n13257), .B(n13258), .ZN(
        n13338) );
  MUX2_X1 U15421 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13338), .S(n14908), .Z(
        P2_U3530) );
  OAI211_X1 U15422 ( .C1(n13260), .C2(n14867), .A(n13259), .B(n13258), .ZN(
        n13339) );
  MUX2_X1 U15423 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13339), .S(n14908), .Z(
        P2_U3529) );
  AOI21_X1 U15424 ( .B1(n14879), .B2(n13263), .A(n13262), .ZN(n13264) );
  MUX2_X1 U15425 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13340), .S(n14908), .Z(
        P2_U3528) );
  MUX2_X1 U15426 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13341), .S(n14908), .Z(
        P2_U3527) );
  AOI21_X1 U15427 ( .B1(n14879), .B2(n13271), .A(n13270), .ZN(n13272) );
  OAI211_X1 U15428 ( .C1(n13274), .C2(n13337), .A(n13273), .B(n13272), .ZN(
        n13342) );
  MUX2_X1 U15429 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13342), .S(n14908), .Z(
        P2_U3526) );
  AOI21_X1 U15430 ( .B1(n14879), .B2(n13276), .A(n13275), .ZN(n13277) );
  OAI211_X1 U15431 ( .C1(n13279), .C2(n13337), .A(n13278), .B(n13277), .ZN(
        n13343) );
  MUX2_X1 U15432 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13343), .S(n14908), .Z(
        P2_U3525) );
  INV_X1 U15433 ( .A(n13280), .ZN(n13281) );
  AOI21_X1 U15434 ( .B1(n14879), .B2(n13282), .A(n13281), .ZN(n13283) );
  OAI211_X1 U15435 ( .C1(n13285), .C2(n13337), .A(n13284), .B(n13283), .ZN(
        n13344) );
  MUX2_X1 U15436 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13344), .S(n14908), .Z(
        P2_U3524) );
  AOI21_X1 U15437 ( .B1(n14879), .B2(n13287), .A(n13286), .ZN(n13288) );
  OAI211_X1 U15438 ( .C1(n13290), .C2(n13337), .A(n13289), .B(n13288), .ZN(
        n13345) );
  MUX2_X1 U15439 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13345), .S(n14908), .Z(
        P2_U3523) );
  AOI21_X1 U15440 ( .B1(n14879), .B2(n13292), .A(n13291), .ZN(n13293) );
  OAI211_X1 U15441 ( .C1(n13337), .C2(n13295), .A(n13294), .B(n13293), .ZN(
        n13346) );
  MUX2_X1 U15442 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13346), .S(n14908), .Z(
        P2_U3522) );
  OAI211_X1 U15443 ( .C1(n13298), .C2(n14867), .A(n13297), .B(n13296), .ZN(
        n13299) );
  AOI21_X1 U15444 ( .B1(n13300), .B2(n14850), .A(n13299), .ZN(n13301) );
  INV_X1 U15445 ( .A(n13301), .ZN(n13347) );
  MUX2_X1 U15446 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13347), .S(n14908), .Z(
        P2_U3521) );
  AOI211_X1 U15447 ( .C1(n14879), .C2(n13304), .A(n13303), .B(n13302), .ZN(
        n13305) );
  OAI21_X1 U15448 ( .B1(n13337), .B2(n13306), .A(n13305), .ZN(n13348) );
  MUX2_X1 U15449 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13348), .S(n14908), .Z(
        P2_U3520) );
  AOI211_X1 U15450 ( .C1(n14879), .C2(n13309), .A(n13308), .B(n13307), .ZN(
        n13310) );
  OAI21_X1 U15451 ( .B1(n13337), .B2(n13311), .A(n13310), .ZN(n13349) );
  MUX2_X1 U15452 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13349), .S(n14908), .Z(
        P2_U3519) );
  AOI211_X1 U15453 ( .C1(n14879), .C2(n7148), .A(n13313), .B(n13312), .ZN(
        n13314) );
  OAI21_X1 U15454 ( .B1(n13337), .B2(n13315), .A(n13314), .ZN(n13350) );
  MUX2_X1 U15455 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13350), .S(n14908), .Z(
        P2_U3518) );
  AOI211_X1 U15456 ( .C1(n14879), .C2(n13318), .A(n13317), .B(n13316), .ZN(
        n13319) );
  OAI21_X1 U15457 ( .B1(n13337), .B2(n13320), .A(n13319), .ZN(n13351) );
  MUX2_X1 U15458 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13351), .S(n14908), .Z(
        P2_U3517) );
  AOI211_X1 U15459 ( .C1(n14879), .C2(n13323), .A(n13322), .B(n13321), .ZN(
        n13324) );
  OAI21_X1 U15460 ( .B1(n13337), .B2(n13325), .A(n13324), .ZN(n13352) );
  MUX2_X1 U15461 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13352), .S(n14908), .Z(
        P2_U3516) );
  AOI211_X1 U15462 ( .C1(n14879), .C2(n13328), .A(n13327), .B(n13326), .ZN(
        n13329) );
  OAI21_X1 U15463 ( .B1(n13337), .B2(n13330), .A(n13329), .ZN(n13353) );
  MUX2_X1 U15464 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13353), .S(n14908), .Z(
        P2_U3515) );
  AOI22_X1 U15465 ( .A1(n13333), .A2(n13332), .B1(n14879), .B2(n13331), .ZN(
        n13334) );
  OAI211_X1 U15466 ( .C1(n13337), .C2(n13336), .A(n13335), .B(n13334), .ZN(
        n13354) );
  MUX2_X1 U15467 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13354), .S(n14908), .Z(
        P2_U3514) );
  MUX2_X1 U15468 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13338), .S(n14887), .Z(
        P2_U3498) );
  MUX2_X1 U15469 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13339), .S(n14887), .Z(
        P2_U3497) );
  MUX2_X1 U15470 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13340), .S(n14887), .Z(
        P2_U3496) );
  MUX2_X1 U15471 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13342), .S(n14887), .Z(
        P2_U3494) );
  MUX2_X1 U15472 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13343), .S(n14887), .Z(
        P2_U3493) );
  MUX2_X1 U15473 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13344), .S(n14887), .Z(
        P2_U3492) );
  MUX2_X1 U15474 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13345), .S(n14887), .Z(
        P2_U3491) );
  MUX2_X1 U15475 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13346), .S(n14887), .Z(
        P2_U3490) );
  MUX2_X1 U15476 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13347), .S(n14887), .Z(
        P2_U3489) );
  MUX2_X1 U15477 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13348), .S(n14887), .Z(
        P2_U3488) );
  MUX2_X1 U15478 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13349), .S(n14887), .Z(
        P2_U3487) );
  MUX2_X1 U15479 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13350), .S(n14887), .Z(
        P2_U3486) );
  MUX2_X1 U15480 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13351), .S(n14887), .Z(
        P2_U3484) );
  MUX2_X1 U15481 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13352), .S(n14887), .Z(
        P2_U3481) );
  MUX2_X1 U15482 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13353), .S(n14887), .Z(
        P2_U3478) );
  MUX2_X1 U15483 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13354), .S(n14887), .Z(
        P2_U3475) );
  INV_X1 U15484 ( .A(n14216), .ZN(n13359) );
  NOR4_X1 U15485 ( .A1(n13355), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7012), .A4(
        P2_U3088), .ZN(n13357) );
  AOI21_X1 U15486 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13361), .A(n13357), 
        .ZN(n13358) );
  OAI21_X1 U15487 ( .B1(n13359), .B2(n13366), .A(n13358), .ZN(P2_U3296) );
  AOI21_X1 U15488 ( .B1(n13361), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13360), 
        .ZN(n13362) );
  OAI21_X1 U15489 ( .B1(n13363), .B2(n13366), .A(n13362), .ZN(P2_U3299) );
  INV_X1 U15490 ( .A(n13364), .ZN(n14220) );
  OAI222_X1 U15491 ( .A1(n13368), .A2(n13367), .B1(n13366), .B2(n14220), .C1(
        P2_U3088), .C2(n13365), .ZN(P2_U3300) );
  MUX2_X1 U15492 ( .A(n13369), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15493 ( .A1(n13371), .A2(n14431), .ZN(n13376) );
  NOR2_X1 U15494 ( .A1(n14436), .A2(n13851), .ZN(n13374) );
  OAI22_X1 U15495 ( .A1(n13372), .A2(n14426), .B1(n14427), .B2(n13421), .ZN(
        n13373) );
  AOI211_X1 U15496 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n13374), 
        .B(n13373), .ZN(n13375) );
  OAI211_X1 U15497 ( .C1(n14066), .C2(n14423), .A(n13376), .B(n13375), .ZN(
        P1_U3214) );
  INV_X1 U15498 ( .A(n13428), .ZN(n13380) );
  NOR3_X1 U15499 ( .A1(n13458), .A2(n13378), .A3(n13377), .ZN(n13379) );
  OAI21_X1 U15500 ( .B1(n13380), .B2(n13379), .A(n14431), .ZN(n13386) );
  NAND2_X1 U15501 ( .A1(n13717), .A2(n14683), .ZN(n13382) );
  NAND2_X1 U15502 ( .A1(n13924), .A2(n14635), .ZN(n13381) );
  NAND2_X1 U15503 ( .A1(n13382), .A2(n13381), .ZN(n14089) );
  AOI22_X1 U15504 ( .A1(n14387), .A2(n14089), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13383) );
  OAI21_X1 U15505 ( .B1(n13919), .B2(n14436), .A(n13383), .ZN(n13384) );
  AOI21_X1 U15506 ( .B1(n13918), .B2(n14415), .A(n13384), .ZN(n13385) );
  NAND2_X1 U15507 ( .A1(n13386), .A2(n13385), .ZN(P1_U3216) );
  AOI21_X1 U15508 ( .B1(n13388), .B2(n13387), .A(n14410), .ZN(n13390) );
  NAND2_X1 U15509 ( .A1(n13390), .A2(n13389), .ZN(n13396) );
  NAND2_X1 U15510 ( .A1(n13729), .A2(n14635), .ZN(n13392) );
  NAND2_X1 U15511 ( .A1(n14636), .A2(n14683), .ZN(n13391) );
  NAND2_X1 U15512 ( .A1(n13392), .A2(n13391), .ZN(n14597) );
  AOI22_X1 U15513 ( .A1(n14387), .A2(n14597), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13395) );
  NAND2_X1 U15514 ( .A1(n14415), .A2(n14602), .ZN(n13394) );
  NAND2_X1 U15515 ( .A1(n13474), .A2(n9587), .ZN(n13393) );
  NAND4_X1 U15516 ( .A1(n13396), .A2(n13395), .A3(n13394), .A4(n13393), .ZN(
        P1_U3218) );
  INV_X1 U15517 ( .A(n13981), .ZN(n14117) );
  AND2_X1 U15518 ( .A1(n13467), .A2(n13397), .ZN(n13400) );
  OAI211_X1 U15519 ( .C1(n13400), .C2(n13399), .A(n14431), .B(n13398), .ZN(
        n13405) );
  AOI22_X1 U15520 ( .A1(n13719), .A2(n14635), .B1(n14683), .B2(n13720), .ZN(
        n14116) );
  OAI21_X1 U15521 ( .B1(n14116), .B2(n13462), .A(n13401), .ZN(n13402) );
  AOI21_X1 U15522 ( .B1(n13403), .B2(n13474), .A(n13402), .ZN(n13404) );
  OAI211_X1 U15523 ( .C1(n14117), .C2(n14423), .A(n13405), .B(n13404), .ZN(
        P1_U3219) );
  INV_X1 U15524 ( .A(n13950), .ZN(n14192) );
  OAI21_X1 U15525 ( .B1(n13407), .B2(n13406), .A(n13456), .ZN(n13408) );
  NAND2_X1 U15526 ( .A1(n13408), .A2(n14431), .ZN(n13414) );
  INV_X1 U15527 ( .A(n13409), .ZN(n13949) );
  AND2_X1 U15528 ( .A1(n13717), .A2(n14635), .ZN(n13410) );
  AOI21_X1 U15529 ( .B1(n13719), .B2(n14683), .A(n13410), .ZN(n14102) );
  INV_X1 U15530 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13411) );
  OAI22_X1 U15531 ( .A1(n14102), .A2(n13462), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13411), .ZN(n13412) );
  AOI21_X1 U15532 ( .B1(n13949), .B2(n13474), .A(n13412), .ZN(n13413) );
  OAI211_X1 U15533 ( .C1(n14192), .C2(n14423), .A(n13414), .B(n13413), .ZN(
        P1_U3223) );
  INV_X1 U15534 ( .A(n13415), .ZN(n13419) );
  NOR3_X1 U15535 ( .A1(n13430), .A2(n13417), .A3(n13416), .ZN(n13418) );
  OAI21_X1 U15536 ( .B1(n13419), .B2(n13418), .A(n14431), .ZN(n13425) );
  OAI22_X1 U15537 ( .A1(n13421), .A2(n14426), .B1(n14427), .B2(n13420), .ZN(
        n13423) );
  NOR2_X1 U15538 ( .A1(n14436), .A2(n13883), .ZN(n13422) );
  AOI211_X1 U15539 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n13423), 
        .B(n13422), .ZN(n13424) );
  OAI211_X1 U15540 ( .C1(n7208), .C2(n14423), .A(n13425), .B(n13424), .ZN(
        P1_U3225) );
  INV_X1 U15541 ( .A(n13903), .ZN(n14181) );
  AND3_X1 U15542 ( .A1(n13428), .A2(n13427), .A3(n13426), .ZN(n13429) );
  OAI21_X1 U15543 ( .B1(n13430), .B2(n13429), .A(n14431), .ZN(n13436) );
  OAI22_X1 U15544 ( .A1(n13432), .A2(n14426), .B1(n14427), .B2(n13431), .ZN(
        n13434) );
  NOR2_X1 U15545 ( .A1(n14436), .A2(n13904), .ZN(n13433) );
  AOI211_X1 U15546 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n13434), 
        .B(n13433), .ZN(n13435) );
  OAI211_X1 U15547 ( .C1(n14181), .C2(n14423), .A(n13436), .B(n13435), .ZN(
        P1_U3229) );
  XNOR2_X1 U15548 ( .A(n13438), .B(n13437), .ZN(n13445) );
  NOR2_X1 U15549 ( .A1(n14436), .A2(n13969), .ZN(n13441) );
  NAND2_X1 U15550 ( .A1(n13718), .A2(n14635), .ZN(n13962) );
  OAI22_X1 U15551 ( .A1(n13462), .A2(n13962), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13439), .ZN(n13440) );
  AOI211_X1 U15552 ( .C1(n13442), .C2(n13994), .A(n13441), .B(n13440), .ZN(
        n13444) );
  NAND2_X1 U15553 ( .A1(n13973), .A2(n14415), .ZN(n13443) );
  OAI211_X1 U15554 ( .C1(n13445), .C2(n14410), .A(n13444), .B(n13443), .ZN(
        P1_U3233) );
  NAND2_X1 U15555 ( .A1(n14387), .A2(n13446), .ZN(n13447) );
  NAND2_X1 U15556 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14519)
         );
  OAI211_X1 U15557 ( .C1(n14436), .C2(n13448), .A(n13447), .B(n14519), .ZN(
        n13452) );
  AOI211_X1 U15558 ( .C1(n13450), .C2(n13449), .A(n14410), .B(n6612), .ZN(
        n13451) );
  AOI211_X1 U15559 ( .C1(n13550), .C2(n14415), .A(n13452), .B(n13451), .ZN(
        n13453) );
  INV_X1 U15560 ( .A(n13453), .ZN(P1_U3234) );
  AND3_X1 U15561 ( .A1(n13456), .A2(n13455), .A3(n13454), .ZN(n13457) );
  OAI21_X1 U15562 ( .B1(n13458), .B2(n13457), .A(n14431), .ZN(n13466) );
  INV_X1 U15563 ( .A(n13937), .ZN(n13464) );
  NAND2_X1 U15564 ( .A1(n13718), .A2(n14683), .ZN(n13460) );
  NAND2_X1 U15565 ( .A1(n13894), .A2(n14635), .ZN(n13459) );
  AND2_X1 U15566 ( .A1(n13460), .A2(n13459), .ZN(n14096) );
  INV_X1 U15567 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13461) );
  OAI22_X1 U15568 ( .A1(n13462), .A2(n14096), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13461), .ZN(n13463) );
  AOI21_X1 U15569 ( .B1(n13464), .B2(n13474), .A(n13463), .ZN(n13465) );
  OAI211_X1 U15570 ( .C1(n14423), .C2(n14188), .A(n13466), .B(n13465), .ZN(
        P1_U3235) );
  OAI21_X1 U15571 ( .B1(n13469), .B2(n13468), .A(n13467), .ZN(n13470) );
  NAND2_X1 U15572 ( .A1(n13470), .A2(n14431), .ZN(n13476) );
  INV_X1 U15573 ( .A(n13471), .ZN(n13995) );
  NAND2_X1 U15574 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14555)
         );
  INV_X1 U15575 ( .A(n14555), .ZN(n13473) );
  OAI22_X1 U15576 ( .A1(n14124), .A2(n14426), .B1(n14427), .B2(n14123), .ZN(
        n13472) );
  AOI211_X1 U15577 ( .C1(n13474), .C2(n13995), .A(n13473), .B(n13472), .ZN(
        n13475) );
  OAI211_X1 U15578 ( .C1(n14201), .C2(n14423), .A(n13476), .B(n13475), .ZN(
        P1_U3238) );
  OAI21_X1 U15579 ( .B1(n13479), .B2(n13478), .A(n13477), .ZN(n13485) );
  NAND2_X1 U15580 ( .A1(n14174), .A2(n14415), .ZN(n13483) );
  NAND2_X1 U15581 ( .A1(n13820), .A2(n14635), .ZN(n13481) );
  NAND2_X1 U15582 ( .A1(n13895), .A2(n14683), .ZN(n13480) );
  NAND2_X1 U15583 ( .A1(n13481), .A2(n13480), .ZN(n13863) );
  AOI22_X1 U15584 ( .A1(n14387), .A2(n13863), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13482) );
  OAI211_X1 U15585 ( .C1(n14436), .C2(n13868), .A(n13483), .B(n13482), .ZN(
        n13484) );
  AOI21_X1 U15586 ( .B1(n13485), .B2(n14431), .A(n13484), .ZN(n13486) );
  INV_X1 U15587 ( .A(n13486), .ZN(P1_U3240) );
  NAND2_X1 U15588 ( .A1(n13732), .A2(n14618), .ZN(n13671) );
  NAND2_X1 U15589 ( .A1(n13671), .A2(n13487), .ZN(n13488) );
  MUX2_X1 U15590 ( .A(n13494), .B(n13493), .S(n6465), .Z(n13491) );
  NAND2_X1 U15591 ( .A1(n13492), .A2(n13491), .ZN(n13497) );
  MUX2_X1 U15592 ( .A(n13494), .B(n13493), .S(n13520), .Z(n13495) );
  AND2_X1 U15593 ( .A1(n14636), .A2(n6465), .ZN(n13500) );
  NOR2_X1 U15594 ( .A1(n14636), .A2(n6465), .ZN(n13499) );
  INV_X1 U15595 ( .A(n13501), .ZN(n13503) );
  AND2_X1 U15596 ( .A1(n13730), .A2(n13520), .ZN(n13505) );
  NOR2_X1 U15597 ( .A1(n13730), .A2(n13520), .ZN(n13504) );
  MUX2_X1 U15598 ( .A(n13505), .B(n13504), .S(n14602), .Z(n13506) );
  INV_X1 U15599 ( .A(n13506), .ZN(n13507) );
  MUX2_X1 U15600 ( .A(n14662), .B(n13729), .S(n6465), .Z(n13508) );
  INV_X1 U15601 ( .A(n13508), .ZN(n13510) );
  MUX2_X1 U15602 ( .A(n14662), .B(n13729), .S(n13520), .Z(n13509) );
  MUX2_X1 U15603 ( .A(n13511), .B(n13728), .S(n13520), .Z(n13513) );
  MUX2_X1 U15604 ( .A(n13511), .B(n13728), .S(n6465), .Z(n13512) );
  MUX2_X1 U15605 ( .A(n13515), .B(n13727), .S(n6465), .Z(n13518) );
  MUX2_X1 U15606 ( .A(n13515), .B(n13727), .S(n13520), .Z(n13516) );
  INV_X1 U15607 ( .A(n13518), .ZN(n13519) );
  MUX2_X1 U15608 ( .A(n14682), .B(n14585), .S(n6465), .Z(n13524) );
  NAND2_X1 U15609 ( .A1(n13523), .A2(n13524), .ZN(n13522) );
  MUX2_X1 U15610 ( .A(n14682), .B(n14585), .S(n13520), .Z(n13521) );
  MUX2_X1 U15611 ( .A(n13726), .B(n14684), .S(n13520), .Z(n13526) );
  MUX2_X1 U15612 ( .A(n13726), .B(n14684), .S(n6465), .Z(n13525) );
  MUX2_X1 U15613 ( .A(n13725), .B(n14570), .S(n6465), .Z(n13528) );
  MUX2_X1 U15614 ( .A(n13725), .B(n14570), .S(n13520), .Z(n13527) );
  MUX2_X1 U15615 ( .A(n13724), .B(n14702), .S(n13520), .Z(n13530) );
  MUX2_X1 U15616 ( .A(n13724), .B(n14702), .S(n6465), .Z(n13529) );
  INV_X1 U15617 ( .A(n13530), .ZN(n13531) );
  MUX2_X1 U15618 ( .A(n13723), .B(n14416), .S(n6465), .Z(n13535) );
  MUX2_X1 U15619 ( .A(n13723), .B(n14416), .S(n13520), .Z(n13532) );
  INV_X1 U15620 ( .A(n13534), .ZN(n13537) );
  INV_X1 U15621 ( .A(n13535), .ZN(n13536) );
  MUX2_X1 U15622 ( .A(n13722), .B(n13538), .S(n13520), .Z(n13540) );
  MUX2_X1 U15623 ( .A(n13722), .B(n13538), .S(n6465), .Z(n13539) );
  NAND2_X1 U15624 ( .A1(n13576), .A2(n14134), .ZN(n13541) );
  OR2_X1 U15625 ( .A1(n14437), .A2(n13520), .ZN(n13543) );
  AOI21_X1 U15626 ( .B1(n13541), .B2(n13543), .A(n14440), .ZN(n13547) );
  NAND2_X1 U15627 ( .A1(n13576), .A2(n14123), .ZN(n13542) );
  OR2_X1 U15628 ( .A1(n14390), .A2(n6465), .ZN(n13568) );
  AOI21_X1 U15629 ( .B1(n13542), .B2(n13568), .A(n7206), .ZN(n13546) );
  NAND2_X1 U15630 ( .A1(n14134), .A2(n13520), .ZN(n13569) );
  OR2_X1 U15631 ( .A1(n14390), .A2(n13569), .ZN(n13545) );
  INV_X1 U15632 ( .A(n13543), .ZN(n13572) );
  NAND2_X1 U15633 ( .A1(n14123), .A2(n13572), .ZN(n13544) );
  NAND2_X1 U15634 ( .A1(n13545), .A2(n13544), .ZN(n13575) );
  AND2_X1 U15635 ( .A1(n13562), .A2(n13548), .ZN(n13554) );
  AND2_X1 U15636 ( .A1(n13563), .A2(n13549), .ZN(n13560) );
  MUX2_X1 U15637 ( .A(n14446), .B(n13550), .S(n6465), .Z(n13555) );
  NOR2_X1 U15638 ( .A1(n14446), .A2(n13520), .ZN(n13553) );
  NOR2_X1 U15639 ( .A1(n13550), .A2(n6465), .ZN(n13556) );
  OR3_X1 U15640 ( .A1(n13555), .A2(n13553), .A3(n13556), .ZN(n13551) );
  AND4_X1 U15641 ( .A1(n13581), .A2(n13554), .A3(n13560), .A4(n13551), .ZN(
        n13552) );
  AOI22_X1 U15642 ( .A1(n13689), .A2(n6465), .B1(n13553), .B2(n13555), .ZN(
        n13567) );
  INV_X1 U15643 ( .A(n13554), .ZN(n13566) );
  INV_X1 U15644 ( .A(n13555), .ZN(n13558) );
  INV_X1 U15645 ( .A(n13556), .ZN(n13557) );
  OAI22_X1 U15646 ( .A1(n13559), .A2(n6465), .B1(n13558), .B2(n13557), .ZN(
        n13561) );
  NAND2_X1 U15647 ( .A1(n13561), .A2(n13560), .ZN(n13565) );
  MUX2_X1 U15648 ( .A(n13563), .B(n13562), .S(n13520), .Z(n13564) );
  OAI211_X1 U15649 ( .C1(n13567), .C2(n13566), .A(n13565), .B(n13564), .ZN(
        n13582) );
  INV_X1 U15650 ( .A(n13568), .ZN(n13571) );
  INV_X1 U15651 ( .A(n13569), .ZN(n13570) );
  AOI21_X1 U15652 ( .B1(n13576), .B2(n13571), .A(n13570), .ZN(n13579) );
  NAND2_X1 U15653 ( .A1(n13576), .A2(n13572), .ZN(n13573) );
  OAI21_X1 U15654 ( .B1(n13520), .B2(n14134), .A(n13573), .ZN(n13574) );
  NAND2_X1 U15655 ( .A1(n13574), .A2(n7206), .ZN(n13578) );
  NAND2_X1 U15656 ( .A1(n13576), .A2(n13575), .ZN(n13577) );
  OAI211_X1 U15657 ( .C1(n13579), .C2(n7206), .A(n13578), .B(n13577), .ZN(
        n13580) );
  AOI21_X1 U15658 ( .B1(n13582), .B2(n13581), .A(n13580), .ZN(n13583) );
  NAND2_X1 U15659 ( .A1(n13584), .A2(n13583), .ZN(n13588) );
  MUX2_X1 U15660 ( .A(n14397), .B(n14201), .S(n13520), .Z(n13585) );
  NAND2_X1 U15661 ( .A1(n13994), .A2(n6465), .ZN(n13590) );
  OR2_X1 U15662 ( .A1(n13994), .A2(n6465), .ZN(n13589) );
  MUX2_X1 U15663 ( .A(n13590), .B(n13589), .S(n13981), .Z(n13591) );
  MUX2_X1 U15664 ( .A(n13592), .B(n14196), .S(n6465), .Z(n13594) );
  MUX2_X1 U15665 ( .A(n13719), .B(n13973), .S(n13520), .Z(n13593) );
  MUX2_X1 U15666 ( .A(n13718), .B(n13950), .S(n13520), .Z(n13597) );
  NAND2_X1 U15667 ( .A1(n13598), .A2(n13597), .ZN(n13596) );
  MUX2_X1 U15668 ( .A(n13718), .B(n13950), .S(n6465), .Z(n13595) );
  NAND2_X1 U15669 ( .A1(n13596), .A2(n13595), .ZN(n13600) );
  MUX2_X1 U15670 ( .A(n13717), .B(n13601), .S(n6465), .Z(n13603) );
  MUX2_X1 U15671 ( .A(n13717), .B(n13601), .S(n13520), .Z(n13602) );
  MUX2_X1 U15672 ( .A(n13894), .B(n13918), .S(n13520), .Z(n13605) );
  MUX2_X1 U15673 ( .A(n13894), .B(n13918), .S(n6465), .Z(n13604) );
  MUX2_X1 U15674 ( .A(n13924), .B(n13903), .S(n6465), .Z(n13609) );
  MUX2_X1 U15675 ( .A(n13924), .B(n13903), .S(n13520), .Z(n13607) );
  NAND2_X1 U15676 ( .A1(n13608), .A2(n13607), .ZN(n13611) );
  MUX2_X1 U15677 ( .A(n13895), .B(n14078), .S(n6465), .Z(n13612) );
  INV_X1 U15678 ( .A(n13613), .ZN(n13614) );
  MUX2_X1 U15679 ( .A(n13879), .B(n14174), .S(n6465), .Z(n13617) );
  MUX2_X1 U15680 ( .A(n13879), .B(n14174), .S(n13520), .Z(n13615) );
  MUX2_X1 U15681 ( .A(n13820), .B(n13618), .S(n13520), .Z(n13620) );
  MUX2_X1 U15682 ( .A(n13820), .B(n13618), .S(n6465), .Z(n13619) );
  MUX2_X1 U15683 ( .A(n14050), .B(n13830), .S(n6465), .Z(n13624) );
  MUX2_X1 U15684 ( .A(n14050), .B(n13830), .S(n13520), .Z(n13621) );
  NAND2_X1 U15685 ( .A1(n13622), .A2(n13621), .ZN(n13628) );
  INV_X1 U15686 ( .A(n13623), .ZN(n13626) );
  INV_X1 U15687 ( .A(n13624), .ZN(n13625) );
  NAND2_X1 U15688 ( .A1(n13626), .A2(n13625), .ZN(n13627) );
  MUX2_X1 U15689 ( .A(n13821), .B(n13629), .S(n13520), .Z(n13631) );
  NAND2_X1 U15690 ( .A1(n13630), .A2(n13631), .ZN(n13634) );
  MUX2_X1 U15691 ( .A(n13821), .B(n13629), .S(n6465), .Z(n13633) );
  INV_X1 U15692 ( .A(n13631), .ZN(n13632) );
  NAND2_X1 U15693 ( .A1(n13635), .A2(n6468), .ZN(n13637) );
  OR2_X1 U15694 ( .A1(n13653), .A2(n14219), .ZN(n13636) );
  INV_X1 U15695 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14043) );
  OR2_X1 U15696 ( .A1(n6463), .A2(n14043), .ZN(n13642) );
  INV_X1 U15697 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13807) );
  OR2_X1 U15698 ( .A1(n13638), .A2(n13807), .ZN(n13641) );
  INV_X1 U15699 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14157) );
  OR2_X1 U15700 ( .A1(n13639), .A2(n14157), .ZN(n13640) );
  INV_X1 U15701 ( .A(n13643), .ZN(n13644) );
  OAI22_X1 U15702 ( .A1(n13806), .A2(n6465), .B1(n13645), .B2(n13644), .ZN(
        n13646) );
  AOI22_X1 U15703 ( .A1(n13815), .A2(n6465), .B1(n13716), .B2(n13646), .ZN(
        n13650) );
  INV_X1 U15704 ( .A(n13806), .ZN(n13715) );
  OAI21_X1 U15705 ( .B1(n13715), .B2(n13647), .A(n13716), .ZN(n13648) );
  MUX2_X1 U15706 ( .A(n13648), .B(n14163), .S(n13520), .Z(n13652) );
  INV_X1 U15707 ( .A(n13650), .ZN(n13651) );
  NAND2_X1 U15708 ( .A1(n14216), .A2(n6468), .ZN(n13655) );
  INV_X1 U15709 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14211) );
  OR2_X1 U15710 ( .A1(n13653), .A2(n14211), .ZN(n13654) );
  XNOR2_X1 U15711 ( .A(n14040), .B(n13806), .ZN(n13668) );
  NAND2_X1 U15712 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  NAND2_X1 U15713 ( .A1(n13659), .A2(n13658), .ZN(n13661) );
  NAND2_X1 U15714 ( .A1(n13661), .A2(n13660), .ZN(n13702) );
  NOR2_X1 U15715 ( .A1(n14040), .A2(n13806), .ZN(n13663) );
  AND2_X1 U15716 ( .A1(n14040), .A2(n13806), .ZN(n13662) );
  MUX2_X1 U15717 ( .A(n13663), .B(n13662), .S(n13520), .Z(n13705) );
  NAND2_X1 U15718 ( .A1(n13665), .A2(n13664), .ZN(n13700) );
  NAND2_X1 U15719 ( .A1(n13702), .A2(n13700), .ZN(n13703) );
  INV_X1 U15720 ( .A(n13703), .ZN(n13666) );
  INV_X1 U15721 ( .A(n13668), .ZN(n13704) );
  NAND2_X1 U15722 ( .A1(n13670), .A2(n13669), .ZN(n14008) );
  AND2_X1 U15723 ( .A1(n13672), .A2(n13671), .ZN(n14628) );
  NAND4_X1 U15724 ( .A1(n13675), .A2(n14628), .A3(n13674), .A4(n13673), .ZN(
        n13677) );
  NOR4_X1 U15725 ( .A1(n14593), .A2(n13678), .A3(n13677), .A4(n13676), .ZN(
        n13680) );
  NAND4_X1 U15726 ( .A1(n13680), .A2(n14561), .A3(n13679), .A4(n14578), .ZN(
        n13681) );
  NOR4_X1 U15727 ( .A1(n13684), .A2(n13683), .A3(n13682), .A4(n13681), .ZN(
        n13687) );
  NAND4_X1 U15728 ( .A1(n14008), .A2(n13687), .A3(n13686), .A4(n13685), .ZN(
        n13690) );
  NOR3_X1 U15729 ( .A1(n13690), .A2(n13689), .A3(n13688), .ZN(n13691) );
  NAND4_X1 U15730 ( .A1(n13967), .A2(n13691), .A3(n7246), .A4(n13993), .ZN(
        n13692) );
  NOR4_X1 U15731 ( .A1(n13912), .A2(n13930), .A3(n13953), .A4(n13692), .ZN(
        n13693) );
  NAND4_X1 U15732 ( .A1(n13861), .A2(n13693), .A3(n13897), .A4(n13877), .ZN(
        n13694) );
  NOR3_X1 U15733 ( .A1(n13818), .A2(n13695), .A3(n13694), .ZN(n13698) );
  XOR2_X1 U15734 ( .A(n13716), .B(n14163), .Z(n13697) );
  NAND4_X1 U15735 ( .A1(n13704), .A2(n13698), .A3(n13697), .A4(n13696), .ZN(
        n13699) );
  XNOR2_X1 U15736 ( .A(n13699), .B(n14614), .ZN(n13701) );
  NOR2_X1 U15737 ( .A1(n13701), .A2(n13700), .ZN(n13710) );
  INV_X1 U15738 ( .A(n13702), .ZN(n13708) );
  NOR2_X1 U15739 ( .A1(n13704), .A2(n13703), .ZN(n13707) );
  INV_X1 U15740 ( .A(n13705), .ZN(n13706) );
  MUX2_X1 U15741 ( .A(n13708), .B(n13707), .S(n13706), .Z(n13709) );
  NAND3_X1 U15742 ( .A1(n13711), .A2(n7231), .A3(n14683), .ZN(n13712) );
  OAI211_X1 U15743 ( .C1(n14225), .C2(n13714), .A(n13712), .B(P1_B_REG_SCAN_IN), .ZN(n13713) );
  MUX2_X1 U15744 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13715), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15745 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13716), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15746 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13821), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15747 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14050), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15748 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13820), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15749 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13879), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15750 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13895), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15751 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13924), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15752 ( .A(n13894), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13721), .Z(
        P1_U3583) );
  MUX2_X1 U15753 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13717), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15754 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13718), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15755 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13719), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15756 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13994), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15757 ( .A(n13720), .B(P1_DATAO_REG_18__SCAN_IN), .S(n13721), .Z(
        P1_U3578) );
  MUX2_X1 U15758 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14134), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15759 ( .A(n14437), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13721), .Z(
        P1_U3576) );
  MUX2_X1 U15760 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14447), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15761 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14147), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15762 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14446), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15763 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13722), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15764 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13723), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15765 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13724), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15766 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13725), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15767 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13726), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15768 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14682), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15769 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13727), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15770 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13728), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15771 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13729), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15772 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13730), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15773 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14636), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15774 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13731), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15775 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13732), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U15776 ( .C1(n13735), .C2(n13734), .A(n14548), .B(n13733), .ZN(
        n13745) );
  MUX2_X1 U15777 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9074), .S(n13736), .Z(
        n13737) );
  OAI21_X1 U15778 ( .B1(n14495), .B2(n13738), .A(n13737), .ZN(n13739) );
  NAND3_X1 U15779 ( .A1(n14545), .A2(n13740), .A3(n13739), .ZN(n13744) );
  NAND2_X1 U15780 ( .A1(n13797), .A2(n13741), .ZN(n13743) );
  AOI22_X1 U15781 ( .A1(n14517), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13742) );
  NAND4_X1 U15782 ( .A1(n13745), .A2(n13744), .A3(n13743), .A4(n13742), .ZN(
        P1_U3244) );
  OAI22_X1 U15783 ( .A1(n14557), .A2(n14292), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9587), .ZN(n13746) );
  AOI21_X1 U15784 ( .B1(n13747), .B2(n13797), .A(n13746), .ZN(n13760) );
  MUX2_X1 U15785 ( .A(n9297), .B(P1_REG1_REG_3__SCAN_IN), .S(n13747), .Z(
        n13748) );
  NAND3_X1 U15786 ( .A1(n13750), .A2(n13749), .A3(n13748), .ZN(n13751) );
  NAND3_X1 U15787 ( .A1(n14545), .A2(n13752), .A3(n13751), .ZN(n13759) );
  NAND3_X1 U15788 ( .A1(n13755), .A2(n13754), .A3(n13753), .ZN(n13756) );
  NAND3_X1 U15789 ( .A1(n14548), .A2(n13757), .A3(n13756), .ZN(n13758) );
  NAND3_X1 U15790 ( .A1(n13760), .A2(n13759), .A3(n13758), .ZN(P1_U3246) );
  OAI21_X1 U15791 ( .B1(n14557), .B2(n14300), .A(n13761), .ZN(n13762) );
  AOI21_X1 U15792 ( .B1(n13763), .B2(n13797), .A(n13762), .ZN(n13778) );
  OAI21_X1 U15793 ( .B1(n13766), .B2(n13765), .A(n13764), .ZN(n13767) );
  NAND2_X1 U15794 ( .A1(n14545), .A2(n13767), .ZN(n13777) );
  INV_X1 U15795 ( .A(n13768), .ZN(n13772) );
  INV_X1 U15796 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n13770) );
  MUX2_X1 U15797 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n13770), .S(n13769), .Z(
        n13771) );
  NAND3_X1 U15798 ( .A1(n13773), .A2(n13772), .A3(n13771), .ZN(n13774) );
  NAND3_X1 U15799 ( .A1(n14548), .A2(n13775), .A3(n13774), .ZN(n13776) );
  NAND3_X1 U15800 ( .A1(n13778), .A2(n13777), .A3(n13776), .ZN(P1_U3248) );
  OAI21_X1 U15801 ( .B1(n13780), .B2(n13779), .A(n14504), .ZN(n13781) );
  NAND2_X1 U15802 ( .A1(n13781), .A2(n14545), .ZN(n13791) );
  NAND2_X1 U15803 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14417)
         );
  OAI21_X1 U15804 ( .B1(n14557), .B2(n14255), .A(n14417), .ZN(n13782) );
  AOI21_X1 U15805 ( .B1(n13797), .B2(n13783), .A(n13782), .ZN(n13790) );
  OR3_X1 U15806 ( .A1(n13786), .A2(n13785), .A3(n13784), .ZN(n13787) );
  NAND3_X1 U15807 ( .A1(n13788), .A2(n14548), .A3(n13787), .ZN(n13789) );
  NAND3_X1 U15808 ( .A1(n13791), .A2(n13790), .A3(n13789), .ZN(P1_U3254) );
  NAND2_X1 U15809 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14391)
         );
  OAI211_X1 U15810 ( .C1(n13794), .C2(n13793), .A(n13792), .B(n14545), .ZN(
        n13795) );
  AND2_X1 U15811 ( .A1(n14391), .A2(n13795), .ZN(n13803) );
  AOI22_X1 U15812 ( .A1(n13797), .A2(n13796), .B1(n14517), .B2(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n13802) );
  OAI211_X1 U15813 ( .C1(n13800), .C2(n13799), .A(n13798), .B(n14548), .ZN(
        n13801) );
  NAND3_X1 U15814 ( .A1(n13803), .A2(n13802), .A3(n13801), .ZN(P1_U3259) );
  NAND2_X1 U15815 ( .A1(n13804), .A2(n14604), .ZN(n14042) );
  OR2_X1 U15816 ( .A1(n13806), .A2(n13805), .ZN(n14041) );
  INV_X1 U15817 ( .A(n14041), .ZN(n14045) );
  NAND2_X1 U15818 ( .A1(n6464), .A2(n14045), .ZN(n13812) );
  OAI21_X1 U15819 ( .B1(n6464), .B2(n13807), .A(n13812), .ZN(n13808) );
  AOI21_X1 U15820 ( .B1(n14040), .B2(n14601), .A(n13808), .ZN(n13809) );
  OAI21_X1 U15821 ( .B1(n14042), .B2(n14035), .A(n13809), .ZN(P1_U3263) );
  AOI211_X1 U15822 ( .C1(n13815), .C2(n13811), .A(n13980), .B(n13810), .ZN(
        n14046) );
  INV_X1 U15823 ( .A(n14046), .ZN(n13817) );
  OAI21_X1 U15824 ( .B1(n6464), .B2(n13813), .A(n13812), .ZN(n13814) );
  AOI21_X1 U15825 ( .B1(n13815), .B2(n14601), .A(n13814), .ZN(n13816) );
  OAI21_X1 U15826 ( .B1(n13817), .B2(n14035), .A(n13816), .ZN(P1_U3264) );
  INV_X1 U15827 ( .A(n13818), .ZN(n13826) );
  XNOR2_X1 U15828 ( .A(n13819), .B(n13826), .ZN(n13824) );
  AOI22_X1 U15829 ( .A1(n14635), .A2(n13821), .B1(n13820), .B2(n14683), .ZN(
        n13822) );
  INV_X1 U15830 ( .A(n13825), .ZN(n13827) );
  NAND2_X1 U15831 ( .A1(n13827), .A2(n13826), .ZN(n13828) );
  AOI21_X1 U15832 ( .B1(n13850), .B2(n13830), .A(n13980), .ZN(n13832) );
  NAND2_X1 U15833 ( .A1(n14057), .A2(n14609), .ZN(n13836) );
  INV_X1 U15834 ( .A(n13833), .ZN(n13834) );
  AOI22_X1 U15835 ( .A1(n14016), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n13834), 
        .B2(n14621), .ZN(n13835) );
  OAI211_X1 U15836 ( .C1(n14168), .C2(n13982), .A(n13836), .B(n13835), .ZN(
        n13837) );
  AOI21_X1 U15837 ( .B1(n14061), .B2(n14624), .A(n13837), .ZN(n13838) );
  OAI21_X1 U15838 ( .B1(n14059), .B2(n14016), .A(n13838), .ZN(P1_U3265) );
  OAI21_X1 U15839 ( .B1(n13840), .B2(n13843), .A(n13839), .ZN(n13841) );
  NAND2_X1 U15840 ( .A1(n13841), .A2(n14699), .ZN(n13849) );
  AOI22_X1 U15841 ( .A1(n14635), .A2(n14050), .B1(n13879), .B2(n14683), .ZN(
        n13848) );
  NAND2_X1 U15842 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  NAND2_X1 U15843 ( .A1(n13846), .A2(n13845), .ZN(n14063) );
  NAND2_X1 U15844 ( .A1(n14063), .A2(n14598), .ZN(n13847) );
  NAND3_X1 U15845 ( .A1(n13849), .A2(n13848), .A3(n13847), .ZN(n14068) );
  INV_X1 U15846 ( .A(n14068), .ZN(n13857) );
  OAI211_X1 U15847 ( .C1(n14066), .C2(n13867), .A(n14604), .B(n13850), .ZN(
        n14064) );
  NOR2_X1 U15848 ( .A1(n14064), .A2(n14035), .ZN(n13855) );
  INV_X1 U15849 ( .A(n13851), .ZN(n13852) );
  AOI22_X1 U15850 ( .A1(n14016), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13852), 
        .B2(n14621), .ZN(n13853) );
  OAI21_X1 U15851 ( .B1(n14066), .B2(n13982), .A(n13853), .ZN(n13854) );
  AOI211_X1 U15852 ( .C1(n14063), .C2(n14610), .A(n13855), .B(n13854), .ZN(
        n13856) );
  OAI21_X1 U15853 ( .B1(n13857), .B2(n14016), .A(n13856), .ZN(P1_U3266) );
  XNOR2_X1 U15854 ( .A(n13859), .B(n13858), .ZN(n14073) );
  OAI21_X1 U15855 ( .B1(n13862), .B2(n13861), .A(n13860), .ZN(n13864) );
  AOI21_X1 U15856 ( .B1(n13864), .B2(n14699), .A(n13863), .ZN(n14072) );
  INV_X1 U15857 ( .A(n14072), .ZN(n13873) );
  NAND2_X1 U15858 ( .A1(n14174), .A2(n13881), .ZN(n13865) );
  NAND2_X1 U15859 ( .A1(n13865), .A2(n14604), .ZN(n13866) );
  OR2_X1 U15860 ( .A1(n13867), .A2(n13866), .ZN(n14071) );
  INV_X1 U15861 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13869) );
  OAI22_X1 U15862 ( .A1(n6464), .A2(n13869), .B1(n13868), .B2(n14599), .ZN(
        n13870) );
  AOI21_X1 U15863 ( .B1(n14174), .B2(n14601), .A(n13870), .ZN(n13871) );
  OAI21_X1 U15864 ( .B1(n14071), .B2(n14035), .A(n13871), .ZN(n13872) );
  AOI21_X1 U15865 ( .B1(n13873), .B2(n6464), .A(n13872), .ZN(n13874) );
  OAI21_X1 U15866 ( .B1(n14073), .B2(n14004), .A(n13874), .ZN(P1_U3267) );
  AND2_X1 U15867 ( .A1(n13896), .A2(n13875), .ZN(n13878) );
  OAI21_X1 U15868 ( .B1(n13878), .B2(n13877), .A(n13876), .ZN(n13880) );
  AOI222_X1 U15869 ( .A1(n14699), .A2(n13880), .B1(n13924), .B2(n14683), .C1(
        n13879), .C2(n14635), .ZN(n14080) );
  INV_X1 U15870 ( .A(n13881), .ZN(n13882) );
  AOI211_X1 U15871 ( .C1(n14078), .C2(n13901), .A(n13980), .B(n13882), .ZN(
        n14077) );
  INV_X1 U15872 ( .A(n13883), .ZN(n13884) );
  AOI22_X1 U15873 ( .A1(n14016), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n13884), 
        .B2(n14621), .ZN(n13885) );
  OAI21_X1 U15874 ( .B1(n7208), .B2(n13982), .A(n13885), .ZN(n13890) );
  OAI21_X1 U15875 ( .B1(n13888), .B2(n13887), .A(n13886), .ZN(n14081) );
  NOR2_X1 U15876 ( .A1(n14081), .A2(n14004), .ZN(n13889) );
  AOI211_X1 U15877 ( .C1(n14077), .C2(n14609), .A(n13890), .B(n13889), .ZN(
        n13891) );
  OAI21_X1 U15878 ( .B1(n14080), .B2(n14016), .A(n13891), .ZN(P1_U3268) );
  AOI21_X1 U15879 ( .B1(n13897), .B2(n13893), .A(n13892), .ZN(n14082) );
  AOI22_X1 U15880 ( .A1(n14635), .A2(n13895), .B1(n13894), .B2(n14683), .ZN(
        n13900) );
  OAI211_X1 U15881 ( .C1(n13898), .C2(n13897), .A(n14699), .B(n13896), .ZN(
        n13899) );
  OAI211_X1 U15882 ( .C1(n14082), .C2(n14647), .A(n13900), .B(n13899), .ZN(
        n14083) );
  NAND2_X1 U15883 ( .A1(n14083), .A2(n6464), .ZN(n13909) );
  AOI211_X1 U15884 ( .C1(n13903), .C2(n13902), .A(n13980), .B(n7209), .ZN(
        n14084) );
  NOR2_X1 U15885 ( .A1(n14181), .A2(n13982), .ZN(n13907) );
  OAI22_X1 U15886 ( .A1(n6464), .A2(n13905), .B1(n13904), .B2(n14599), .ZN(
        n13906) );
  AOI211_X1 U15887 ( .C1(n14084), .C2(n14609), .A(n13907), .B(n13906), .ZN(
        n13908) );
  OAI211_X1 U15888 ( .C1(n14082), .C2(n13910), .A(n13909), .B(n13908), .ZN(
        P1_U3269) );
  OAI21_X1 U15889 ( .B1(n7685), .B2(n13912), .A(n13911), .ZN(n14088) );
  OAI21_X1 U15890 ( .B1(n13915), .B2(n13914), .A(n13913), .ZN(n13916) );
  AND2_X1 U15891 ( .A1(n13916), .A2(n14699), .ZN(n14092) );
  NAND2_X1 U15892 ( .A1(n14092), .A2(n6464), .ZN(n13928) );
  XNOR2_X1 U15893 ( .A(n13918), .B(n13935), .ZN(n13917) );
  NOR2_X1 U15894 ( .A1(n13917), .A2(n13980), .ZN(n14090) );
  OAI22_X1 U15895 ( .A1(n6464), .A2(n13920), .B1(n13919), .B2(n14599), .ZN(
        n13923) );
  NOR2_X1 U15896 ( .A1(n14029), .A2(n13921), .ZN(n13922) );
  AOI211_X1 U15897 ( .C1(n14032), .C2(n13924), .A(n13923), .B(n13922), .ZN(
        n13925) );
  OAI21_X1 U15898 ( .B1(n7210), .B2(n13982), .A(n13925), .ZN(n13926) );
  AOI21_X1 U15899 ( .B1(n14090), .B2(n14609), .A(n13926), .ZN(n13927) );
  OAI211_X1 U15900 ( .C1(n14088), .C2(n14004), .A(n13928), .B(n13927), .ZN(
        P1_U3270) );
  OAI21_X1 U15901 ( .B1(n13931), .B2(n13930), .A(n13929), .ZN(n13932) );
  INV_X1 U15902 ( .A(n13932), .ZN(n14097) );
  XNOR2_X1 U15903 ( .A(n13934), .B(n13933), .ZN(n14099) );
  NAND2_X1 U15904 ( .A1(n14099), .A2(n14623), .ZN(n13943) );
  INV_X1 U15905 ( .A(n13947), .ZN(n13936) );
  OAI211_X1 U15906 ( .C1(n14188), .C2(n13936), .A(n14604), .B(n13935), .ZN(
        n14095) );
  INV_X1 U15907 ( .A(n14095), .ZN(n13941) );
  OAI22_X1 U15908 ( .A1(n14016), .A2(n14096), .B1(n13937), .B2(n14599), .ZN(
        n13938) );
  AOI21_X1 U15909 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n14016), .A(n13938), 
        .ZN(n13939) );
  OAI21_X1 U15910 ( .B1(n14188), .B2(n13982), .A(n13939), .ZN(n13940) );
  AOI21_X1 U15911 ( .B1(n13941), .B2(n14609), .A(n13940), .ZN(n13942) );
  OAI211_X1 U15912 ( .C1(n14097), .C2(n14004), .A(n13943), .B(n13942), .ZN(
        P1_U3271) );
  XNOR2_X1 U15913 ( .A(n13945), .B(n13944), .ZN(n14105) );
  AOI21_X1 U15914 ( .B1(n13946), .B2(n13950), .A(n13980), .ZN(n13948) );
  NAND2_X1 U15915 ( .A1(n13948), .A2(n13947), .ZN(n14103) );
  AOI22_X1 U15916 ( .A1(n14016), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n13949), 
        .B2(n14621), .ZN(n13952) );
  NAND2_X1 U15917 ( .A1(n13950), .A2(n14601), .ZN(n13951) );
  OAI211_X1 U15918 ( .C1(n14103), .C2(n14035), .A(n13952), .B(n13951), .ZN(
        n13957) );
  XNOR2_X1 U15919 ( .A(n13954), .B(n13953), .ZN(n13955) );
  NAND2_X1 U15920 ( .A1(n13955), .A2(n14699), .ZN(n14107) );
  AOI21_X1 U15921 ( .B1(n14107), .B2(n14102), .A(n14016), .ZN(n13956) );
  AOI211_X1 U15922 ( .C1(n14624), .C2(n14105), .A(n13957), .B(n13956), .ZN(
        n13958) );
  INV_X1 U15923 ( .A(n13958), .ZN(P1_U3272) );
  INV_X1 U15924 ( .A(n13959), .ZN(n13961) );
  OAI211_X1 U15925 ( .C1(n13961), .C2(n13967), .A(n14699), .B(n13960), .ZN(
        n13963) );
  NAND2_X1 U15926 ( .A1(n13963), .A2(n13962), .ZN(n14111) );
  INV_X1 U15927 ( .A(n14111), .ZN(n13977) );
  INV_X1 U15928 ( .A(n13964), .ZN(n13965) );
  AOI21_X1 U15929 ( .B1(n13967), .B2(n13966), .A(n13965), .ZN(n14113) );
  XNOR2_X1 U15930 ( .A(n13979), .B(n13973), .ZN(n13968) );
  NAND2_X1 U15931 ( .A1(n13968), .A2(n14604), .ZN(n14110) );
  NOR2_X1 U15932 ( .A1(n14124), .A2(n14029), .ZN(n13972) );
  OAI22_X1 U15933 ( .A1(n6464), .A2(n13970), .B1(n13969), .B2(n14599), .ZN(
        n13971) );
  AOI211_X1 U15934 ( .C1(n13973), .C2(n14601), .A(n13972), .B(n13971), .ZN(
        n13974) );
  OAI21_X1 U15935 ( .B1(n14110), .B2(n14035), .A(n13974), .ZN(n13975) );
  AOI21_X1 U15936 ( .B1(n14113), .B2(n14624), .A(n13975), .ZN(n13976) );
  OAI21_X1 U15937 ( .B1(n13977), .B2(n14016), .A(n13976), .ZN(P1_U3273) );
  XNOR2_X1 U15938 ( .A(n13978), .B(n7246), .ZN(n14122) );
  AOI211_X1 U15939 ( .C1(n13981), .C2(n13998), .A(n13980), .B(n13979), .ZN(
        n14119) );
  NOR2_X1 U15940 ( .A1(n14117), .A2(n13982), .ZN(n13986) );
  OAI21_X1 U15941 ( .B1(n14599), .B2(n13983), .A(n14116), .ZN(n13984) );
  MUX2_X1 U15942 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13984), .S(n6464), .Z(
        n13985) );
  AOI211_X1 U15943 ( .C1(n14119), .C2(n14609), .A(n13986), .B(n13985), .ZN(
        n13990) );
  XNOR2_X1 U15944 ( .A(n13988), .B(n13987), .ZN(n14120) );
  NAND2_X1 U15945 ( .A1(n14120), .A2(n14624), .ZN(n13989) );
  OAI211_X1 U15946 ( .C1(n14122), .C2(n14038), .A(n13990), .B(n13989), .ZN(
        P1_U3274) );
  XOR2_X1 U15947 ( .A(n13993), .B(n13991), .Z(n14128) );
  XOR2_X1 U15948 ( .A(n13993), .B(n13992), .Z(n14130) );
  NAND2_X1 U15949 ( .A1(n14130), .A2(n14623), .ZN(n14003) );
  NAND2_X1 U15950 ( .A1(n13994), .A2(n14032), .ZN(n13997) );
  AOI22_X1 U15951 ( .A1(n14016), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13995), 
        .B2(n14621), .ZN(n13996) );
  OAI211_X1 U15952 ( .C1(n14123), .C2(n14029), .A(n13997), .B(n13996), .ZN(
        n14000) );
  OAI211_X1 U15953 ( .C1(n14010), .C2(n14201), .A(n14604), .B(n13998), .ZN(
        n14126) );
  NOR2_X1 U15954 ( .A1(n14126), .A2(n14035), .ZN(n13999) );
  AOI211_X1 U15955 ( .C1(n14601), .C2(n14001), .A(n14000), .B(n13999), .ZN(
        n14002) );
  OAI211_X1 U15956 ( .C1(n14128), .C2(n14004), .A(n14003), .B(n14002), .ZN(
        P1_U3275) );
  XOR2_X1 U15957 ( .A(n14008), .B(n14005), .Z(n14006) );
  OAI22_X1 U15958 ( .A1(n14006), .A2(n14629), .B1(n14397), .B2(n14615), .ZN(
        n14441) );
  INV_X1 U15959 ( .A(n14441), .ZN(n14017) );
  XOR2_X1 U15960 ( .A(n14008), .B(n14007), .Z(n14443) );
  OAI21_X1 U15961 ( .B1(n14027), .B2(n14440), .A(n14604), .ZN(n14009) );
  OR2_X1 U15962 ( .A1(n14010), .A2(n14009), .ZN(n14439) );
  NOR2_X1 U15963 ( .A1(n14029), .A2(n14425), .ZN(n14012) );
  OAI22_X1 U15964 ( .A1(n6464), .A2(n10410), .B1(n14403), .B2(n14599), .ZN(
        n14011) );
  AOI211_X1 U15965 ( .C1(n7206), .C2(n14601), .A(n14012), .B(n14011), .ZN(
        n14013) );
  OAI21_X1 U15966 ( .B1(n14439), .B2(n14035), .A(n14013), .ZN(n14014) );
  AOI21_X1 U15967 ( .B1(n14443), .B2(n14624), .A(n14014), .ZN(n14015) );
  OAI21_X1 U15968 ( .B1(n14017), .B2(n14016), .A(n14015), .ZN(P1_U3276) );
  NAND2_X1 U15969 ( .A1(n14018), .A2(n14021), .ZN(n14019) );
  NAND2_X1 U15970 ( .A1(n14020), .A2(n14019), .ZN(n14133) );
  INV_X1 U15971 ( .A(n14133), .ZN(n14039) );
  OR2_X1 U15972 ( .A1(n14022), .A2(n14021), .ZN(n14023) );
  NAND2_X1 U15973 ( .A1(n14024), .A2(n14023), .ZN(n14140) );
  OAI21_X1 U15974 ( .B1(n14025), .B2(n14205), .A(n14604), .ZN(n14026) );
  OR2_X1 U15975 ( .A1(n14027), .A2(n14026), .ZN(n14138) );
  OAI22_X1 U15976 ( .A1(n6464), .A2(n14028), .B1(n14393), .B2(n14599), .ZN(
        n14031) );
  NOR2_X1 U15977 ( .A1(n14029), .A2(n14374), .ZN(n14030) );
  AOI211_X1 U15978 ( .C1(n14032), .C2(n14134), .A(n14031), .B(n14030), .ZN(
        n14034) );
  NAND2_X1 U15979 ( .A1(n14390), .A2(n14601), .ZN(n14033) );
  OAI211_X1 U15980 ( .C1(n14138), .C2(n14035), .A(n14034), .B(n14033), .ZN(
        n14036) );
  AOI21_X1 U15981 ( .B1(n14140), .B2(n14624), .A(n14036), .ZN(n14037) );
  OAI21_X1 U15982 ( .B1(n14039), .B2(n14038), .A(n14037), .ZN(P1_U3277) );
  INV_X1 U15983 ( .A(n14040), .ZN(n14159) );
  MUX2_X1 U15984 ( .A(n14043), .B(n14156), .S(n14730), .Z(n14044) );
  OAI21_X1 U15985 ( .B1(n14159), .B2(n14155), .A(n14044), .ZN(P1_U3559) );
  INV_X1 U15986 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14047) );
  NOR2_X1 U15987 ( .A1(n14046), .A2(n14045), .ZN(n14160) );
  MUX2_X1 U15988 ( .A(n14047), .B(n14160), .S(n14730), .Z(n14048) );
  OAI21_X1 U15989 ( .B1(n14163), .B2(n14155), .A(n14048), .ZN(P1_U3558) );
  AOI21_X1 U15990 ( .B1(n14683), .B2(n14050), .A(n14049), .ZN(n14051) );
  OAI211_X1 U15991 ( .C1(n7198), .C2(n14691), .A(n14052), .B(n14051), .ZN(
        n14053) );
  AOI21_X1 U15992 ( .B1(n14054), .B2(n14699), .A(n14053), .ZN(n14055) );
  OAI21_X1 U15993 ( .B1(n14056), .B2(n14639), .A(n14055), .ZN(n14164) );
  MUX2_X1 U15994 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14164), .S(n14730), .Z(
        P1_U3557) );
  INV_X1 U15995 ( .A(n14057), .ZN(n14058) );
  AOI21_X1 U15996 ( .B1(n14061), .B2(n14708), .A(n14060), .ZN(n14166) );
  NAND2_X1 U15997 ( .A1(n14063), .A2(n14697), .ZN(n14065) );
  OAI211_X1 U15998 ( .C1(n14066), .C2(n14691), .A(n14065), .B(n14064), .ZN(
        n14067) );
  NOR2_X1 U15999 ( .A1(n14068), .A2(n14067), .ZN(n14169) );
  MUX2_X1 U16000 ( .A(n14069), .B(n14169), .S(n14730), .Z(n14070) );
  INV_X1 U16001 ( .A(n14070), .ZN(P1_U3555) );
  INV_X1 U16002 ( .A(n14155), .ZN(n14075) );
  OAI211_X1 U16003 ( .C1(n14639), .C2(n14073), .A(n14072), .B(n14071), .ZN(
        n14172) );
  MUX2_X1 U16004 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14172), .S(n14730), .Z(
        n14074) );
  AOI21_X1 U16005 ( .B1(n14075), .B2(n14174), .A(n14074), .ZN(n14076) );
  INV_X1 U16006 ( .A(n14076), .ZN(P1_U3554) );
  AOI21_X1 U16007 ( .B1(n14078), .B2(n14701), .A(n14077), .ZN(n14079) );
  OAI211_X1 U16008 ( .C1(n14639), .C2(n14081), .A(n14080), .B(n14079), .ZN(
        n14177) );
  MUX2_X1 U16009 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14177), .S(n14730), .Z(
        P1_U3553) );
  INV_X1 U16010 ( .A(n14082), .ZN(n14085) );
  AOI211_X1 U16011 ( .C1(n14697), .C2(n14085), .A(n14084), .B(n14083), .ZN(
        n14178) );
  MUX2_X1 U16012 ( .A(n14086), .B(n14178), .S(n14730), .Z(n14087) );
  OAI21_X1 U16013 ( .B1(n14181), .B2(n14155), .A(n14087), .ZN(P1_U3552) );
  INV_X1 U16014 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n14093) );
  NOR2_X1 U16015 ( .A1(n14088), .A2(n14639), .ZN(n14091) );
  NOR4_X1 U16016 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14182) );
  MUX2_X1 U16017 ( .A(n14093), .B(n14182), .S(n14730), .Z(n14094) );
  OAI21_X1 U16018 ( .B1(n7210), .B2(n14155), .A(n14094), .ZN(P1_U3551) );
  OAI211_X1 U16019 ( .C1(n14097), .C2(n14639), .A(n14096), .B(n14095), .ZN(
        n14098) );
  AOI21_X1 U16020 ( .B1(n14699), .B2(n14099), .A(n14098), .ZN(n14185) );
  MUX2_X1 U16021 ( .A(n14100), .B(n14185), .S(n14730), .Z(n14101) );
  OAI21_X1 U16022 ( .B1(n14155), .B2(n14188), .A(n14101), .ZN(P1_U3550) );
  NAND2_X1 U16023 ( .A1(n14103), .A2(n14102), .ZN(n14104) );
  AOI21_X1 U16024 ( .B1(n14105), .B2(n14708), .A(n14104), .ZN(n14106) );
  AND2_X1 U16025 ( .A1(n14107), .A2(n14106), .ZN(n14190) );
  MUX2_X1 U16026 ( .A(n14108), .B(n14190), .S(n14730), .Z(n14109) );
  OAI21_X1 U16027 ( .B1(n14192), .B2(n14155), .A(n14109), .ZN(P1_U3549) );
  INV_X1 U16028 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14114) );
  OAI21_X1 U16029 ( .B1(n14124), .B2(n14704), .A(n14110), .ZN(n14112) );
  AOI211_X1 U16030 ( .C1(n14113), .C2(n14708), .A(n14112), .B(n14111), .ZN(
        n14193) );
  MUX2_X1 U16031 ( .A(n14114), .B(n14193), .S(n14730), .Z(n14115) );
  OAI21_X1 U16032 ( .B1(n14196), .B2(n14155), .A(n14115), .ZN(P1_U3548) );
  OAI21_X1 U16033 ( .B1(n14117), .B2(n14691), .A(n14116), .ZN(n14118) );
  AOI211_X1 U16034 ( .C1(n14120), .C2(n14708), .A(n14119), .B(n14118), .ZN(
        n14121) );
  OAI21_X1 U16035 ( .B1(n14122), .B2(n14629), .A(n14121), .ZN(n14197) );
  MUX2_X1 U16036 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14197), .S(n14730), .Z(
        P1_U3547) );
  INV_X1 U16037 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14131) );
  OAI22_X1 U16038 ( .A1(n14124), .A2(n14615), .B1(n14123), .B2(n14704), .ZN(
        n14125) );
  INV_X1 U16039 ( .A(n14125), .ZN(n14127) );
  OAI211_X1 U16040 ( .C1(n14128), .C2(n14639), .A(n14127), .B(n14126), .ZN(
        n14129) );
  AOI21_X1 U16041 ( .B1(n14130), .B2(n14699), .A(n14129), .ZN(n14198) );
  MUX2_X1 U16042 ( .A(n14131), .B(n14198), .S(n14730), .Z(n14132) );
  OAI21_X1 U16043 ( .B1(n14201), .B2(n14155), .A(n14132), .ZN(P1_U3546) );
  NAND2_X1 U16044 ( .A1(n14133), .A2(n14699), .ZN(n14142) );
  NAND2_X1 U16045 ( .A1(n14134), .A2(n14635), .ZN(n14136) );
  NAND2_X1 U16046 ( .A1(n14447), .A2(n14683), .ZN(n14135) );
  NAND2_X1 U16047 ( .A1(n14136), .A2(n14135), .ZN(n14388) );
  INV_X1 U16048 ( .A(n14388), .ZN(n14137) );
  NAND2_X1 U16049 ( .A1(n14138), .A2(n14137), .ZN(n14139) );
  AOI21_X1 U16050 ( .B1(n14140), .B2(n14708), .A(n14139), .ZN(n14141) );
  AND2_X1 U16051 ( .A1(n14142), .A2(n14141), .ZN(n14203) );
  MUX2_X1 U16052 ( .A(n14143), .B(n14203), .S(n14730), .Z(n14144) );
  OAI21_X1 U16053 ( .B1(n14205), .B2(n14155), .A(n14144), .ZN(P1_U3544) );
  INV_X1 U16054 ( .A(n14145), .ZN(n14424) );
  NAND2_X1 U16055 ( .A1(n14146), .A2(n14699), .ZN(n14153) );
  AOI22_X1 U16056 ( .A1(n14147), .A2(n14683), .B1(n14437), .B2(n14635), .ZN(
        n14148) );
  NAND2_X1 U16057 ( .A1(n14149), .A2(n14148), .ZN(n14150) );
  AOI21_X1 U16058 ( .B1(n14151), .B2(n14708), .A(n14150), .ZN(n14152) );
  AND2_X1 U16059 ( .A1(n14153), .A2(n14152), .ZN(n14207) );
  MUX2_X1 U16060 ( .A(n10725), .B(n14207), .S(n14730), .Z(n14154) );
  OAI21_X1 U16061 ( .B1(n14424), .B2(n14155), .A(n14154), .ZN(P1_U3543) );
  MUX2_X1 U16062 ( .A(n14157), .B(n14156), .S(n14714), .Z(n14158) );
  OAI21_X1 U16063 ( .B1(n14159), .B2(n14209), .A(n14158), .ZN(P1_U3527) );
  INV_X1 U16064 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14161) );
  MUX2_X1 U16065 ( .A(n14161), .B(n14160), .S(n14714), .Z(n14162) );
  OAI21_X1 U16066 ( .B1(n14163), .B2(n14209), .A(n14162), .ZN(P1_U3526) );
  MUX2_X1 U16067 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14164), .S(n14714), .Z(
        P1_U3525) );
  OAI21_X1 U16068 ( .B1(n14168), .B2(n14209), .A(n14167), .ZN(P1_U3524) );
  MUX2_X1 U16069 ( .A(n14170), .B(n14169), .S(n14714), .Z(n14171) );
  INV_X1 U16070 ( .A(n14171), .ZN(P1_U3523) );
  INV_X1 U16071 ( .A(n14209), .ZN(n14175) );
  MUX2_X1 U16072 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14172), .S(n14714), .Z(
        n14173) );
  AOI21_X1 U16073 ( .B1(n14175), .B2(n14174), .A(n14173), .ZN(n14176) );
  INV_X1 U16074 ( .A(n14176), .ZN(P1_U3522) );
  MUX2_X1 U16075 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14177), .S(n14714), .Z(
        P1_U3521) );
  INV_X1 U16076 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14179) );
  MUX2_X1 U16077 ( .A(n14179), .B(n14178), .S(n14714), .Z(n14180) );
  OAI21_X1 U16078 ( .B1(n14181), .B2(n14209), .A(n14180), .ZN(P1_U3520) );
  MUX2_X1 U16079 ( .A(n14183), .B(n14182), .S(n14714), .Z(n14184) );
  OAI21_X1 U16080 ( .B1(n7210), .B2(n14209), .A(n14184), .ZN(P1_U3519) );
  MUX2_X1 U16081 ( .A(n14186), .B(n14185), .S(n14714), .Z(n14187) );
  OAI21_X1 U16082 ( .B1(n14209), .B2(n14188), .A(n14187), .ZN(P1_U3518) );
  MUX2_X1 U16083 ( .A(n14190), .B(n14189), .S(n14713), .Z(n14191) );
  OAI21_X1 U16084 ( .B1(n14192), .B2(n14209), .A(n14191), .ZN(P1_U3517) );
  INV_X1 U16085 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14194) );
  MUX2_X1 U16086 ( .A(n14194), .B(n14193), .S(n14714), .Z(n14195) );
  OAI21_X1 U16087 ( .B1(n14196), .B2(n14209), .A(n14195), .ZN(P1_U3516) );
  MUX2_X1 U16088 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14197), .S(n14714), .Z(
        P1_U3515) );
  INV_X1 U16089 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14199) );
  MUX2_X1 U16090 ( .A(n14199), .B(n14198), .S(n14714), .Z(n14200) );
  OAI21_X1 U16091 ( .B1(n14201), .B2(n14209), .A(n14200), .ZN(P1_U3513) );
  INV_X1 U16092 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14202) );
  MUX2_X1 U16093 ( .A(n14203), .B(n14202), .S(n14713), .Z(n14204) );
  OAI21_X1 U16094 ( .B1(n14205), .B2(n14209), .A(n14204), .ZN(P1_U3507) );
  INV_X1 U16095 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14206) );
  MUX2_X1 U16096 ( .A(n14207), .B(n14206), .S(n14713), .Z(n14208) );
  OAI21_X1 U16097 ( .B1(n14424), .B2(n14209), .A(n14208), .ZN(P1_U3504) );
  NAND3_X1 U16098 ( .A1(n14210), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14212) );
  OAI22_X1 U16099 ( .A1(n14213), .A2(n14212), .B1(n14211), .B2(n14223), .ZN(
        n14214) );
  AOI21_X1 U16100 ( .B1(n14216), .B2(n14215), .A(n14214), .ZN(n14217) );
  INV_X1 U16101 ( .A(n14217), .ZN(P1_U3324) );
  OAI222_X1 U16102 ( .A1(n14223), .A2(n14219), .B1(n14221), .B2(n14218), .C1(
        n9054), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U16103 ( .A1(n14223), .A2(n14222), .B1(n14221), .B2(n14220), .C1(
        P1_U3086), .C2(n14496), .ZN(P1_U3328) );
  MUX2_X1 U16104 ( .A(n14225), .B(n14224), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16105 ( .A(n14226), .ZN(n14227) );
  MUX2_X1 U16106 ( .A(n14227), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NAND2_X1 U16107 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14228), .ZN(n14264) );
  INV_X1 U16108 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14229) );
  AOI22_X1 U16109 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14229), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n14228), .ZN(n14272) );
  INV_X1 U16110 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14230) );
  XOR2_X1 U16111 ( .A(n14261), .B(n14230), .Z(n14274) );
  INV_X1 U16112 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14516) );
  XOR2_X1 U16113 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .Z(n14317) );
  XNOR2_X1 U16114 ( .A(n14251), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n14313) );
  XNOR2_X1 U16115 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14279) );
  XNOR2_X1 U16116 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14283) );
  NAND2_X1 U16117 ( .A1(n14286), .A2(n14285), .ZN(n14231) );
  NAND2_X1 U16118 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14234), .ZN(n14235) );
  NAND2_X1 U16119 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14236), .ZN(n14238) );
  NAND2_X1 U16120 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14239), .ZN(n14241) );
  NAND2_X1 U16121 ( .A1(n14299), .A2(n14300), .ZN(n14240) );
  INV_X1 U16122 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14244) );
  NAND2_X1 U16123 ( .A1(n14245), .A2(n14244), .ZN(n14247) );
  XNOR2_X1 U16124 ( .A(n14245), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U16125 ( .A1(n14307), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U16126 ( .A1(n14247), .A2(n14246), .ZN(n14280) );
  NAND2_X1 U16127 ( .A1(n14279), .A2(n14280), .ZN(n14248) );
  NAND2_X1 U16128 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14277), .ZN(n14253) );
  NOR2_X1 U16129 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14277), .ZN(n14252) );
  XOR2_X1 U16130 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n14255), .Z(n14275) );
  NAND2_X1 U16131 ( .A1(n14276), .A2(n14275), .ZN(n14254) );
  INV_X1 U16132 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14257) );
  NOR2_X1 U16133 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14257), .ZN(n14259) );
  NOR2_X1 U16134 ( .A1(n14274), .A2(n14273), .ZN(n14260) );
  AOI21_X1 U16135 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14261), .A(n14260), 
        .ZN(n14326) );
  NAND2_X1 U16136 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14324), .ZN(n14262) );
  NOR2_X1 U16137 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14324), .ZN(n14323) );
  AOI21_X1 U16138 ( .B1(n14326), .B2(n14262), .A(n14323), .ZN(n14271) );
  NAND2_X1 U16139 ( .A1(n14272), .A2(n14271), .ZN(n14263) );
  NAND2_X1 U16140 ( .A1(n14264), .A2(n14263), .ZN(n14265) );
  NOR2_X1 U16141 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14265), .ZN(n14267) );
  INV_X1 U16142 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14270) );
  XNOR2_X1 U16143 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14265), .ZN(n14269) );
  NOR2_X1 U16144 ( .A1(n14270), .A2(n14269), .ZN(n14266) );
  NOR2_X1 U16145 ( .A1(n14267), .A2(n14266), .ZN(n15189) );
  INV_X1 U16146 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14558) );
  NAND2_X1 U16147 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n14558), .ZN(n15188) );
  OAI21_X1 U16148 ( .B1(n14558), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n15188), 
        .ZN(n14268) );
  XOR2_X1 U16149 ( .A(n15189), .B(n14268), .Z(n15183) );
  XNOR2_X1 U16150 ( .A(n14270), .B(n14269), .ZN(n14329) );
  INV_X1 U16151 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14493) );
  XNOR2_X1 U16152 ( .A(n14272), .B(n14271), .ZN(n14327) );
  INV_X1 U16153 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14483) );
  XOR2_X1 U16154 ( .A(n14274), .B(n14273), .Z(n14481) );
  INV_X1 U16155 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14478) );
  XOR2_X1 U16156 ( .A(n14276), .B(n14275), .Z(n14470) );
  XOR2_X1 U16157 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14277), .Z(n14278) );
  XNOR2_X1 U16158 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14278), .ZN(n14344) );
  XOR2_X1 U16159 ( .A(n14280), .B(n14279), .Z(n14311) );
  NAND2_X1 U16160 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14282), .ZN(n14298) );
  XOR2_X1 U16161 ( .A(n14282), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15382) );
  INV_X1 U16162 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14336) );
  XNOR2_X1 U16163 ( .A(n14284), .B(n14283), .ZN(n14334) );
  XNOR2_X1 U16164 ( .A(n14286), .B(n14285), .ZN(n14288) );
  NAND2_X1 U16165 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14288), .ZN(n14289) );
  AOI21_X1 U16166 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14287), .A(n14286), .ZN(
        n15385) );
  INV_X1 U16167 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15384) );
  NOR2_X1 U16168 ( .A1(n15385), .A2(n15384), .ZN(n15390) );
  NAND2_X1 U16169 ( .A1(n14334), .A2(n14335), .ZN(n14290) );
  XNOR2_X1 U16170 ( .A(n14292), .B(n14291), .ZN(n14293) );
  NAND2_X1 U16171 ( .A1(n14294), .A2(n14293), .ZN(n14296) );
  XOR2_X1 U16172 ( .A(n14294), .B(n14293), .Z(n15388) );
  NAND2_X1 U16173 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15388), .ZN(n14295) );
  NAND2_X1 U16174 ( .A1(n14296), .A2(n14295), .ZN(n15381) );
  NAND2_X1 U16175 ( .A1(n15382), .A2(n15381), .ZN(n14297) );
  XNOR2_X1 U16176 ( .A(n14300), .B(n14299), .ZN(n14301) );
  NAND2_X1 U16177 ( .A1(n14303), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14306) );
  XNOR2_X1 U16178 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14305) );
  XNOR2_X1 U16179 ( .A(n14305), .B(n14304), .ZN(n14338) );
  NAND2_X1 U16180 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14308), .ZN(n14310) );
  XOR2_X1 U16181 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14307), .Z(n15387) );
  NAND2_X1 U16182 ( .A1(n15387), .A2(n15386), .ZN(n14309) );
  XNOR2_X1 U16183 ( .A(n14313), .B(n14312), .ZN(n14314) );
  NAND2_X1 U16184 ( .A1(n6523), .A2(n14314), .ZN(n14315) );
  XOR2_X1 U16185 ( .A(n14317), .B(n14316), .Z(n14319) );
  XOR2_X1 U16186 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .Z(n14320) );
  XNOR2_X1 U16187 ( .A(n14321), .B(n14320), .ZN(n14477) );
  NAND2_X1 U16188 ( .A1(n14476), .A2(n14477), .ZN(n14322) );
  NOR2_X1 U16189 ( .A1(n14476), .A2(n14477), .ZN(n14475) );
  AOI21_X1 U16190 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n14324), .A(n14323), 
        .ZN(n14325) );
  XNOR2_X1 U16191 ( .A(n14326), .B(n14325), .ZN(n14487) );
  NAND2_X1 U16192 ( .A1(n14328), .A2(n14327), .ZN(n14491) );
  INV_X1 U16193 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14350) );
  NAND2_X1 U16194 ( .A1(n14330), .A2(n14329), .ZN(n14349) );
  NAND2_X1 U16195 ( .A1(n14350), .A2(n14349), .ZN(n14346) );
  AOI21_X1 U16196 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14331) );
  OAI21_X1 U16197 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14331), 
        .ZN(U28) );
  AOI21_X1 U16198 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14332) );
  OAI21_X1 U16199 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14332), 
        .ZN(U29) );
  AOI21_X1 U16200 ( .B1(n14335), .B2(n14334), .A(n14333), .ZN(n14337) );
  XNOR2_X1 U16201 ( .A(n14337), .B(n14336), .ZN(SUB_1596_U61) );
  XOR2_X1 U16202 ( .A(n14339), .B(n14338), .Z(SUB_1596_U57) );
  XNOR2_X1 U16203 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14340), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16204 ( .A(n14341), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  OAI21_X1 U16205 ( .B1(n14344), .B2(n14343), .A(n14342), .ZN(n14345) );
  XNOR2_X1 U16206 ( .A(n14345), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI222_X1 U16207 ( .A1(n14350), .A2(n14349), .B1(n14350), .B2(n14348), .C1(
        n14347), .C2(n14346), .ZN(SUB_1596_U63) );
  XOR2_X1 U16208 ( .A(n14352), .B(n14351), .Z(n14364) );
  XNOR2_X1 U16209 ( .A(n14353), .B(n14352), .ZN(n14354) );
  OAI222_X1 U16210 ( .A1(n15072), .A2(n14356), .B1(n15096), .B2(n14355), .C1(
        n14354), .C2(n15075), .ZN(n14362) );
  AOI21_X1 U16211 ( .B1(n14364), .B2(n15034), .A(n14362), .ZN(n14361) );
  NOR2_X1 U16212 ( .A1(n14357), .A2(n15131), .ZN(n14363) );
  AOI22_X1 U16213 ( .A1(n14363), .A2(n15064), .B1(n15102), .B2(n14358), .ZN(
        n14359) );
  OAI221_X1 U16214 ( .B1(n15068), .B2(n14361), .C1(n15107), .C2(n14360), .A(
        n14359), .ZN(P3_U3220) );
  AOI211_X1 U16215 ( .C1(n14364), .C2(n15160), .A(n14363), .B(n14362), .ZN(
        n14371) );
  AOI22_X1 U16216 ( .A1(n15181), .A2(n14371), .B1(n14365), .B2(n6961), .ZN(
        P3_U3472) );
  NOR2_X1 U16217 ( .A1(n14366), .A2(n15131), .ZN(n14368) );
  AOI211_X1 U16218 ( .C1(n15160), .C2(n14369), .A(n14368), .B(n14367), .ZN(
        n14373) );
  AOI22_X1 U16219 ( .A1(n15181), .A2(n14373), .B1(n12244), .B2(n6961), .ZN(
        P3_U3471) );
  INV_X1 U16220 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14370) );
  AOI22_X1 U16221 ( .A1(n15164), .A2(n14371), .B1(n14370), .B2(n15162), .ZN(
        P3_U3429) );
  INV_X1 U16222 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U16223 ( .A1(n15164), .A2(n14373), .B1(n14372), .B2(n15162), .ZN(
        P3_U3426) );
  OAI22_X1 U16224 ( .A1(n14375), .A2(n14427), .B1(n14426), .B2(n14374), .ZN(
        n14381) );
  OAI21_X1 U16225 ( .B1(n6612), .B2(n14377), .A(n14376), .ZN(n14378) );
  AOI21_X1 U16226 ( .B1(n14379), .B2(n14378), .A(n14410), .ZN(n14380) );
  AOI211_X1 U16227 ( .C1(n14445), .C2(n14415), .A(n14381), .B(n14380), .ZN(
        n14383) );
  OAI211_X1 U16228 ( .C1(n14436), .C2(n14384), .A(n14383), .B(n14382), .ZN(
        P1_U3215) );
  XNOR2_X1 U16229 ( .A(n14385), .B(n14386), .ZN(n14389) );
  AOI222_X1 U16230 ( .A1(n14415), .A2(n14390), .B1(n14431), .B2(n14389), .C1(
        n14388), .C2(n14387), .ZN(n14392) );
  OAI211_X1 U16231 ( .C1(n14436), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        P1_U3226) );
  NAND2_X1 U16232 ( .A1(n6629), .A2(n14394), .ZN(n14395) );
  XNOR2_X1 U16233 ( .A(n14396), .B(n14395), .ZN(n14400) );
  NOR2_X1 U16234 ( .A1(n14440), .A2(n14423), .ZN(n14399) );
  OAI22_X1 U16235 ( .A1(n14425), .A2(n14427), .B1(n14426), .B2(n14397), .ZN(
        n14398) );
  AOI211_X1 U16236 ( .C1(n14400), .C2(n14431), .A(n14399), .B(n14398), .ZN(
        n14402) );
  OAI211_X1 U16237 ( .C1(n14436), .C2(n14403), .A(n14402), .B(n14401), .ZN(
        P1_U3228) );
  OAI22_X1 U16238 ( .A1(n14405), .A2(n14426), .B1(n14427), .B2(n14404), .ZN(
        n14414) );
  AOI21_X1 U16239 ( .B1(n14408), .B2(n14407), .A(n14406), .ZN(n14409) );
  INV_X1 U16240 ( .A(n14409), .ZN(n14412) );
  AOI21_X1 U16241 ( .B1(n14412), .B2(n14411), .A(n14410), .ZN(n14413) );
  AOI211_X1 U16242 ( .C1(n14416), .C2(n14415), .A(n14414), .B(n14413), .ZN(
        n14418) );
  OAI211_X1 U16243 ( .C1(n14436), .C2(n14419), .A(n14418), .B(n14417), .ZN(
        P1_U3236) );
  OAI21_X1 U16244 ( .B1(n14422), .B2(n14421), .A(n14420), .ZN(n14432) );
  NOR2_X1 U16245 ( .A1(n14424), .A2(n14423), .ZN(n14430) );
  OAI22_X1 U16246 ( .A1(n14428), .A2(n14427), .B1(n14426), .B2(n14425), .ZN(
        n14429) );
  AOI211_X1 U16247 ( .C1(n14432), .C2(n14431), .A(n14430), .B(n14429), .ZN(
        n14434) );
  NAND2_X1 U16248 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14541)
         );
  OAI211_X1 U16249 ( .C1(n14436), .C2(n14435), .A(n14434), .B(n14541), .ZN(
        P1_U3241) );
  NAND2_X1 U16250 ( .A1(n14437), .A2(n14683), .ZN(n14438) );
  OAI211_X1 U16251 ( .C1(n14440), .C2(n14691), .A(n14439), .B(n14438), .ZN(
        n14442) );
  AOI211_X1 U16252 ( .C1(n14443), .C2(n14708), .A(n14442), .B(n14441), .ZN(
        n14463) );
  AOI22_X1 U16253 ( .A1(n14730), .A2(n14463), .B1(n14444), .B2(n14727), .ZN(
        P1_U3545) );
  INV_X1 U16254 ( .A(n14445), .ZN(n14450) );
  AOI22_X1 U16255 ( .A1(n14635), .A2(n14447), .B1(n14446), .B2(n14683), .ZN(
        n14448) );
  OAI211_X1 U16256 ( .C1(n14450), .C2(n14691), .A(n14449), .B(n14448), .ZN(
        n14453) );
  INV_X1 U16257 ( .A(n14451), .ZN(n14452) );
  AOI211_X1 U16258 ( .C1(n14454), .C2(n14708), .A(n14453), .B(n14452), .ZN(
        n14465) );
  AOI22_X1 U16259 ( .A1(n14730), .A2(n14465), .B1(n14455), .B2(n14727), .ZN(
        P1_U3542) );
  OAI21_X1 U16260 ( .B1(n14457), .B2(n14691), .A(n14456), .ZN(n14459) );
  AOI211_X1 U16261 ( .C1(n14460), .C2(n14708), .A(n14459), .B(n14458), .ZN(
        n14467) );
  AOI22_X1 U16262 ( .A1(n14730), .A2(n14467), .B1(n14461), .B2(n14727), .ZN(
        P1_U3539) );
  INV_X1 U16263 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14462) );
  AOI22_X1 U16264 ( .A1(n14714), .A2(n14463), .B1(n14462), .B2(n14713), .ZN(
        P1_U3510) );
  INV_X1 U16265 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14464) );
  AOI22_X1 U16266 ( .A1(n14714), .A2(n14465), .B1(n14464), .B2(n14713), .ZN(
        P1_U3501) );
  INV_X1 U16267 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U16268 ( .A1(n14714), .A2(n14467), .B1(n14466), .B2(n14713), .ZN(
        P1_U3492) );
  AOI21_X1 U16269 ( .B1(n14470), .B2(n14469), .A(n14468), .ZN(n14471) );
  XOR2_X1 U16270 ( .A(n14471), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  NOR2_X1 U16271 ( .A1(n14473), .A2(n14472), .ZN(n14474) );
  XOR2_X1 U16272 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14474), .Z(SUB_1596_U68)
         );
  AOI21_X1 U16273 ( .B1(n14477), .B2(n14476), .A(n14475), .ZN(n14479) );
  XNOR2_X1 U16274 ( .A(n14479), .B(n14478), .ZN(SUB_1596_U67) );
  AOI21_X1 U16275 ( .B1(n14482), .B2(n14481), .A(n14480), .ZN(n14484) );
  XNOR2_X1 U16276 ( .A(n14484), .B(n14483), .ZN(SUB_1596_U66) );
  OAI21_X1 U16277 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n14488) );
  XNOR2_X1 U16278 ( .A(n14488), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  INV_X1 U16279 ( .A(n14491), .ZN(n14490) );
  OAI222_X1 U16280 ( .A1(n14493), .A2(n14492), .B1(n14493), .B2(n14491), .C1(
        n14490), .C2(n14489), .ZN(SUB_1596_U64) );
  AOI21_X1 U16281 ( .B1(n14496), .B2(n14495), .A(n14494), .ZN(n14497) );
  XNOR2_X1 U16282 ( .A(n14497), .B(P1_IR_REG_0__SCAN_IN), .ZN(n14500) );
  AOI22_X1 U16283 ( .A1(n14517), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14498) );
  OAI21_X1 U16284 ( .B1(n14500), .B2(n14499), .A(n14498), .ZN(P1_U3243) );
  INV_X1 U16285 ( .A(n14501), .ZN(n14506) );
  NAND3_X1 U16286 ( .A1(n14504), .A2(n14503), .A3(n14502), .ZN(n14505) );
  AOI21_X1 U16287 ( .B1(n14506), .B2(n14505), .A(n14538), .ZN(n14513) );
  AOI21_X1 U16288 ( .B1(n14509), .B2(n14508), .A(n14507), .ZN(n14511) );
  OAI22_X1 U16289 ( .A1(n14511), .A2(n14536), .B1(n14510), .B2(n14553), .ZN(
        n14512) );
  NOR2_X1 U16290 ( .A1(n14513), .A2(n14512), .ZN(n14515) );
  OAI211_X1 U16291 ( .C1(n14516), .C2(n14557), .A(n14515), .B(n14514), .ZN(
        P1_U3255) );
  NAND2_X1 U16292 ( .A1(n14517), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14518) );
  OAI211_X1 U16293 ( .C1(n14553), .C2(n14520), .A(n14519), .B(n14518), .ZN(
        n14521) );
  INV_X1 U16294 ( .A(n14521), .ZN(n14530) );
  OAI211_X1 U16295 ( .C1(n14524), .C2(n14523), .A(n14545), .B(n14522), .ZN(
        n14529) );
  OAI211_X1 U16296 ( .C1(n14527), .C2(n14526), .A(n14548), .B(n14525), .ZN(
        n14528) );
  NAND3_X1 U16297 ( .A1(n14530), .A2(n14529), .A3(n14528), .ZN(P1_U3256) );
  INV_X1 U16298 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14543) );
  AOI21_X1 U16299 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14532), .A(n14531), 
        .ZN(n14537) );
  AOI21_X1 U16300 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14534), .A(n14533), 
        .ZN(n14535) );
  OAI222_X1 U16301 ( .A1(n14553), .A2(n14539), .B1(n14538), .B2(n14537), .C1(
        n14536), .C2(n14535), .ZN(n14540) );
  INV_X1 U16302 ( .A(n14540), .ZN(n14542) );
  OAI211_X1 U16303 ( .C1(n14543), .C2(n14557), .A(n14542), .B(n14541), .ZN(
        P1_U3258) );
  OAI211_X1 U16304 ( .C1(n14546), .C2(P1_REG1_REG_18__SCAN_IN), .A(n14545), 
        .B(n14544), .ZN(n14551) );
  OAI211_X1 U16305 ( .C1(n14549), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14548), 
        .B(n14547), .ZN(n14550) );
  OAI211_X1 U16306 ( .C1(n14553), .C2(n14552), .A(n14551), .B(n14550), .ZN(
        n14554) );
  INV_X1 U16307 ( .A(n14554), .ZN(n14556) );
  OAI211_X1 U16308 ( .C1(n14558), .C2(n14557), .A(n14556), .B(n14555), .ZN(
        P1_U3261) );
  OAI21_X1 U16309 ( .B1(n14560), .B2(n14561), .A(n14559), .ZN(n14565) );
  XNOR2_X1 U16310 ( .A(n14562), .B(n14561), .ZN(n14568) );
  NOR2_X1 U16311 ( .A1(n14568), .A2(n14647), .ZN(n14563) );
  AOI211_X1 U16312 ( .C1(n14699), .C2(n14565), .A(n14564), .B(n14563), .ZN(
        n14693) );
  INV_X1 U16313 ( .A(n14566), .ZN(n14567) );
  AOI222_X1 U16314 ( .A1(n14570), .A2(n14601), .B1(P1_REG2_REG_9__SCAN_IN), 
        .B2(n14016), .C1(n14621), .C2(n14567), .ZN(n14575) );
  INV_X1 U16315 ( .A(n14568), .ZN(n14696) );
  INV_X1 U16316 ( .A(n14569), .ZN(n14572) );
  INV_X1 U16317 ( .A(n14570), .ZN(n14692) );
  OAI211_X1 U16318 ( .C1(n14572), .C2(n14692), .A(n14604), .B(n14571), .ZN(
        n14690) );
  INV_X1 U16319 ( .A(n14690), .ZN(n14573) );
  AOI22_X1 U16320 ( .A1(n14696), .A2(n14610), .B1(n14609), .B2(n14573), .ZN(
        n14574) );
  OAI211_X1 U16321 ( .C1(n14016), .C2(n14693), .A(n14575), .B(n14574), .ZN(
        P1_U3284) );
  XNOR2_X1 U16322 ( .A(n14577), .B(n14576), .ZN(n14680) );
  XNOR2_X1 U16323 ( .A(n14579), .B(n14578), .ZN(n14580) );
  NOR2_X1 U16324 ( .A1(n14580), .A2(n14629), .ZN(n14581) );
  AOI211_X1 U16325 ( .C1(n14598), .C2(n14680), .A(n14582), .B(n14581), .ZN(
        n14677) );
  INV_X1 U16326 ( .A(n14583), .ZN(n14584) );
  AOI222_X1 U16327 ( .A1(n14585), .A2(n14601), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n14016), .C1(n14621), .C2(n14584), .ZN(n14591) );
  INV_X1 U16328 ( .A(n14586), .ZN(n14587) );
  OAI211_X1 U16329 ( .C1(n14676), .C2(n14588), .A(n14587), .B(n14604), .ZN(
        n14675) );
  INV_X1 U16330 ( .A(n14675), .ZN(n14589) );
  AOI22_X1 U16331 ( .A1(n14680), .A2(n14610), .B1(n14609), .B2(n14589), .ZN(
        n14590) );
  OAI211_X1 U16332 ( .C1(n14016), .C2(n14677), .A(n14591), .B(n14590), .ZN(
        P1_U3286) );
  XNOR2_X1 U16333 ( .A(n14592), .B(n14593), .ZN(n14659) );
  XNOR2_X1 U16334 ( .A(n14594), .B(n14593), .ZN(n14595) );
  NOR2_X1 U16335 ( .A1(n14595), .A2(n14629), .ZN(n14596) );
  AOI211_X1 U16336 ( .C1(n14598), .C2(n14659), .A(n14597), .B(n14596), .ZN(
        n14656) );
  OAI22_X1 U16337 ( .A1(n6464), .A2(n8804), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n14599), .ZN(n14600) );
  AOI21_X1 U16338 ( .B1(n14601), .B2(n14602), .A(n14600), .ZN(n14612) );
  NAND2_X1 U16339 ( .A1(n14603), .A2(n14602), .ZN(n14605) );
  NAND2_X1 U16340 ( .A1(n14605), .A2(n14604), .ZN(n14607) );
  OR2_X1 U16341 ( .A1(n14607), .A2(n14606), .ZN(n14654) );
  INV_X1 U16342 ( .A(n14654), .ZN(n14608) );
  AOI22_X1 U16343 ( .A1(n14659), .A2(n14610), .B1(n14609), .B2(n14608), .ZN(
        n14611) );
  OAI211_X1 U16344 ( .C1(n14016), .C2(n14656), .A(n14612), .B(n14611), .ZN(
        P1_U3290) );
  AOI21_X1 U16345 ( .B1(n14633), .B2(n14614), .A(n14613), .ZN(n14619) );
  NOR2_X1 U16346 ( .A1(n14616), .A2(n14615), .ZN(n14631) );
  INV_X1 U16347 ( .A(n14631), .ZN(n14617) );
  OAI21_X1 U16348 ( .B1(n14619), .B2(n14618), .A(n14617), .ZN(n14620) );
  AOI22_X1 U16349 ( .A1(n14621), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n6464), .B2(
        n14620), .ZN(n14626) );
  INV_X1 U16350 ( .A(n14628), .ZN(n14622) );
  OAI21_X1 U16351 ( .B1(n14624), .B2(n14623), .A(n14622), .ZN(n14625) );
  OAI211_X1 U16352 ( .C1(n6464), .C2(n9056), .A(n14626), .B(n14625), .ZN(
        P1_U3293) );
  AND2_X1 U16353 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14627), .ZN(P1_U3294) );
  AND2_X1 U16354 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14627), .ZN(P1_U3295) );
  AND2_X1 U16355 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14627), .ZN(P1_U3296) );
  AND2_X1 U16356 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14627), .ZN(P1_U3297) );
  AND2_X1 U16357 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14627), .ZN(P1_U3298) );
  AND2_X1 U16358 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14627), .ZN(P1_U3299) );
  AND2_X1 U16359 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14627), .ZN(P1_U3300) );
  AND2_X1 U16360 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14627), .ZN(P1_U3301) );
  AND2_X1 U16361 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14627), .ZN(P1_U3302) );
  AND2_X1 U16362 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14627), .ZN(P1_U3303) );
  AND2_X1 U16363 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14627), .ZN(P1_U3304) );
  AND2_X1 U16364 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14627), .ZN(P1_U3305) );
  AND2_X1 U16365 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14627), .ZN(P1_U3306) );
  AND2_X1 U16366 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14627), .ZN(P1_U3307) );
  AND2_X1 U16367 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14627), .ZN(P1_U3308) );
  AND2_X1 U16368 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14627), .ZN(P1_U3309) );
  AND2_X1 U16369 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14627), .ZN(P1_U3310) );
  AND2_X1 U16370 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14627), .ZN(P1_U3311) );
  AND2_X1 U16371 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14627), .ZN(P1_U3312) );
  AND2_X1 U16372 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14627), .ZN(P1_U3313) );
  AND2_X1 U16373 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14627), .ZN(P1_U3314) );
  AND2_X1 U16374 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14627), .ZN(P1_U3315) );
  AND2_X1 U16375 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14627), .ZN(P1_U3316) );
  AND2_X1 U16376 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14627), .ZN(P1_U3317) );
  AND2_X1 U16377 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14627), .ZN(P1_U3318) );
  AND2_X1 U16378 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14627), .ZN(P1_U3319) );
  AND2_X1 U16379 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14627), .ZN(P1_U3320) );
  AND2_X1 U16380 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14627), .ZN(P1_U3321) );
  AND2_X1 U16381 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14627), .ZN(P1_U3322) );
  AND2_X1 U16382 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14627), .ZN(P1_U3323) );
  AOI21_X1 U16383 ( .B1(n14639), .B2(n14629), .A(n14628), .ZN(n14630) );
  AOI211_X1 U16384 ( .C1(n14633), .C2(n14632), .A(n14631), .B(n14630), .ZN(
        n14715) );
  INV_X1 U16385 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U16386 ( .A1(n14714), .A2(n14715), .B1(n14634), .B2(n14713), .ZN(
        P1_U3459) );
  AOI22_X1 U16387 ( .A1(n14636), .A2(n14635), .B1(n6668), .B2(n14701), .ZN(
        n14638) );
  OAI211_X1 U16388 ( .C1(n14640), .C2(n14639), .A(n14638), .B(n14637), .ZN(
        n14643) );
  INV_X1 U16389 ( .A(n14641), .ZN(n14642) );
  NOR2_X1 U16390 ( .A1(n14643), .A2(n14642), .ZN(n14716) );
  INV_X1 U16391 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14644) );
  AOI22_X1 U16392 ( .A1(n14714), .A2(n14716), .B1(n14644), .B2(n14713), .ZN(
        P1_U3462) );
  AOI21_X1 U16393 ( .B1(n14647), .B2(n14646), .A(n14645), .ZN(n14652) );
  OAI21_X1 U16394 ( .B1(n14649), .B2(n14691), .A(n14648), .ZN(n14650) );
  NOR3_X1 U16395 ( .A1(n14652), .A2(n14651), .A3(n14650), .ZN(n14717) );
  INV_X1 U16396 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14653) );
  AOI22_X1 U16397 ( .A1(n14714), .A2(n14717), .B1(n14653), .B2(n14713), .ZN(
        P1_U3465) );
  OAI21_X1 U16398 ( .B1(n14655), .B2(n14691), .A(n14654), .ZN(n14658) );
  INV_X1 U16399 ( .A(n14656), .ZN(n14657) );
  AOI211_X1 U16400 ( .C1(n14697), .C2(n14659), .A(n14658), .B(n14657), .ZN(
        n14718) );
  INV_X1 U16401 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14660) );
  AOI22_X1 U16402 ( .A1(n14714), .A2(n14718), .B1(n14660), .B2(n14713), .ZN(
        P1_U3468) );
  NAND2_X1 U16403 ( .A1(n14661), .A2(n14708), .ZN(n14666) );
  NAND2_X1 U16404 ( .A1(n14662), .A2(n14701), .ZN(n14663) );
  NAND4_X1 U16405 ( .A1(n14666), .A2(n14665), .A3(n14664), .A4(n14663), .ZN(
        n14667) );
  AOI21_X1 U16406 ( .B1(n14699), .B2(n14668), .A(n14667), .ZN(n14720) );
  INV_X1 U16407 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14669) );
  AOI22_X1 U16408 ( .A1(n14714), .A2(n14720), .B1(n14669), .B2(n14713), .ZN(
        P1_U3471) );
  OAI21_X1 U16409 ( .B1(n14671), .B2(n14691), .A(n14670), .ZN(n14673) );
  AOI211_X1 U16410 ( .C1(n14697), .C2(n14674), .A(n14673), .B(n14672), .ZN(
        n14722) );
  AOI22_X1 U16411 ( .A1(n14714), .A2(n14722), .B1(n9608), .B2(n14713), .ZN(
        P1_U3474) );
  OAI21_X1 U16412 ( .B1(n14676), .B2(n14691), .A(n14675), .ZN(n14679) );
  INV_X1 U16413 ( .A(n14677), .ZN(n14678) );
  AOI211_X1 U16414 ( .C1(n14697), .C2(n14680), .A(n14679), .B(n14678), .ZN(
        n14723) );
  INV_X1 U16415 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U16416 ( .A1(n14714), .A2(n14723), .B1(n14681), .B2(n14713), .ZN(
        P1_U3480) );
  AOI22_X1 U16417 ( .A1(n14684), .A2(n14701), .B1(n14683), .B2(n14682), .ZN(
        n14685) );
  NAND2_X1 U16418 ( .A1(n14686), .A2(n14685), .ZN(n14688) );
  AOI211_X1 U16419 ( .C1(n14689), .C2(n14708), .A(n14688), .B(n14687), .ZN(
        n14724) );
  AOI22_X1 U16420 ( .A1(n14714), .A2(n14724), .B1(n9980), .B2(n14713), .ZN(
        P1_U3483) );
  OAI21_X1 U16421 ( .B1(n14692), .B2(n14691), .A(n14690), .ZN(n14695) );
  INV_X1 U16422 ( .A(n14693), .ZN(n14694) );
  AOI211_X1 U16423 ( .C1(n14697), .C2(n14696), .A(n14695), .B(n14694), .ZN(
        n14726) );
  INV_X1 U16424 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14698) );
  AOI22_X1 U16425 ( .A1(n14714), .A2(n14726), .B1(n14698), .B2(n14713), .ZN(
        P1_U3486) );
  NAND2_X1 U16426 ( .A1(n14700), .A2(n14699), .ZN(n14712) );
  NAND2_X1 U16427 ( .A1(n14702), .A2(n14701), .ZN(n14703) );
  OAI21_X1 U16428 ( .B1(n14705), .B2(n14704), .A(n14703), .ZN(n14706) );
  NOR2_X1 U16429 ( .A1(n14707), .A2(n14706), .ZN(n14711) );
  NAND2_X1 U16430 ( .A1(n14709), .A2(n14708), .ZN(n14710) );
  AOI22_X1 U16431 ( .A1(n14714), .A2(n14729), .B1(n10339), .B2(n14713), .ZN(
        P1_U3489) );
  AOI22_X1 U16432 ( .A1(n14730), .A2(n14715), .B1(n14495), .B2(n14727), .ZN(
        P1_U3528) );
  AOI22_X1 U16433 ( .A1(n14730), .A2(n14716), .B1(n9074), .B2(n14727), .ZN(
        P1_U3529) );
  AOI22_X1 U16434 ( .A1(n14730), .A2(n14717), .B1(n9128), .B2(n14727), .ZN(
        P1_U3530) );
  AOI22_X1 U16435 ( .A1(n14730), .A2(n14718), .B1(n9297), .B2(n14727), .ZN(
        P1_U3531) );
  AOI22_X1 U16436 ( .A1(n14730), .A2(n14720), .B1(n14719), .B2(n14727), .ZN(
        P1_U3532) );
  AOI22_X1 U16437 ( .A1(n14730), .A2(n14722), .B1(n14721), .B2(n14727), .ZN(
        P1_U3533) );
  AOI22_X1 U16438 ( .A1(n14730), .A2(n14723), .B1(n9849), .B2(n14727), .ZN(
        P1_U3535) );
  AOI22_X1 U16439 ( .A1(n14730), .A2(n14724), .B1(n9984), .B2(n14727), .ZN(
        P1_U3536) );
  AOI22_X1 U16440 ( .A1(n14730), .A2(n14726), .B1(n14725), .B2(n14727), .ZN(
        P1_U3537) );
  AOI22_X1 U16441 ( .A1(n14730), .A2(n14729), .B1(n14728), .B2(n14727), .ZN(
        P1_U3538) );
  NOR2_X1 U16442 ( .A1(n14784), .A2(P2_U3947), .ZN(P2_U3087) );
  INV_X1 U16443 ( .A(n14731), .ZN(n14732) );
  AOI21_X1 U16444 ( .B1(n14785), .B2(P2_REG1_REG_0__SCAN_IN), .A(n14732), .ZN(
        n14737) );
  AOI22_X1 U16445 ( .A1(n14784), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14736) );
  OAI22_X1 U16446 ( .A1(n14733), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14742), .ZN(n14734) );
  OAI21_X1 U16447 ( .B1(n14790), .B2(n14734), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14735) );
  OAI211_X1 U16448 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14737), .A(n14736), .B(
        n14735), .ZN(P2_U3214) );
  AOI22_X1 U16449 ( .A1(n14784), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14750) );
  OAI211_X1 U16450 ( .C1(n14740), .C2(n14739), .A(n14738), .B(n14791), .ZN(
        n14749) );
  AOI211_X1 U16451 ( .C1(n14744), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        n14745) );
  INV_X1 U16452 ( .A(n14745), .ZN(n14748) );
  NAND2_X1 U16453 ( .A1(n14790), .A2(n14746), .ZN(n14747) );
  NAND4_X1 U16454 ( .A1(n14750), .A2(n14749), .A3(n14748), .A4(n14747), .ZN(
        P2_U3227) );
  INV_X1 U16455 ( .A(n14751), .ZN(n14753) );
  OAI21_X1 U16456 ( .B1(n14753), .B2(n14752), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14754) );
  OAI21_X1 U16457 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14754), .ZN(n14763) );
  OAI211_X1 U16458 ( .C1(n14756), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14755), 
        .B(n14791), .ZN(n14762) );
  NAND2_X1 U16459 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n14784), .ZN(n14761) );
  XOR2_X1 U16460 ( .A(n14758), .B(n14757), .Z(n14759) );
  NAND2_X1 U16461 ( .A1(n14759), .A2(n14785), .ZN(n14760) );
  NAND4_X1 U16462 ( .A1(n14763), .A2(n14762), .A3(n14761), .A4(n14760), .ZN(
        P2_U3228) );
  AOI22_X1 U16463 ( .A1(n14784), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14772) );
  NAND2_X1 U16464 ( .A1(n14790), .A2(n14764), .ZN(n14771) );
  OAI211_X1 U16465 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14766), .A(n14791), 
        .B(n14765), .ZN(n14770) );
  OAI211_X1 U16466 ( .C1(n14768), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14785), 
        .B(n14767), .ZN(n14769) );
  NAND4_X1 U16467 ( .A1(n14772), .A2(n14771), .A3(n14770), .A4(n14769), .ZN(
        P2_U3229) );
  AOI22_X1 U16468 ( .A1(n14784), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n14783) );
  NAND2_X1 U16469 ( .A1(n14790), .A2(n14773), .ZN(n14782) );
  OAI211_X1 U16470 ( .C1(n14776), .C2(n14775), .A(n14774), .B(n14791), .ZN(
        n14781) );
  XNOR2_X1 U16471 ( .A(n14778), .B(n14777), .ZN(n14779) );
  NAND2_X1 U16472 ( .A1(n14779), .A2(n14785), .ZN(n14780) );
  NAND4_X1 U16473 ( .A1(n14783), .A2(n14782), .A3(n14781), .A4(n14780), .ZN(
        P2_U3230) );
  AOI22_X1 U16474 ( .A1(n14784), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14798) );
  OAI211_X1 U16475 ( .C1(n14788), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n14797) );
  NAND2_X1 U16476 ( .A1(n14790), .A2(n14789), .ZN(n14796) );
  OAI211_X1 U16477 ( .C1(n14794), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        n14795) );
  NAND4_X1 U16478 ( .A1(n14798), .A2(n14797), .A3(n14796), .A4(n14795), .ZN(
        P2_U3231) );
  INV_X1 U16479 ( .A(n14799), .ZN(n14800) );
  AND2_X1 U16480 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14801), .ZN(P2_U3266) );
  AND2_X1 U16481 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14801), .ZN(P2_U3267) );
  AND2_X1 U16482 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14801), .ZN(P2_U3268) );
  AND2_X1 U16483 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14801), .ZN(P2_U3269) );
  AND2_X1 U16484 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14801), .ZN(P2_U3270) );
  AND2_X1 U16485 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14801), .ZN(P2_U3271) );
  AND2_X1 U16486 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14801), .ZN(P2_U3272) );
  AND2_X1 U16487 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14801), .ZN(P2_U3273) );
  AND2_X1 U16488 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14801), .ZN(P2_U3274) );
  AND2_X1 U16489 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14801), .ZN(P2_U3275) );
  AND2_X1 U16490 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14801), .ZN(P2_U3276) );
  AND2_X1 U16491 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14801), .ZN(P2_U3277) );
  AND2_X1 U16492 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14801), .ZN(P2_U3278) );
  AND2_X1 U16493 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14801), .ZN(P2_U3279) );
  AND2_X1 U16494 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14801), .ZN(P2_U3280) );
  AND2_X1 U16495 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14801), .ZN(P2_U3281) );
  AND2_X1 U16496 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14801), .ZN(P2_U3282) );
  AND2_X1 U16497 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14801), .ZN(P2_U3283) );
  AND2_X1 U16498 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14801), .ZN(P2_U3284) );
  AND2_X1 U16499 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14801), .ZN(P2_U3285) );
  AND2_X1 U16500 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14801), .ZN(P2_U3286) );
  AND2_X1 U16501 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14801), .ZN(P2_U3287) );
  AND2_X1 U16502 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14801), .ZN(P2_U3288) );
  AND2_X1 U16503 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14801), .ZN(P2_U3289) );
  AND2_X1 U16504 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14801), .ZN(P2_U3290) );
  AND2_X1 U16505 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14801), .ZN(P2_U3291) );
  AND2_X1 U16506 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14801), .ZN(P2_U3292) );
  AND2_X1 U16507 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14801), .ZN(P2_U3293) );
  AND2_X1 U16508 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14801), .ZN(P2_U3294) );
  AND2_X1 U16509 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14801), .ZN(P2_U3295) );
  AOI22_X1 U16510 ( .A1(n14805), .A2(n14802), .B1(n8882), .B2(n14803), .ZN(
        P2_U3416) );
  AOI22_X1 U16511 ( .A1(n14805), .A2(n14804), .B1(n8885), .B2(n14803), .ZN(
        P2_U3417) );
  INV_X1 U16512 ( .A(n14806), .ZN(n14810) );
  INV_X1 U16513 ( .A(n14807), .ZN(n14808) );
  AOI211_X1 U16514 ( .C1(n14875), .C2(n14810), .A(n14809), .B(n14808), .ZN(
        n14888) );
  INV_X1 U16515 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14811) );
  AOI22_X1 U16516 ( .A1(n14887), .A2(n14888), .B1(n14811), .B2(n14886), .ZN(
        P2_U3430) );
  INV_X1 U16517 ( .A(n14812), .ZN(n14818) );
  INV_X1 U16518 ( .A(n14819), .ZN(n14816) );
  AOI21_X1 U16519 ( .B1(n14879), .B2(n14814), .A(n14813), .ZN(n14815) );
  OAI21_X1 U16520 ( .B1(n14816), .B2(n14871), .A(n14815), .ZN(n14817) );
  AOI211_X1 U16521 ( .C1(n14875), .C2(n14819), .A(n14818), .B(n14817), .ZN(
        n14890) );
  INV_X1 U16522 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14820) );
  AOI22_X1 U16523 ( .A1(n14887), .A2(n14890), .B1(n14820), .B2(n14886), .ZN(
        P2_U3433) );
  OAI21_X1 U16524 ( .B1(n14822), .B2(n14867), .A(n14821), .ZN(n14823) );
  AOI21_X1 U16525 ( .B1(n14824), .B2(n14875), .A(n14823), .ZN(n14825) );
  AND2_X1 U16526 ( .A1(n14826), .A2(n14825), .ZN(n14892) );
  AOI22_X1 U16527 ( .A1(n14887), .A2(n14892), .B1(n8957), .B2(n14886), .ZN(
        P2_U3436) );
  INV_X1 U16528 ( .A(n14827), .ZN(n14828) );
  OAI21_X1 U16529 ( .B1(n14829), .B2(n14867), .A(n14828), .ZN(n14831) );
  AOI211_X1 U16530 ( .C1(n14875), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        n14894) );
  INV_X1 U16531 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14833) );
  AOI22_X1 U16532 ( .A1(n14887), .A2(n14894), .B1(n14833), .B2(n14886), .ZN(
        P2_U3442) );
  OAI211_X1 U16533 ( .C1(n14836), .C2(n14867), .A(n14835), .B(n14834), .ZN(
        n14837) );
  AOI21_X1 U16534 ( .B1(n14850), .B2(n14838), .A(n14837), .ZN(n14895) );
  AOI22_X1 U16535 ( .A1(n14887), .A2(n14895), .B1(n9338), .B2(n14886), .ZN(
        P2_U3445) );
  AOI21_X1 U16536 ( .B1(n14871), .B2(n14881), .A(n14839), .ZN(n14844) );
  OAI21_X1 U16537 ( .B1(n14841), .B2(n14867), .A(n14840), .ZN(n14842) );
  NOR3_X1 U16538 ( .A1(n14844), .A2(n14843), .A3(n14842), .ZN(n14897) );
  AOI22_X1 U16539 ( .A1(n14887), .A2(n14897), .B1(n9548), .B2(n14886), .ZN(
        P2_U3448) );
  INV_X1 U16540 ( .A(n14845), .ZN(n14851) );
  OAI21_X1 U16541 ( .B1(n14847), .B2(n14867), .A(n14846), .ZN(n14849) );
  AOI211_X1 U16542 ( .C1(n14851), .C2(n14850), .A(n14849), .B(n14848), .ZN(
        n14898) );
  AOI22_X1 U16543 ( .A1(n14887), .A2(n14898), .B1(n9533), .B2(n14886), .ZN(
        P2_U3451) );
  OAI21_X1 U16544 ( .B1(n14853), .B2(n14867), .A(n14852), .ZN(n14857) );
  OAI21_X1 U16545 ( .B1(n14871), .B2(n14855), .A(n14854), .ZN(n14856) );
  AOI211_X1 U16546 ( .C1(n14875), .C2(n14858), .A(n14857), .B(n14856), .ZN(
        n14900) );
  AOI22_X1 U16547 ( .A1(n14887), .A2(n14900), .B1(n9649), .B2(n14886), .ZN(
        P2_U3454) );
  INV_X1 U16548 ( .A(n14862), .ZN(n14865) );
  AOI21_X1 U16549 ( .B1(n14879), .B2(n14860), .A(n14859), .ZN(n14861) );
  OAI21_X1 U16550 ( .B1(n14862), .B2(n14881), .A(n14861), .ZN(n14864) );
  AOI211_X1 U16551 ( .C1(n14885), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        n14902) );
  AOI22_X1 U16552 ( .A1(n14887), .A2(n14902), .B1(n9661), .B2(n14886), .ZN(
        P2_U3457) );
  OAI21_X1 U16553 ( .B1(n14868), .B2(n14867), .A(n14866), .ZN(n14873) );
  OAI21_X1 U16554 ( .B1(n14871), .B2(n14870), .A(n14869), .ZN(n14872) );
  AOI211_X1 U16555 ( .C1(n14875), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14904) );
  AOI22_X1 U16556 ( .A1(n14887), .A2(n14904), .B1(n9669), .B2(n14886), .ZN(
        P2_U3460) );
  INV_X1 U16557 ( .A(n14882), .ZN(n14884) );
  AOI211_X1 U16558 ( .C1(n14879), .C2(n14878), .A(n14877), .B(n14876), .ZN(
        n14880) );
  OAI21_X1 U16559 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14883) );
  AOI21_X1 U16560 ( .B1(n14885), .B2(n14884), .A(n14883), .ZN(n14907) );
  AOI22_X1 U16561 ( .A1(n14887), .A2(n14907), .B1(n10181), .B2(n14886), .ZN(
        P2_U3463) );
  AOI22_X1 U16562 ( .A1(n14908), .A2(n14888), .B1(n8623), .B2(n14905), .ZN(
        P2_U3499) );
  AOI22_X1 U16563 ( .A1(n14908), .A2(n14890), .B1(n14889), .B2(n14905), .ZN(
        P2_U3500) );
  AOI22_X1 U16564 ( .A1(n14908), .A2(n14892), .B1(n14891), .B2(n14905), .ZN(
        P2_U3501) );
  AOI22_X1 U16565 ( .A1(n14908), .A2(n14894), .B1(n14893), .B2(n14905), .ZN(
        P2_U3503) );
  AOI22_X1 U16566 ( .A1(n14908), .A2(n14895), .B1(n9333), .B2(n14905), .ZN(
        P2_U3504) );
  AOI22_X1 U16567 ( .A1(n14908), .A2(n14897), .B1(n14896), .B2(n14905), .ZN(
        P2_U3505) );
  AOI22_X1 U16568 ( .A1(n14908), .A2(n14898), .B1(n9531), .B2(n14905), .ZN(
        P2_U3506) );
  AOI22_X1 U16569 ( .A1(n14908), .A2(n14900), .B1(n14899), .B2(n14905), .ZN(
        P2_U3507) );
  AOI22_X1 U16570 ( .A1(n14908), .A2(n14902), .B1(n14901), .B2(n14905), .ZN(
        P2_U3508) );
  AOI22_X1 U16571 ( .A1(n14908), .A2(n14904), .B1(n14903), .B2(n14905), .ZN(
        P2_U3509) );
  AOI22_X1 U16572 ( .A1(n14908), .A2(n14907), .B1(n14906), .B2(n14905), .ZN(
        P2_U3510) );
  NOR2_X1 U16573 ( .A1(P3_U3897), .A2(n14996), .ZN(P3_U3150) );
  AOI22_X1 U16574 ( .A1(n15005), .A2(n14910), .B1(n14997), .B2(n14909), .ZN(
        n14919) );
  AOI22_X1 U16575 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n14996), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n14918) );
  NAND3_X1 U16576 ( .A1(n14990), .A2(n14977), .A3(n14911), .ZN(n14913) );
  NAND3_X1 U16577 ( .A1(n15007), .A2(n14915), .A3(n14914), .ZN(n14916) );
  NAND4_X1 U16578 ( .A1(n14919), .A2(n14918), .A3(n14917), .A4(n14916), .ZN(
        P3_U3182) );
  AOI21_X1 U16579 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(n14996), .A(n14920), .ZN(
        n14934) );
  OAI21_X1 U16580 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14925) );
  AOI22_X1 U16581 ( .A1(n14925), .A2(n15007), .B1(n14924), .B2(n14983), .ZN(
        n14933) );
  XNOR2_X1 U16582 ( .A(n14926), .B(n15169), .ZN(n14927) );
  NAND2_X1 U16583 ( .A1(n15005), .A2(n14927), .ZN(n14932) );
  OAI221_X1 U16584 ( .B1(n14930), .B2(n14929), .C1(n14930), .C2(n14928), .A(
        n14997), .ZN(n14931) );
  NAND4_X1 U16585 ( .A1(n14934), .A2(n14933), .A3(n14932), .A4(n14931), .ZN(
        P3_U3185) );
  AOI21_X1 U16586 ( .B1(P3_ADDR_REG_5__SCAN_IN), .B2(n14996), .A(n14935), .ZN(
        n14950) );
  OAI21_X1 U16587 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n14939) );
  AOI22_X1 U16588 ( .A1(n14983), .A2(n14940), .B1(n14939), .B2(n15007), .ZN(
        n14949) );
  OAI221_X1 U16589 ( .B1(n14943), .B2(n14942), .C1(n14943), .C2(n14941), .A(
        n14997), .ZN(n14948) );
  AOI21_X1 U16590 ( .B1(n14945), .B2(n15172), .A(n14944), .ZN(n14946) );
  OR2_X1 U16591 ( .A1(n14977), .A2(n14946), .ZN(n14947) );
  NAND4_X1 U16592 ( .A1(n14950), .A2(n14949), .A3(n14948), .A4(n14947), .ZN(
        P3_U3187) );
  AOI21_X1 U16593 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(n14996), .A(n14951), .ZN(
        n14966) );
  OAI21_X1 U16594 ( .B1(n14954), .B2(n14953), .A(n14952), .ZN(n14955) );
  AOI22_X1 U16595 ( .A1(n14983), .A2(n14956), .B1(n14955), .B2(n15007), .ZN(
        n14965) );
  AOI21_X1 U16596 ( .B1(n14958), .B2(n15175), .A(n14957), .ZN(n14959) );
  OR2_X1 U16597 ( .A1(n14959), .A2(n14977), .ZN(n14964) );
  OAI221_X1 U16598 ( .B1(n14962), .B2(n14961), .C1(n14962), .C2(n14960), .A(
        n14997), .ZN(n14963) );
  NAND4_X1 U16599 ( .A1(n14966), .A2(n14965), .A3(n14964), .A4(n14963), .ZN(
        P3_U3189) );
  INV_X1 U16600 ( .A(n14967), .ZN(n14968) );
  AOI21_X1 U16601 ( .B1(n14970), .B2(n14969), .A(n14968), .ZN(n14991) );
  INV_X1 U16602 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14973) );
  INV_X1 U16603 ( .A(n14971), .ZN(n14972) );
  OAI21_X1 U16604 ( .B1(n14974), .B2(n14973), .A(n14972), .ZN(n14981) );
  NAND2_X1 U16605 ( .A1(n14976), .A2(n14975), .ZN(n14978) );
  AOI21_X1 U16606 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n14980) );
  AOI211_X1 U16607 ( .C1(n14983), .C2(n14982), .A(n14981), .B(n14980), .ZN(
        n14989) );
  NOR2_X1 U16608 ( .A1(n14985), .A2(n14984), .ZN(n14986) );
  OAI21_X1 U16609 ( .B1(n14987), .B2(n14986), .A(n15007), .ZN(n14988) );
  OAI211_X1 U16610 ( .C1(n14991), .C2(n14990), .A(n14989), .B(n14988), .ZN(
        P3_U3192) );
  NOR2_X1 U16611 ( .A1(n14993), .A2(n14992), .ZN(n14994) );
  AOI211_X1 U16612 ( .C1(n14996), .C2(P3_ADDR_REG_12__SCAN_IN), .A(n14995), 
        .B(n14994), .ZN(n15014) );
  OAI221_X1 U16613 ( .B1(n15000), .B2(n14999), .C1(n15000), .C2(n14998), .A(
        n14997), .ZN(n15013) );
  INV_X1 U16614 ( .A(n15001), .ZN(n15004) );
  OAI21_X1 U16615 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15006) );
  NAND2_X1 U16616 ( .A1(n15006), .A2(n15005), .ZN(n15012) );
  OAI211_X1 U16617 ( .C1(n15010), .C2(n15009), .A(n15008), .B(n15007), .ZN(
        n15011) );
  NAND4_X1 U16618 ( .A1(n15014), .A2(n15013), .A3(n15012), .A4(n15011), .ZN(
        P3_U3194) );
  XNOR2_X1 U16619 ( .A(n15016), .B(n15015), .ZN(n15161) );
  OR2_X1 U16620 ( .A1(n15037), .A2(n15017), .ZN(n15020) );
  AND2_X1 U16621 ( .A1(n15020), .A2(n15018), .ZN(n15023) );
  NAND2_X1 U16622 ( .A1(n15020), .A2(n15019), .ZN(n15021) );
  OAI211_X1 U16623 ( .C1(n15023), .C2(n15022), .A(n15021), .B(n15099), .ZN(
        n15027) );
  AOI22_X1 U16624 ( .A1(n15025), .A2(n15045), .B1(n15093), .B2(n15024), .ZN(
        n15026) );
  NAND2_X1 U16625 ( .A1(n15027), .A2(n15026), .ZN(n15158) );
  AOI21_X1 U16626 ( .B1(n15161), .B2(n15080), .A(n15158), .ZN(n15033) );
  AOI22_X1 U16627 ( .A1(n15068), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15102), 
        .B2(n15028), .ZN(n15032) );
  NOR2_X1 U16628 ( .A1(n15029), .A2(n15131), .ZN(n15159) );
  AOI22_X1 U16629 ( .A1(n15161), .A2(n15030), .B1(n15064), .B2(n15159), .ZN(
        n15031) );
  OAI211_X1 U16630 ( .C1(n15068), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        P3_U3223) );
  INV_X1 U16631 ( .A(n15034), .ZN(n15105) );
  XNOR2_X1 U16632 ( .A(n15035), .B(n15042), .ZN(n15155) );
  OR2_X1 U16633 ( .A1(n15037), .A2(n15036), .ZN(n15040) );
  AND2_X1 U16634 ( .A1(n15040), .A2(n15038), .ZN(n15043) );
  NAND2_X1 U16635 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  OAI211_X1 U16636 ( .C1(n15043), .C2(n15042), .A(n15041), .B(n15099), .ZN(
        n15047) );
  AOI22_X1 U16637 ( .A1(n8302), .A2(n15045), .B1(n15093), .B2(n15044), .ZN(
        n15046) );
  AND2_X1 U16638 ( .A1(n15047), .A2(n15046), .ZN(n15154) );
  OAI21_X1 U16639 ( .B1(n15105), .B2(n15155), .A(n15154), .ZN(n15051) );
  OAI22_X1 U16640 ( .A1(n15049), .A2(n15048), .B1(n10228), .B2(n15107), .ZN(
        n15050) );
  AOI21_X1 U16641 ( .B1(n15051), .B2(n15107), .A(n15050), .ZN(n15052) );
  OAI21_X1 U16642 ( .B1(n15054), .B2(n15053), .A(n15052), .ZN(P3_U3224) );
  AOI21_X1 U16643 ( .B1(n6632), .B2(n15061), .A(n15075), .ZN(n15059) );
  OAI22_X1 U16644 ( .A1(n15056), .A2(n15096), .B1(n15055), .B2(n15072), .ZN(
        n15057) );
  AOI21_X1 U16645 ( .B1(n15059), .B2(n15058), .A(n15057), .ZN(n15137) );
  AOI22_X1 U16646 ( .A1(n15068), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n15102), 
        .B2(n15060), .ZN(n15067) );
  XNOR2_X1 U16647 ( .A(n15062), .B(n15061), .ZN(n15140) );
  NOR2_X1 U16648 ( .A1(n15063), .A2(n15131), .ZN(n15139) );
  AOI22_X1 U16649 ( .A1(n15140), .A2(n15065), .B1(n15064), .B2(n15139), .ZN(
        n15066) );
  OAI211_X1 U16650 ( .C1(n15068), .C2(n15137), .A(n15067), .B(n15066), .ZN(
        P3_U3227) );
  OAI21_X1 U16651 ( .B1(n15070), .B2(n15074), .A(n15069), .ZN(n15118) );
  OAI22_X1 U16652 ( .A1(n7018), .A2(n15072), .B1(n15071), .B2(n15096), .ZN(
        n15079) );
  NAND3_X1 U16653 ( .A1(n15092), .A2(n15074), .A3(n15073), .ZN(n15076) );
  AOI21_X1 U16654 ( .B1(n15077), .B2(n15076), .A(n15075), .ZN(n15078) );
  AOI211_X1 U16655 ( .C1(n15080), .C2(n15118), .A(n15079), .B(n15078), .ZN(
        n15081) );
  INV_X1 U16656 ( .A(n15081), .ZN(n15116) );
  NOR2_X1 U16657 ( .A1(n15082), .A2(n15131), .ZN(n15117) );
  AOI22_X1 U16658 ( .A1(n15118), .A2(n15083), .B1(n15117), .B2(n15103), .ZN(
        n15084) );
  INV_X1 U16659 ( .A(n15084), .ZN(n15085) );
  AOI211_X1 U16660 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15102), .A(n15116), .B(
        n15085), .ZN(n15086) );
  AOI22_X1 U16661 ( .A1(n15068), .A2(n15087), .B1(n15086), .B2(n15107), .ZN(
        P3_U3231) );
  XNOR2_X1 U16662 ( .A(n15090), .B(n15088), .ZN(n15110) );
  OR2_X1 U16663 ( .A1(n15090), .A2(n15089), .ZN(n15091) );
  NAND2_X1 U16664 ( .A1(n15092), .A2(n15091), .ZN(n15100) );
  NAND2_X1 U16665 ( .A1(n15094), .A2(n15093), .ZN(n15095) );
  OAI21_X1 U16666 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n15098) );
  AOI21_X1 U16667 ( .B1(n15100), .B2(n15099), .A(n15098), .ZN(n15114) );
  AND2_X1 U16668 ( .A1(n15101), .A2(n15151), .ZN(n15111) );
  AOI22_X1 U16669 ( .A1(n15111), .A2(n15103), .B1(n15102), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n15104) );
  OAI211_X1 U16670 ( .C1(n15105), .C2(n15110), .A(n15114), .B(n15104), .ZN(
        n15106) );
  INV_X1 U16671 ( .A(n15106), .ZN(n15108) );
  AOI22_X1 U16672 ( .A1(n15068), .A2(n15109), .B1(n15108), .B2(n15107), .ZN(
        P3_U3232) );
  OR2_X1 U16673 ( .A1(n15110), .A2(n15156), .ZN(n15113) );
  INV_X1 U16674 ( .A(n15111), .ZN(n15112) );
  AND3_X1 U16675 ( .A1(n15114), .A2(n15113), .A3(n15112), .ZN(n15166) );
  INV_X1 U16676 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15115) );
  AOI22_X1 U16677 ( .A1(n15164), .A2(n15166), .B1(n15115), .B2(n15162), .ZN(
        P3_U3393) );
  AOI211_X1 U16678 ( .C1(n15148), .C2(n15118), .A(n15117), .B(n15116), .ZN(
        n15168) );
  INV_X1 U16679 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15119) );
  AOI22_X1 U16680 ( .A1(n15164), .A2(n15168), .B1(n15119), .B2(n15162), .ZN(
        P3_U3396) );
  NOR2_X1 U16681 ( .A1(n15120), .A2(n15131), .ZN(n15122) );
  AOI211_X1 U16682 ( .C1(n15148), .C2(n15123), .A(n15122), .B(n15121), .ZN(
        n15170) );
  INV_X1 U16683 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15124) );
  AOI22_X1 U16684 ( .A1(n15164), .A2(n15170), .B1(n15124), .B2(n15162), .ZN(
        P3_U3399) );
  INV_X1 U16685 ( .A(n15125), .ZN(n15129) );
  INV_X1 U16686 ( .A(n15126), .ZN(n15127) );
  AOI211_X1 U16687 ( .C1(n15129), .C2(n15148), .A(n15128), .B(n15127), .ZN(
        n15171) );
  INV_X1 U16688 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15130) );
  AOI22_X1 U16689 ( .A1(n15164), .A2(n15171), .B1(n15130), .B2(n15162), .ZN(
        P3_U3402) );
  NOR2_X1 U16690 ( .A1(n15132), .A2(n15131), .ZN(n15134) );
  AOI211_X1 U16691 ( .C1(n15148), .C2(n15135), .A(n15134), .B(n15133), .ZN(
        n15173) );
  INV_X1 U16692 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15136) );
  AOI22_X1 U16693 ( .A1(n15164), .A2(n15173), .B1(n15136), .B2(n15162), .ZN(
        P3_U3405) );
  INV_X1 U16694 ( .A(n15137), .ZN(n15138) );
  AOI211_X1 U16695 ( .C1(n15140), .C2(n15160), .A(n15139), .B(n15138), .ZN(
        n15174) );
  INV_X1 U16696 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15141) );
  AOI22_X1 U16697 ( .A1(n15164), .A2(n15174), .B1(n15141), .B2(n15162), .ZN(
        P3_U3408) );
  AOI211_X1 U16698 ( .C1(n15148), .C2(n15144), .A(n15143), .B(n15142), .ZN(
        n15176) );
  INV_X1 U16699 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15145) );
  AOI22_X1 U16700 ( .A1(n15164), .A2(n15176), .B1(n15145), .B2(n15162), .ZN(
        P3_U3411) );
  AOI211_X1 U16701 ( .C1(n15149), .C2(n15148), .A(n15147), .B(n15146), .ZN(
        n15177) );
  INV_X1 U16702 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15150) );
  AOI22_X1 U16703 ( .A1(n15164), .A2(n15177), .B1(n15150), .B2(n15162), .ZN(
        P3_U3414) );
  NAND2_X1 U16704 ( .A1(n15152), .A2(n15151), .ZN(n15153) );
  OAI211_X1 U16705 ( .C1(n15156), .C2(n15155), .A(n15154), .B(n15153), .ZN(
        n15178) );
  OAI22_X1 U16706 ( .A1(n15162), .A2(n15178), .B1(P3_REG0_REG_9__SCAN_IN), 
        .B2(n15164), .ZN(n15157) );
  INV_X1 U16707 ( .A(n15157), .ZN(P3_U3417) );
  AOI211_X1 U16708 ( .C1(n15161), .C2(n15160), .A(n15159), .B(n15158), .ZN(
        n15180) );
  INV_X1 U16709 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15163) );
  AOI22_X1 U16710 ( .A1(n15164), .A2(n15180), .B1(n15163), .B2(n15162), .ZN(
        P3_U3420) );
  INV_X1 U16711 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15165) );
  AOI22_X1 U16712 ( .A1(n15181), .A2(n15166), .B1(n15165), .B2(n6961), .ZN(
        P3_U3460) );
  AOI22_X1 U16713 ( .A1(n15181), .A2(n15168), .B1(n15167), .B2(n6961), .ZN(
        P3_U3461) );
  AOI22_X1 U16714 ( .A1(n15181), .A2(n15170), .B1(n15169), .B2(n6961), .ZN(
        P3_U3462) );
  AOI22_X1 U16715 ( .A1(n15181), .A2(n15171), .B1(n9161), .B2(n6961), .ZN(
        P3_U3463) );
  AOI22_X1 U16716 ( .A1(n15181), .A2(n15173), .B1(n15172), .B2(n6961), .ZN(
        P3_U3464) );
  AOI22_X1 U16717 ( .A1(n15181), .A2(n15174), .B1(n9501), .B2(n6961), .ZN(
        P3_U3465) );
  AOI22_X1 U16718 ( .A1(n15181), .A2(n15176), .B1(n15175), .B2(n6961), .ZN(
        P3_U3466) );
  AOI22_X1 U16719 ( .A1(n15181), .A2(n15177), .B1(n9884), .B2(n6961), .ZN(
        P3_U3467) );
  OAI22_X1 U16720 ( .A1(n6961), .A2(n15178), .B1(P3_REG1_REG_9__SCAN_IN), .B2(
        n15181), .ZN(n15179) );
  INV_X1 U16721 ( .A(n15179), .ZN(P3_U3468) );
  AOI22_X1 U16722 ( .A1(n15181), .A2(n15180), .B1(n10573), .B2(n6961), .ZN(
        P3_U3469) );
  XNOR2_X1 U16723 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15185) );
  XNOR2_X1 U16724 ( .A(n15185), .B(n15184), .ZN(n15186) );
  AOI22_X1 U16725 ( .A1(n15189), .A2(n15188), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n15187), .ZN(n15380) );
  AOI22_X1 U16726 ( .A1(SI_9_), .A2(keyinput_f23), .B1(SI_16_), .B2(
        keyinput_f16), .ZN(n15190) );
  OAI221_X1 U16727 ( .B1(SI_9_), .B2(keyinput_f23), .C1(SI_16_), .C2(
        keyinput_f16), .A(n15190), .ZN(n15197) );
  AOI22_X1 U16728 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n15191) );
  OAI221_X1 U16729 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n15191), .ZN(n15196)
         );
  AOI22_X1 U16730 ( .A1(SI_24_), .A2(keyinput_f8), .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n15192) );
  OAI221_X1 U16731 ( .B1(SI_24_), .B2(keyinput_f8), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n15192), .ZN(n15195)
         );
  AOI22_X1 U16732 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n15193) );
  OAI221_X1 U16733 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_f56), .A(n15193), .ZN(n15194)
         );
  NOR4_X1 U16734 ( .A1(n15197), .A2(n15196), .A3(n15195), .A4(n15194), .ZN(
        n15226) );
  XNOR2_X1 U16735 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_f42), .ZN(n15205)
         );
  AOI22_X1 U16736 ( .A1(SI_14_), .A2(keyinput_f18), .B1(n15199), .B2(
        keyinput_f41), .ZN(n15198) );
  OAI221_X1 U16737 ( .B1(SI_14_), .B2(keyinput_f18), .C1(n15199), .C2(
        keyinput_f41), .A(n15198), .ZN(n15204) );
  AOI22_X1 U16738 ( .A1(SI_23_), .A2(keyinput_f9), .B1(SI_10_), .B2(
        keyinput_f22), .ZN(n15200) );
  OAI221_X1 U16739 ( .B1(SI_23_), .B2(keyinput_f9), .C1(SI_10_), .C2(
        keyinput_f22), .A(n15200), .ZN(n15203) );
  AOI22_X1 U16740 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n15201) );
  OAI221_X1 U16741 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n15201), .ZN(n15202)
         );
  NOR4_X1 U16742 ( .A1(n15205), .A2(n15204), .A3(n15203), .A4(n15202), .ZN(
        n15225) );
  AOI22_X1 U16743 ( .A1(SI_26_), .A2(keyinput_f6), .B1(SI_13_), .B2(
        keyinput_f19), .ZN(n15206) );
  OAI221_X1 U16744 ( .B1(SI_26_), .B2(keyinput_f6), .C1(SI_13_), .C2(
        keyinput_f19), .A(n15206), .ZN(n15214) );
  AOI22_X1 U16745 ( .A1(SI_5_), .A2(keyinput_f27), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n15207) );
  OAI221_X1 U16746 ( .B1(SI_5_), .B2(keyinput_f27), .C1(P3_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n15207), .ZN(n15213) );
  AOI22_X1 U16747 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_f57), .B1(
        n15209), .B2(keyinput_f47), .ZN(n15208) );
  OAI221_X1 U16748 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .C1(
        n15209), .C2(keyinput_f47), .A(n15208), .ZN(n15212) );
  AOI22_X1 U16749 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(keyinput_f44), .ZN(n15210) );
  OAI221_X1 U16750 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P3_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n15210), .ZN(n15211) );
  NOR4_X1 U16751 ( .A1(n15214), .A2(n15213), .A3(n15212), .A4(n15211), .ZN(
        n15224) );
  AOI22_X1 U16752 ( .A1(SI_4_), .A2(keyinput_f28), .B1(SI_15_), .B2(
        keyinput_f17), .ZN(n15215) );
  OAI221_X1 U16753 ( .B1(SI_4_), .B2(keyinput_f28), .C1(SI_15_), .C2(
        keyinput_f17), .A(n15215), .ZN(n15222) );
  AOI22_X1 U16754 ( .A1(keyinput_f0), .A2(P3_WR_REG_SCAN_IN), .B1(keyinput_f33), .B2(P3_RD_REG_SCAN_IN), .ZN(n15216) );
  OAI221_X1 U16755 ( .B1(keyinput_f0), .B2(P3_WR_REG_SCAN_IN), .C1(
        keyinput_f33), .C2(P3_RD_REG_SCAN_IN), .A(n15216), .ZN(n15221) );
  AOI22_X1 U16756 ( .A1(SI_8_), .A2(keyinput_f24), .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n15217) );
  OAI221_X1 U16757 ( .B1(SI_8_), .B2(keyinput_f24), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n15217), .ZN(n15220)
         );
  AOI22_X1 U16758 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n15218) );
  OAI221_X1 U16759 ( .B1(SI_25_), .B2(keyinput_f7), .C1(
        P3_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n15218), .ZN(n15219)
         );
  NOR4_X1 U16760 ( .A1(n15222), .A2(n15221), .A3(n15220), .A4(n15219), .ZN(
        n15223) );
  NAND4_X1 U16761 ( .A1(n15226), .A2(n15225), .A3(n15224), .A4(n15223), .ZN(
        n15281) );
  AOI22_X1 U16762 ( .A1(n15228), .A2(keyinput_f10), .B1(n15347), .B2(
        keyinput_f5), .ZN(n15227) );
  OAI221_X1 U16763 ( .B1(n15228), .B2(keyinput_f10), .C1(n15347), .C2(
        keyinput_f5), .A(n15227), .ZN(n15239) );
  AOI22_X1 U16764 ( .A1(n15230), .A2(keyinput_f52), .B1(n15348), .B2(
        keyinput_f43), .ZN(n15229) );
  OAI221_X1 U16765 ( .B1(n15230), .B2(keyinput_f52), .C1(n15348), .C2(
        keyinput_f43), .A(n15229), .ZN(n15238) );
  AOI22_X1 U16766 ( .A1(n15232), .A2(keyinput_f20), .B1(n15363), .B2(
        keyinput_f39), .ZN(n15231) );
  OAI221_X1 U16767 ( .B1(n15232), .B2(keyinput_f20), .C1(n15363), .C2(
        keyinput_f39), .A(n15231), .ZN(n15237) );
  INV_X1 U16768 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15235) );
  INV_X1 U16769 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U16770 ( .A1(n15235), .A2(keyinput_f55), .B1(keyinput_f54), .B2(
        n15234), .ZN(n15233) );
  OAI221_X1 U16771 ( .B1(n15235), .B2(keyinput_f55), .C1(n15234), .C2(
        keyinput_f54), .A(n15233), .ZN(n15236) );
  NOR4_X1 U16772 ( .A1(n15239), .A2(n15238), .A3(n15237), .A4(n15236), .ZN(
        n15279) );
  INV_X1 U16773 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15241) );
  AOI22_X1 U16774 ( .A1(n15345), .A2(keyinput_f58), .B1(n15241), .B2(
        keyinput_f60), .ZN(n15240) );
  OAI221_X1 U16775 ( .B1(n15345), .B2(keyinput_f58), .C1(n15241), .C2(
        keyinput_f60), .A(n15240), .ZN(n15251) );
  AOI22_X1 U16776 ( .A1(n15244), .A2(keyinput_f37), .B1(keyinput_f4), .B2(
        n15243), .ZN(n15242) );
  OAI221_X1 U16777 ( .B1(n15244), .B2(keyinput_f37), .C1(n15243), .C2(
        keyinput_f4), .A(n15242), .ZN(n15250) );
  XNOR2_X1 U16778 ( .A(SI_0_), .B(keyinput_f32), .ZN(n15248) );
  XNOR2_X1 U16779 ( .A(P3_REG3_REG_21__SCAN_IN), .B(keyinput_f45), .ZN(n15247)
         );
  XNOR2_X1 U16780 ( .A(SI_1_), .B(keyinput_f31), .ZN(n15246) );
  XNOR2_X1 U16781 ( .A(SI_3_), .B(keyinput_f29), .ZN(n15245) );
  NAND4_X1 U16782 ( .A1(n15248), .A2(n15247), .A3(n15246), .A4(n15245), .ZN(
        n15249) );
  NOR3_X1 U16783 ( .A1(n15251), .A2(n15250), .A3(n15249), .ZN(n15278) );
  AOI22_X1 U16784 ( .A1(P3_U3151), .A2(keyinput_f34), .B1(keyinput_f59), .B2(
        n15253), .ZN(n15252) );
  OAI221_X1 U16785 ( .B1(P3_U3151), .B2(keyinput_f34), .C1(n15253), .C2(
        keyinput_f59), .A(n15252), .ZN(n15264) );
  AOI22_X1 U16786 ( .A1(n15255), .A2(keyinput_f50), .B1(keyinput_f3), .B2(
        n15364), .ZN(n15254) );
  OAI221_X1 U16787 ( .B1(n15255), .B2(keyinput_f50), .C1(n15364), .C2(
        keyinput_f3), .A(n15254), .ZN(n15263) );
  AOI22_X1 U16788 ( .A1(n15258), .A2(keyinput_f30), .B1(n15257), .B2(
        keyinput_f15), .ZN(n15256) );
  OAI221_X1 U16789 ( .B1(n15258), .B2(keyinput_f30), .C1(n15257), .C2(
        keyinput_f15), .A(n15256), .ZN(n15262) );
  XNOR2_X1 U16790 ( .A(SI_7_), .B(keyinput_f25), .ZN(n15260) );
  XNOR2_X1 U16791 ( .A(SI_21_), .B(keyinput_f11), .ZN(n15259) );
  NAND2_X1 U16792 ( .A1(n15260), .A2(n15259), .ZN(n15261) );
  NOR4_X1 U16793 ( .A1(n15264), .A2(n15263), .A3(n15262), .A4(n15261), .ZN(
        n15277) );
  AOI22_X1 U16794 ( .A1(n15344), .A2(keyinput_f14), .B1(n7852), .B2(
        keyinput_f49), .ZN(n15265) );
  OAI221_X1 U16795 ( .B1(n15344), .B2(keyinput_f14), .C1(n7852), .C2(
        keyinput_f49), .A(n15265), .ZN(n15275) );
  AOI22_X1 U16796 ( .A1(n7912), .A2(keyinput_f53), .B1(keyinput_f13), .B2(
        n15267), .ZN(n15266) );
  OAI221_X1 U16797 ( .B1(n7912), .B2(keyinput_f53), .C1(n15267), .C2(
        keyinput_f13), .A(n15266), .ZN(n15274) );
  INV_X1 U16798 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15269) );
  AOI22_X1 U16799 ( .A1(n15325), .A2(keyinput_f12), .B1(n15269), .B2(
        keyinput_f48), .ZN(n15268) );
  OAI221_X1 U16800 ( .B1(n15325), .B2(keyinput_f12), .C1(n15269), .C2(
        keyinput_f48), .A(n15268), .ZN(n15273) );
  XOR2_X1 U16801 ( .A(n15338), .B(keyinput_f35), .Z(n15271) );
  XNOR2_X1 U16802 ( .A(SI_6_), .B(keyinput_f26), .ZN(n15270) );
  NAND2_X1 U16803 ( .A1(n15271), .A2(n15270), .ZN(n15272) );
  NOR4_X1 U16804 ( .A1(n15275), .A2(n15274), .A3(n15273), .A4(n15272), .ZN(
        n15276) );
  NAND4_X1 U16805 ( .A1(n15279), .A2(n15278), .A3(n15277), .A4(n15276), .ZN(
        n15280) );
  OAI22_X1 U16806 ( .A1(n15281), .A2(n15280), .B1(keyinput_f21), .B2(SI_11_), 
        .ZN(n15282) );
  AOI21_X1 U16807 ( .B1(keyinput_f21), .B2(SI_11_), .A(n15282), .ZN(n15378) );
  AOI22_X1 U16808 ( .A1(SI_7_), .A2(keyinput_g25), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n15283) );
  OAI221_X1 U16809 ( .B1(SI_7_), .B2(keyinput_g25), .C1(SI_22_), .C2(
        keyinput_g10), .A(n15283), .ZN(n15290) );
  AOI22_X1 U16810 ( .A1(SI_30_), .A2(keyinput_g2), .B1(SI_17_), .B2(
        keyinput_g15), .ZN(n15284) );
  OAI221_X1 U16811 ( .B1(SI_30_), .B2(keyinput_g2), .C1(SI_17_), .C2(
        keyinput_g15), .A(n15284), .ZN(n15289) );
  AOI22_X1 U16812 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n15285) );
  OAI221_X1 U16813 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_g51), .A(n15285), .ZN(n15288)
         );
  AOI22_X1 U16814 ( .A1(SI_10_), .A2(keyinput_g22), .B1(SI_1_), .B2(
        keyinput_g31), .ZN(n15286) );
  OAI221_X1 U16815 ( .B1(SI_10_), .B2(keyinput_g22), .C1(SI_1_), .C2(
        keyinput_g31), .A(n15286), .ZN(n15287) );
  NOR4_X1 U16816 ( .A1(n15290), .A2(n15289), .A3(n15288), .A4(n15287), .ZN(
        n15317) );
  XOR2_X1 U16817 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_g52), .Z(n15297) );
  AOI22_X1 U16818 ( .A1(SI_12_), .A2(keyinput_g20), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n15291) );
  OAI221_X1 U16819 ( .B1(SI_12_), .B2(keyinput_g20), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n15291), .ZN(n15296)
         );
  AOI22_X1 U16820 ( .A1(SI_25_), .A2(keyinput_g7), .B1(P3_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n15292) );
  OAI221_X1 U16821 ( .B1(SI_25_), .B2(keyinput_g7), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n15292), .ZN(n15295)
         );
  AOI22_X1 U16822 ( .A1(SI_23_), .A2(keyinput_g9), .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .ZN(n15293) );
  OAI221_X1 U16823 ( .B1(SI_23_), .B2(keyinput_g9), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n15293), .ZN(n15294)
         );
  NOR4_X1 U16824 ( .A1(n15297), .A2(n15296), .A3(n15295), .A4(n15294), .ZN(
        n15316) );
  AOI22_X1 U16825 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(SI_13_), .B2(keyinput_g19), .ZN(n15298) );
  OAI221_X1 U16826 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        SI_13_), .C2(keyinput_g19), .A(n15298), .ZN(n15305) );
  AOI22_X1 U16827 ( .A1(SI_3_), .A2(keyinput_g29), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_g53), .ZN(n15299) );
  OAI221_X1 U16828 ( .B1(SI_3_), .B2(keyinput_g29), .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_g53), .A(n15299), .ZN(n15304) );
  AOI22_X1 U16829 ( .A1(SI_19_), .A2(keyinput_g13), .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n15300) );
  OAI221_X1 U16830 ( .B1(SI_19_), .B2(keyinput_g13), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n15300), .ZN(n15303) );
  AOI22_X1 U16831 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n15301) );
  OAI221_X1 U16832 ( .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n15301), .ZN(n15302)
         );
  NOR4_X1 U16833 ( .A1(n15305), .A2(n15304), .A3(n15303), .A4(n15302), .ZN(
        n15315) );
  AOI22_X1 U16834 ( .A1(SI_28_), .A2(keyinput_g4), .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n15306) );
  OAI221_X1 U16835 ( .B1(SI_28_), .B2(keyinput_g4), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n15306), .ZN(n15313)
         );
  AOI22_X1 U16836 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n15307) );
  OAI221_X1 U16837 ( .B1(P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n15307), .ZN(n15312)
         );
  AOI22_X1 U16838 ( .A1(SI_6_), .A2(keyinput_g26), .B1(SI_24_), .B2(
        keyinput_g8), .ZN(n15308) );
  OAI221_X1 U16839 ( .B1(SI_6_), .B2(keyinput_g26), .C1(SI_24_), .C2(
        keyinput_g8), .A(n15308), .ZN(n15311) );
  AOI22_X1 U16840 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P3_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .ZN(n15309) );
  OAI221_X1 U16841 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_g38), .A(n15309), .ZN(n15310)
         );
  NOR4_X1 U16842 ( .A1(n15313), .A2(n15312), .A3(n15311), .A4(n15310), .ZN(
        n15314) );
  NAND4_X1 U16843 ( .A1(n15317), .A2(n15316), .A3(n15315), .A4(n15314), .ZN(
        n15376) );
  INV_X1 U16844 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15319) );
  AOI22_X1 U16845 ( .A1(n15320), .A2(keyinput_g63), .B1(keyinput_g0), .B2(
        n15319), .ZN(n15318) );
  OAI221_X1 U16846 ( .B1(n15320), .B2(keyinput_g63), .C1(n15319), .C2(
        keyinput_g0), .A(n15318), .ZN(n15331) );
  AOI22_X1 U16847 ( .A1(n7689), .A2(keyinput_g56), .B1(keyinput_g18), .B2(
        n15322), .ZN(n15321) );
  OAI221_X1 U16848 ( .B1(n7689), .B2(keyinput_g56), .C1(n15322), .C2(
        keyinput_g18), .A(n15321), .ZN(n15330) );
  AOI22_X1 U16849 ( .A1(n15325), .A2(keyinput_g12), .B1(n15324), .B2(
        keyinput_g36), .ZN(n15323) );
  OAI221_X1 U16850 ( .B1(n15325), .B2(keyinput_g12), .C1(n15324), .C2(
        keyinput_g36), .A(n15323), .ZN(n15329) );
  XNOR2_X1 U16851 ( .A(SI_4_), .B(keyinput_g28), .ZN(n15327) );
  XNOR2_X1 U16852 ( .A(SI_15_), .B(keyinput_g17), .ZN(n15326) );
  NAND2_X1 U16853 ( .A1(n15327), .A2(n15326), .ZN(n15328) );
  NOR4_X1 U16854 ( .A1(n15331), .A2(n15330), .A3(n15329), .A4(n15328), .ZN(
        n15374) );
  AOI22_X1 U16855 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(
        P3_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n15332) );
  OAI221_X1 U16856 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        P3_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n15332), .ZN(n15342) );
  AOI22_X1 U16857 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n15333) );
  OAI221_X1 U16858 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n15333), .ZN(n15341)
         );
  AOI22_X1 U16859 ( .A1(n15336), .A2(keyinput_g16), .B1(keyinput_g23), .B2(
        n15335), .ZN(n15334) );
  OAI221_X1 U16860 ( .B1(n15336), .B2(keyinput_g16), .C1(n15335), .C2(
        keyinput_g23), .A(n15334), .ZN(n15340) );
  AOI22_X1 U16861 ( .A1(P3_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(n15338), 
        .B2(keyinput_g35), .ZN(n15337) );
  OAI221_X1 U16862 ( .B1(P3_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(n15338), 
        .C2(keyinput_g35), .A(n15337), .ZN(n15339) );
  NOR4_X1 U16863 ( .A1(n15342), .A2(n15341), .A3(n15340), .A4(n15339), .ZN(
        n15373) );
  AOI22_X1 U16864 ( .A1(n15345), .A2(keyinput_g58), .B1(keyinput_g14), .B2(
        n15344), .ZN(n15343) );
  OAI221_X1 U16865 ( .B1(n15345), .B2(keyinput_g58), .C1(n15344), .C2(
        keyinput_g14), .A(n15343), .ZN(n15355) );
  AOI22_X1 U16866 ( .A1(n15348), .A2(keyinput_g43), .B1(keyinput_g5), .B2(
        n15347), .ZN(n15346) );
  OAI221_X1 U16867 ( .B1(n15348), .B2(keyinput_g43), .C1(n15347), .C2(
        keyinput_g5), .A(n15346), .ZN(n15354) );
  XNOR2_X1 U16868 ( .A(SI_0_), .B(keyinput_g32), .ZN(n15352) );
  XNOR2_X1 U16869 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_g46), .ZN(n15351)
         );
  XNOR2_X1 U16870 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_g44), .ZN(n15350)
         );
  XNOR2_X1 U16871 ( .A(SI_5_), .B(keyinput_g27), .ZN(n15349) );
  NAND4_X1 U16872 ( .A1(n15352), .A2(n15351), .A3(n15350), .A4(n15349), .ZN(
        n15353) );
  NOR3_X1 U16873 ( .A1(n15355), .A2(n15354), .A3(n15353), .ZN(n15372) );
  INV_X1 U16874 ( .A(SI_31_), .ZN(n15357) );
  AOI22_X1 U16875 ( .A1(n15358), .A2(keyinput_g6), .B1(keyinput_g1), .B2(
        n15357), .ZN(n15356) );
  OAI221_X1 U16876 ( .B1(n15358), .B2(keyinput_g6), .C1(n15357), .C2(
        keyinput_g1), .A(n15356), .ZN(n15370) );
  AOI22_X1 U16877 ( .A1(n15361), .A2(keyinput_g11), .B1(n15360), .B2(
        keyinput_g40), .ZN(n15359) );
  OAI221_X1 U16878 ( .B1(n15361), .B2(keyinput_g11), .C1(n15360), .C2(
        keyinput_g40), .A(n15359), .ZN(n15369) );
  AOI22_X1 U16879 ( .A1(n15364), .A2(keyinput_g3), .B1(n15363), .B2(
        keyinput_g39), .ZN(n15362) );
  OAI221_X1 U16880 ( .B1(n15364), .B2(keyinput_g3), .C1(n15363), .C2(
        keyinput_g39), .A(n15362), .ZN(n15368) );
  XNOR2_X1 U16881 ( .A(SI_2_), .B(keyinput_g30), .ZN(n15366) );
  XNOR2_X1 U16882 ( .A(SI_8_), .B(keyinput_g24), .ZN(n15365) );
  NAND2_X1 U16883 ( .A1(n15366), .A2(n15365), .ZN(n15367) );
  NOR4_X1 U16884 ( .A1(n15370), .A2(n15369), .A3(n15368), .A4(n15367), .ZN(
        n15371) );
  NAND4_X1 U16885 ( .A1(n15374), .A2(n15373), .A3(n15372), .A4(n15371), .ZN(
        n15375) );
  OAI22_X1 U16886 ( .A1(SI_11_), .A2(keyinput_g21), .B1(n15376), .B2(n15375), 
        .ZN(n15377) );
  AOI211_X1 U16887 ( .C1(SI_11_), .C2(keyinput_g21), .A(n15378), .B(n15377), 
        .ZN(n15379) );
  XOR2_X1 U16888 ( .A(n15382), .B(n15381), .Z(SUB_1596_U59) );
  XNOR2_X1 U16889 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15383), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16890 ( .B1(n15385), .B2(n15384), .A(n15390), .ZN(SUB_1596_U53) );
  XOR2_X1 U16891 ( .A(n15387), .B(n15386), .Z(SUB_1596_U56) );
  XOR2_X1 U16892 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15388), .Z(SUB_1596_U60) );
  XOR2_X1 U16893 ( .A(n15390), .B(n15389), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7217 ( .A(n11051), .Z(n6477) );
  CLKBUF_X1 U7258 ( .A(n11100), .Z(n7010) );
  CLKBUF_X1 U7881 ( .A(n8948), .Z(n11959) );
endmodule

