

module b17_C_SARLock_k_64_9 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820;

  XNOR2_X1 U11023 ( .A(n10730), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14273) );
  INV_X1 U11024 ( .A(n14873), .ZN(n14840) );
  AOI21_X1 U11025 ( .B1(n14609), .B2(n15710), .A(n11529), .ZN(n15708) );
  NAND3_X1 U11026 ( .A1(n13699), .A2(n13700), .A3(n11680), .ZN(n13769) );
  INV_X2 U11027 ( .A(n13108), .ZN(n18810) );
  CLKBUF_X2 U11029 ( .A(n10739), .Z(n10844) );
  INV_X1 U11030 ( .A(n19232), .ZN(n19230) );
  OR2_X1 U11031 ( .A1(n10226), .A2(n10225), .ZN(n10449) );
  OR2_X1 U11032 ( .A1(n10207), .A2(n14217), .ZN(n10384) );
  OR2_X1 U11033 ( .A1(n10207), .A2(n13533), .ZN(n10380) );
  CLKBUF_X2 U11034 ( .A(n12251), .Z(n16917) );
  INV_X2 U11036 ( .A(n15453), .ZN(n16915) );
  CLKBUF_X2 U11038 ( .A(n11277), .Z(n12072) );
  CLKBUF_X2 U11039 ( .A(n11989), .Z(n11369) );
  CLKBUF_X2 U11040 ( .A(n11292), .Z(n12044) );
  CLKBUF_X1 U11041 ( .A(n11251), .Z(n14796) );
  AND2_X1 U11042 ( .A1(n12941), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10249) );
  AND2_X1 U11043 ( .A1(n9591), .A2(n10023), .ZN(n12748) );
  AND2_X1 U11044 ( .A1(n10033), .A2(n10023), .ZN(n12749) );
  AND2_X1 U11045 ( .A1(n12940), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10250) );
  CLKBUF_X1 U11046 ( .A(n10302), .Z(n12697) );
  INV_X1 U11047 ( .A(n10179), .ZN(n10739) );
  INV_X1 U11048 ( .A(n19979), .ZN(n11253) );
  CLKBUF_X1 U11049 ( .A(n11249), .Z(n19994) );
  CLKBUF_X2 U11050 ( .A(n12154), .Z(n9586) );
  CLKBUF_X2 U11051 ( .A(n12154), .Z(n9585) );
  INV_X1 U11052 ( .A(n16840), .ZN(n15473) );
  BUF_X1 U11053 ( .A(n12207), .Z(n16922) );
  BUF_X2 U11054 ( .A(n12149), .Z(n16916) );
  CLKBUF_X1 U11055 ( .A(n12251), .Z(n16942) );
  CLKBUF_X1 U11056 ( .A(n12250), .Z(n16683) );
  CLKBUF_X1 U11057 ( .A(n12149), .Z(n16943) );
  INV_X4 U11058 ( .A(n12127), .ZN(n9594) );
  CLKBUF_X3 U11059 ( .A(n12142), .Z(n9602) );
  NAND4_X2 U11060 ( .A1(n11239), .A2(n11238), .A3(n11237), .A4(n11236), .ZN(
        n19979) );
  CLKBUF_X2 U11061 ( .A(n11326), .Z(n11275) );
  NAND2_X1 U11062 ( .A1(n9633), .A2(n9627), .ZN(n10127) );
  OR2_X1 U11063 ( .A1(n10136), .A2(n9598), .ZN(n10143) );
  AND2_X1 U11065 ( .A1(n13669), .A2(n13418), .ZN(n11292) );
  CLKBUF_X1 U11066 ( .A(n10144), .Z(n13785) );
  AND2_X2 U11067 ( .A1(n11111), .A2(n13418), .ZN(n11363) );
  NAND2_X1 U11068 ( .A1(n10078), .A2(n10077), .ZN(n11055) );
  INV_X2 U11070 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16054) );
  OR2_X1 U11071 ( .A1(n10835), .A2(n10128), .ZN(n10129) );
  BUF_X2 U11072 ( .A(n10025), .Z(n10102) );
  AND2_X2 U11073 ( .A1(n10624), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9592) );
  AND2_X1 U11074 ( .A1(n10421), .A2(n10420), .ZN(n10469) );
  INV_X1 U11075 ( .A(n11180), .ZN(n11242) );
  INV_X1 U11076 ( .A(n19983), .ZN(n9599) );
  NAND2_X1 U11077 ( .A1(n10519), .A2(n9996), .ZN(n10531) );
  INV_X1 U11078 ( .A(n10339), .ZN(n9930) );
  AND2_X1 U11079 ( .A1(n12940), .A2(n10023), .ZN(n10917) );
  NAND2_X1 U11081 ( .A1(n11055), .A2(n9598), .ZN(n10644) );
  AND2_X1 U11082 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10624) );
  NAND2_X1 U11083 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18580), .ZN(
        n12119) );
  NOR2_X1 U11084 ( .A1(n19983), .A2(n19987), .ZN(n11258) );
  AOI21_X1 U11085 ( .B1(n14251), .B2(n14698), .A(n13064), .ZN(n14533) );
  AND4_X1 U11086 ( .A1(n11147), .A2(n11146), .A3(n11145), .A4(n11144), .ZN(
        n11158) );
  INV_X2 U11087 ( .A(n10155), .ZN(n10848) );
  AND2_X1 U11088 ( .A1(n10270), .A2(n10269), .ZN(n9867) );
  INV_X1 U11089 ( .A(n10449), .ZN(n14044) );
  OR2_X1 U11090 ( .A1(n10223), .A2(n10225), .ZN(n19232) );
  INV_X1 U11091 ( .A(n12163), .ZN(n15453) );
  INV_X2 U11092 ( .A(n12258), .ZN(n9595) );
  INV_X1 U11093 ( .A(n11528), .ZN(n15702) );
  NAND2_X1 U11094 ( .A1(n10118), .A2(n10119), .ZN(n10854) );
  NAND2_X1 U11095 ( .A1(n10566), .A2(n10565), .ZN(n15013) );
  XNOR2_X1 U11096 ( .A(n10193), .B(n10192), .ZN(n10201) );
  AND3_X1 U11097 ( .A1(n9695), .A2(n12975), .A3(n9578), .ZN(n15500) );
  NAND2_X1 U11098 ( .A1(n9859), .A2(n10215), .ZN(n19132) );
  INV_X2 U11099 ( .A(n9627), .ZN(n10121) );
  INV_X1 U11100 ( .A(n17465), .ZN(n17450) );
  INV_X1 U11101 ( .A(n15655), .ZN(n19809) );
  INV_X1 U11102 ( .A(n15677), .ZN(n15623) );
  NAND2_X1 U11103 ( .A1(n11536), .A2(n14581), .ZN(n14251) );
  NAND2_X1 U11104 ( .A1(n10127), .A2(n10661), .ZN(n11054) );
  NOR2_X1 U11105 ( .A1(n14876), .A2(n14863), .ZN(n14864) );
  NOR2_X1 U11106 ( .A1(n15359), .A2(n9708), .ZN(n15313) );
  BUF_X1 U11107 ( .A(n12618), .Z(n13444) );
  NAND2_X1 U11109 ( .A1(n10729), .A2(n10728), .ZN(n14972) );
  XNOR2_X1 U11110 ( .A(n10195), .B(n10194), .ZN(n10198) );
  INV_X1 U11111 ( .A(n17960), .ZN(n18605) );
  AOI221_X1 U11112 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17362), 
        .C1(n17723), .C2(n17381), .A(n17348), .ZN(n17349) );
  NAND2_X1 U11113 ( .A1(n17923), .A2(n18424), .ZN(n17882) );
  OR2_X1 U11114 ( .A1(n13210), .A2(n13212), .ZN(n15172) );
  NAND2_X1 U11115 ( .A1(n10196), .A2(n10189), .ZN(n15399) );
  NOR2_X1 U11116 ( .A1(n16770), .A2(n16794), .ZN(n16783) );
  AND2_X1 U11117 ( .A1(n11423), .A2(n11422), .ZN(n11454) );
  AND2_X1 U11118 ( .A1(n13738), .A2(n11056), .ZN(n9578) );
  AND2_X1 U11119 ( .A1(n9679), .A2(n13533), .ZN(n9579) );
  XOR2_X1 U11120 ( .A(n9798), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n9580)
         );
  AND2_X1 U11121 ( .A1(n15708), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9581) );
  XOR2_X1 U11122 ( .A(n19909), .B(n9604), .Z(n9582) );
  NAND2_X1 U11123 ( .A1(n10853), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10179) );
  NOR2_X2 U11124 ( .A1(n12120), .A2(n12119), .ZN(n12163) );
  OR2_X1 U11125 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  NAND2_X1 U11126 ( .A1(n18573), .A2(n18562), .ZN(n12118) );
  OAI21_X2 U11128 ( .B1(n18694), .B2(n10894), .A(n15065), .ZN(n15061) );
  NOR2_X1 U11129 ( .A1(n12117), .A2(n12119), .ZN(n12154) );
  BUF_X2 U11130 ( .A(n13716), .Z(n9587) );
  XNOR2_X1 U11131 ( .A(n10201), .B(n10197), .ZN(n13716) );
  NOR4_X1 U11133 ( .A1(n17960), .A2(n16612), .A3(n15604), .A4(n18452), .ZN(
        n16990) );
  INV_X2 U11134 ( .A(n9580), .ZN(n9589) );
  AND2_X1 U11135 ( .A1(n12778), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9590) );
  AND2_X1 U11136 ( .A1(n12778), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10294) );
  OAI211_X2 U11137 ( .C1(n9654), .C2(n13714), .A(n10157), .B(n10178), .ZN(
        n10186) );
  NOR2_X2 U11138 ( .A1(n17348), .A2(n12239), .ZN(n17300) );
  OR2_X2 U11139 ( .A1(n17348), .A2(n17337), .ZN(n17383) );
  OAI21_X2 U11140 ( .B1(n15079), .B2(n15080), .A(n12491), .ZN(n15025) );
  NOR2_X1 U11141 ( .A1(n17989), .A2(n17955), .ZN(n12340) );
  AND2_X2 U11142 ( .A1(n10624), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9591) );
  AND2_X1 U11143 ( .A1(n10624), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10236) );
  OR2_X1 U11144 ( .A1(n15167), .A2(n16040), .ZN(n9991) );
  XNOR2_X1 U11145 ( .A(n14950), .B(n14949), .ZN(n14963) );
  INV_X1 U11146 ( .A(n9884), .ZN(n14941) );
  NAND2_X1 U11147 ( .A1(n14960), .A2(n14959), .ZN(n15167) );
  NAND2_X1 U11148 ( .A1(n12470), .A2(n9723), .ZN(n15298) );
  NAND2_X1 U11149 ( .A1(n14050), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14049) );
  NAND2_X1 U11150 ( .A1(n9781), .A2(n9784), .ZN(n14050) );
  AND2_X1 U11151 ( .A1(n10712), .A2(n9782), .ZN(n9781) );
  NAND2_X1 U11152 ( .A1(n14334), .A2(n14323), .ZN(n14322) );
  OR2_X1 U11153 ( .A1(n14925), .A2(n14926), .ZN(n9671) );
  AND2_X2 U11154 ( .A1(n9645), .A2(n9646), .ZN(n15757) );
  NAND2_X1 U11155 ( .A1(n11665), .A2(n11664), .ZN(n13700) );
  AND2_X1 U11156 ( .A1(n13443), .A2(n13442), .ZN(n19678) );
  INV_X1 U11157 ( .A(n15702), .ZN(n15735) );
  OR2_X1 U11158 ( .A1(n11528), .A2(n15814), .ZN(n14625) );
  XNOR2_X1 U11159 ( .A(n9668), .B(n11503), .ZN(n11654) );
  XNOR2_X1 U11160 ( .A(n11491), .B(n11487), .ZN(n11643) );
  NAND2_X1 U11161 ( .A1(n13588), .A2(n13590), .ZN(n13589) );
  NAND2_X1 U11162 ( .A1(n11454), .A2(n11453), .ZN(n11491) );
  NOR2_X1 U11163 ( .A1(n10212), .A2(n13533), .ZN(n10199) );
  OAI21_X1 U11164 ( .B1(n15399), .B2(n12990), .A(n12637), .ZN(n15405) );
  INV_X2 U11165 ( .A(n9589), .ZN(n16599) );
  NOR2_X1 U11166 ( .A1(n16931), .A2(n16956), .ZN(n16953) );
  NOR2_X1 U11167 ( .A1(n14171), .A2(n15517), .ZN(n15494) );
  NOR2_X2 U11168 ( .A1(n17108), .A2(n16158), .ZN(n17518) );
  NAND2_X1 U11169 ( .A1(n11260), .A2(n11259), .ZN(n13019) );
  INV_X1 U11171 ( .A(n13778), .ZN(n9598) );
  NAND2_X1 U11172 ( .A1(n12502), .A2(n12501), .ZN(n12583) );
  INV_X1 U11173 ( .A(n12501), .ZN(n12997) );
  NOR2_X2 U11174 ( .A1(n12257), .A2(n12256), .ZN(n17960) );
  INV_X1 U11175 ( .A(n11612), .ZN(n9593) );
  NOR2_X1 U11176 ( .A1(n11206), .A2(n11205), .ZN(n11217) );
  AND4_X1 U11177 ( .A1(n11151), .A2(n11150), .A3(n11149), .A4(n11148), .ZN(
        n11157) );
  AND4_X1 U11178 ( .A1(n11155), .A2(n11154), .A3(n11153), .A4(n11152), .ZN(
        n11156) );
  CLKBUF_X3 U11179 ( .A(n12177), .Z(n16934) );
  CLKBUF_X2 U11181 ( .A(n12935), .Z(n12929) );
  CLKBUF_X2 U11182 ( .A(n12172), .Z(n16900) );
  CLKBUF_X3 U11183 ( .A(n12155), .Z(n9601) );
  BUF_X2 U11184 ( .A(n11278), .Z(n12071) );
  CLKBUF_X2 U11185 ( .A(n11327), .Z(n12074) );
  BUF_X2 U11186 ( .A(n11223), .Z(n12076) );
  BUF_X2 U11187 ( .A(n12064), .Z(n12043) );
  NOR2_X2 U11188 ( .A1(n18412), .A2(n12117), .ZN(n12207) );
  CLKBUF_X2 U11189 ( .A(n11298), .Z(n12065) );
  AND2_X2 U11190 ( .A1(n11104), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11112) );
  AND2_X1 U11191 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13669) );
  INV_X1 U11192 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18562) );
  NOR2_X1 U11193 ( .A1(n9880), .A2(n9881), .ZN(n15158) );
  NAND2_X1 U11194 ( .A1(n14941), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10730) );
  NAND2_X1 U11195 ( .A1(n14948), .A2(n14947), .ZN(n14950) );
  NOR2_X1 U11196 ( .A1(n12485), .A2(n9686), .ZN(n9785) );
  OAI21_X1 U11197 ( .B1(n9788), .B2(n9787), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9786) );
  OAI21_X1 U11198 ( .B1(n9778), .B2(n9908), .A(n9907), .ZN(n9909) );
  OR2_X1 U11199 ( .A1(n12474), .A2(n9789), .ZN(n9788) );
  OAI21_X1 U11200 ( .B1(n14250), .B2(n15655), .A(n9834), .ZN(n9833) );
  OR2_X1 U11201 ( .A1(n12889), .A2(n9961), .ZN(n9960) );
  AND2_X1 U11202 ( .A1(n14513), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9677) );
  NOR2_X1 U11203 ( .A1(n15298), .A2(n12472), .ZN(n15084) );
  AOI211_X1 U11204 ( .C1(n15731), .C2(n14549), .A(n14548), .B(n14547), .ZN(
        n14550) );
  XNOR2_X1 U11205 ( .A(n9657), .B(n12098), .ZN(n12500) );
  NOR2_X1 U11206 ( .A1(n14523), .A2(n9649), .ZN(n14513) );
  XNOR2_X1 U11207 ( .A(n14308), .B(n9987), .ZN(n14521) );
  AOI21_X1 U11208 ( .B1(n14962), .B2(n16001), .A(n14961), .ZN(n9873) );
  AND2_X1 U11209 ( .A1(n9962), .A2(n14811), .ZN(n9959) );
  XNOR2_X1 U11210 ( .A(n12987), .B(n10852), .ZN(n14271) );
  NOR2_X1 U11211 ( .A1(n15157), .A2(n9887), .ZN(n9886) );
  AND2_X1 U11212 ( .A1(n9945), .A2(n9699), .ZN(n15003) );
  OR2_X1 U11213 ( .A1(n12866), .A2(n12865), .ZN(n9962) );
  OR2_X1 U11214 ( .A1(n14335), .A2(n9989), .ZN(n14309) );
  NOR2_X1 U11215 ( .A1(n14335), .A2(n9988), .ZN(n14308) );
  CLKBUF_X1 U11216 ( .A(n14348), .Z(n14349) );
  OAI21_X1 U11217 ( .B1(n15102), .B2(n12489), .A(n15100), .ZN(n15094) );
  NAND2_X1 U11218 ( .A1(n11537), .A2(n14543), .ZN(n14535) );
  CLKBUF_X1 U11219 ( .A(n14376), .Z(n14377) );
  AND2_X1 U11220 ( .A1(n14827), .A2(n9742), .ZN(n14813) );
  NAND2_X1 U11221 ( .A1(n14831), .A2(n12815), .ZN(n12839) );
  NOR2_X2 U11222 ( .A1(n14835), .A2(n14826), .ZN(n14827) );
  AND2_X1 U11223 ( .A1(n9852), .A2(n9851), .ZN(n16154) );
  OAI21_X2 U11224 ( .B1(n14588), .B2(n9725), .A(n15702), .ZN(n14581) );
  NAND2_X1 U11225 ( .A1(n14582), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11536) );
  NAND2_X1 U11226 ( .A1(n14834), .A2(n10824), .ZN(n14835) );
  OAI21_X1 U11227 ( .B1(n14587), .B2(n11533), .A(n14633), .ZN(n14582) );
  OR2_X1 U11228 ( .A1(n17257), .A2(n16166), .ZN(n9852) );
  NAND2_X1 U11229 ( .A1(n10001), .A2(n10713), .ZN(n9784) );
  NOR2_X1 U11230 ( .A1(n17258), .A2(n9847), .ZN(n17257) );
  NAND2_X1 U11231 ( .A1(n14604), .A2(n9659), .ZN(n14587) );
  NOR3_X1 U11232 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17518), .A3(
        n12418), .ZN(n15530) );
  INV_X1 U11233 ( .A(n14604), .ZN(n9596) );
  AND2_X1 U11234 ( .A1(n10477), .A2(n9949), .ZN(n9948) );
  AOI21_X1 U11235 ( .B1(n16995), .B2(P3_EAX_REG_30__SCAN_IN), .A(n9726), .ZN(
        n16996) );
  NOR2_X1 U11236 ( .A1(n14911), .A2(n14905), .ZN(n14898) );
  NOR2_X1 U11237 ( .A1(n14284), .A2(n12956), .ZN(n12955) );
  NOR2_X1 U11238 ( .A1(n13213), .A2(n14882), .ZN(n14881) );
  XNOR2_X1 U11239 ( .A(n9836), .B(n13094), .ZN(n14659) );
  NAND2_X1 U11240 ( .A1(n14648), .A2(n11520), .ZN(n14608) );
  NAND2_X1 U11241 ( .A1(n9606), .A2(n9684), .ZN(n14648) );
  INV_X1 U11242 ( .A(n13093), .ZN(n9836) );
  AND2_X1 U11243 ( .A1(n17267), .A2(n12243), .ZN(n12244) );
  OAI211_X1 U11244 ( .C1(n9610), .C2(n15744), .A(n9607), .B(n11518), .ZN(n9606) );
  NOR2_X1 U11245 ( .A1(n9581), .A2(n9614), .ZN(n9613) );
  AND2_X1 U11246 ( .A1(n10717), .A2(n10724), .ZN(n15989) );
  AND2_X1 U11247 ( .A1(n9674), .A2(n12785), .ZN(n12761) );
  NAND2_X1 U11248 ( .A1(n10348), .A2(n13619), .ZN(n13762) );
  OR2_X1 U11249 ( .A1(n10707), .A2(n10716), .ZN(n10724) );
  AND2_X1 U11250 ( .A1(n11532), .A2(n9612), .ZN(n9611) );
  NOR2_X2 U11251 ( .A1(n19172), .A2(n19312), .ZN(n19157) );
  AND3_X2 U11252 ( .A1(n9630), .A2(n9867), .A3(n10699), .ZN(n10470) );
  AND2_X1 U11253 ( .A1(n10469), .A2(n10711), .ZN(n9934) );
  OR2_X1 U11254 ( .A1(n15244), .A2(n15245), .ZN(n15233) );
  NAND2_X1 U11255 ( .A1(n11645), .A2(n11644), .ZN(n13595) );
  AND2_X1 U11256 ( .A1(n10468), .A2(n10467), .ZN(n10711) );
  NOR2_X1 U11257 ( .A1(n17017), .A2(n17150), .ZN(n17011) );
  OR2_X1 U11258 ( .A1(n11531), .A2(n14623), .ZN(n14610) );
  NAND2_X1 U11259 ( .A1(n9614), .A2(n11522), .ZN(n9612) );
  INV_X1 U11260 ( .A(n14633), .ZN(n9614) );
  NOR2_X1 U11261 ( .A1(n15283), .A2(n14139), .ZN(n14138) );
  INV_X1 U11262 ( .A(n13564), .ZN(n9735) );
  INV_X1 U11263 ( .A(n15702), .ZN(n14633) );
  AND2_X1 U11264 ( .A1(n11499), .A2(n11498), .ZN(n15751) );
  INV_X1 U11265 ( .A(n15702), .ZN(n9597) );
  OAI211_X1 U11266 ( .C1(n10402), .C2(n12881), .A(n10404), .B(n10403), .ZN(
        n10405) );
  NAND2_X1 U11267 ( .A1(n11493), .A2(n11492), .ZN(n11653) );
  NAND2_X1 U11268 ( .A1(n14444), .A2(n14441), .ZN(n14440) );
  AND2_X1 U11269 ( .A1(n12625), .A2(n13575), .ZN(n13440) );
  OR2_X1 U11270 ( .A1(n12645), .A2(n12624), .ZN(n12625) );
  NOR2_X2 U11271 ( .A1(n14454), .A2(n14445), .ZN(n14444) );
  NAND2_X1 U11272 ( .A1(n11452), .A2(n11425), .ZN(n11624) );
  NOR2_X1 U11273 ( .A1(n17158), .A2(n17031), .ZN(n17030) );
  NAND2_X1 U11274 ( .A1(n12623), .A2(n12622), .ZN(n12645) );
  NAND2_X1 U11275 ( .A1(n12631), .A2(n12632), .ZN(n12643) );
  NOR3_X1 U11276 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n12231), .ZN(n17419) );
  OAI21_X1 U11277 ( .B1(n13690), .B2(n11752), .A(n11603), .ZN(n9958) );
  CLKBUF_X1 U11278 ( .A(n12461), .Z(n14510) );
  INV_X1 U11279 ( .A(n11424), .ZN(n11423) );
  NOR2_X1 U11280 ( .A1(n12230), .A2(n9847), .ZN(n9845) );
  INV_X2 U11281 ( .A(n17806), .ZN(n18384) );
  AND2_X1 U11282 ( .A1(n14227), .A2(n9714), .ZN(n15372) );
  NOR2_X1 U11283 ( .A1(n10218), .A2(n9858), .ZN(n9857) );
  NOR2_X1 U11284 ( .A1(n17080), .A2(n17256), .ZN(n17073) );
  INV_X1 U11285 ( .A(n13716), .ZN(n10212) );
  AND2_X1 U11286 ( .A1(n11421), .A2(n11420), .ZN(n19961) );
  NAND2_X1 U11287 ( .A1(n17960), .A2(n12363), .ZN(n17806) );
  XNOR2_X1 U11288 ( .A(n15405), .B(n12638), .ZN(n13287) );
  OR2_X1 U11289 ( .A1(n10485), .A2(n9930), .ZN(n10591) );
  INV_X2 U11290 ( .A(n17079), .ZN(n17131) );
  AOI21_X1 U11291 ( .B1(n9648), .B2(n20790), .A(n9994), .ZN(n11386) );
  NOR2_X2 U11292 ( .A1(n18385), .A2(n18409), .ZN(n17923) );
  OAI21_X1 U11293 ( .B1(n10184), .B2(n10190), .A(n10191), .ZN(n10174) );
  AND2_X1 U11294 ( .A1(n10482), .A2(n9693), .ZN(n10494) );
  XNOR2_X1 U11295 ( .A(n10734), .B(n10735), .ZN(n10733) );
  NAND2_X1 U11296 ( .A1(n12527), .A2(n10005), .ZN(n13704) );
  NAND2_X1 U11297 ( .A1(n9957), .A2(n11380), .ZN(n11389) );
  AND2_X1 U11298 ( .A1(n10472), .A2(n10473), .ZN(n10482) );
  NOR2_X1 U11299 ( .A1(n13517), .A2(n10875), .ZN(n13621) );
  NAND2_X1 U11300 ( .A1(n11323), .A2(n11322), .ZN(n20009) );
  NOR3_X2 U11301 ( .A1(n12350), .A2(n12349), .A3(n15489), .ZN(n18398) );
  NAND2_X1 U11302 ( .A1(n11406), .A2(n11405), .ZN(n20113) );
  AOI221_X2 U11303 ( .B1(n17960), .B2(n18408), .C1(n15493), .C2(n18408), .A(
        n15496), .ZN(n15606) );
  AOI21_X1 U11304 ( .B1(n9698), .B2(n10891), .A(n9904), .ZN(n9903) );
  INV_X1 U11305 ( .A(n18411), .ZN(n18413) );
  NOR2_X1 U11306 ( .A1(n10376), .A2(n10375), .ZN(n10423) );
  AND2_X1 U11307 ( .A1(n11321), .A2(n11320), .ZN(n11324) );
  NOR2_X1 U11308 ( .A1(n13569), .A2(n13568), .ZN(n15874) );
  NAND2_X1 U11309 ( .A1(n10349), .A2(n10347), .ZN(n10376) );
  NOR2_X2 U11310 ( .A1(n10350), .A2(n10355), .ZN(n10349) );
  NAND2_X1 U11311 ( .A1(n9933), .A2(n10161), .ZN(n10853) );
  NAND2_X1 U11312 ( .A1(n17569), .A2(n17570), .ZN(n17568) );
  OAI211_X1 U11313 ( .C1(n18599), .C2(n17960), .A(n17208), .B(n17207), .ZN(
        n17252) );
  NAND2_X1 U11314 ( .A1(n11318), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11348) );
  OR2_X1 U11315 ( .A1(n13556), .A2(n13555), .ZN(n13569) );
  XNOR2_X1 U11316 ( .A(n9672), .B(n13102), .ZN(n14269) );
  NAND2_X1 U11317 ( .A1(n10338), .A2(n10337), .ZN(n10350) );
  INV_X1 U11318 ( .A(n10835), .ZN(n10847) );
  AND2_X1 U11319 ( .A1(n11265), .A2(n11252), .ZN(n13038) );
  NOR2_X1 U11320 ( .A1(n18402), .A2(n17965), .ZN(n16277) );
  NAND2_X1 U11321 ( .A1(n9687), .A2(n12951), .ZN(n10155) );
  NAND4_X1 U11322 ( .A1(n10126), .A2(n10125), .A3(n11054), .A4(n11061), .ZN(
        n10161) );
  OR2_X1 U11323 ( .A1(n12330), .A2(n12343), .ZN(n18402) );
  CLKBUF_X1 U11324 ( .A(n10628), .Z(n16070) );
  AND2_X1 U11325 ( .A1(n11061), .A2(n13785), .ZN(n9932) );
  AOI21_X1 U11326 ( .B1(n12347), .B2(n17977), .A(n15512), .ZN(n12335) );
  AND2_X1 U11327 ( .A1(n10143), .A2(n10122), .ZN(n10126) );
  NAND2_X1 U11328 ( .A1(n10091), .A2(n10141), .ZN(n10138) );
  OAI21_X1 U11329 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(n12586), .A(n12505), .ZN(
        n12509) );
  AND2_X1 U11330 ( .A1(n10340), .A2(n10867), .ZN(n10355) );
  AND2_X1 U11331 ( .A1(n11247), .A2(n11254), .ZN(n11267) );
  NOR2_X1 U11332 ( .A1(n11309), .A2(n20790), .ZN(n11512) );
  AND2_X1 U11333 ( .A1(n14305), .A2(n12565), .ZN(n13249) );
  NAND2_X1 U11334 ( .A1(n14302), .A2(n13089), .ZN(n13386) );
  AND2_X1 U11335 ( .A1(n14156), .A2(n11256), .ZN(n11257) );
  AND2_X1 U11336 ( .A1(n11195), .A2(n11194), .ZN(n11196) );
  OR2_X1 U11337 ( .A1(n12565), .A2(n12520), .ZN(n12586) );
  NAND4_X1 U11338 ( .A1(n12957), .A2(n11056), .A3(n9656), .A4(n13785), .ZN(
        n11059) );
  OR2_X1 U11339 ( .A1(n10646), .A2(n13754), .ZN(n10648) );
  INV_X1 U11340 ( .A(n15510), .ZN(n17973) );
  OR2_X1 U11341 ( .A1(n10308), .A2(n10307), .ZN(n10345) );
  NAND3_X1 U11342 ( .A1(n12278), .A2(n12277), .A3(n12276), .ZN(n15509) );
  OR2_X1 U11343 ( .A1(n10268), .A2(n10267), .ZN(n9912) );
  OR2_X1 U11344 ( .A1(n10256), .A2(n10255), .ZN(n10687) );
  AND2_X1 U11345 ( .A1(n11258), .A2(n11255), .ZN(n13089) );
  NAND4_X2 U11346 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10478) );
  NAND3_X1 U11347 ( .A1(n12268), .A2(n12267), .A3(n12266), .ZN(n17955) );
  XNOR2_X1 U11348 ( .A(n12394), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17599) );
  AOI211_X1 U11349 ( .C1(n9595), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n12265), .B(n12264), .ZN(n12266) );
  CLKBUF_X2 U11350 ( .A(n9593), .Z(n11270) );
  AND2_X2 U11351 ( .A1(n12501), .A2(n19979), .ZN(n13410) );
  OR2_X1 U11352 ( .A1(n11291), .A2(n11290), .ZN(n11515) );
  OR2_X1 U11353 ( .A1(n11306), .A2(n11305), .ZN(n11395) );
  NOR2_X2 U11354 ( .A1(n17351), .A2(n17350), .ZN(n17325) );
  CLKBUF_X1 U11355 ( .A(n11242), .Z(n11243) );
  NAND2_X1 U11356 ( .A1(n10065), .A2(n10064), .ZN(n13754) );
  NAND2_X1 U11357 ( .A1(n10053), .A2(n10052), .ZN(n10144) );
  NAND2_X2 U11358 ( .A1(n10014), .A2(n9675), .ZN(n11254) );
  AND4_X1 U11359 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n10070) );
  INV_X2 U11360 ( .A(U214), .ZN(n16224) );
  AND2_X2 U11361 ( .A1(n11119), .A2(n11118), .ZN(n11612) );
  NAND4_X2 U11362 ( .A1(n11139), .A2(n11138), .A3(n11137), .A4(n11136), .ZN(
        n11249) );
  AND4_X1 U11363 ( .A1(n11131), .A2(n11130), .A3(n11129), .A4(n11128), .ZN(
        n11137) );
  AND4_X1 U11364 ( .A1(n11117), .A2(n11116), .A3(n11115), .A4(n11114), .ZN(
        n11118) );
  AND4_X1 U11365 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n11138) );
  AND4_X1 U11366 ( .A1(n11108), .A2(n11107), .A3(n11106), .A4(n11105), .ZN(
        n11119) );
  AND4_X1 U11367 ( .A1(n11123), .A2(n11122), .A3(n11121), .A4(n11120), .ZN(
        n11139) );
  INV_X2 U11368 ( .A(n16262), .ZN(U215) );
  AND4_X1 U11369 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(
        n11216) );
  AND4_X1 U11370 ( .A1(n11235), .A2(n11234), .A3(n11233), .A4(n11232), .ZN(
        n11236) );
  AND4_X1 U11371 ( .A1(n11167), .A2(n11166), .A3(n11165), .A4(n11164), .ZN(
        n9675) );
  AND4_X1 U11372 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n11237) );
  AND4_X1 U11373 ( .A1(n11201), .A2(n11200), .A3(n11199), .A4(n11198), .ZN(
        n11218) );
  AND4_X1 U11374 ( .A1(n11143), .A2(n11142), .A3(n11141), .A4(n11140), .ZN(
        n11159) );
  AND4_X1 U11375 ( .A1(n11135), .A2(n11134), .A3(n11133), .A4(n11132), .ZN(
        n11136) );
  AND4_X1 U11376 ( .A1(n11222), .A2(n11221), .A3(n11220), .A4(n11219), .ZN(
        n11239) );
  AND4_X1 U11377 ( .A1(n11191), .A2(n11190), .A3(n11189), .A4(n11188), .ZN(
        n11192) );
  AND4_X1 U11378 ( .A1(n11227), .A2(n11226), .A3(n11225), .A4(n11224), .ZN(
        n11238) );
  NAND2_X2 U11379 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19736), .ZN(n19656) );
  NAND2_X2 U11380 ( .A1(n19736), .A2(n19608), .ZN(n19655) );
  INV_X2 U11381 ( .A(n19853), .ZN(n19873) );
  BUF_X2 U11382 ( .A(n11276), .Z(n12066) );
  BUF_X2 U11383 ( .A(n12207), .Z(n16935) );
  BUF_X2 U11384 ( .A(n12250), .Z(n16944) );
  BUF_X2 U11385 ( .A(n12172), .Z(n16877) );
  NAND2_X2 U11386 ( .A1(n18543), .A2(n18482), .ZN(n18540) );
  BUF_X2 U11387 ( .A(n11325), .Z(n11368) );
  INV_X2 U11388 ( .A(n19942), .ZN(n12105) );
  AND2_X2 U11389 ( .A1(n11110), .A2(n13669), .ZN(n11326) );
  INV_X2 U11390 ( .A(n16266), .ZN(n16268) );
  OR2_X1 U11391 ( .A1(n12115), .A2(n12116), .ZN(n12127) );
  BUF_X2 U11392 ( .A(n11300), .Z(n12075) );
  AND2_X2 U11393 ( .A1(n11112), .A2(n13682), .ZN(n11276) );
  AND2_X2 U11394 ( .A1(n11110), .A2(n11112), .ZN(n11277) );
  AND2_X2 U11395 ( .A1(n11109), .A2(n11111), .ZN(n11278) );
  AND2_X1 U11396 ( .A1(n11112), .A2(n13418), .ZN(n11989) );
  NOR2_X1 U11397 ( .A1(n18566), .A2(n18464), .ZN(n18600) );
  NAND4_X1 U11398 ( .A1(n18608), .A2(n18617), .A3(n16275), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18460) );
  NOR2_X1 U11399 ( .A1(n18412), .A2(n12120), .ZN(n12110) );
  NAND2_X1 U11400 ( .A1(n18573), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12116) );
  NAND3_X1 U11401 ( .A1(n15797), .A2(n11521), .A3(n12552), .ZN(n11522) );
  INV_X1 U11402 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9634) );
  INV_X1 U11403 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11263) );
  INV_X1 U11404 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9635) );
  NOR2_X2 U11405 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11111) );
  AND2_X2 U11406 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13418) );
  INV_X1 U11407 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19729) );
  AND2_X1 U11408 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13448) );
  INV_X1 U11409 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19064) );
  INV_X1 U11410 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U11411 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18412) );
  INV_X1 U11412 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10228) );
  INV_X1 U11413 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12766) );
  NAND2_X1 U11414 ( .A1(n9603), .A2(n11451), .ZN(n9646) );
  INV_X1 U11415 ( .A(n9604), .ZN(n9603) );
  XNOR2_X1 U11416 ( .A(n11450), .B(n19922), .ZN(n9604) );
  XNOR2_X1 U11417 ( .A(n11473), .B(n20699), .ZN(n15756) );
  NAND2_X1 U11418 ( .A1(n9605), .A2(n11472), .ZN(n11473) );
  NAND2_X1 U11419 ( .A1(n11643), .A2(n11511), .ZN(n9605) );
  INV_X1 U11420 ( .A(n15746), .ZN(n9609) );
  NAND2_X1 U11421 ( .A1(n9609), .A2(n15745), .ZN(n9607) );
  NAND2_X1 U11422 ( .A1(n9608), .A2(n15745), .ZN(n14002) );
  NAND2_X1 U11423 ( .A1(n15744), .A2(n15746), .ZN(n9608) );
  INV_X1 U11424 ( .A(n15745), .ZN(n9610) );
  OAI21_X2 U11425 ( .B1(n14608), .B2(n9613), .A(n9611), .ZN(n14604) );
  AND2_X4 U11426 ( .A1(n11109), .A2(n13669), .ZN(n11332) );
  AND2_X2 U11427 ( .A1(n11263), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11109) );
  OAI21_X2 U11428 ( .B1(n9624), .B2(n11361), .A(n9615), .ZN(n13417) );
  NOR2_X1 U11429 ( .A1(n9615), .A2(n20360), .ZN(n13405) );
  XNOR2_X1 U11430 ( .A(n9615), .B(n20113), .ZN(n20233) );
  NAND2_X2 U11431 ( .A1(n11362), .A2(n11361), .ZN(n9615) );
  OR2_X2 U11432 ( .A1(n11178), .A2(n11179), .ZN(n19987) );
  NAND2_X1 U11433 ( .A1(n10162), .A2(n9619), .ZN(n9616) );
  AND2_X1 U11434 ( .A1(n9616), .A2(n9617), .ZN(n10185) );
  OR2_X1 U11435 ( .A1(n9618), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9617) );
  INV_X1 U11436 ( .A(n10163), .ZN(n9618) );
  AND2_X1 U11437 ( .A1(n10161), .A2(n10163), .ZN(n9619) );
  NOR2_X1 U11438 ( .A1(n10116), .A2(n10115), .ZN(n10117) );
  OR2_X1 U11439 ( .A1(n10110), .A2(n10109), .ZN(n10116) );
  INV_X1 U11440 ( .A(n12939), .ZN(n9620) );
  NOR2_X2 U11441 ( .A1(n16483), .A2(n16835), .ZN(n16811) );
  NOR2_X2 U11442 ( .A1(n16729), .A2(n15410), .ZN(n16715) );
  NAND2_X1 U11443 ( .A1(n13589), .A2(n11401), .ZN(n11432) );
  NAND2_X1 U11444 ( .A1(n11340), .A2(n11257), .ZN(n9621) );
  NAND2_X1 U11445 ( .A1(n11340), .A2(n11257), .ZN(n13393) );
  NAND2_X1 U11446 ( .A1(n9679), .A2(n10227), .ZN(n19280) );
  CLKBUF_X1 U11447 ( .A(n13989), .Z(n9622) );
  NOR2_X2 U11448 ( .A1(n10531), .A2(n10530), .ZN(n10522) );
  NOR2_X2 U11449 ( .A1(n10528), .A2(n10526), .ZN(n10519) );
  NAND2_X1 U11450 ( .A1(n14535), .A2(n11538), .ZN(n14523) );
  BUF_X2 U11451 ( .A(n9670), .Z(n10402) );
  NOR2_X2 U11453 ( .A1(n14404), .A2(n14387), .ZN(n14373) );
  NOR2_X4 U11454 ( .A1(n14105), .A2(n12551), .ZN(n14154) );
  INV_X2 U11455 ( .A(n13410), .ZN(n12520) );
  INV_X2 U11456 ( .A(n10339), .ZN(n9656) );
  NAND2_X1 U11457 ( .A1(n11353), .A2(n11352), .ZN(n9624) );
  INV_X1 U11458 ( .A(n9596), .ZN(n9625) );
  NAND2_X1 U11459 ( .A1(n14002), .A2(n11518), .ZN(n9626) );
  NAND2_X1 U11460 ( .A1(n11353), .A2(n11352), .ZN(n11362) );
  MUX2_X2 U11461 ( .A(n9628), .B(n9629), .S(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n9627) );
  NAND4_X1 U11462 ( .A1(n10095), .A2(n10094), .A3(n10093), .A4(n10092), .ZN(
        n9628) );
  NAND4_X1 U11463 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n9629) );
  NAND2_X1 U11464 ( .A1(n10024), .A2(n10023), .ZN(n10032) );
  INV_X1 U11465 ( .A(n10661), .ZN(n16067) );
  INV_X1 U11466 ( .A(n10311), .ZN(n9630) );
  OR2_X1 U11467 ( .A1(n10206), .A2(n10205), .ZN(n10211) );
  NAND2_X1 U11468 ( .A1(n9579), .A2(n9587), .ZN(n9631) );
  NAND2_X1 U11470 ( .A1(n12437), .A2(n12444), .ZN(n13013) );
  NOR2_X2 U11471 ( .A1(n12918), .A2(n12917), .ZN(n12928) );
  NAND2_X1 U11472 ( .A1(n9579), .A2(n10212), .ZN(n9670) );
  INV_X1 U11473 ( .A(n10854), .ZN(n9633) );
  NOR2_X2 U11474 ( .A1(n13021), .A2(n11246), .ZN(n11265) );
  NAND2_X2 U11475 ( .A1(n10186), .A2(n10185), .ZN(n10184) );
  NOR2_X1 U11476 ( .A1(n16055), .A2(n9583), .ZN(n18942) );
  NAND2_X2 U11477 ( .A1(n9679), .A2(n10199), .ZN(n10392) );
  AND2_X2 U11478 ( .A1(n12618), .A2(n15399), .ZN(n9679) );
  NOR2_X1 U11479 ( .A1(n9636), .A2(n9637), .ZN(n9639) );
  OR2_X1 U11480 ( .A1(n11244), .A2(n12501), .ZN(n9636) );
  NAND2_X1 U11481 ( .A1(n11195), .A2(n9638), .ZN(n9637) );
  NAND2_X1 U11482 ( .A1(n11244), .A2(n19983), .ZN(n9638) );
  NAND2_X1 U11483 ( .A1(n11197), .A2(n11196), .ZN(n9640) );
  INV_X1 U11484 ( .A(n9640), .ZN(n13040) );
  NOR2_X2 U11485 ( .A1(n17733), .A2(n17511), .ZN(n17391) );
  AOI22_X1 U11486 ( .A1(n17805), .A2(n17601), .B1(n17520), .B2(n17808), .ZN(
        n17511) );
  NAND2_X1 U11487 ( .A1(n13600), .A2(n13602), .ZN(n9641) );
  NAND2_X1 U11488 ( .A1(n13600), .A2(n13602), .ZN(n13601) );
  OR2_X2 U11489 ( .A1(n11491), .A2(n11489), .ZN(n9668) );
  NAND2_X1 U11490 ( .A1(n11423), .A2(n11422), .ZN(n11452) );
  XNOR2_X1 U11491 ( .A(n11452), .B(n11453), .ZN(n11599) );
  NOR2_X1 U11492 ( .A1(n13595), .A2(n13709), .ZN(n9642) );
  NOR2_X2 U11493 ( .A1(n13769), .A2(n9643), .ZN(n13967) );
  OR2_X1 U11494 ( .A1(n13943), .A2(n9644), .ZN(n9643) );
  INV_X1 U11495 ( .A(n13970), .ZN(n9644) );
  NOR2_X2 U11496 ( .A1(n13595), .A2(n13709), .ZN(n13699) );
  NAND2_X1 U11497 ( .A1(n13601), .A2(n9647), .ZN(n9645) );
  AND2_X1 U11498 ( .A1(n11433), .A2(n11451), .ZN(n9647) );
  NOR2_X2 U11499 ( .A1(n12501), .A2(n19979), .ZN(n14302) );
  INV_X1 U11500 ( .A(n9648), .ZN(n13694) );
  OR2_X1 U11501 ( .A1(n11244), .A2(n13022), .ZN(n13385) );
  AND2_X2 U11502 ( .A1(n20009), .A2(n11353), .ZN(n9648) );
  XNOR2_X1 U11503 ( .A(n9650), .B(n9649), .ZN(n14677) );
  INV_X1 U11504 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9649) );
  NOR2_X1 U11505 ( .A1(n14525), .A2(n14524), .ZN(n9650) );
  NOR2_X2 U11506 ( .A1(n18605), .A2(n16279), .ZN(n17601) );
  AND2_X2 U11507 ( .A1(n9639), .A2(n11197), .ZN(n12492) );
  NAND2_X1 U11509 ( .A1(n9641), .A2(n11433), .ZN(n19909) );
  OR2_X1 U11510 ( .A1(n13023), .A2(n11180), .ZN(n12998) );
  OAI211_X2 U11511 ( .C1(n15028), .C2(n15027), .A(n15049), .B(n15061), .ZN(
        n15040) );
  NOR2_X2 U11512 ( .A1(n14020), .A2(n14019), .ZN(n14018) );
  AOI21_X2 U11513 ( .B1(n11251), .B2(n19987), .A(n11181), .ZN(n11197) );
  OR2_X1 U11514 ( .A1(n12618), .A2(n13533), .ZN(n10226) );
  NOR2_X1 U11515 ( .A1(n13769), .A2(n13943), .ZN(n13942) );
  AOI211_X2 U11516 ( .C1(n15731), .C2(n14326), .A(n14264), .B(n14263), .ZN(
        n14265) );
  NOR2_X2 U11517 ( .A1(n12488), .A2(n15110), .ZN(n15102) );
  NAND4_X4 U11518 ( .A1(n11159), .A2(n11158), .A3(n11157), .A4(n11156), .ZN(
        n11180) );
  AND2_X1 U11519 ( .A1(n11112), .A2(n13418), .ZN(n9652) );
  AND2_X1 U11520 ( .A1(n11112), .A2(n13418), .ZN(n9653) );
  XNOR2_X2 U11521 ( .A(n11378), .B(n11377), .ZN(n11392) );
  OAI22_X2 U11522 ( .A1(n13417), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11426), 
        .B2(n11408), .ZN(n11378) );
  XNOR2_X1 U11523 ( .A(n13433), .B(n11345), .ZN(n13489) );
  NAND2_X2 U11524 ( .A1(n9668), .A2(n11513), .ZN(n11528) );
  NAND2_X2 U11525 ( .A1(n11392), .A2(n11391), .ZN(n11424) );
  OR2_X2 U11526 ( .A1(n11392), .A2(n11391), .ZN(n11393) );
  NAND2_X1 U11527 ( .A1(n20071), .A2(n11324), .ZN(n11353) );
  NAND2_X2 U11528 ( .A1(n12492), .A2(n11253), .ZN(n12437) );
  NAND2_X1 U11529 ( .A1(n10853), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9654) );
  XNOR2_X1 U11530 ( .A(n11432), .B(n19933), .ZN(n13600) );
  AOI21_X1 U11531 ( .B1(n11604), .B2(n11386), .A(n11390), .ZN(n11391) );
  XNOR2_X1 U11532 ( .A(n11400), .B(n19954), .ZN(n13588) );
  NAND2_X1 U11533 ( .A1(n13490), .A2(n11347), .ZN(n11400) );
  INV_X1 U11534 ( .A(n10339), .ZN(n9655) );
  NOR2_X2 U11535 ( .A1(n18619), .A2(n14171), .ZN(n18385) );
  NAND2_X1 U11536 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9871) );
  NAND2_X1 U11537 ( .A1(n9779), .A2(n10584), .ZN(n9778) );
  NAND2_X1 U11538 ( .A1(n10583), .A2(n11090), .ZN(n9779) );
  AND4_X1 U11539 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10330) );
  AND4_X1 U11540 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10329) );
  AND4_X1 U11541 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10331) );
  NAND2_X1 U11542 ( .A1(n10858), .A2(n10339), .ZN(n11005) );
  NOR3_X1 U11543 ( .A1(n17983), .A2(n15509), .A3(n18399), .ZN(n14173) );
  NOR2_X1 U11544 ( .A1(n9762), .A2(n9759), .ZN(n9758) );
  INV_X1 U11545 ( .A(n10616), .ZN(n9759) );
  NAND2_X1 U11546 ( .A1(n10135), .A2(n10134), .ZN(n10137) );
  AND2_X1 U11547 ( .A1(n10133), .A2(n9627), .ZN(n10134) );
  NAND2_X1 U11548 ( .A1(n11059), .A2(n9598), .ZN(n10133) );
  INV_X1 U11549 ( .A(n10178), .ZN(n10164) );
  OR2_X1 U11550 ( .A1(n12359), .A2(n12360), .ZN(n12352) );
  NAND3_X1 U11551 ( .A1(n11180), .A2(n12501), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11575) );
  OR2_X1 U11552 ( .A1(n12501), .A2(n20790), .ZN(n11407) );
  NOR2_X1 U11553 ( .A1(n10620), .A2(n10618), .ZN(n10668) );
  OR2_X1 U11554 ( .A1(n10835), .A2(n10168), .ZN(n10170) );
  AND2_X1 U11555 ( .A1(n9965), .A2(n9964), .ZN(n9963) );
  INV_X1 U11556 ( .A(n14390), .ZN(n9964) );
  OR2_X1 U11557 ( .A1(n11338), .A2(n11337), .ZN(n11394) );
  OR2_X1 U11558 ( .A1(n11180), .A2(n20790), .ZN(n11408) );
  OAI21_X1 U11559 ( .B1(n13688), .B2(n14789), .A(n20623), .ZN(n19963) );
  NOR2_X1 U11560 ( .A1(n10017), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10018) );
  INV_X1 U11561 ( .A(n9663), .ZN(n9976) );
  INV_X1 U11563 ( .A(n15328), .ZN(n9893) );
  INV_X1 U11564 ( .A(n10183), .ZN(n10735) );
  OAI21_X1 U11565 ( .B1(n9651), .B2(n16047), .A(n10182), .ZN(n10183) );
  NOR2_X1 U11566 ( .A1(n10514), .A2(n9776), .ZN(n9775) );
  INV_X1 U11567 ( .A(n10506), .ZN(n9776) );
  NOR2_X1 U11568 ( .A1(n10127), .A2(n19729), .ZN(n9864) );
  NAND2_X1 U11569 ( .A1(n12630), .A2(n12629), .ZN(n12631) );
  AND2_X1 U11570 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19450), .ZN(
        n12626) );
  NOR2_X1 U11571 ( .A1(n12118), .A2(n18412), .ZN(n12149) );
  OAI21_X1 U11572 ( .B1(n12348), .B2(n12347), .A(n12346), .ZN(n15489) );
  OR2_X1 U11573 ( .A1(n14295), .A2(n14301), .ZN(n13401) );
  NAND2_X1 U11574 ( .A1(n11253), .A2(n12501), .ZN(n13251) );
  INV_X1 U11575 ( .A(n13857), .ZN(n9905) );
  INV_X1 U11576 ( .A(n12985), .ZN(n10846) );
  NAND2_X1 U11577 ( .A1(n14953), .A2(n15164), .ZN(n9910) );
  NAND2_X1 U11578 ( .A1(n10686), .A2(n10685), .ZN(n11075) );
  AND2_X1 U11579 ( .A1(n10675), .A2(n10674), .ZN(n16055) );
  OR2_X1 U11580 ( .A1(n18946), .A2(n10673), .ZN(n10674) );
  OR2_X1 U11581 ( .A1(n13152), .A2(n19504), .ZN(n18631) );
  NAND2_X1 U11582 ( .A1(n12331), .A2(n12348), .ZN(n15493) );
  AND2_X1 U11583 ( .A1(n16369), .A2(n9589), .ZN(n16358) );
  AOI21_X1 U11584 ( .B1(n14173), .B2(n14172), .A(n15494), .ZN(n15604) );
  NAND2_X1 U11585 ( .A1(n17579), .A2(n12220), .ZN(n17569) );
  INV_X1 U11586 ( .A(n16165), .ZN(n9851) );
  NOR2_X1 U11587 ( .A1(n18617), .A2(n18455), .ZN(n18603) );
  INV_X1 U11588 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n9858) );
  CLKBUF_X1 U11589 ( .A(n11363), .Z(n12073) );
  AOI22_X1 U11590 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11326), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U11591 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11332), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11105) );
  AND2_X1 U11592 ( .A1(n11486), .A2(n11485), .ZN(n11492) );
  AND2_X2 U11593 ( .A1(n11358), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11113) );
  AOI21_X1 U11594 ( .B1(n11551), .B2(n11550), .A(n11547), .ZN(n11579) );
  NOR2_X1 U11595 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n11548), .ZN(
        n11578) );
  OR2_X1 U11596 ( .A1(n13193), .A2(n10576), .ZN(n10577) );
  AND4_X1 U11597 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10324), .ZN(
        n10328) );
  AND2_X1 U11598 ( .A1(n10148), .A2(n11065), .ZN(n10149) );
  OAI211_X1 U11599 ( .C1(n12954), .C2(n11056), .A(n10648), .B(n13800), .ZN(
        n11052) );
  INV_X1 U11600 ( .A(n10214), .ZN(n10221) );
  AND2_X1 U11601 ( .A1(n18869), .A2(n10201), .ZN(n10214) );
  AOI22_X1 U11602 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U11603 ( .A1(n10371), .A2(n10370), .ZN(n10620) );
  OR2_X1 U11604 ( .A1(n10369), .A2(n10368), .ZN(n10371) );
  NAND2_X1 U11605 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16073), .ZN(
        n10618) );
  NAND2_X1 U11606 ( .A1(n17973), .A2(n17983), .ZN(n12347) );
  AOI21_X1 U11607 ( .B1(n12998), .B2(n14796), .A(n11258), .ZN(n11252) );
  NAND2_X1 U11608 ( .A1(n14261), .A2(n9990), .ZN(n9989) );
  INV_X1 U11609 ( .A(n14337), .ZN(n9990) );
  NAND2_X1 U11610 ( .A1(n11803), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12059) );
  NOR2_X1 U11611 ( .A1(n11907), .A2(n9967), .ZN(n9966) );
  INV_X1 U11612 ( .A(n14443), .ZN(n9967) );
  NOR2_X1 U11613 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  INV_X1 U11614 ( .A(n14461), .ZN(n9970) );
  AND2_X1 U11615 ( .A1(n11592), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11637) );
  OR2_X1 U11616 ( .A1(n11254), .A2(n20640), .ZN(n12090) );
  NAND2_X1 U11617 ( .A1(n9596), .A2(n11534), .ZN(n14588) );
  NOR2_X1 U11618 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11534) );
  NOR2_X1 U11619 ( .A1(n9831), .A2(n9830), .ZN(n9829) );
  INV_X1 U11620 ( .A(n14458), .ZN(n9831) );
  INV_X1 U11621 ( .A(n14153), .ZN(n9830) );
  NAND2_X1 U11622 ( .A1(n13410), .A2(n12565), .ZN(n12580) );
  AND3_X1 U11623 ( .A1(n11540), .A2(n11340), .A3(n11539), .ZN(n13015) );
  NAND2_X1 U11624 ( .A1(n19994), .A2(n19979), .ZN(n11541) );
  AND2_X1 U11625 ( .A1(n11379), .A2(n20790), .ZN(n9744) );
  NAND2_X1 U11626 ( .A1(n11308), .A2(n9747), .ZN(n9746) );
  NAND2_X1 U11627 ( .A1(n9749), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9747) );
  INV_X1 U11628 ( .A(n11376), .ZN(n11426) );
  AND3_X1 U11629 ( .A1(n11385), .A2(n11384), .A3(n11383), .ZN(n11387) );
  INV_X1 U11630 ( .A(n11185), .ZN(n11186) );
  NOR2_X1 U11631 ( .A1(n11575), .A2(n11541), .ZN(n11577) );
  NAND2_X1 U11632 ( .A1(n11408), .A2(n11407), .ZN(n11555) );
  OAI21_X1 U11633 ( .B1(n9912), .B2(n10127), .A(n10336), .ZN(n10630) );
  OR2_X1 U11634 ( .A1(n10332), .A2(n10335), .ZN(n10336) );
  OR2_X1 U11635 ( .A1(n10594), .A2(n9906), .ZN(n10611) );
  INV_X1 U11636 ( .A(n10591), .ZN(n9906) );
  NAND2_X1 U11637 ( .A1(n10568), .A2(n9913), .ZN(n10593) );
  AND2_X1 U11638 ( .A1(n9718), .A2(n14838), .ZN(n9913) );
  NAND2_X1 U11639 ( .A1(n10567), .A2(n10591), .ZN(n10568) );
  NAND2_X1 U11640 ( .A1(n10481), .A2(n9929), .ZN(n9928) );
  INV_X1 U11641 ( .A(n10483), .ZN(n9929) );
  NAND2_X1 U11642 ( .A1(n14823), .A2(n12842), .ZN(n12866) );
  INV_X1 U11643 ( .A(n14860), .ZN(n9977) );
  AND2_X1 U11644 ( .A1(n13812), .A2(n12670), .ZN(n13890) );
  INV_X1 U11645 ( .A(n11005), .ZN(n10962) );
  OR2_X1 U11646 ( .A1(n9822), .A2(n18753), .ZN(n9821) );
  NAND2_X1 U11647 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U11648 ( .A1(n14049), .A2(n10715), .ZN(n10720) );
  NAND2_X1 U11649 ( .A1(n9899), .A2(n14897), .ZN(n9898) );
  NOR2_X1 U11650 ( .A1(n9900), .A2(n14912), .ZN(n9899) );
  INV_X1 U11651 ( .A(n13215), .ZN(n9900) );
  NAND2_X1 U11652 ( .A1(n15925), .A2(n10478), .ZN(n10587) );
  OR2_X1 U11653 ( .A1(n15933), .A2(n10894), .ZN(n10602) );
  INV_X1 U11654 ( .A(n15002), .ZN(n9937) );
  AND2_X1 U11655 ( .A1(n14016), .A2(n14088), .ZN(n9739) );
  NAND2_X1 U11656 ( .A1(n9895), .A2(n10966), .ZN(n9894) );
  INV_X1 U11657 ( .A(n15342), .ZN(n9895) );
  INV_X1 U11658 ( .A(n13565), .ZN(n9737) );
  INV_X1 U11659 ( .A(n14219), .ZN(n9949) );
  INV_X1 U11660 ( .A(n10000), .ZN(n9783) );
  NAND2_X1 U11661 ( .A1(n13990), .A2(n13991), .ZN(n10713) );
  INV_X1 U11662 ( .A(n13584), .ZN(n10743) );
  INV_X1 U11663 ( .A(n9772), .ZN(n9771) );
  INV_X1 U11664 ( .A(n9770), .ZN(n9769) );
  OAI21_X1 U11665 ( .B1(n9773), .B2(n9771), .A(n13907), .ZN(n9770) );
  XNOR2_X1 U11666 ( .A(n10698), .B(n10699), .ZN(n10701) );
  NOR2_X1 U11667 ( .A1(n13533), .A2(n9587), .ZN(n10227) );
  AOI22_X1 U11668 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U11669 ( .A1(n10051), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10052) );
  NAND2_X1 U11670 ( .A1(n10046), .A2(n10023), .ZN(n10053) );
  OAI21_X1 U11671 ( .B1(n10620), .B2(n10619), .A(n10618), .ZN(n10673) );
  AND2_X1 U11672 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15603), .ZN(
        n10619) );
  AND3_X1 U11673 ( .A1(n11056), .A2(n11055), .A3(n13778), .ZN(n10141) );
  NOR2_X1 U11674 ( .A1(n15492), .A2(n12342), .ZN(n15488) );
  NOR2_X1 U11675 ( .A1(n16651), .A2(n12117), .ZN(n12142) );
  NOR3_X1 U11676 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18562), .A3(
        n18419), .ZN(n12245) );
  NOR2_X1 U11677 ( .A1(n16651), .A2(n12116), .ZN(n12155) );
  NOR2_X1 U11678 ( .A1(n17312), .A2(n17310), .ZN(n9799) );
  XNOR2_X1 U11679 ( .A(n17129), .B(n12394), .ZN(n12215) );
  NOR2_X1 U11680 ( .A1(n17115), .A2(n12198), .ZN(n12197) );
  INV_X1 U11681 ( .A(n18383), .ZN(n12333) );
  NAND2_X1 U11682 ( .A1(n17528), .A2(n12229), .ZN(n12382) );
  AOI21_X1 U11683 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18437), .A(
        n12354), .ZN(n12366) );
  OAI211_X1 U11684 ( .C1(n12360), .C2(n12359), .A(n12361), .B(n12358), .ZN(
        n12367) );
  NAND2_X1 U11685 ( .A1(n12335), .A2(n12334), .ZN(n15491) );
  INV_X1 U11686 ( .A(n16277), .ZN(n15492) );
  OR2_X1 U11687 ( .A1(n20645), .A2(n12498), .ZN(n14405) );
  INV_X1 U11688 ( .A(n19740), .ZN(n14307) );
  AND2_X1 U11689 ( .A1(n20640), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12095) );
  OR2_X1 U11690 ( .A1(n9989), .A2(n14310), .ZN(n9988) );
  NOR2_X1 U11691 ( .A1(n12039), .A2(n14260), .ZN(n12040) );
  INV_X1 U11692 ( .A(n14514), .ZN(n9955) );
  OAI21_X1 U11693 ( .B1(n14514), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n13424), .ZN(n9953) );
  NOR2_X1 U11694 ( .A1(n9824), .A2(n14351), .ZN(n9823) );
  INV_X1 U11695 ( .A(n9825), .ZN(n9824) );
  NAND2_X1 U11696 ( .A1(n14154), .A2(n9827), .ZN(n14454) );
  NOR2_X1 U11697 ( .A1(n9828), .A2(n14452), .ZN(n9827) );
  INV_X1 U11698 ( .A(n9829), .ZN(n9828) );
  NAND2_X1 U11699 ( .A1(n14154), .A2(n9829), .ZN(n14460) );
  OR2_X1 U11700 ( .A1(n13704), .A2(n9838), .ZN(n15838) );
  AND2_X1 U11701 ( .A1(n13043), .A2(n14764), .ZN(n15848) );
  NAND2_X1 U11702 ( .A1(n12583), .A2(n12565), .ZN(n13413) );
  XNOR2_X1 U11703 ( .A(n11389), .B(n11387), .ZN(n11604) );
  AND2_X1 U11704 ( .A1(n13402), .A2(n13401), .ZN(n13684) );
  AND2_X1 U11705 ( .A1(n20445), .A2(n19965), .ZN(n20294) );
  NOR2_X1 U11706 ( .A1(n20288), .A2(n20119), .ZN(n20452) );
  OR2_X1 U11707 ( .A1(n13691), .A2(n11611), .ZN(n20422) );
  OR2_X1 U11708 ( .A1(n13690), .A2(n19961), .ZN(n20444) );
  NAND2_X1 U11709 ( .A1(n11611), .A2(n13691), .ZN(n20443) );
  NOR2_X1 U11710 ( .A1(n10593), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10594) );
  OR2_X1 U11711 ( .A1(n9808), .A2(n18656), .ZN(n9807) );
  OR2_X1 U11712 ( .A1(n18669), .A2(n9710), .ZN(n9806) );
  OR2_X1 U11713 ( .A1(n18669), .A2(n18670), .ZN(n9809) );
  NOR2_X1 U11714 ( .A1(n9928), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n9927) );
  AND2_X1 U11715 ( .A1(n10797), .A2(n10796), .ZN(n12477) );
  AND2_X1 U11716 ( .A1(n9981), .A2(n13514), .ZN(n9980) );
  NAND2_X1 U11717 ( .A1(n12866), .A2(n12865), .ZN(n12869) );
  INV_X1 U11718 ( .A(n16027), .ZN(n9890) );
  AND3_X1 U11719 ( .A1(n10886), .A2(n10885), .A3(n10884), .ZN(n13857) );
  AND2_X1 U11720 ( .A1(n10123), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13278) );
  AND2_X1 U11721 ( .A1(n10862), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U11722 ( .A1(n13100), .A2(n9812), .ZN(n9811) );
  NAND2_X1 U11723 ( .A1(n10793), .A2(n10792), .ZN(n13933) );
  AND2_X1 U11724 ( .A1(n15021), .A2(n10564), .ZN(n10565) );
  AND2_X1 U11725 ( .A1(n10563), .A2(n15038), .ZN(n10564) );
  INV_X1 U11726 ( .A(n16014), .ZN(n11094) );
  NAND2_X1 U11727 ( .A1(n10108), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10119) );
  NAND2_X1 U11728 ( .A1(n10117), .A2(n10023), .ZN(n10118) );
  NOR2_X1 U11729 ( .A1(n10107), .A2(n9868), .ZN(n10108) );
  OR2_X1 U11730 ( .A1(n13760), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9773) );
  NAND2_X1 U11731 ( .A1(n13760), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9772) );
  NOR2_X1 U11732 ( .A1(n19678), .A2(n18873), .ZN(n13832) );
  NAND2_X1 U11733 ( .A1(n13855), .A2(n18873), .ZN(n19199) );
  INV_X1 U11734 ( .A(n14039), .ZN(n19083) );
  INV_X1 U11735 ( .A(n19312), .ZN(n19358) );
  AND2_X1 U11736 ( .A1(n12628), .A2(n12627), .ZN(n19390) );
  AOI21_X2 U11737 ( .B1(n19729), .B2(n16049), .A(n13730), .ZN(n19392) );
  AND2_X1 U11738 ( .A1(n19678), .A2(n18873), .ZN(n19428) );
  AND2_X1 U11739 ( .A1(n19678), .A2(n19698), .ZN(n19449) );
  AND2_X1 U11740 ( .A1(n12626), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19517) );
  NOR2_X1 U11741 ( .A1(n15488), .A2(n17208), .ZN(n18383) );
  BUF_X1 U11742 ( .A(n12245), .Z(n15475) );
  NAND2_X1 U11743 ( .A1(n16119), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9798) );
  AND2_X1 U11744 ( .A1(n17479), .A2(n9795), .ZN(n17364) );
  AND2_X1 U11745 ( .A1(n9796), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9795) );
  NAND2_X1 U11746 ( .A1(n12197), .A2(n17111), .ZN(n16158) );
  NAND2_X1 U11747 ( .A1(n9840), .A2(n9843), .ZN(n17267) );
  AND2_X1 U11748 ( .A1(n17284), .A2(n9841), .ZN(n9840) );
  NOR2_X1 U11749 ( .A1(n9842), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9841) );
  INV_X1 U11750 ( .A(n9700), .ZN(n9842) );
  NAND2_X1 U11751 ( .A1(n12241), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9843) );
  AOI211_X1 U11752 ( .C1(n16917), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n12275), .B(n12274), .ZN(n12276) );
  NAND2_X1 U11753 ( .A1(n17568), .A2(n9848), .ZN(n17558) );
  AND2_X1 U11754 ( .A1(n9849), .A2(n12221), .ZN(n9848) );
  INV_X1 U11755 ( .A(n12217), .ZN(n12218) );
  NAND2_X1 U11756 ( .A1(n18411), .A2(n13178), .ZN(n18408) );
  AND2_X1 U11757 ( .A1(n14248), .A2(n14249), .ZN(n9835) );
  NAND2_X1 U11758 ( .A1(n12606), .A2(n12605), .ZN(n19825) );
  AND2_X1 U11759 ( .A1(n12606), .A2(n12595), .ZN(n19828) );
  INV_X1 U11760 ( .A(n14521), .ZN(n14250) );
  INV_X1 U11761 ( .A(n14482), .ZN(n14506) );
  AND2_X1 U11762 ( .A1(n13291), .A2(n13290), .ZN(n19854) );
  NAND2_X1 U11763 ( .A1(n13042), .A2(n15550), .ZN(n14761) );
  OR2_X1 U11764 ( .A1(n20207), .A2(n20327), .ZN(n20215) );
  NAND2_X1 U11765 ( .A1(n12978), .A2(n13154), .ZN(n18633) );
  NOR2_X1 U11766 ( .A1(n18704), .A2(n18691), .ZN(n18690) );
  NAND2_X1 U11767 ( .A1(n18922), .A2(n12958), .ZN(n14928) );
  OR2_X1 U11768 ( .A1(n13464), .A2(n12952), .ZN(n12953) );
  NOR2_X1 U11769 ( .A1(n15156), .A2(n15164), .ZN(n9885) );
  NAND2_X1 U11770 ( .A1(n14959), .A2(n15156), .ZN(n9883) );
  INV_X1 U11771 ( .A(n15167), .ZN(n9875) );
  INV_X1 U11772 ( .A(n19057), .ZN(n16001) );
  INV_X1 U11773 ( .A(n19049), .ZN(n15144) );
  OR2_X1 U11774 ( .A1(n18633), .A2(n9583), .ZN(n15995) );
  NAND2_X1 U11775 ( .A1(n19061), .A2(n19688), .ZN(n19057) );
  INV_X1 U11776 ( .A(n15995), .ZN(n19050) );
  NAND2_X1 U11777 ( .A1(n9757), .A2(n9755), .ZN(n14272) );
  AOI21_X1 U11778 ( .B1(n15890), .B2(n15354), .A(n11074), .ZN(n11099) );
  XNOR2_X1 U11779 ( .A(n12983), .B(n12982), .ZN(n13082) );
  INV_X1 U11780 ( .A(n15154), .ZN(n9888) );
  INV_X1 U11781 ( .A(n9790), .ZN(n9789) );
  AOI21_X1 U11782 ( .B1(n15090), .B2(n12475), .A(n15321), .ZN(n9790) );
  NAND2_X1 U11783 ( .A1(n10853), .A2(n11075), .ZN(n16008) );
  AND2_X1 U11784 ( .A1(n11075), .A2(n19707), .ZN(n16044) );
  NOR2_X2 U11785 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19681) );
  NAND2_X1 U11786 ( .A1(n17002), .A2(n17128), .ZN(n17001) );
  INV_X1 U11787 ( .A(n17008), .ZN(n17003) );
  NAND2_X1 U11788 ( .A1(n17003), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n17002) );
  NAND2_X1 U11789 ( .A1(n17077), .A2(n16992), .ZN(n17128) );
  INV_X1 U11790 ( .A(n17138), .ZN(n17126) );
  INV_X1 U11791 ( .A(n9852), .ZN(n12371) );
  OAI22_X1 U11792 ( .A1(n16154), .A2(n9705), .B1(n17669), .B2(n9850), .ZN(
        n16152) );
  OR2_X1 U11793 ( .A1(n17922), .A2(n16151), .ZN(n9850) );
  INV_X1 U11794 ( .A(n10380), .ZN(n9765) );
  AOI21_X1 U11795 ( .B1(n10654), .B2(n10621), .A(n10333), .ZN(n10342) );
  INV_X1 U11796 ( .A(n12941), .ZN(n12728) );
  INV_X1 U11797 ( .A(n12939), .ZN(n12724) );
  INV_X1 U11798 ( .A(n12940), .ZN(n12729) );
  INV_X1 U11799 ( .A(n12938), .ZN(n12725) );
  NAND2_X1 U11800 ( .A1(n9859), .A2(n9857), .ZN(n10279) );
  XNOR2_X1 U11801 ( .A(n10023), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10368) );
  OR2_X1 U11802 ( .A1(n11464), .A2(n11463), .ZN(n11494) );
  OR2_X1 U11803 ( .A1(n11443), .A2(n11442), .ZN(n11468) );
  OR3_X1 U11804 ( .A1(n11572), .A2(n11571), .A3(n12439), .ZN(n11573) );
  CLKBUF_X1 U11805 ( .A(n12729), .Z(n12905) );
  CLKBUF_X1 U11806 ( .A(n12728), .Z(n12902) );
  CLKBUF_X1 U11807 ( .A(n12725), .Z(n12907) );
  OR2_X1 U11808 ( .A1(n10466), .A2(n10465), .ZN(n10471) );
  OR2_X1 U11809 ( .A1(n10419), .A2(n10418), .ZN(n10422) );
  INV_X1 U11810 ( .A(n10144), .ZN(n10123) );
  OAI21_X1 U11811 ( .B1(n15002), .B2(n9938), .A(n10577), .ZN(n9942) );
  AND2_X1 U11812 ( .A1(n9943), .A2(n9699), .ZN(n9938) );
  AOI22_X1 U11813 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10054) );
  INV_X1 U11814 ( .A(n10071), .ZN(n10072) );
  AOI22_X1 U11815 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10019) );
  AND2_X1 U11816 ( .A1(n12365), .A2(n12364), .ZN(n12351) );
  NOR2_X1 U11817 ( .A1(n17955), .A2(n15512), .ZN(n12344) );
  NAND2_X1 U11818 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18562), .ZN(
        n12117) );
  AND2_X1 U11819 ( .A1(n9966), .A2(n14400), .ZN(n9965) );
  INV_X1 U11820 ( .A(n12059), .ZN(n12085) );
  NAND2_X1 U11821 ( .A1(n9972), .A2(n11791), .ZN(n9971) );
  INV_X1 U11822 ( .A(n14149), .ZN(n9972) );
  AND2_X1 U11823 ( .A1(n11756), .A2(n9986), .ZN(n9985) );
  OR2_X1 U11824 ( .A1(n14092), .A2(n14065), .ZN(n9986) );
  AND2_X1 U11825 ( .A1(n14103), .A2(n14095), .ZN(n11756) );
  NAND2_X1 U11826 ( .A1(n11681), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11696) );
  AND2_X1 U11827 ( .A1(n11646), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11656) );
  AND2_X1 U11828 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11591), .ZN(
        n11592) );
  AND2_X1 U11829 ( .A1(n11259), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11633) );
  NOR2_X1 U11830 ( .A1(n14362), .A2(n9826), .ZN(n9825) );
  INV_X1 U11831 ( .A(n14375), .ZN(n9826) );
  OR2_X1 U11832 ( .A1(n13703), .A2(n9839), .ZN(n9838) );
  INV_X1 U11833 ( .A(n13827), .ZN(n9839) );
  AND2_X1 U11834 ( .A1(n11500), .A2(n15756), .ZN(n9750) );
  NAND2_X1 U11835 ( .A1(n11500), .A2(n9754), .ZN(n9751) );
  INV_X1 U11836 ( .A(n11474), .ZN(n9754) );
  OR2_X1 U11837 ( .A1(n11484), .A2(n11483), .ZN(n11505) );
  NAND2_X1 U11838 ( .A1(n11488), .A2(n11487), .ZN(n11489) );
  INV_X1 U11839 ( .A(n11492), .ZN(n11488) );
  INV_X1 U11840 ( .A(n12586), .ZN(n12577) );
  OR2_X1 U11841 ( .A1(n11419), .A2(n11418), .ZN(n11467) );
  INV_X1 U11842 ( .A(n11575), .ZN(n11581) );
  OR2_X1 U11843 ( .A1(n11357), .A2(n11104), .ZN(n11406) );
  NAND2_X1 U11844 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11210) );
  AND2_X1 U11845 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11206) );
  AND2_X1 U11846 ( .A1(n10568), .A2(n9718), .ZN(n10588) );
  NOR2_X1 U11847 ( .A1(n10573), .A2(n9916), .ZN(n9915) );
  INV_X1 U11848 ( .A(n10569), .ZN(n9916) );
  OR2_X1 U11849 ( .A1(n10543), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U11850 ( .A1(n9920), .A2(n9919), .ZN(n10543) );
  NOR2_X1 U11851 ( .A1(n9921), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n9919) );
  INV_X1 U11852 ( .A(n10531), .ZN(n9920) );
  OR2_X1 U11853 ( .A1(n9923), .A2(n9922), .ZN(n9921) );
  INV_X1 U11854 ( .A(n10517), .ZN(n9922) );
  NAND2_X1 U11855 ( .A1(n9924), .A2(n10523), .ZN(n9923) );
  INV_X1 U11856 ( .A(n10530), .ZN(n9924) );
  NOR2_X1 U11857 ( .A1(n10508), .A2(n9918), .ZN(n9917) );
  INV_X1 U11858 ( .A(n10501), .ZN(n9918) );
  INV_X1 U11859 ( .A(n10482), .ZN(n9926) );
  NAND2_X1 U11860 ( .A1(n10630), .A2(n10339), .ZN(n10338) );
  OR2_X1 U11861 ( .A1(n12813), .A2(n12814), .ZN(n12815) );
  INV_X1 U11862 ( .A(n14869), .ZN(n9979) );
  INV_X1 U11863 ( .A(n14053), .ZN(n9904) );
  INV_X1 U11864 ( .A(n12863), .ZN(n13574) );
  AND2_X1 U11865 ( .A1(n10123), .A2(n10339), .ZN(n10136) );
  NOR2_X1 U11866 ( .A1(n9813), .A2(n15004), .ZN(n9812) );
  INV_X1 U11867 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U11868 ( .A1(n13118), .A2(n9810), .ZN(n13101) );
  INV_X1 U11869 ( .A(n9812), .ZN(n9810) );
  AND2_X1 U11870 ( .A1(n9715), .A2(n9815), .ZN(n9814) );
  NOR2_X1 U11871 ( .A1(n13126), .A2(n9816), .ZN(n9815) );
  OAI21_X1 U11872 ( .B1(n10178), .B2(n10023), .A(n10177), .ZN(n10734) );
  INV_X1 U11873 ( .A(n9912), .ZN(n10872) );
  AND2_X1 U11874 ( .A1(n13211), .A2(n14815), .ZN(n9742) );
  NAND2_X1 U11875 ( .A1(n12470), .A2(n9722), .ZN(n14971) );
  AND2_X1 U11876 ( .A1(n9681), .A2(n9775), .ZN(n9774) );
  NOR2_X1 U11877 ( .A1(n15303), .A2(n12480), .ZN(n9892) );
  NAND2_X1 U11878 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n9872) );
  NAND2_X1 U11879 ( .A1(n12940), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9870) );
  NAND2_X1 U11880 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n9869) );
  NOR2_X1 U11881 ( .A1(n9793), .A2(n9792), .ZN(n9791) );
  NAND2_X1 U11882 ( .A1(n9866), .A2(n10311), .ZN(n9780) );
  INV_X1 U11883 ( .A(n12954), .ZN(n10864) );
  AND2_X1 U11884 ( .A1(n19729), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12635) );
  INV_X1 U11885 ( .A(n10190), .ZN(n10193) );
  INV_X1 U11886 ( .A(n10191), .ZN(n10192) );
  AND3_X1 U11887 ( .A1(n11054), .A2(n10126), .A3(n10125), .ZN(n13717) );
  NOR2_X1 U11888 ( .A1(n12863), .A2(n13853), .ZN(n12632) );
  NAND2_X1 U11889 ( .A1(n13574), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12638) );
  INV_X1 U11890 ( .A(n9583), .ZN(n10208) );
  AOI22_X1 U11891 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10028) );
  AND2_X1 U11892 ( .A1(n10669), .A2(n10673), .ZN(n10670) );
  NAND2_X1 U11893 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12120) );
  INV_X1 U11894 ( .A(n12162), .ZN(n16840) );
  NAND2_X1 U11895 ( .A1(n18586), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12115) );
  NAND2_X1 U11896 ( .A1(n9799), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16300) );
  NOR2_X1 U11897 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18586), .ZN(
        n12364) );
  INV_X1 U11898 ( .A(n17965), .ZN(n15512) );
  AND2_X1 U11899 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18401) );
  NOR2_X1 U11900 ( .A1(n18581), .A2(n18461), .ZN(n17954) );
  OAI21_X1 U11901 ( .B1(n15488), .B2(n15487), .A(n18604), .ZN(n17142) );
  AND2_X1 U11902 ( .A1(n12492), .A2(n12493), .ZN(n14303) );
  AND2_X1 U11903 ( .A1(n11811), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U11904 ( .A1(n14405), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13863) );
  AND2_X1 U11905 ( .A1(n12539), .A2(n12538), .ZN(n14080) );
  AND2_X1 U11906 ( .A1(n11864), .A2(n11863), .ZN(n14443) );
  AND2_X1 U11907 ( .A1(n11255), .A2(n11254), .ZN(n14156) );
  NAND2_X1 U11908 ( .A1(n12003), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12004) );
  INV_X1 U11909 ( .A(n12000), .ZN(n12003) );
  OR2_X1 U11910 ( .A1(n11967), .A2(n14366), .ZN(n12000) );
  NAND2_X1 U11911 ( .A1(n11922), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11923) );
  OR2_X1 U11912 ( .A1(n11923), .A2(n14392), .ZN(n11963) );
  AND2_X1 U11913 ( .A1(n11880), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11881) );
  INV_X1 U11914 ( .A(n11904), .ZN(n11880) );
  NAND2_X1 U11915 ( .A1(n11881), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11921) );
  NOR2_X1 U11916 ( .A1(n11861), .A2(n14601), .ZN(n11862) );
  NAND2_X1 U11917 ( .A1(n11828), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11861) );
  INV_X1 U11918 ( .A(n14451), .ZN(n11845) );
  NAND2_X1 U11919 ( .A1(n11774), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11792) );
  INV_X1 U11920 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15664) );
  NOR2_X1 U11921 ( .A1(n11757), .A2(n14108), .ZN(n11774) );
  CLKBUF_X1 U11922 ( .A(n14071), .Z(n14072) );
  AND2_X1 U11923 ( .A1(n11712), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11713) );
  CLKBUF_X1 U11924 ( .A(n13967), .Z(n13968) );
  AND2_X1 U11925 ( .A1(n11656), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11681) );
  INV_X1 U11926 ( .A(n11663), .ZN(n11664) );
  CLKBUF_X1 U11927 ( .A(n13539), .Z(n13540) );
  OAI21_X1 U11928 ( .B1(n13690), .B2(n11541), .A(n11399), .ZN(n13590) );
  INV_X1 U11929 ( .A(n13502), .ZN(n11621) );
  NOR2_X1 U11930 ( .A1(n13424), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9954) );
  OAI21_X1 U11931 ( .B1(n14552), .B2(n14254), .A(n15702), .ZN(n14543) );
  NAND2_X1 U11932 ( .A1(n14373), .A2(n14375), .ZN(n14374) );
  NAND2_X1 U11933 ( .A1(n14373), .A2(n9825), .ZN(n14364) );
  INV_X1 U11934 ( .A(n14610), .ZN(n11532) );
  AND2_X1 U11935 ( .A1(n12557), .A2(n12556), .ZN(n14458) );
  OR2_X1 U11936 ( .A1(n14127), .A2(n14106), .ZN(n14105) );
  AND2_X1 U11937 ( .A1(n14081), .A2(n14080), .ZN(n14125) );
  NAND2_X1 U11938 ( .A1(n14125), .A2(n14124), .ZN(n14127) );
  CLKBUF_X1 U11939 ( .A(n14648), .Z(n14649) );
  INV_X1 U11940 ( .A(n15876), .ZN(n12527) );
  NOR2_X1 U11941 ( .A1(n13704), .A2(n13703), .ZN(n13828) );
  NAND2_X1 U11942 ( .A1(n12515), .A2(n12514), .ZN(n13556) );
  INV_X1 U11943 ( .A(n13504), .ZN(n12514) );
  INV_X1 U11944 ( .A(n13505), .ZN(n12515) );
  INV_X1 U11945 ( .A(n19940), .ZN(n15850) );
  AND2_X1 U11946 ( .A1(n13042), .A2(n13036), .ZN(n14763) );
  NAND2_X1 U11947 ( .A1(n13042), .A2(n13039), .ZN(n19936) );
  OAI21_X1 U11948 ( .B1(n11308), .B2(n11379), .A(n9746), .ZN(n9745) );
  NAND2_X1 U11949 ( .A1(n11308), .A2(n9749), .ZN(n9748) );
  OAI211_X1 U11950 ( .C1(n19964), .C2(n12104), .A(n11360), .B(n11359), .ZN(
        n11361) );
  OR2_X1 U11951 ( .A1(n11357), .A2(n11358), .ZN(n11360) );
  NAND2_X1 U11952 ( .A1(n11624), .A2(n13690), .ZN(n20076) );
  OR2_X1 U11953 ( .A1(n11624), .A2(n20230), .ZN(n20334) );
  NOR2_X1 U11954 ( .A1(n11187), .A2(n11186), .ZN(n11193) );
  AND3_X1 U11955 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20790), .A3(n19963), 
        .ZN(n20002) );
  INV_X1 U11956 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20416) );
  INV_X1 U11957 ( .A(n11324), .ZN(n11322) );
  AOI21_X1 U11958 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20416), .A(n20119), 
        .ZN(n20499) );
  INV_X1 U11959 ( .A(n20418), .ZN(n20493) );
  NAND2_X1 U11960 ( .A1(n11590), .A2(n11589), .ZN(n14301) );
  INV_X1 U11961 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20363) );
  INV_X1 U11962 ( .A(n15884), .ZN(n14789) );
  OR2_X1 U11963 ( .A1(n11049), .A2(n11048), .ZN(n16060) );
  NOR2_X1 U11964 ( .A1(n10599), .A2(n10598), .ZN(n10608) );
  NAND2_X1 U11965 ( .A1(n10611), .A2(n10595), .ZN(n10599) );
  NOR2_X1 U11966 ( .A1(n10611), .A2(n10586), .ZN(n15925) );
  OAI21_X1 U11967 ( .B1(n15945), .B2(n9717), .A(n9817), .ZN(n15937) );
  OR2_X1 U11968 ( .A1(n9808), .A2(n15938), .ZN(n9817) );
  OR2_X1 U11969 ( .A1(n15945), .A2(n15946), .ZN(n9818) );
  NAND2_X1 U11970 ( .A1(n10568), .A2(n9915), .ZN(n10585) );
  AND2_X1 U11971 ( .A1(n11015), .A2(n11014), .ZN(n14139) );
  INV_X1 U11972 ( .A(n10519), .ZN(n10520) );
  INV_X1 U11973 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13126) );
  AND2_X1 U11974 ( .A1(n10498), .A2(n9917), .ZN(n10537) );
  NAND2_X1 U11975 ( .A1(n10498), .A2(n10501), .ZN(n10509) );
  INV_X1 U11976 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13530) );
  INV_X1 U11977 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13638) );
  NOR2_X1 U11978 ( .A1(n13255), .A2(n13155), .ZN(n18847) );
  NAND2_X1 U11979 ( .A1(n14827), .A2(n9741), .ZN(n12985) );
  AND2_X1 U11980 ( .A1(n9742), .A2(n12921), .ZN(n9741) );
  AND2_X1 U11981 ( .A1(n13813), .A2(n13811), .ZN(n13812) );
  AND2_X1 U11982 ( .A1(n13819), .A2(n13613), .ZN(n13811) );
  XNOR2_X1 U11983 ( .A(n12839), .B(n12840), .ZN(n14825) );
  NAND2_X1 U11984 ( .A1(n14825), .A2(n14824), .ZN(n14823) );
  AND2_X1 U11985 ( .A1(n11029), .A2(n11028), .ZN(n14905) );
  NOR2_X1 U11986 ( .A1(n14842), .A2(n14844), .ZN(n14843) );
  NAND2_X1 U11987 ( .A1(n9978), .A2(n9976), .ZN(n9975) );
  NOR2_X1 U11988 ( .A1(n9976), .A2(n9978), .ZN(n9974) );
  NAND2_X1 U11989 ( .A1(n14084), .A2(n9697), .ZN(n14867) );
  NAND2_X1 U11990 ( .A1(n9983), .A2(n9706), .ZN(n14020) );
  AND2_X1 U11991 ( .A1(n12671), .A2(n13938), .ZN(n12672) );
  AND3_X1 U11992 ( .A1(n10912), .A2(n10911), .A3(n10910), .ZN(n16027) );
  AOI211_X1 U11993 ( .C1(n10860), .C2(n10962), .A(n10870), .B(n10859), .ZN(
        n13281) );
  INV_X1 U11994 ( .A(n12968), .ZN(n18892) );
  OAI21_X1 U11995 ( .B1(n12967), .B2(n12966), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12968) );
  NAND2_X1 U11996 ( .A1(n9820), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9819) );
  INV_X1 U11997 ( .A(n9821), .ZN(n9820) );
  NAND2_X1 U11998 ( .A1(n10720), .A2(n10719), .ZN(n15986) );
  NOR2_X1 U11999 ( .A1(n18821), .A2(n9802), .ZN(n9801) );
  NOR2_X1 U12000 ( .A1(n13135), .A2(n18821), .ZN(n13136) );
  INV_X1 U12001 ( .A(n14937), .ZN(n9761) );
  INV_X1 U12002 ( .A(n12981), .ZN(n9760) );
  AND2_X1 U12003 ( .A1(n9764), .A2(n14938), .ZN(n9763) );
  OR2_X1 U12004 ( .A1(n11073), .A2(n11072), .ZN(n11074) );
  OR2_X1 U12005 ( .A1(n13208), .A2(n10894), .ZN(n14951) );
  INV_X1 U12006 ( .A(n15912), .ZN(n10601) );
  INV_X1 U12007 ( .A(n14951), .ZN(n14949) );
  AOI21_X1 U12008 ( .B1(n15189), .B2(n10587), .A(n10604), .ZN(n14974) );
  AND2_X1 U12009 ( .A1(n10603), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14983) );
  NAND2_X1 U12010 ( .A1(n9937), .A2(n15014), .ZN(n9940) );
  INV_X1 U12011 ( .A(n15013), .ZN(n9941) );
  NOR2_X1 U12012 ( .A1(n9876), .A2(n9879), .ZN(n15000) );
  INV_X1 U12013 ( .A(n12470), .ZN(n9876) );
  AND2_X1 U12014 ( .A1(n11021), .A2(n11020), .ZN(n15231) );
  AND2_X1 U12015 ( .A1(n10809), .A2(n10808), .ZN(n14863) );
  AND2_X1 U12016 ( .A1(n11019), .A2(n11018), .ZN(n14926) );
  NAND2_X1 U12017 ( .A1(n12478), .A2(n9664), .ZN(n14876) );
  AND2_X1 U12018 ( .A1(n11013), .A2(n11012), .ZN(n15280) );
  NAND2_X1 U12019 ( .A1(n9892), .A2(n9891), .ZN(n15283) );
  INV_X1 U12020 ( .A(n15280), .ZN(n9891) );
  INV_X1 U12021 ( .A(n9892), .ZN(n15281) );
  AND2_X1 U12022 ( .A1(n12478), .A2(n14016), .ZN(n14089) );
  AND2_X1 U12023 ( .A1(n9777), .A2(n9775), .ZN(n12488) );
  AND3_X1 U12024 ( .A1(n10979), .A2(n10978), .A3(n10977), .ZN(n15342) );
  NOR2_X1 U12025 ( .A1(n9736), .A2(n13608), .ZN(n9733) );
  INV_X1 U12026 ( .A(n16007), .ZN(n9889) );
  NOR2_X1 U12027 ( .A1(n13564), .A2(n13565), .ZN(n13659) );
  NAND2_X1 U12028 ( .A1(n9950), .A2(n9948), .ZN(n15141) );
  AND2_X1 U12029 ( .A1(n18813), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14219) );
  NAND3_X1 U12030 ( .A1(n10738), .A2(n9740), .A3(n9676), .ZN(n13653) );
  INV_X1 U12031 ( .A(n13632), .ZN(n9740) );
  NOR2_X2 U12032 ( .A1(n13653), .A2(n13652), .ZN(n14225) );
  AOI21_X1 U12033 ( .B1(n9769), .B2(n9771), .A(n9709), .ZN(n9766) );
  INV_X1 U12034 ( .A(n10701), .ZN(n10702) );
  NAND2_X1 U12035 ( .A1(n9780), .A2(n10698), .ZN(n13759) );
  INV_X1 U12036 ( .A(n9861), .ZN(n10157) );
  OAI211_X1 U12037 ( .C1(n10835), .C2(n10156), .A(n9863), .B(n9862), .ZN(n9861) );
  NOR2_X1 U12038 ( .A1(n11071), .A2(n9707), .ZN(n9862) );
  NAND2_X1 U12039 ( .A1(n12619), .A2(n19697), .ZN(n12636) );
  INV_X1 U12040 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13714) );
  NAND2_X1 U12041 ( .A1(n9584), .A2(n10121), .ZN(n10661) );
  INV_X1 U12042 ( .A(n13832), .ZN(n19172) );
  NAND2_X1 U12043 ( .A1(n19171), .A2(n19692), .ZN(n19670) );
  OR2_X1 U12044 ( .A1(n19171), .A2(n19689), .ZN(n19312) );
  NAND2_X1 U12045 ( .A1(n10088), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10089) );
  NAND2_X1 U12046 ( .A1(n10083), .A2(n10023), .ZN(n10090) );
  NOR2_X2 U12047 ( .A1(n18892), .A2(n13734), .ZN(n13795) );
  NOR2_X2 U12048 ( .A1(n18891), .A2(n13734), .ZN(n13796) );
  NAND2_X1 U12049 ( .A1(n9856), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9855) );
  NAND2_X1 U12050 ( .A1(n9854), .A2(n10023), .ZN(n9853) );
  INV_X1 U12051 ( .A(n13750), .ZN(n13799) );
  INV_X1 U12052 ( .A(n13796), .ZN(n13798) );
  AND2_X1 U12053 ( .A1(n10384), .A2(n19505), .ZN(n19512) );
  INV_X1 U12054 ( .A(n18472), .ZN(n18604) );
  AND2_X1 U12055 ( .A1(n16333), .A2(n9589), .ZN(n16323) );
  INV_X1 U12056 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16337) );
  NAND2_X1 U12057 ( .A1(n9794), .A2(n16310), .ZN(n16369) );
  AND2_X1 U12058 ( .A1(n16400), .A2(n9589), .ZN(n16393) );
  AND2_X1 U12059 ( .A1(n16423), .A2(n9589), .ZN(n16415) );
  NOR2_X1 U12060 ( .A1(n17329), .A2(n16415), .ZN(n16414) );
  OR2_X1 U12061 ( .A1(n16425), .A2(n17344), .ZN(n16423) );
  NOR2_X1 U12062 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16603), .ZN(n16588) );
  INV_X1 U12063 ( .A(n18620), .ZN(n13180) );
  NOR2_X1 U12064 ( .A1(n16955), .A2(n16964), .ZN(n16959) );
  NOR2_X1 U12065 ( .A1(n12171), .A2(n12170), .ZN(n12175) );
  INV_X1 U12066 ( .A(n12169), .ZN(n12170) );
  NOR2_X1 U12067 ( .A1(n17143), .A2(n17142), .ZN(n17173) );
  NOR2_X1 U12068 ( .A1(n18452), .A2(n15508), .ZN(n17207) );
  NOR2_X2 U12069 ( .A1(n16337), .A2(n16120), .ZN(n16119) );
  AND2_X1 U12070 ( .A1(n17618), .A2(n15524), .ZN(n15506) );
  NOR2_X2 U12071 ( .A1(n16308), .A2(n16309), .ZN(n16307) );
  INV_X1 U12072 ( .A(n9799), .ZN(n17288) );
  INV_X1 U12073 ( .A(n16300), .ZN(n17280) );
  AND2_X1 U12074 ( .A1(n9660), .A2(n17408), .ZN(n9796) );
  AND2_X1 U12075 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17567) );
  NOR2_X1 U12076 ( .A1(n18394), .A2(n18452), .ZN(n12373) );
  INV_X1 U12077 ( .A(n17882), .ZN(n12363) );
  OR2_X1 U12078 ( .A1(n17402), .A2(n17294), .ZN(n12238) );
  NOR2_X1 U12079 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17338), .ZN(
        n17332) );
  NOR2_X1 U12080 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17388), .ZN(
        n17387) );
  NOR2_X1 U12081 ( .A1(n17487), .A2(n17846), .ZN(n17808) );
  NAND2_X1 U12082 ( .A1(n12409), .A2(n17851), .ZN(n17805) );
  INV_X1 U12083 ( .A(n17400), .ZN(n9846) );
  INV_X1 U12084 ( .A(n12228), .ZN(n12226) );
  NAND2_X1 U12085 ( .A1(n17529), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17528) );
  INV_X1 U12086 ( .A(n18391), .ZN(n16156) );
  NOR2_X1 U12087 ( .A1(n18402), .A2(n15489), .ZN(n13178) );
  NAND2_X1 U12088 ( .A1(n18586), .A2(n18580), .ZN(n16651) );
  AND2_X1 U12089 ( .A1(n18383), .A2(n9731), .ZN(n18411) );
  NAND2_X1 U12090 ( .A1(n12332), .A2(n12340), .ZN(n9731) );
  INV_X1 U12091 ( .A(n18401), .ZN(n18419) );
  NOR2_X1 U12092 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17954), .ZN(n18290) );
  NOR2_X1 U12093 ( .A1(n12329), .A2(n12328), .ZN(n17969) );
  INV_X1 U12094 ( .A(n15509), .ZN(n17977) );
  NOR2_X2 U12095 ( .A1(n12299), .A2(n12298), .ZN(n17983) );
  NOR2_X1 U12096 ( .A1(n12319), .A2(n12318), .ZN(n17989) );
  INV_X1 U12097 ( .A(n18290), .ZN(n18147) );
  NAND2_X1 U12098 ( .A1(n15583), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19740) );
  NAND2_X1 U12099 ( .A1(n14292), .A2(n14293), .ZN(n20645) );
  INV_X1 U12100 ( .A(n19820), .ZN(n19775) );
  NAND2_X1 U12101 ( .A1(n14405), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19769) );
  INV_X1 U12102 ( .A(n19825), .ZN(n19797) );
  INV_X1 U12103 ( .A(n19769), .ZN(n19823) );
  NAND2_X1 U12104 ( .A1(n12606), .A2(n12604), .ZN(n15677) );
  NAND2_X1 U12105 ( .A1(n12592), .A2(n12591), .ZN(n12594) );
  OR2_X1 U12106 ( .A1(n14334), .A2(n14333), .ZN(n14692) );
  NAND2_X1 U12107 ( .A1(n19851), .A2(n13095), .ZN(n14465) );
  INV_X1 U12108 ( .A(n19851), .ZN(n14446) );
  INV_X1 U12109 ( .A(n14484), .ZN(n14507) );
  NAND2_X1 U12110 ( .A1(n13399), .A2(n14307), .ZN(n12449) );
  OR2_X1 U12111 ( .A1(n14506), .A2(n13357), .ZN(n14137) );
  XNOR2_X1 U12112 ( .A(n12103), .B(n12607), .ZN(n13866) );
  INV_X1 U12113 ( .A(n12097), .ZN(n12098) );
  INV_X1 U12114 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14601) );
  OR2_X1 U12115 ( .A1(n15564), .A2(n19740), .ZN(n19746) );
  NOR2_X2 U12116 ( .A1(n19908), .A2(n13471), .ZN(n15731) );
  INV_X1 U12117 ( .A(n19908), .ZN(n14653) );
  INV_X1 U12118 ( .A(n19911), .ZN(n19960) );
  INV_X1 U12119 ( .A(n19746), .ZN(n19912) );
  OAI211_X1 U12120 ( .C1(n9677), .C2(n9953), .A(n9952), .B(n9951), .ZN(n13018)
         );
  NAND2_X1 U12121 ( .A1(n9955), .A2(n9954), .ZN(n9951) );
  NAND2_X1 U12122 ( .A1(n9677), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9952) );
  NOR2_X1 U12123 ( .A1(n15872), .A2(n13063), .ZN(n14734) );
  OAI21_X1 U12124 ( .B1(n19950), .B2(n19936), .A(n15853), .ZN(n19928) );
  NOR2_X1 U12125 ( .A1(n15850), .A2(n13493), .ZN(n19935) );
  OR2_X1 U12126 ( .A1(n13059), .A2(n14763), .ZN(n19940) );
  NOR2_X1 U12127 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13059), .ZN(
        n13493) );
  AND2_X1 U12128 ( .A1(n13042), .A2(n13017), .ZN(n19929) );
  AND2_X1 U12129 ( .A1(n14737), .A2(n19936), .ZN(n13436) );
  INV_X1 U12130 ( .A(n19929), .ZN(n19946) );
  INV_X1 U12131 ( .A(n11386), .ZN(n11605) );
  OAI21_X1 U12132 ( .B1(n13689), .B2(n15888), .A(n20119), .ZN(n19956) );
  AND2_X1 U12133 ( .A1(n13040), .A2(n13041), .ZN(n15550) );
  NOR2_X1 U12134 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14800) );
  OR2_X1 U12135 ( .A1(n20076), .A2(n20327), .ZN(n20100) );
  OR2_X1 U12136 ( .A1(n20076), .A2(n20443), .ZN(n20106) );
  OAI211_X1 U12137 ( .C1(n20255), .C2(n20371), .A(n20294), .B(n20240), .ZN(
        n20258) );
  INV_X1 U12138 ( .A(n20215), .ZN(n20257) );
  OR2_X1 U12139 ( .A1(n20334), .A2(n20443), .ZN(n20320) );
  OAI211_X1 U12140 ( .C1(n20297), .C2(n20296), .A(n20295), .B(n20294), .ZN(
        n20323) );
  INV_X1 U12141 ( .A(n20320), .ZN(n20353) );
  OAI211_X1 U12142 ( .C1(n20483), .C2(n20453), .A(n20452), .B(n20451), .ZN(
        n20486) );
  INV_X1 U12143 ( .A(n20364), .ZN(n20495) );
  INV_X1 U12144 ( .A(n20377), .ZN(n20506) );
  INV_X1 U12145 ( .A(n20387), .ZN(n20518) );
  INV_X1 U12146 ( .A(n20392), .ZN(n20524) );
  INV_X1 U12147 ( .A(n20402), .ZN(n20536) );
  INV_X1 U12148 ( .A(n19966), .ZN(n20547) );
  NAND2_X1 U12149 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n14301), .ZN(n20623) );
  INV_X1 U12150 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20553) );
  INV_X2 U12151 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20640) );
  NAND2_X1 U12152 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20647) );
  INV_X1 U12153 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n18626) );
  OR2_X1 U12154 ( .A1(n14277), .A2(n18858), .ZN(n13166) );
  NOR2_X1 U12155 ( .A1(n18810), .A2(n15914), .ZN(n15902) );
  NOR2_X1 U12156 ( .A1(n15937), .A2(n18810), .ZN(n15923) );
  NOR2_X1 U12157 ( .A1(n18810), .A2(n13190), .ZN(n15945) );
  INV_X1 U12158 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15004) );
  AND2_X1 U12159 ( .A1(n9806), .A2(n9712), .ZN(n15540) );
  AND2_X1 U12160 ( .A1(n9809), .A2(n9808), .ZN(n18655) );
  NAND2_X1 U12161 ( .A1(n9806), .A2(n9807), .ZN(n18654) );
  AND2_X1 U12162 ( .A1(n9685), .A2(n13108), .ZN(n18704) );
  NOR2_X1 U12163 ( .A1(n13142), .A2(n18733), .ZN(n18720) );
  INV_X1 U12164 ( .A(n18871), .ZN(n18842) );
  AND2_X1 U12165 ( .A1(n19724), .A2(n16050), .ZN(n18859) );
  NOR2_X1 U12166 ( .A1(n18781), .A2(n18779), .ZN(n18772) );
  NAND2_X1 U12167 ( .A1(n10482), .A2(n9927), .ZN(n10493) );
  NOR2_X1 U12168 ( .A1(n18826), .A2(n18824), .ZN(n18809) );
  OR3_X1 U12169 ( .A1(n19724), .A2(n18838), .A3(n13153), .ZN(n18845) );
  INV_X1 U12170 ( .A(n18845), .ZN(n18862) );
  INV_X1 U12171 ( .A(n19678), .ZN(n13855) );
  INV_X1 U12172 ( .A(n19582), .ZN(n18838) );
  INV_X1 U12173 ( .A(n18868), .ZN(n18858) );
  AOI22_X1 U12174 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19729), .ZN(n18878) );
  NOR2_X1 U12175 ( .A1(n12646), .A2(n9982), .ZN(n9981) );
  INV_X1 U12176 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U12177 ( .A1(n14840), .A2(n13800), .ZN(n14880) );
  NAND2_X1 U12178 ( .A1(n13462), .A2(n13454), .ZN(n12919) );
  INV_X1 U12179 ( .A(n15910), .ZN(n15155) );
  NOR2_X1 U12180 ( .A1(n14820), .A2(n14819), .ZN(n14818) );
  NAND2_X1 U12181 ( .A1(n9962), .A2(n12869), .ZN(n14820) );
  AND2_X1 U12182 ( .A1(n13275), .A2(n18891), .ZN(n18884) );
  AND2_X1 U12183 ( .A1(n14227), .A2(n9701), .ZN(n15386) );
  OAI21_X1 U12184 ( .B1(n13622), .B2(n9698), .A(n10891), .ZN(n14054) );
  NOR2_X1 U12185 ( .A1(n13622), .A2(n13857), .ZN(n13995) );
  NOR2_X1 U12186 ( .A1(n18890), .A2(n18932), .ZN(n18920) );
  NAND2_X1 U12187 ( .A1(n13276), .A2(n14928), .ZN(n18913) );
  AND2_X1 U12188 ( .A1(n18922), .A2(n12957), .ZN(n18932) );
  NOR2_X1 U12189 ( .A1(n15405), .A2(n13279), .ZN(n18873) );
  INV_X1 U12190 ( .A(n18936), .ZN(n18890) );
  INV_X1 U12191 ( .A(n18922), .ZN(n18931) );
  INV_X1 U12192 ( .A(n18913), .ZN(n18940) );
  NOR2_X1 U12193 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16095), .ZN(n19008) );
  INV_X1 U12194 ( .A(n18943), .ZN(n19043) );
  NAND2_X1 U12195 ( .A1(n13256), .A2(n19586), .ZN(n19046) );
  CLKBUF_X1 U12196 ( .A(n19016), .Z(n19044) );
  INV_X1 U12197 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18753) );
  INV_X1 U12198 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18799) );
  INV_X1 U12199 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20762) );
  NAND2_X1 U12200 ( .A1(n10738), .A2(n10737), .ZN(n13585) );
  NAND2_X1 U12201 ( .A1(n18633), .A2(n12988), .ZN(n19061) );
  AND2_X1 U12202 ( .A1(n19061), .A2(n13236), .ZN(n19049) );
  INV_X1 U12203 ( .A(n19061), .ZN(n15105) );
  AND2_X1 U12204 ( .A1(n15200), .A2(n11093), .ZN(n15174) );
  INV_X1 U12205 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15173) );
  NAND2_X1 U12206 ( .A1(n15013), .A2(n15014), .ZN(n9945) );
  NAND2_X1 U12207 ( .A1(n13762), .A2(n9773), .ZN(n9768) );
  INV_X1 U12208 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16047) );
  INV_X1 U12209 ( .A(n16008), .ZN(n16038) );
  INV_X1 U12210 ( .A(n18873), .ZN(n19698) );
  INV_X1 U12211 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19687) );
  INV_X1 U12212 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19680) );
  INV_X1 U12213 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15603) );
  NAND2_X1 U12214 ( .A1(n13837), .A2(n13836), .ZN(n19076) );
  INV_X1 U12215 ( .A(n19095), .ZN(n19104) );
  OAI21_X1 U12216 ( .B1(n19102), .B2(n19697), .A(n19086), .ZN(n19105) );
  INV_X1 U12217 ( .A(n19126), .ZN(n19108) );
  NAND2_X1 U12218 ( .A1(n9860), .A2(n19697), .ZN(n19136) );
  NOR2_X1 U12219 ( .A1(n19670), .A2(n19172), .ZN(n19274) );
  OAI21_X1 U12220 ( .B1(n19305), .B2(n19283), .A(n19515), .ZN(n19308) );
  NAND2_X1 U12221 ( .A1(n19449), .A2(n19083), .ZN(n19311) );
  AND2_X1 U12222 ( .A1(n19428), .A2(n19083), .ZN(n19343) );
  INV_X1 U12223 ( .A(n19327), .ZN(n19344) );
  OAI22_X1 U12224 ( .A1(n16191), .A2(n13798), .B1(n17038), .B2(n13797), .ZN(
        n19408) );
  OAI21_X1 U12225 ( .B1(n19413), .B2(n19697), .A(n19395), .ZN(n19416) );
  INV_X1 U12226 ( .A(n19411), .ZN(n19415) );
  INV_X1 U12227 ( .A(n19437), .ZN(n19445) );
  INV_X1 U12228 ( .A(n19522), .ZN(n19465) );
  INV_X1 U12229 ( .A(n19530), .ZN(n19470) );
  INV_X1 U12230 ( .A(n19529), .ZN(n19469) );
  INV_X1 U12231 ( .A(n19542), .ZN(n19474) );
  INV_X1 U12232 ( .A(n19536), .ZN(n19473) );
  INV_X1 U12233 ( .A(n19544), .ZN(n19481) );
  INV_X1 U12234 ( .A(n19551), .ZN(n19488) );
  INV_X1 U12235 ( .A(n19550), .ZN(n19486) );
  INV_X1 U12236 ( .A(n19560), .ZN(n19493) );
  INV_X1 U12237 ( .A(n19559), .ZN(n19492) );
  OAI21_X1 U12238 ( .B1(n19461), .B2(n19460), .A(n19459), .ZN(n19499) );
  AND2_X1 U12239 ( .A1(n19428), .A2(n19427), .ZN(n19498) );
  INV_X1 U12240 ( .A(n19485), .ZN(n19546) );
  INV_X1 U12241 ( .A(n19576), .ZN(n19554) );
  INV_X1 U12242 ( .A(n19412), .ZN(n19562) );
  INV_X1 U12243 ( .A(n19408), .ZN(n19565) );
  NAND2_X1 U12244 ( .A1(n19428), .A2(n19673), .ZN(n19576) );
  AND2_X1 U12245 ( .A1(n19449), .A2(n19673), .ZN(n19572) );
  INV_X1 U12246 ( .A(n18631), .ZN(n19720) );
  NOR3_X1 U12247 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19597), .A3(n19600), 
        .ZN(n19730) );
  AOI21_X1 U12248 ( .B1(n18383), .B2(n18408), .A(n17143), .ZN(n18620) );
  INV_X1 U12249 ( .A(n15493), .ZN(n17208) );
  INV_X1 U12250 ( .A(n17207), .ZN(n17143) );
  INV_X1 U12251 ( .A(n12373), .ZN(n16279) );
  NOR2_X1 U12252 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16408), .ZN(n16391) );
  NOR2_X1 U12253 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16436), .ZN(n16431) );
  AND2_X1 U12254 ( .A1(n9589), .A2(n9797), .ZN(n13177) );
  NAND2_X1 U12255 ( .A1(n13176), .A2(n16466), .ZN(n9797) );
  NOR2_X1 U12256 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16481), .ZN(n16469) );
  NOR2_X1 U12257 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16539), .ZN(n16538) );
  NOR2_X1 U12258 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16579), .ZN(n16560) );
  NOR2_X2 U12259 ( .A1(n18555), .A2(n16653), .ZN(n16610) );
  INV_X1 U12260 ( .A(n16659), .ZN(n16648) );
  INV_X1 U12261 ( .A(n16669), .ZN(n16653) );
  INV_X1 U12262 ( .A(n16665), .ZN(n16654) );
  NAND4_X1 U12263 ( .A1(n17930), .A2(n13180), .A3(n18460), .A4(n18450), .ZN(
        n16669) );
  AND2_X1 U12264 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16743), .ZN(n16728) );
  NOR2_X1 U12265 ( .A1(n16730), .A2(n16729), .ZN(n16743) );
  NOR2_X1 U12266 ( .A1(n15409), .A2(n16766), .ZN(n16754) );
  INV_X1 U12267 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U12268 ( .A1(n17020), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n17017) );
  NOR2_X1 U12269 ( .A1(n9673), .A2(n17154), .ZN(n17020) );
  NAND2_X1 U12270 ( .A1(n9730), .A2(n9728), .ZN(n17031) );
  NOR2_X1 U12271 ( .A1(n17036), .A2(n9729), .ZN(n9728) );
  INV_X1 U12272 ( .A(n17069), .ZN(n9730) );
  NAND2_X1 U12273 ( .A1(n17073), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17069) );
  NOR2_X1 U12274 ( .A1(n12137), .A2(n12136), .ZN(n17115) );
  NOR2_X1 U12275 ( .A1(n12148), .A2(n12147), .ZN(n17123) );
  NOR3_X1 U12276 ( .A1(n17200), .A2(n17137), .A3(n17126), .ZN(n17133) );
  NAND2_X1 U12277 ( .A1(n18423), .A2(n17095), .ZN(n17134) );
  INV_X1 U12278 ( .A(n12394), .ZN(n17141) );
  OAI21_X1 U12279 ( .B1(n15606), .B2(n15605), .A(n18603), .ZN(n17135) );
  INV_X1 U12280 ( .A(n17135), .ZN(n16992) );
  INV_X1 U12281 ( .A(n17134), .ZN(n17136) );
  NOR2_X1 U12282 ( .A1(n18423), .A2(n17135), .ZN(n17079) );
  CLKBUF_X1 U12283 ( .A(n17190), .Z(n17202) );
  NOR2_X1 U12286 ( .A1(n17245), .A2(n17960), .ZN(n17253) );
  NAND2_X1 U12287 ( .A1(n17325), .A2(n10008), .ZN(n17312) );
  NAND2_X1 U12288 ( .A1(n17364), .A2(n10007), .ZN(n17351) );
  NAND2_X1 U12289 ( .A1(n17479), .A2(n9796), .ZN(n17390) );
  NOR2_X2 U12290 ( .A1(n18566), .A2(n17604), .ZN(n17465) );
  OR2_X1 U12291 ( .A1(n18287), .A2(n18147), .ZN(n17980) );
  NAND2_X1 U12292 ( .A1(n17479), .A2(n10009), .ZN(n17429) );
  NOR2_X1 U12293 ( .A1(n16527), .A2(n16537), .ZN(n12374) );
  NOR2_X2 U12294 ( .A1(n17108), .A2(n17612), .ZN(n17519) );
  INV_X1 U12295 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20724) );
  NAND3_X1 U12296 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17553) );
  INV_X2 U12297 ( .A(n17980), .ZN(n18329) );
  INV_X1 U12298 ( .A(n17603), .ZN(n17593) );
  NAND2_X1 U12299 ( .A1(n17609), .A2(n17566), .ZN(n17604) );
  NAND2_X1 U12300 ( .A1(n17354), .A2(n17450), .ZN(n17603) );
  OAI21_X2 U12301 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18602), .A(n16279), 
        .ZN(n17609) );
  INV_X1 U12302 ( .A(n17601), .ZN(n17613) );
  INV_X1 U12303 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18566) );
  NAND2_X1 U12304 ( .A1(n9843), .A2(n9844), .ZN(n17269) );
  AND2_X1 U12305 ( .A1(n17284), .A2(n9700), .ZN(n9844) );
  INV_X1 U12306 ( .A(n17681), .ZN(n17752) );
  INV_X1 U12307 ( .A(n17807), .ZN(n17839) );
  NOR2_X1 U12308 ( .A1(n17400), .A2(n12230), .ZN(n17840) );
  OAI21_X2 U12309 ( .B1(n15520), .B2(n15519), .A(n18603), .ZN(n17922) );
  NAND2_X1 U12310 ( .A1(n16156), .A2(n17928), .ZN(n17934) );
  INV_X1 U12311 ( .A(n17921), .ZN(n17936) );
  NOR2_X1 U12312 ( .A1(n13178), .A2(n18413), .ZN(n18424) );
  INV_X1 U12313 ( .A(n17922), .ZN(n17928) );
  INV_X1 U12314 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18437) );
  AND2_X2 U12315 ( .A1(n12460), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19957)
         );
  OAI21_X1 U12317 ( .B1(n14659), .B2(n19793), .A(n9832), .ZN(P1_U2810) );
  INV_X1 U12318 ( .A(n9833), .ZN(n9832) );
  NOR2_X1 U12319 ( .A1(n14247), .A2(n9835), .ZN(n9834) );
  OAI21_X1 U12320 ( .B1(n15906), .B2(n14873), .A(n12922), .ZN(n12923) );
  AOI21_X1 U12321 ( .B1(n14272), .B2(n19050), .A(n14270), .ZN(n9732) );
  NAND2_X1 U12322 ( .A1(n13082), .A2(n19050), .ZN(n12995) );
  OAI211_X1 U12323 ( .C1(n15171), .C2(n15995), .A(n9874), .B(n9873), .ZN(
        P2_U2986) );
  NAND2_X1 U12324 ( .A1(n9875), .A2(n19052), .ZN(n9874) );
  INV_X1 U12325 ( .A(n11100), .ZN(n11101) );
  INV_X1 U12326 ( .A(n13080), .ZN(n13085) );
  NOR2_X1 U12327 ( .A1(n15910), .A2(n16036), .ZN(n9881) );
  NAND2_X1 U12328 ( .A1(n9882), .A2(n9886), .ZN(n9880) );
  NAND2_X1 U12329 ( .A1(n9786), .A2(n9785), .ZN(P2_U3029) );
  NOR2_X1 U12330 ( .A1(n13344), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9787) );
  INV_X1 U12331 ( .A(n9788), .ZN(n15312) );
  AOI21_X1 U12332 ( .B1(n17001), .B2(n9720), .A(n9727), .ZN(n9726) );
  NOR2_X1 U12333 ( .A1(n12414), .A2(n9999), .ZN(n12415) );
  NOR2_X1 U12334 ( .A1(n12115), .A2(n12117), .ZN(n12250) );
  NOR2_X2 U12335 ( .A1(n12118), .A2(n12119), .ZN(n12177) );
  NAND2_X1 U12336 ( .A1(n9625), .A2(n14603), .ZN(n14605) );
  INV_X1 U12337 ( .A(n11037), .ZN(n11041) );
  INV_X1 U12338 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10017) );
  NAND2_X1 U12339 ( .A1(n14442), .A2(n14443), .ZN(n14434) );
  OR3_X1 U12340 ( .A1(n14335), .A2(n9987), .A3(n9988), .ZN(n9657) );
  NAND2_X1 U12341 ( .A1(n14442), .A2(n9965), .ZN(n14389) );
  OR2_X1 U12342 ( .A1(n13131), .A2(n9822), .ZN(n9658) );
  NOR2_X1 U12343 ( .A1(n14070), .A2(n9971), .ZN(n14148) );
  NAND2_X1 U12344 ( .A1(n13127), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13125) );
  INV_X1 U12345 ( .A(n12980), .ZN(n9764) );
  AND2_X1 U12346 ( .A1(n14603), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9659) );
  AND2_X1 U12347 ( .A1(n10009), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9660) );
  AND2_X1 U12348 ( .A1(n9701), .A2(n15387), .ZN(n9661) );
  NOR2_X1 U12349 ( .A1(n13198), .A2(n9719), .ZN(n13214) );
  NOR2_X1 U12350 ( .A1(n9838), .A2(n15837), .ZN(n9662) );
  OAI22_X2 U12351 ( .A1(n14269), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19729), 
        .B2(n13103), .ZN(n13108) );
  AND2_X1 U12352 ( .A1(n9983), .A2(n9984), .ZN(n13649) );
  NOR2_X1 U12353 ( .A1(n13120), .A2(n18659), .ZN(n13119) );
  NOR2_X1 U12354 ( .A1(n13118), .A2(n15004), .ZN(n13116) );
  AND2_X1 U12355 ( .A1(n13127), .A2(n9713), .ZN(n13121) );
  AND2_X1 U12356 ( .A1(n9697), .A2(n9977), .ZN(n9663) );
  NOR2_X1 U12357 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11071) );
  AND2_X1 U12358 ( .A1(n9739), .A2(n9738), .ZN(n9664) );
  OR2_X1 U12359 ( .A1(n15359), .A2(n15360), .ZN(n9665) );
  AND2_X1 U12360 ( .A1(n9818), .A2(n9808), .ZN(n9666) );
  NAND2_X1 U12361 ( .A1(n14225), .A2(n14224), .ZN(n13509) );
  AND2_X1 U12362 ( .A1(n10726), .A2(n9724), .ZN(n9667) );
  AND2_X2 U12363 ( .A1(n12941), .A2(n10023), .ZN(n10361) );
  INV_X2 U12364 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U12365 ( .A1(n12470), .A2(n10726), .ZN(n15010) );
  AND2_X1 U12366 ( .A1(n10033), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10296) );
  AND2_X2 U12367 ( .A1(n12939), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10301) );
  NAND2_X1 U12368 ( .A1(n12470), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9669) );
  NAND2_X1 U12369 ( .A1(n10499), .A2(n10591), .ZN(n10498) );
  INV_X1 U12370 ( .A(n11379), .ZN(n9749) );
  INV_X1 U12371 ( .A(n9778), .ZN(n14973) );
  OR2_X1 U12372 ( .A1(n13118), .A2(n9811), .ZN(n9672) );
  INV_X1 U12373 ( .A(n17518), .ZN(n9847) );
  NAND2_X1 U12374 ( .A1(n13967), .A2(n14065), .ZN(n14064) );
  NOR2_X1 U12375 ( .A1(n10531), .A2(n9921), .ZN(n10542) );
  AND2_X1 U12376 ( .A1(n12951), .A2(n10332), .ZN(n10158) );
  NOR2_X1 U12377 ( .A1(n13137), .A2(n20762), .ZN(n13138) );
  NOR2_X1 U12378 ( .A1(n13133), .A2(n18799), .ZN(n13134) );
  NOR2_X1 U12379 ( .A1(n13131), .A2(n18787), .ZN(n13132) );
  AND2_X1 U12380 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13139) );
  OR2_X1 U12381 ( .A1(n17025), .A2(n17156), .ZN(n9673) );
  AND2_X1 U12382 ( .A1(n14084), .A2(n9663), .ZN(n9674) );
  AND2_X1 U12383 ( .A1(n10743), .A2(n10737), .ZN(n9676) );
  INV_X1 U12384 ( .A(n10127), .ZN(n10332) );
  NAND2_X1 U12385 ( .A1(n15118), .A2(n10504), .ZN(n9777) );
  AND2_X1 U12386 ( .A1(n14442), .A2(n9966), .ZN(n14399) );
  AND2_X1 U12387 ( .A1(n12470), .A2(n9791), .ZN(n9678) );
  NOR2_X1 U12388 ( .A1(n14843), .A2(n12789), .ZN(n12813) );
  OR2_X1 U12389 ( .A1(n13280), .A2(n10868), .ZN(n9680) );
  INV_X1 U12390 ( .A(n15014), .ZN(n9943) );
  NAND2_X1 U12391 ( .A1(n9777), .A2(n10506), .ZN(n15109) );
  AND3_X1 U12392 ( .A1(n10546), .A2(n15037), .A3(n15022), .ZN(n9681) );
  OR2_X1 U12393 ( .A1(n9761), .A2(n9760), .ZN(n9682) );
  OR2_X1 U12394 ( .A1(n11528), .A2(n14025), .ZN(n9683) );
  AND2_X1 U12395 ( .A1(n11519), .A2(n9683), .ZN(n9684) );
  NAND2_X1 U12396 ( .A1(n18706), .A2(n18705), .ZN(n9685) );
  NOR2_X1 U12397 ( .A1(n15078), .A2(n16034), .ZN(n9686) );
  INV_X1 U12398 ( .A(n9877), .ZN(n15012) );
  NAND2_X1 U12399 ( .A1(n12470), .A2(n9667), .ZN(n9877) );
  AND2_X1 U12400 ( .A1(n10332), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9687) );
  INV_X1 U12401 ( .A(n9897), .ZN(n14911) );
  NOR2_X1 U12402 ( .A1(n13198), .A2(n14912), .ZN(n9897) );
  NOR3_X1 U12403 ( .A1(n13198), .A2(n14905), .A3(n9898), .ZN(n9896) );
  NAND2_X1 U12404 ( .A1(n10090), .A2(n10089), .ZN(n13778) );
  INV_X1 U12405 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17428) );
  INV_X1 U12406 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12775) );
  NAND2_X1 U12407 ( .A1(n10894), .A2(n10711), .ZN(n9688) );
  AND2_X1 U12408 ( .A1(n14827), .A2(n13211), .ZN(n13210) );
  OR2_X1 U12409 ( .A1(n19057), .A2(n14271), .ZN(n9689) );
  NAND2_X1 U12410 ( .A1(n10568), .A2(n10569), .ZN(n10572) );
  AND2_X1 U12411 ( .A1(n9682), .A2(n10616), .ZN(n9690) );
  AND2_X1 U12412 ( .A1(n10469), .A2(n10894), .ZN(n9691) );
  AND2_X1 U12413 ( .A1(n14974), .A2(n14981), .ZN(n9692) );
  AND2_X1 U12414 ( .A1(n9927), .A2(n9925), .ZN(n9693) );
  AND2_X1 U12415 ( .A1(n9884), .A2(n9883), .ZN(n9694) );
  INV_X1 U12416 ( .A(n11307), .ZN(n11308) );
  AND2_X1 U12417 ( .A1(n9598), .A2(n10339), .ZN(n9695) );
  NAND2_X1 U12418 ( .A1(n14951), .A2(n15173), .ZN(n9696) );
  INV_X1 U12419 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17389) );
  AND2_X1 U12420 ( .A1(n9983), .A2(n9980), .ZN(n13611) );
  INV_X1 U12421 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11358) );
  INV_X1 U12422 ( .A(n10861), .ZN(n11024) );
  INV_X1 U12423 ( .A(n11024), .ZN(n11030) );
  NOR2_X1 U12424 ( .A1(n9583), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U12425 ( .A1(n9968), .A2(n11791), .ZN(n14116) );
  NAND2_X1 U12426 ( .A1(n14084), .A2(n14874), .ZN(n14866) );
  NAND2_X1 U12427 ( .A1(n9735), .A2(n9734), .ZN(n13607) );
  AND2_X1 U12428 ( .A1(n14373), .A2(n9823), .ZN(n14331) );
  NOR2_X1 U12429 ( .A1(n13131), .A2(n9821), .ZN(n13130) );
  NAND2_X1 U12430 ( .A1(n14138), .A2(n15254), .ZN(n14925) );
  NAND2_X1 U12431 ( .A1(n9735), .A2(n9733), .ZN(n13609) );
  NAND2_X1 U12432 ( .A1(n9584), .A2(n19697), .ZN(n10863) );
  INV_X1 U12433 ( .A(n13086), .ZN(n9987) );
  AND2_X1 U12434 ( .A1(n9979), .A2(n14874), .ZN(n9697) );
  AND2_X1 U12435 ( .A1(n10423), .A2(n10424), .ZN(n10472) );
  NAND2_X1 U12436 ( .A1(n13996), .A2(n9905), .ZN(n9698) );
  NOR2_X1 U12437 ( .A1(n15359), .A2(n9894), .ZN(n15327) );
  NOR2_X1 U12438 ( .A1(n9671), .A2(n15231), .ZN(n13199) );
  OR3_X1 U12439 ( .A1(n15543), .A2(n10894), .A3(n15234), .ZN(n9699) );
  NAND2_X1 U12440 ( .A1(n13127), .A2(n9814), .ZN(n13122) );
  NAND2_X1 U12441 ( .A1(n9642), .A2(n13700), .ZN(n13698) );
  INV_X1 U12442 ( .A(n10138), .ZN(n9865) );
  AND2_X1 U12443 ( .A1(n17479), .A2(n9660), .ZN(n13174) );
  OR2_X1 U12444 ( .A1(n9847), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9700) );
  NAND2_X1 U12445 ( .A1(n9767), .A2(n9766), .ZN(n13988) );
  NAND2_X1 U12446 ( .A1(n9768), .A2(n9772), .ZN(n13906) );
  NAND2_X1 U12447 ( .A1(n9626), .A2(n11519), .ZN(n14024) );
  NAND2_X1 U12448 ( .A1(n9950), .A2(n10477), .ZN(n14218) );
  NAND2_X1 U12449 ( .A1(n15755), .A2(n11474), .ZN(n15750) );
  AND2_X1 U12450 ( .A1(n13128), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13127) );
  AND2_X1 U12451 ( .A1(n14864), .A2(n14858), .ZN(n13195) );
  AND2_X1 U12452 ( .A1(n9890), .A2(n14226), .ZN(n9701) );
  AND2_X1 U12453 ( .A1(n12641), .A2(n12640), .ZN(n9702) );
  AND2_X1 U12454 ( .A1(n13127), .A2(n9815), .ZN(n9703) );
  AND2_X1 U12455 ( .A1(n9599), .A2(n19987), .ZN(n11340) );
  NOR2_X1 U12456 ( .A1(n13131), .A2(n9819), .ZN(n13128) );
  OR2_X1 U12457 ( .A1(n9926), .A2(n9928), .ZN(n9704) );
  NOR2_X1 U12458 ( .A1(n14853), .A2(n12761), .ZN(n14842) );
  NOR2_X1 U12459 ( .A1(n13609), .A2(n13821), .ZN(n13808) );
  NOR2_X1 U12460 ( .A1(n13933), .A2(n12477), .ZN(n12478) );
  OR2_X1 U12461 ( .A1(n17934), .A2(n9847), .ZN(n9705) );
  OR2_X1 U12462 ( .A1(n10367), .A2(n10366), .ZN(n10699) );
  INV_X1 U12463 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17602) );
  AND2_X1 U12464 ( .A1(n14154), .A2(n14153), .ZN(n14151) );
  AND2_X1 U12465 ( .A1(n12672), .A2(n9980), .ZN(n9706) );
  AND2_X1 U12466 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n9707) );
  INV_X1 U12467 ( .A(n9736), .ZN(n9734) );
  NAND2_X1 U12468 ( .A1(n9737), .A2(n13658), .ZN(n9736) );
  INV_X1 U12469 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13123) );
  OR2_X1 U12470 ( .A1(n9894), .A2(n9893), .ZN(n9708) );
  AND2_X1 U12471 ( .A1(n18848), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9709) );
  NAND2_X1 U12472 ( .A1(n12478), .A2(n9739), .ZN(n14087) );
  OR2_X1 U12473 ( .A1(n18656), .A2(n18670), .ZN(n9710) );
  AND2_X1 U12474 ( .A1(n9917), .A2(n10535), .ZN(n9711) );
  AND2_X1 U12475 ( .A1(n9807), .A2(n9808), .ZN(n9712) );
  AND2_X1 U12476 ( .A1(n9814), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9713) );
  AND2_X1 U12477 ( .A1(n9661), .A2(n9889), .ZN(n9714) );
  AND2_X1 U12478 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9715) );
  NAND2_X2 U12479 ( .A1(n12919), .A2(n19720), .ZN(n14873) );
  NOR2_X1 U12480 ( .A1(n13654), .A2(n14225), .ZN(n9716) );
  INV_X1 U12481 ( .A(n15354), .ZN(n16036) );
  NAND2_X1 U12482 ( .A1(n14227), .A2(n14226), .ZN(n14228) );
  NAND2_X1 U12483 ( .A1(n14227), .A2(n9661), .ZN(n15388) );
  NAND2_X1 U12484 ( .A1(n10738), .A2(n9676), .ZN(n13583) );
  INV_X1 U12485 ( .A(n12785), .ZN(n9978) );
  INV_X1 U12486 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9802) );
  INV_X1 U12487 ( .A(n11752), .ZN(n11783) );
  INV_X1 U12488 ( .A(n15991), .ZN(n9947) );
  INV_X1 U12489 ( .A(n14875), .ZN(n9738) );
  OR2_X1 U12490 ( .A1(n15938), .A2(n15946), .ZN(n9717) );
  AND2_X1 U12491 ( .A1(n9915), .A2(n9914), .ZN(n9718) );
  OR3_X1 U12492 ( .A1(n14905), .A2(n9901), .A3(n14912), .ZN(n9719) );
  AND2_X1 U12493 ( .A1(n9983), .A2(n9981), .ZN(n13513) );
  INV_X1 U12494 ( .A(n14897), .ZN(n9901) );
  INV_X1 U12495 ( .A(n13509), .ZN(n10758) );
  OR2_X1 U12496 ( .A1(n17126), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9720) );
  AND2_X1 U12497 ( .A1(n10101), .A2(n10640), .ZN(n9721) );
  INV_X1 U12498 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n9792) );
  NOR2_X2 U12499 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13682) );
  INV_X1 U12500 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n9925) );
  OR2_X1 U12501 ( .A1(n18633), .A2(n10208), .ZN(n15996) );
  AND2_X1 U12502 ( .A1(n9878), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9722) );
  INV_X1 U12503 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9816) );
  AND3_X1 U12504 ( .A1(n10965), .A2(n10964), .A3(n10963), .ZN(n15360) );
  INV_X1 U12505 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n9914) );
  INV_X1 U12506 ( .A(n17553), .ZN(n16598) );
  AND2_X1 U12507 ( .A1(n9791), .A2(n15296), .ZN(n9723) );
  AND2_X1 U12508 ( .A1(n10727), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9724) );
  NOR2_X1 U12509 ( .A1(n17476), .A2(n20724), .ZN(n16526) );
  NAND2_X1 U12510 ( .A1(n14743), .A2(n14751), .ZN(n9725) );
  INV_X1 U12511 ( .A(n9879), .ZN(n9878) );
  NAND2_X1 U12512 ( .A1(n9667), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9879) );
  INV_X1 U12513 ( .A(n12646), .ZN(n9984) );
  INV_X1 U12514 ( .A(n15376), .ZN(n9793) );
  INV_X1 U12515 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19504) );
  OAI221_X1 U12516 ( .B1(n20136), .B2(n20371), .C1(n20136), .C2(n20120), .A(
        n20452), .ZN(n20138) );
  AOI22_X2 U12517 ( .A1(DATAI_16_), .A2(n19958), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20001), .ZN(n20457) );
  NOR3_X2 U12518 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18456), .A3(
        n18165), .ZN(n18139) );
  INV_X1 U12519 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18617) );
  AOI22_X2 U12520 ( .A1(DATAI_17_), .A2(n19958), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20001), .ZN(n20461) );
  NOR2_X2 U12521 ( .A1(n19960), .A2(n19959), .ZN(n20001) );
  NOR3_X2 U12522 ( .A1(n18456), .A2(n18428), .A3(n18077), .ZN(n18049) );
  NAND3_X1 U12523 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_22__SCAN_IN), .ZN(n9729) );
  INV_X2 U12524 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18573) );
  INV_X2 U12525 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18580) );
  NAND3_X1 U12526 ( .A1(n14274), .A2(n9732), .A3(n9689), .ZN(P2_U2983) );
  NAND2_X1 U12527 ( .A1(n11614), .A2(n9744), .ZN(n9743) );
  XNOR2_X2 U12528 ( .A(n11321), .B(n11274), .ZN(n11614) );
  OAI211_X1 U12529 ( .C1(n11614), .C2(n9748), .A(n9745), .B(n9743), .ZN(n11611) );
  NAND2_X1 U12530 ( .A1(n15757), .A2(n9750), .ZN(n9753) );
  AND2_X1 U12531 ( .A1(n11502), .A2(n9751), .ZN(n9752) );
  NAND2_X1 U12532 ( .A1(n15757), .A2(n15756), .ZN(n15755) );
  NAND2_X1 U12533 ( .A1(n9753), .A2(n9752), .ZN(n15744) );
  NAND2_X1 U12534 ( .A1(n14939), .A2(n14938), .ZN(n12979) );
  NAND2_X1 U12535 ( .A1(n14939), .A2(n9763), .ZN(n9762) );
  NAND2_X1 U12536 ( .A1(n14272), .A2(n16044), .ZN(n11103) );
  NAND2_X1 U12537 ( .A1(n9762), .A2(n9756), .ZN(n9755) );
  NOR2_X1 U12538 ( .A1(n9682), .A2(n10616), .ZN(n9756) );
  NOR2_X1 U12539 ( .A1(n9758), .A2(n9690), .ZN(n9757) );
  NAND2_X1 U12540 ( .A1(n9765), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10209) );
  NAND2_X1 U12541 ( .A1(n12618), .A2(n10215), .ZN(n10207) );
  XNOR2_X2 U12542 ( .A(n10732), .B(n10733), .ZN(n12618) );
  NAND2_X1 U12543 ( .A1(n13762), .A2(n9769), .ZN(n9767) );
  NAND2_X1 U12544 ( .A1(n9777), .A2(n9774), .ZN(n10566) );
  NAND3_X1 U12545 ( .A1(n9780), .A2(n10698), .A3(n10894), .ZN(n10348) );
  NAND2_X1 U12546 ( .A1(n9630), .A2(n9867), .ZN(n10698) );
  NAND3_X1 U12547 ( .A1(n13990), .A2(n13991), .A3(n9783), .ZN(n9782) );
  XNOR2_X2 U12548 ( .A(n10470), .B(n10469), .ZN(n10706) );
  NOR2_X1 U12549 ( .A1(n16358), .A2(n16359), .ZN(n16357) );
  INV_X1 U12550 ( .A(n16371), .ZN(n9794) );
  NOR2_X2 U12551 ( .A1(n16300), .A2(n17290), .ZN(n16298) );
  INV_X1 U12552 ( .A(n13135), .ZN(n9800) );
  NAND2_X1 U12553 ( .A1(n9800), .A2(n9801), .ZN(n13133) );
  NAND2_X1 U12554 ( .A1(n9803), .A2(n13168), .ZN(P2_U2825) );
  NAND2_X1 U12555 ( .A1(n9804), .A2(n18838), .ZN(n9803) );
  XNOR2_X1 U12556 ( .A(n9805), .B(n15897), .ZN(n9804) );
  NOR2_X1 U12557 ( .A1(n15900), .A2(n18810), .ZN(n9805) );
  INV_X1 U12558 ( .A(n9809), .ZN(n18668) );
  INV_X1 U12559 ( .A(n18810), .ZN(n9808) );
  INV_X1 U12560 ( .A(n13101), .ZN(n13104) );
  NOR2_X1 U12561 ( .A1(n18810), .A2(n18690), .ZN(n18680) );
  INV_X1 U12562 ( .A(n9818), .ZN(n15944) );
  INV_X1 U12563 ( .A(n13704), .ZN(n9837) );
  NAND2_X1 U12564 ( .A1(n9837), .A2(n9662), .ZN(n15840) );
  INV_X1 U12565 ( .A(n12241), .ZN(n17285) );
  NAND2_X1 U12566 ( .A1(n17517), .A2(n12231), .ZN(n17420) );
  NAND2_X1 U12567 ( .A1(n9846), .A2(n9845), .ZN(n17517) );
  NOR2_X1 U12568 ( .A1(n17420), .A2(n17733), .ZN(n12234) );
  NAND2_X1 U12569 ( .A1(n17568), .A2(n12221), .ZN(n12223) );
  INV_X1 U12570 ( .A(n12222), .ZN(n9849) );
  INV_X2 U12571 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18586) );
  INV_X1 U12572 ( .A(n13800), .ZN(n12957) );
  NAND2_X2 U12573 ( .A1(n9855), .A2(n9853), .ZN(n13800) );
  NAND4_X1 U12574 ( .A1(n10037), .A2(n10034), .A3(n10035), .A4(n10036), .ZN(
        n9854) );
  NAND4_X1 U12575 ( .A1(n10041), .A2(n10038), .A3(n10040), .A4(n10039), .ZN(
        n9856) );
  AND3_X4 U12576 ( .A1(n9634), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10033) );
  INV_X1 U12577 ( .A(n10226), .ZN(n9859) );
  NAND2_X1 U12578 ( .A1(n19132), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n9860) );
  NAND3_X1 U12579 ( .A1(n9687), .A2(n12951), .A3(P2_EBX_REG_0__SCAN_IN), .ZN(
        n9863) );
  NAND2_X4 U12580 ( .A1(n9865), .A2(n9864), .ZN(n10835) );
  INV_X1 U12581 ( .A(n9867), .ZN(n9866) );
  NAND4_X1 U12582 ( .A1(n9872), .A2(n9871), .A3(n9870), .A4(n9869), .ZN(n9868)
         );
  NAND2_X1 U12583 ( .A1(n14964), .A2(n9885), .ZN(n9884) );
  NAND3_X1 U12584 ( .A1(n9884), .A2(n9883), .A3(n10731), .ZN(n9882) );
  NAND2_X1 U12585 ( .A1(n14964), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14959) );
  OAI21_X1 U12586 ( .B1(n15165), .B2(n15156), .A(n9888), .ZN(n9887) );
  INV_X1 U12587 ( .A(n9896), .ZN(n13213) );
  NAND2_X1 U12588 ( .A1(n13622), .A2(n10891), .ZN(n9902) );
  NAND2_X1 U12589 ( .A1(n9902), .A2(n9903), .ZN(n10896) );
  OR2_X1 U12590 ( .A1(n14953), .A2(n9911), .ZN(n9907) );
  NAND3_X1 U12591 ( .A1(n14974), .A2(n9696), .A3(n14981), .ZN(n9908) );
  NAND2_X1 U12592 ( .A1(n9909), .A2(n9910), .ZN(n10605) );
  NAND2_X1 U12593 ( .A1(n14973), .A2(n9692), .ZN(n14948) );
  AND2_X1 U12594 ( .A1(n15164), .A2(n15173), .ZN(n9911) );
  NAND2_X1 U12595 ( .A1(n10498), .A2(n9711), .ZN(n10528) );
  NOR2_X1 U12596 ( .A1(n10531), .A2(n9923), .ZN(n10525) );
  NAND2_X1 U12597 ( .A1(n10482), .A2(n10481), .ZN(n10485) );
  NAND2_X1 U12598 ( .A1(n9655), .A2(n13800), .ZN(n10120) );
  NAND2_X1 U12599 ( .A1(n10165), .A2(n9584), .ZN(n9933) );
  NAND3_X1 U12600 ( .A1(n10101), .A2(n9931), .A3(n10640), .ZN(n10165) );
  NAND3_X1 U12601 ( .A1(n9932), .A2(n12958), .A3(n16067), .ZN(n9931) );
  NAND2_X1 U12602 ( .A1(n9934), .A2(n10470), .ZN(n10707) );
  AND2_X1 U12603 ( .A1(n10470), .A2(n10469), .ZN(n10708) );
  NAND2_X1 U12604 ( .A1(n9935), .A2(n10707), .ZN(n10475) );
  NAND2_X1 U12605 ( .A1(n9688), .A2(n9936), .ZN(n9935) );
  NAND2_X1 U12606 ( .A1(n10470), .A2(n9691), .ZN(n9936) );
  OAI21_X1 U12607 ( .B1(n15002), .B2(n9699), .A(n10577), .ZN(n9944) );
  OAI21_X2 U12608 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n14994) );
  INV_X1 U12609 ( .A(n9944), .ZN(n9939) );
  OAI211_X1 U12610 ( .C1(n15013), .C2(n9944), .A(n9942), .B(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10582) );
  NAND2_X1 U12611 ( .A1(n14051), .A2(n14052), .ZN(n9950) );
  NAND2_X1 U12612 ( .A1(n9946), .A2(n10489), .ZN(n15118) );
  NAND3_X1 U12613 ( .A1(n9950), .A2(n9947), .A3(n9948), .ZN(n9946) );
  NAND2_X2 U12614 ( .A1(n11393), .A2(n11424), .ZN(n13690) );
  OAI21_X1 U12615 ( .B1(n13018), .B2(n19946), .A(n13071), .ZN(P1_U3000) );
  OAI21_X1 U12616 ( .B1(n11614), .B2(n11307), .A(n9956), .ZN(n9957) );
  AOI21_X1 U12617 ( .B1(n11308), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9749), 
        .ZN(n9956) );
  NAND3_X1 U12618 ( .A1(n11536), .A2(n14581), .A3(n11535), .ZN(n14552) );
  AND2_X2 U12619 ( .A1(n11314), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11110) );
  INV_X1 U12620 ( .A(n13503), .ZN(n11622) );
  NAND2_X1 U12621 ( .A1(n9958), .A2(n11623), .ZN(n13503) );
  NAND2_X1 U12622 ( .A1(n9960), .A2(n9959), .ZN(n12918) );
  INV_X1 U12623 ( .A(n14819), .ZN(n9961) );
  AND2_X2 U12624 ( .A1(n14442), .A2(n9963), .ZN(n14376) );
  INV_X1 U12625 ( .A(n14070), .ZN(n9968) );
  NAND2_X1 U12626 ( .A1(n9968), .A2(n9969), .ZN(n14448) );
  NAND2_X1 U12627 ( .A1(n14084), .A2(n9974), .ZN(n9973) );
  OAI211_X1 U12628 ( .C1(n14084), .C2(n12785), .A(n9975), .B(n9973), .ZN(
        n14852) );
  NAND2_X1 U12629 ( .A1(n13442), .A2(n13577), .ZN(n9983) );
  NAND2_X1 U12630 ( .A1(n13967), .A2(n9985), .ZN(n14071) );
  INV_X1 U12631 ( .A(n14071), .ZN(n11773) );
  NOR2_X1 U12632 ( .A1(n14335), .A2(n14337), .ZN(n14336) );
  INV_X1 U12633 ( .A(n10608), .ZN(n10600) );
  AOI21_X1 U12634 ( .B1(n11653), .B2(n11783), .A(n11652), .ZN(n13709) );
  NAND2_X1 U12635 ( .A1(n12920), .A2(n10010), .ZN(n12925) );
  CLKBUF_X1 U12636 ( .A(n14971), .Z(n14991) );
  INV_X1 U12637 ( .A(n14971), .ZN(n10729) );
  NAND2_X1 U12638 ( .A1(n10896), .A2(n10895), .ZN(n14227) );
  OR2_X1 U12639 ( .A1(n13081), .A2(n15996), .ZN(n12996) );
  OAI22_X1 U12640 ( .A1(n14659), .A2(n14465), .B1(n19851), .B2(n14246), .ZN(
        n13096) );
  OR2_X1 U12641 ( .A1(n14318), .A2(n14317), .ZN(n14674) );
  OAI22_X1 U12642 ( .A1(n14318), .A2(n12565), .B1(n13092), .B2(n14322), .ZN(
        n13093) );
  NAND2_X1 U12643 ( .A1(n14318), .A2(n13094), .ZN(n12591) );
  OR2_X1 U12644 ( .A1(n14318), .A2(n12589), .ZN(n12592) );
  OR2_X1 U12645 ( .A1(n13441), .A2(n13440), .ZN(n13443) );
  AND2_X1 U12646 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19696), .ZN(
        n10333) );
  NOR2_X2 U12647 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13918) );
  XNOR2_X1 U12648 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11550) );
  NOR2_X2 U12650 ( .A1(n13393), .A2(n12997), .ZN(n12494) );
  NAND2_X1 U12651 ( .A1(n12494), .A2(n19979), .ZN(n12444) );
  INV_X1 U12652 ( .A(n12494), .ZN(n14300) );
  NAND2_X1 U12653 ( .A1(n11169), .A2(n11168), .ZN(n11251) );
  INV_X1 U12654 ( .A(n11266), .ZN(n11169) );
  AND2_X1 U12655 ( .A1(n11180), .A2(n11254), .ZN(n11168) );
  NAND2_X1 U12656 ( .A1(n13440), .A2(n13441), .ZN(n13442) );
  NAND2_X1 U12657 ( .A1(n12644), .A2(n12643), .ZN(n13441) );
  AND2_X4 U12658 ( .A1(n11112), .A2(n11109), .ZN(n11297) );
  NAND2_X1 U12659 ( .A1(n10160), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10178) );
  NAND2_X1 U12660 ( .A1(n11242), .A2(n11612), .ZN(n11248) );
  OAI21_X2 U12661 ( .B1(n15094), .B2(n12490), .A(n15092), .ZN(n15079) );
  NAND2_X1 U12662 ( .A1(n11622), .A2(n11621), .ZN(n13500) );
  XNOR2_X1 U12663 ( .A(n10339), .B(n10144), .ZN(n10646) );
  AND2_X2 U12664 ( .A1(n11113), .A2(n11110), .ZN(n11327) );
  AND2_X2 U12665 ( .A1(n11110), .A2(n11111), .ZN(n11325) );
  INV_X1 U12666 ( .A(n11604), .ZN(n11606) );
  NAND2_X1 U12667 ( .A1(n11052), .A2(n13778), .ZN(n10135) );
  XNOR2_X1 U12668 ( .A(n13383), .B(n9702), .ZN(n19171) );
  OAI22_X2 U12669 ( .A1(n13759), .A2(n13758), .B1(n10697), .B2(n16047), .ZN(
        n10700) );
  OAI21_X1 U12670 ( .B1(n12632), .B2(n12631), .A(n12643), .ZN(n13383) );
  INV_X1 U12671 ( .A(n12110), .ZN(n12258) );
  NOR2_X1 U12672 ( .A1(n18412), .A2(n12116), .ZN(n12251) );
  AND2_X1 U12673 ( .A1(n13079), .A2(n13078), .ZN(n9992) );
  AND2_X1 U12674 ( .A1(n12935), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10293) );
  NAND2_X1 U12675 ( .A1(n20790), .A2(n19963), .ZN(n20119) );
  AND2_X1 U12676 ( .A1(n19851), .A2(n11254), .ZN(n19847) );
  NAND2_X2 U12677 ( .A1(n14482), .A2(n13357), .ZN(n14493) );
  INV_X1 U12678 ( .A(n12496), .ZN(n12087) );
  AND2_X1 U12679 ( .A1(n11249), .A2(n9593), .ZN(n9993) );
  AND2_X1 U12680 ( .A1(n11339), .A2(n11394), .ZN(n9994) );
  AND2_X1 U12681 ( .A1(n15283), .A2(n15282), .ZN(n9995) );
  OR2_X1 U12682 ( .A1(n10339), .A2(n10790), .ZN(n9996) );
  AND4_X1 U12683 ( .A1(n12167), .A2(n12166), .A3(n12165), .A4(n12164), .ZN(
        n9997) );
  AND2_X1 U12684 ( .A1(n10511), .A2(n15126), .ZN(n15122) );
  INV_X1 U12685 ( .A(n15122), .ZN(n10512) );
  OR2_X1 U12686 ( .A1(n18467), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18615) );
  OR2_X1 U12687 ( .A1(n14633), .A2(n14678), .ZN(n9998) );
  AND3_X1 U12688 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17264), .A3(
        n16153), .ZN(n9999) );
  AND2_X1 U12689 ( .A1(n10707), .A2(n10709), .ZN(n10000) );
  AND2_X1 U12690 ( .A1(n10000), .A2(n13992), .ZN(n10001) );
  INV_X1 U12691 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15686) );
  INV_X1 U12692 ( .A(n16987), .ZN(n16972) );
  INV_X1 U12693 ( .A(n16987), .ZN(n16975) );
  INV_X1 U12694 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11535) );
  NOR2_X1 U12695 ( .A1(n11040), .A2(n14882), .ZN(n10002) );
  INV_X1 U12696 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11314) );
  INV_X1 U12697 ( .A(n11092), .ZN(n10728) );
  AND2_X1 U12698 ( .A1(n12977), .A2(n12976), .ZN(n10003) );
  OR2_X1 U12699 ( .A1(n15135), .A2(n15371), .ZN(n10004) );
  OR2_X1 U12700 ( .A1(n12526), .A2(n12525), .ZN(n10005) );
  AND4_X1 U12701 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10006) );
  INV_X1 U12702 ( .A(n13004), .ZN(n11259) );
  INV_X1 U12703 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11548) );
  INV_X1 U12704 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15558) );
  INV_X1 U12705 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14108) );
  INV_X1 U12706 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12240) );
  AND2_X1 U12707 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10007) );
  AND2_X1 U12708 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10008) );
  OR2_X1 U12709 ( .A1(n19587), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19737) );
  AND2_X1 U12710 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10009) );
  AND2_X1 U12711 ( .A1(n14281), .A2(n14870), .ZN(n10010) );
  NAND2_X1 U12712 ( .A1(n10599), .A2(n10598), .ZN(n10011) );
  AND3_X1 U12713 ( .A1(n10239), .A2(n10238), .A3(n10237), .ZN(n10012) );
  INV_X1 U12714 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19696) );
  AND3_X1 U12715 ( .A1(n12435), .A2(n12434), .A3(n12433), .ZN(n10013) );
  AOI21_X1 U12716 ( .B1(n9587), .B2(n12635), .A(n12634), .ZN(n13286) );
  AND2_X1 U12717 ( .A1(n19681), .A2(n11071), .ZN(n15127) );
  INV_X1 U12718 ( .A(n10198), .ZN(n14217) );
  AND2_X2 U12719 ( .A1(n11113), .A2(n13418), .ZN(n11223) );
  AND4_X1 U12720 ( .A1(n11163), .A2(n11162), .A3(n11161), .A4(n11160), .ZN(
        n10014) );
  AND4_X1 U12721 ( .A1(n11273), .A2(n11272), .A3(n11271), .A4(n13034), .ZN(
        n10015) );
  NAND2_X1 U12722 ( .A1(n19987), .A2(n19979), .ZN(n13022) );
  INV_X1 U12723 ( .A(n12565), .ZN(n12589) );
  INV_X1 U12724 ( .A(n11244), .ZN(n11245) );
  INV_X1 U12725 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10200) );
  INV_X1 U12726 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11542) );
  OAI22_X1 U12727 ( .A1(n19280), .A2(n12827), .B1(n10392), .B2(n10281), .ZN(
        n10282) );
  INV_X1 U12728 ( .A(n19203), .ZN(n10444) );
  AOI22_X1 U12729 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10049) );
  INV_X1 U12730 ( .A(n11487), .ZN(n11490) );
  AOI22_X1 U12731 ( .A1(n11276), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11223), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11114) );
  INV_X1 U12732 ( .A(n10353), .ZN(n10621) );
  INV_X1 U12733 ( .A(n10660), .ZN(n10335) );
  INV_X1 U12734 ( .A(n12840), .ZN(n12841) );
  INV_X1 U12735 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12774) );
  INV_X1 U12736 ( .A(n10374), .ZN(n10375) );
  NAND2_X1 U12737 ( .A1(n9930), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10337) );
  NOR2_X1 U12738 ( .A1(n10072), .A2(n10023), .ZN(n10076) );
  INV_X1 U12739 ( .A(n11556), .ZN(n11552) );
  NAND2_X1 U12740 ( .A1(n11546), .A2(n11545), .ZN(n11551) );
  INV_X1 U12741 ( .A(n11921), .ZN(n11922) );
  OAI21_X1 U12742 ( .B1(n12090), .B2(n11662), .A(n11661), .ZN(n11663) );
  OR2_X1 U12743 ( .A1(n11375), .A2(n11374), .ZN(n11376) );
  INV_X1 U12744 ( .A(n19961), .ZN(n11422) );
  NAND2_X1 U12745 ( .A1(n12839), .A2(n12841), .ZN(n12842) );
  AND2_X1 U12746 ( .A1(n12938), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10262) );
  OAI21_X1 U12747 ( .B1(n13075), .B2(n11070), .A(n13074), .ZN(n13076) );
  INV_X1 U12748 ( .A(n14992), .ZN(n10581) );
  INV_X1 U12749 ( .A(n10644), .ZN(n11061) );
  AOI22_X1 U12750 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U12751 ( .A1(n10070), .A2(n10023), .ZN(n10078) );
  AND2_X1 U12752 ( .A1(n11579), .A2(n11578), .ZN(n12441) );
  INV_X1 U12753 ( .A(n11320), .ZN(n11274) );
  OR2_X1 U12754 ( .A1(n11995), .A2(n11994), .ZN(n12016) );
  NAND2_X1 U12755 ( .A1(n11966), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11967) );
  OR2_X1 U12756 ( .A1(n14435), .A2(n14439), .ZN(n11907) );
  INV_X1 U12757 ( .A(n14073), .ZN(n11772) );
  INV_X1 U12758 ( .A(n13770), .ZN(n11680) );
  OAI211_X1 U12759 ( .C1(n11575), .C2(n11311), .A(n11310), .B(n11309), .ZN(
        n11379) );
  INV_X1 U12760 ( .A(n11248), .ZN(n11256) );
  NAND2_X1 U12761 ( .A1(n13278), .A2(n10208), .ZN(n12863) );
  INV_X1 U12762 ( .A(n10990), .ZN(n11027) );
  OR2_X1 U12763 ( .A1(n10831), .A2(n13106), .ZN(n13105) );
  INV_X1 U12764 ( .A(n14837), .ZN(n10824) );
  NAND2_X1 U12765 ( .A1(n10513), .A2(n10512), .ZN(n10514) );
  AND2_X1 U12766 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n15989), .ZN(
        n10723) );
  AOI21_X1 U12767 ( .B1(n10164), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10151), .ZN(n10152) );
  AND2_X1 U12768 ( .A1(n19678), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19511) );
  INV_X1 U12769 ( .A(n17315), .ZN(n16305) );
  AOI21_X1 U12770 ( .B1(n18428), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12351), .ZN(n12360) );
  INV_X1 U12771 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20774) );
  INV_X1 U12772 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16813) );
  AOI21_X1 U12773 ( .B1(n11579), .B2(n11549), .A(n11578), .ZN(n12443) );
  AND2_X1 U12774 ( .A1(n13866), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13867) );
  INV_X1 U12775 ( .A(n11249), .ZN(n11255) );
  OR2_X1 U12776 ( .A1(n12102), .A2(n14519), .ZN(n12103) );
  OR2_X1 U12777 ( .A1(n12004), .A2(n14341), .ZN(n12039) );
  INV_X1 U12778 ( .A(n12090), .ZN(n12096) );
  OR2_X1 U12779 ( .A1(n11270), .A2(n20640), .ZN(n11752) );
  AND4_X1 U12780 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n13770) );
  AND2_X1 U12781 ( .A1(n20328), .A2(n11356), .ZN(n19964) );
  AND2_X1 U12783 ( .A1(n10827), .A2(n10826), .ZN(n14826) );
  INV_X1 U12784 ( .A(n13935), .ZN(n10792) );
  INV_X1 U12785 ( .A(n13608), .ZN(n10775) );
  INV_X1 U12786 ( .A(n12932), .ZN(n12942) );
  OR2_X1 U12787 ( .A1(n12836), .A2(n12838), .ZN(n12864) );
  AND2_X1 U12788 ( .A1(n13936), .A2(n13890), .ZN(n13938) );
  INV_X1 U12789 ( .A(n15360), .ZN(n10966) );
  AND2_X1 U12790 ( .A1(n10876), .A2(n12954), .ZN(n10870) );
  OR2_X1 U12791 ( .A1(n18673), .A2(n10894), .ZN(n10561) );
  XNOR2_X1 U12792 ( .A(n10720), .B(n10718), .ZN(n14222) );
  NAND2_X1 U12793 ( .A1(n10703), .A2(n10702), .ZN(n13898) );
  OR2_X2 U12794 ( .A1(n10223), .A2(n10222), .ZN(n19170) );
  AND2_X1 U12795 ( .A1(n10380), .A2(n19348), .ZN(n19353) );
  OR2_X1 U12796 ( .A1(n15491), .A2(n18400), .ZN(n14171) );
  NOR2_X1 U12797 ( .A1(n12344), .A2(n15509), .ZN(n12348) );
  NAND2_X1 U12798 ( .A1(n17932), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n12410) );
  INV_X1 U12799 ( .A(n17289), .ZN(n17446) );
  NOR2_X1 U12800 ( .A1(n18464), .A2(n17596), .ZN(n17353) );
  NAND2_X1 U12801 ( .A1(n12242), .A2(n17518), .ZN(n12243) );
  AND2_X1 U12802 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  OR2_X1 U12803 ( .A1(n17531), .A2(n17532), .ZN(n12404) );
  OAI21_X2 U12804 ( .B1(n18399), .B2(n18413), .A(n18398), .ZN(n18409) );
  INV_X1 U12805 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14392) );
  AND2_X1 U12806 ( .A1(n12561), .A2(n12560), .ZN(n14452) );
  INV_X1 U12807 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19768) );
  NOR2_X1 U12808 ( .A1(n13863), .A2(n12997), .ZN(n12606) );
  OAI21_X1 U12809 ( .B1(n12437), .B2(n12447), .A(n12446), .ZN(n13399) );
  INV_X1 U12810 ( .A(n20647), .ZN(n13250) );
  INV_X1 U12811 ( .A(n11963), .ZN(n11966) );
  NOR2_X1 U12812 ( .A1(n11792), .A2(n15664), .ZN(n11811) );
  OR2_X1 U12813 ( .A1(n11740), .A2(n15686), .ZN(n11757) );
  NOR2_X1 U12814 ( .A1(n11696), .A2(n19768), .ZN(n11712) );
  AND2_X1 U12815 ( .A1(n11637), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11646) );
  AND2_X1 U12816 ( .A1(n15577), .A2(n12101), .ZN(n13471) );
  INV_X1 U12817 ( .A(n14761), .ZN(n13059) );
  AND2_X1 U12818 ( .A1(n20074), .A2(n20105), .ZN(n20080) );
  OR2_X1 U12819 ( .A1(n20334), .A2(n20422), .ZN(n20306) );
  INV_X1 U12820 ( .A(n11611), .ZN(n19962) );
  OR2_X1 U12821 ( .A1(n20444), .A2(n20327), .ZN(n19966) );
  INV_X1 U12822 ( .A(n20643), .ZN(n13688) );
  INV_X1 U12823 ( .A(n10678), .ZN(n16063) );
  INV_X1 U12824 ( .A(n13162), .ZN(n13163) );
  NAND2_X1 U12825 ( .A1(n10600), .A2(n10011), .ZN(n15912) );
  NOR2_X1 U12826 ( .A1(n18810), .A2(n18679), .ZN(n18669) );
  AND2_X1 U12827 ( .A1(n11011), .A2(n11010), .ZN(n12480) );
  INV_X1 U12828 ( .A(n12814), .ZN(n12810) );
  AND2_X1 U12829 ( .A1(n18922), .A2(n12975), .ZN(n13275) );
  AND2_X1 U12830 ( .A1(n13278), .A2(n13277), .ZN(n13279) );
  OR2_X1 U12831 ( .A1(n13222), .A2(n9583), .ZN(n13255) );
  AND2_X1 U12832 ( .A1(n10779), .A2(n10778), .ZN(n13821) );
  OR2_X1 U12833 ( .A1(n18813), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15140) );
  AND2_X1 U12834 ( .A1(n14204), .A2(n13344), .ZN(n16014) );
  AND2_X1 U12835 ( .A1(n11076), .A2(n13343), .ZN(n14204) );
  OR2_X1 U12836 ( .A1(n10627), .A2(n19700), .ZN(n19712) );
  AND2_X1 U12837 ( .A1(n16093), .A2(n16095), .ZN(n13730) );
  INV_X1 U12838 ( .A(n19427), .ZN(n19422) );
  OR2_X1 U12839 ( .A1(n19171), .A2(n19692), .ZN(n14039) );
  OR2_X1 U12840 ( .A1(n19353), .A2(n19351), .ZN(n19381) );
  NAND2_X1 U12841 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19515), .ZN(n13750) );
  INV_X1 U12842 ( .A(n13795), .ZN(n13797) );
  NAND3_X1 U12843 ( .A1(n19681), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19515), 
        .ZN(n13734) );
  NOR2_X1 U12844 ( .A1(n16394), .A2(n16393), .ZN(n16392) );
  NOR2_X1 U12845 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16460), .ZN(n16445) );
  NOR2_X1 U12846 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16504), .ZN(n16489) );
  NOR2_X1 U12847 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16533), .ZN(n16515) );
  INV_X1 U12848 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16581) );
  NAND2_X1 U12849 ( .A1(n13183), .A2(n13182), .ZN(n16659) );
  INV_X1 U12850 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16483) );
  NAND2_X1 U12851 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12173) );
  INV_X1 U12852 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17310) );
  INV_X1 U12853 ( .A(n13175), .ZN(n17408) );
  INV_X1 U12854 ( .A(n16526), .ZN(n17525) );
  INV_X1 U12855 ( .A(n17567), .ZN(n16614) );
  NOR2_X1 U12856 ( .A1(n17387), .A2(n17518), .ZN(n17348) );
  INV_X1 U12857 ( .A(n17682), .ZN(n17760) );
  OAI21_X1 U12858 ( .B1(n12368), .B2(n12367), .A(n12366), .ZN(n15508) );
  INV_X1 U12859 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18428) );
  NOR2_X2 U12860 ( .A1(n12309), .A2(n12308), .ZN(n17965) );
  AOI22_X1 U12861 ( .A1(n18384), .A2(n18386), .B1(n16156), .B2(n18390), .ZN(
        n18394) );
  NOR2_X2 U12862 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20418) );
  OAI21_X1 U12863 ( .B1(n14419), .B2(n19793), .A(n12614), .ZN(n12615) );
  INV_X1 U12864 ( .A(n19821), .ZN(n19766) );
  NOR2_X1 U12865 ( .A1(n13866), .A2(n20553), .ZN(n12499) );
  OR2_X1 U12866 ( .A1(n13401), .A2(n19740), .ZN(n13091) );
  INV_X1 U12867 ( .A(n14465), .ZN(n19846) );
  OR2_X1 U12868 ( .A1(n13386), .A2(n13087), .ZN(n12448) );
  INV_X1 U12869 ( .A(n13318), .ZN(n19890) );
  NAND2_X1 U12870 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n11862), .ZN(
        n11904) );
  NAND2_X1 U12871 ( .A1(n11713), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11740) );
  AND2_X1 U12872 ( .A1(n19746), .A2(n12100), .ZN(n19908) );
  AND2_X1 U12873 ( .A1(n12099), .A2(n20418), .ZN(n19911) );
  OR2_X1 U12874 ( .A1(n14718), .A2(n13052), .ZN(n14711) );
  NAND2_X1 U12875 ( .A1(n14800), .A2(n20790), .ZN(n12104) );
  AND2_X1 U12876 ( .A1(n13012), .A2(n14307), .ZN(n13042) );
  NAND2_X1 U12877 ( .A1(n13436), .A2(n14761), .ZN(n15854) );
  INV_X1 U12878 ( .A(n15848), .ZN(n19938) );
  INV_X1 U12879 ( .A(n19945), .ZN(n19925) );
  INV_X1 U12880 ( .A(n20029), .ZN(n20032) );
  OAI22_X1 U12881 ( .A1(n20042), .A2(n20041), .B1(n20236), .B2(n20171), .ZN(
        n20066) );
  INV_X1 U12882 ( .A(n20100), .ZN(n20137) );
  INV_X1 U12883 ( .A(n20200), .ZN(n20161) );
  INV_X1 U12884 ( .A(n20207), .ZN(n20112) );
  OAI22_X1 U12885 ( .A1(n20173), .A2(n20172), .B1(n20171), .B2(n20445), .ZN(
        n20196) );
  OR2_X1 U12886 ( .A1(n13690), .A2(n11422), .ZN(n20207) );
  INV_X1 U12887 ( .A(n20357), .ZN(n20231) );
  INV_X1 U12888 ( .A(n20306), .ZN(n20322) );
  AND2_X1 U12889 ( .A1(n20330), .A2(n9648), .ZN(n20296) );
  NAND2_X1 U12890 ( .A1(n13691), .A2(n19962), .ZN(n20327) );
  INV_X1 U12891 ( .A(n20373), .ZN(n20410) );
  OR2_X1 U12892 ( .A1(n13691), .A2(n19962), .ZN(n20357) );
  NOR2_X2 U12893 ( .A1(n20444), .A2(n20422), .ZN(n20485) );
  INV_X1 U12894 ( .A(n20382), .ZN(n20512) );
  INV_X1 U12895 ( .A(n20397), .ZN(n20530) );
  INV_X1 U12896 ( .A(n20408), .ZN(n20542) );
  AND2_X1 U12897 ( .A1(n20553), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15583) );
  INV_X1 U12898 ( .A(n20606), .ZN(n20609) );
  INV_X1 U12899 ( .A(n16056), .ZN(n13221) );
  NOR2_X1 U12900 ( .A1(n10121), .A2(n18631), .ZN(n13154) );
  XNOR2_X1 U12901 ( .A(n13149), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15897) );
  INV_X1 U12902 ( .A(n18847), .ZN(n18865) );
  OR2_X1 U12903 ( .A1(n12703), .A2(n12702), .ZN(n14874) );
  OR2_X1 U12904 ( .A1(n10909), .A2(n10908), .ZN(n13514) );
  INV_X1 U12905 ( .A(n14880), .ZN(n14870) );
  OR2_X1 U12906 ( .A1(n12692), .A2(n12691), .ZN(n14086) );
  AND2_X1 U12907 ( .A1(n13275), .A2(n18892), .ZN(n18883) );
  AND2_X1 U12908 ( .A1(n18945), .A2(n19730), .ZN(n18978) );
  INV_X1 U12909 ( .A(n19046), .ZN(n13271) );
  INV_X1 U12910 ( .A(n14056), .ZN(n15392) );
  INV_X1 U12911 ( .A(n15996), .ZN(n19052) );
  OAI211_X1 U12912 ( .C1(n16008), .C2(n15921), .A(n15168), .B(n9991), .ZN(
        n15169) );
  AND2_X1 U12913 ( .A1(n11075), .A2(n11047), .ZN(n15354) );
  NOR2_X1 U12914 ( .A1(n19728), .A2(n16070), .ZN(n19708) );
  NOR2_X1 U12915 ( .A1(n16055), .A2(n19697), .ZN(n16049) );
  OAI21_X1 U12916 ( .B1(n13845), .B2(n13844), .A(n13843), .ZN(n19075) );
  NOR2_X2 U12917 ( .A1(n14039), .A2(n19199), .ZN(n19126) );
  OAI21_X1 U12918 ( .B1(n19139), .B2(n19138), .A(n19137), .ZN(n19159) );
  NOR2_X2 U12919 ( .A1(n19199), .A2(n19312), .ZN(n19195) );
  NOR2_X1 U12920 ( .A1(n19172), .A2(n19422), .ZN(n19225) );
  NOR2_X1 U12921 ( .A1(n19199), .A2(n19422), .ZN(n19254) );
  INV_X1 U12922 ( .A(n19311), .ZN(n19299) );
  INV_X1 U12923 ( .A(n19302), .ZN(n19306) );
  OAI21_X1 U12924 ( .B1(n13749), .B2(n13748), .A(n13747), .ZN(n13804) );
  INV_X1 U12925 ( .A(n19392), .ZN(n19515) );
  NOR2_X1 U12926 ( .A1(n19313), .A2(n19312), .ZN(n19383) );
  AND2_X1 U12927 ( .A1(n19171), .A2(n19689), .ZN(n19427) );
  INV_X1 U12928 ( .A(n19509), .ZN(n19462) );
  AND2_X1 U12929 ( .A1(n13754), .A2(n13799), .ZN(n19479) );
  INV_X1 U12930 ( .A(n19566), .ZN(n19497) );
  INV_X1 U12931 ( .A(n19491), .ZN(n19553) );
  INV_X1 U12932 ( .A(n19670), .ZN(n19673) );
  INV_X1 U12933 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19608) );
  INV_X1 U12934 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19587) );
  NAND2_X1 U12935 ( .A1(n12363), .A2(n15507), .ZN(n18391) );
  NOR2_X1 U12936 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16385), .ZN(n16368) );
  NOR2_X1 U12937 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16430), .ZN(n16413) );
  INV_X1 U12938 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17350) );
  NOR2_X1 U12939 ( .A1(n17352), .A2(n13177), .ZN(n16302) );
  INV_X1 U12940 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16534) );
  NOR2_X1 U12941 ( .A1(n13180), .A2(n16612), .ZN(n13182) );
  INV_X1 U12942 ( .A(n16666), .ZN(n16646) );
  NAND2_X1 U12943 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16754), .ZN(n16729) );
  NAND2_X1 U12944 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16953), .ZN(n16929) );
  INV_X1 U12945 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16968) );
  INV_X1 U12946 ( .A(n17955), .ZN(n16612) );
  INV_X1 U12947 ( .A(n17072), .ZN(n17061) );
  NOR2_X1 U12948 ( .A1(n17183), .A2(n17099), .ZN(n17094) );
  INV_X1 U12949 ( .A(n17989), .ZN(n17077) );
  OR2_X1 U12950 ( .A1(n12413), .A2(n12412), .ZN(n12414) );
  INV_X1 U12951 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17794) );
  INV_X1 U12952 ( .A(n17609), .ZN(n17596) );
  INV_X1 U12953 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17668) );
  INV_X1 U12954 ( .A(n17841), .ZN(n17903) );
  INV_X1 U12955 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17771) );
  INV_X1 U12956 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17822) );
  NOR2_X2 U12957 ( .A1(n17108), .A2(n17934), .ZN(n17850) );
  NOR2_X1 U12958 ( .A1(n17627), .A2(n17928), .ZN(n17924) );
  NOR2_X1 U12959 ( .A1(n16272), .A2(n16275), .ZN(n18191) );
  INV_X1 U12960 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18583) );
  NOR2_X1 U12961 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18555), .ZN(
        n18581) );
  INV_X1 U12962 ( .A(n18053), .ZN(n18046) );
  INV_X1 U12963 ( .A(n18075), .ZN(n18068) );
  INV_X1 U12964 ( .A(n18098), .ZN(n18087) );
  NOR2_X1 U12965 ( .A1(n18436), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18213) );
  INV_X1 U12966 ( .A(n18248), .ZN(n18254) );
  INV_X1 U12967 ( .A(n18293), .ZN(n18317) );
  INV_X1 U12968 ( .A(n20812), .ZN(n18353) );
  INV_X1 U12969 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18467) );
  INV_X2 U12970 ( .A(n18892), .ZN(n18891) );
  NOR2_X1 U12971 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13173), .ZN(n16249)
         );
  NAND3_X1 U12972 ( .A1(n12494), .A2(n14307), .A3(n14301), .ZN(n14293) );
  INV_X1 U12973 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20641) );
  INV_X1 U12974 ( .A(n12615), .ZN(n12616) );
  INV_X1 U12975 ( .A(n19828), .ZN(n19793) );
  NAND2_X1 U12976 ( .A1(n14405), .A2(n12499), .ZN(n15655) );
  NAND2_X2 U12977 ( .A1(n13091), .A2(n13090), .ZN(n19851) );
  AND2_X1 U12978 ( .A1(n13332), .A2(n13331), .ZN(n19998) );
  NAND2_X1 U12979 ( .A1(n12449), .A2(n12448), .ZN(n14482) );
  INV_X1 U12980 ( .A(n19854), .ZN(n19875) );
  NOR2_X1 U12981 ( .A1(n14293), .A2(n13252), .ZN(n13317) );
  INV_X1 U12982 ( .A(n12107), .ZN(n12108) );
  INV_X1 U12983 ( .A(n15731), .ZN(n19916) );
  OR2_X1 U12984 ( .A1(n12104), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19942) );
  NAND2_X1 U12985 ( .A1(n13042), .A2(n13020), .ZN(n19945) );
  NAND2_X1 U12986 ( .A1(n13060), .A2(n19928), .ZN(n15872) );
  INV_X1 U12987 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19941) );
  OR2_X1 U12988 ( .A1(n20076), .A2(n20357), .ZN(n20029) );
  OR2_X1 U12989 ( .A1(n20076), .A2(n20422), .ZN(n20064) );
  AOI22_X1 U12990 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20078), .B1(n20081), 
        .B2(n20075), .ZN(n20111) );
  NAND2_X1 U12991 ( .A1(n20112), .A2(n20231), .ZN(n20165) );
  OR2_X1 U12992 ( .A1(n20207), .A2(n20422), .ZN(n20200) );
  OR2_X1 U12993 ( .A1(n20207), .A2(n20443), .ZN(n20229) );
  NAND2_X1 U12994 ( .A1(n20232), .A2(n20231), .ZN(n20285) );
  AOI22_X1 U12995 ( .A1(n20291), .A2(n20296), .B1(n20289), .B2(n20288), .ZN(
        n20326) );
  OR2_X1 U12996 ( .A1(n20334), .A2(n20327), .ZN(n20373) );
  AOI22_X1 U12997 ( .A1(n20369), .A2(n20366), .B1(n20362), .B2(n20361), .ZN(
        n20415) );
  OR2_X1 U12998 ( .A1(n20444), .A2(n20357), .ZN(n20442) );
  OR2_X1 U12999 ( .A1(n20444), .A2(n20443), .ZN(n20551) );
  INV_X2 U13000 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20790) );
  INV_X1 U13001 ( .A(n20621), .ZN(n20556) );
  INV_X1 U13002 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20570) );
  OR2_X1 U13003 ( .A1(n20650), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20603) );
  NOR2_X1 U13004 ( .A1(n16065), .A2(n18631), .ZN(n19724) );
  INV_X1 U13005 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19668) );
  AND2_X1 U13006 ( .A1(n13167), .A2(n13166), .ZN(n13168) );
  NAND2_X1 U13007 ( .A1(n18845), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18871) );
  INV_X1 U13008 ( .A(n18859), .ZN(n18841) );
  INV_X1 U13009 ( .A(n12923), .ZN(n12924) );
  OR2_X1 U13010 ( .A1(n13888), .A2(n13810), .ZN(n18740) );
  INV_X1 U13011 ( .A(n19692), .ZN(n19689) );
  AND2_X1 U13012 ( .A1(n12953), .A2(n19720), .ZN(n18922) );
  NAND2_X1 U13013 ( .A1(n12954), .A2(n18922), .ZN(n18936) );
  NAND2_X1 U13014 ( .A1(n18978), .A2(n18947), .ZN(n18976) );
  INV_X1 U13015 ( .A(n18978), .ZN(n19010) );
  OR2_X1 U13016 ( .A1(n13222), .A2(n10208), .ZN(n18943) );
  INV_X1 U13017 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18787) );
  INV_X1 U13018 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18821) );
  INV_X1 U13019 ( .A(n16044), .ZN(n16034) );
  NAND2_X1 U13020 ( .A1(n11075), .A2(n19708), .ZN(n16040) );
  INV_X1 U13021 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19703) );
  INV_X1 U13022 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16073) );
  INV_X1 U13023 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13853) );
  NAND2_X1 U13024 ( .A1(n19083), .A2(n13832), .ZN(n19095) );
  NOR2_X1 U13025 ( .A1(n14043), .A2(n19392), .ZN(n19130) );
  AOI21_X1 U13026 ( .B1(n19134), .B2(n19138), .A(n19133), .ZN(n19162) );
  INV_X1 U13027 ( .A(n19195), .ZN(n19190) );
  INV_X1 U13028 ( .A(n19225), .ZN(n19223) );
  INV_X1 U13029 ( .A(n19254), .ZN(n19249) );
  INV_X1 U13030 ( .A(n19274), .ZN(n19270) );
  OR2_X1 U13031 ( .A1(n19199), .A2(n19670), .ZN(n19302) );
  NOR2_X1 U13032 ( .A1(n13744), .A2(n13743), .ZN(n13807) );
  INV_X1 U13033 ( .A(n19343), .ZN(n19336) );
  INV_X1 U13034 ( .A(n19383), .ZN(n19376) );
  NAND2_X1 U13035 ( .A1(n19428), .A2(n19358), .ZN(n19411) );
  NAND2_X1 U13036 ( .A1(n19449), .A2(n19427), .ZN(n19437) );
  INV_X1 U13037 ( .A(n19498), .ZN(n19484) );
  INV_X1 U13038 ( .A(n19572), .ZN(n19557) );
  INV_X1 U13039 ( .A(n19667), .ZN(n19585) );
  NAND2_X1 U13040 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18566), .ZN(n18455) );
  AOI211_X1 U13041 ( .C1(n16328), .C2(n16655), .A(n16327), .B(n16326), .ZN(
        n16331) );
  INV_X1 U13042 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16537) );
  INV_X1 U13043 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20743) );
  INV_X1 U13044 ( .A(n16610), .ZN(n16656) );
  AND2_X1 U13045 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16728), .ZN(n16723) );
  INV_X1 U13046 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20785) );
  AND2_X1 U13047 ( .A1(n17077), .A2(n9588), .ZN(n16987) );
  INV_X1 U13048 ( .A(n17128), .ZN(n17095) );
  NOR2_X2 U13049 ( .A1(n12126), .A2(n12125), .ZN(n17108) );
  NOR2_X1 U13050 ( .A1(n18600), .A2(n17173), .ZN(n17190) );
  INV_X1 U13051 ( .A(n17173), .ZN(n17205) );
  INV_X1 U13052 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17693) );
  INV_X1 U13053 ( .A(n17519), .ZN(n17498) );
  NAND2_X1 U13054 ( .A1(n12373), .A2(n18605), .ZN(n17612) );
  INV_X1 U13055 ( .A(n17850), .ZN(n17827) );
  INV_X1 U13056 ( .A(n17924), .ZN(n17915) );
  INV_X1 U13057 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18433) );
  OAI211_X1 U13058 ( .C1(n18452), .C2(n18431), .A(n17953), .B(n15497), .ZN(
        n18584) );
  INV_X1 U13059 ( .A(n18111), .ZN(n18120) );
  INV_X1 U13060 ( .A(n18140), .ZN(n18136) );
  INV_X1 U13061 ( .A(n20808), .ZN(n18163) );
  INV_X1 U13062 ( .A(n18179), .ZN(n20811) );
  INV_X1 U13063 ( .A(n18205), .ZN(n18212) );
  INV_X1 U13064 ( .A(n18281), .ZN(n18277) );
  INV_X1 U13065 ( .A(n18377), .ZN(n18334) );
  INV_X1 U13066 ( .A(n18603), .ZN(n18452) );
  INV_X1 U13067 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18555) );
  INV_X1 U13068 ( .A(n18552), .ZN(n18465) );
  INV_X1 U13069 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18480) );
  INV_X1 U13070 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18506) );
  INV_X1 U13071 ( .A(n16225), .ZN(n16229) );
  INV_X1 U13072 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19611) );
  NAND2_X1 U13073 ( .A1(n13098), .A2(n13097), .ZN(P1_U2842) );
  OR4_X1 U13074 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n13202), .ZN(
        P2_U2832) );
  NAND2_X1 U13075 ( .A1(n12925), .A2(n12924), .ZN(P2_U2858) );
  OR4_X1 U13076 ( .A1(n13189), .A2(n13188), .A3(n13187), .A4(n13186), .ZN(
        P3_U2651) );
  NAND2_X1 U13077 ( .A1(n12416), .A2(n12415), .ZN(P3_U2802) );
  INV_X1 U13078 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10016) );
  AND2_X2 U13079 ( .A1(n10017), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13720) );
  AND2_X2 U13080 ( .A1(n13720), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10025) );
  BUF_X4 U13081 ( .A(n10025), .Z(n10235) );
  AND2_X4 U13082 ( .A1(n13720), .A2(n16054), .ZN(n12935) );
  AOI22_X1 U13083 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10022) );
  AND2_X4 U13084 ( .A1(n13918), .A2(n9635), .ZN(n12938) );
  AND3_X4 U13085 ( .A1(n9635), .A2(n10016), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U13086 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10021) );
  AND2_X4 U13087 ( .A1(n13448), .A2(n16054), .ZN(n12941) );
  AND2_X4 U13088 ( .A1(n10018), .A2(n9635), .ZN(n12939) );
  AOI22_X1 U13089 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10020) );
  NAND4_X1 U13090 ( .A1(n10022), .A2(n10021), .A3(n10020), .A4(n10019), .ZN(
        n10024) );
  AOI22_X1 U13091 ( .A1(n10102), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10029) );
  AOI22_X1 U13092 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U13093 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10026) );
  NAND4_X1 U13094 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10030) );
  NAND2_X2 U13095 ( .A1(n10030), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10031) );
  NAND2_X4 U13096 ( .A1(n10032), .A2(n10031), .ZN(n10339) );
  AOI22_X1 U13097 ( .A1(n10102), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10037) );
  AOI22_X1 U13098 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U13099 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12939), .B1(
        n12941), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10035) );
  AOI22_X1 U13100 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10034) );
  AOI22_X1 U13101 ( .A1(n10102), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U13102 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U13103 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10039) );
  AOI22_X1 U13104 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U13105 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10045) );
  AOI22_X1 U13106 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U13107 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10043) );
  AOI22_X1 U13108 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10042) );
  NAND4_X1 U13109 ( .A1(n10045), .A2(n10044), .A3(n10043), .A4(n10042), .ZN(
        n10046) );
  AOI22_X1 U13110 ( .A1(n10102), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U13111 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10048) );
  AOI22_X1 U13112 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10047) );
  NAND4_X1 U13113 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10051) );
  NOR2_X1 U13114 ( .A1(n10120), .A2(n13785), .ZN(n10091) );
  AOI22_X1 U13115 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U13116 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U13117 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10055) );
  NAND4_X1 U13118 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n10058) );
  NAND2_X1 U13119 ( .A1(n10058), .A2(n10023), .ZN(n10065) );
  AOI22_X1 U13120 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10062) );
  AOI22_X1 U13121 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10060) );
  AOI22_X1 U13122 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10059) );
  NAND4_X1 U13123 ( .A1(n10062), .A2(n10061), .A3(n10060), .A4(n10059), .ZN(
        n10063) );
  NAND2_X1 U13124 ( .A1(n10063), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10064) );
  INV_X2 U13125 ( .A(n13754), .ZN(n11056) );
  AOI22_X1 U13126 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10069) );
  AOI22_X1 U13127 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10068) );
  AOI22_X1 U13128 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U13129 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10066) );
  AOI22_X1 U13130 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10071) );
  AOI22_X1 U13131 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U13132 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10074) );
  AOI22_X1 U13133 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10073) );
  NAND4_X1 U13134 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10077) );
  AOI22_X1 U13135 ( .A1(n10102), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10082) );
  AOI22_X1 U13136 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U13137 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10080) );
  NAND4_X1 U13138 ( .A1(n10082), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n10083) );
  AOI22_X1 U13139 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U13140 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10086) );
  AOI22_X1 U13141 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10085) );
  NAND4_X1 U13142 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        n10088) );
  INV_X1 U13143 ( .A(n10138), .ZN(n10100) );
  AOI22_X1 U13144 ( .A1(n10102), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U13145 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U13146 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U13147 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U13148 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U13149 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10098) );
  AOI22_X1 U13150 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10097) );
  AOI22_X1 U13151 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U13152 ( .A1(n10100), .A2(n9627), .ZN(n10101) );
  NAND2_X1 U13153 ( .A1(n10144), .A2(n13800), .ZN(n10139) );
  INV_X1 U13154 ( .A(n10139), .ZN(n12975) );
  INV_X2 U13155 ( .A(n11055), .ZN(n13738) );
  NAND4_X1 U13156 ( .A1(n12975), .A2(n9695), .A3(n13738), .A4(n11056), .ZN(
        n10145) );
  NAND2_X1 U13157 ( .A1(n10121), .A2(n15500), .ZN(n10640) );
  NAND2_X1 U13158 ( .A1(n10102), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10106) );
  NAND2_X1 U13159 ( .A1(n12935), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10105) );
  NAND2_X1 U13160 ( .A1(n9592), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10104) );
  NAND2_X1 U13161 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10103) );
  NAND4_X1 U13162 ( .A1(n10106), .A2(n10105), .A3(n10104), .A4(n10103), .ZN(
        n10107) );
  OAI22_X1 U13163 ( .A1(n12725), .A2(n19064), .B1(n12729), .B2(n12766), .ZN(
        n10110) );
  OAI22_X1 U13164 ( .A1(n9620), .A2(n10228), .B1(n12728), .B2(n10216), .ZN(
        n10109) );
  NAND2_X1 U13165 ( .A1(n10235), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10114) );
  NAND2_X1 U13166 ( .A1(n12935), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10113) );
  NAND2_X1 U13167 ( .A1(n9591), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10112) );
  NAND2_X1 U13168 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10111) );
  NAND4_X1 U13169 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10115) );
  INV_X1 U13170 ( .A(n10855), .ZN(n12958) );
  AND2_X1 U13171 ( .A1(n13754), .A2(n13800), .ZN(n10122) );
  NAND3_X1 U13172 ( .A1(n9584), .A2(n10123), .A3(n9656), .ZN(n10124) );
  NAND2_X1 U13173 ( .A1(n10124), .A2(n9598), .ZN(n10125) );
  NOR2_X2 U13174 ( .A1(n11059), .A2(n10644), .ZN(n12951) );
  INV_X1 U13175 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U13176 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10130) );
  INV_X1 U13177 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10128) );
  OAI211_X1 U13178 ( .C1(n10155), .C2(n10131), .A(n10130), .B(n10129), .ZN(
        n10132) );
  AOI21_X1 U13179 ( .B1(n10739), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10132), .ZN(n10153) );
  NAND2_X1 U13180 ( .A1(n10864), .A2(n9583), .ZN(n11058) );
  NAND2_X1 U13181 ( .A1(n10137), .A2(n11058), .ZN(n10150) );
  NOR2_X1 U13182 ( .A1(n10139), .A2(n9656), .ZN(n10140) );
  NAND2_X1 U13183 ( .A1(n10141), .A2(n10140), .ZN(n10628) );
  NOR2_X1 U13184 ( .A1(n13738), .A2(n9583), .ZN(n10142) );
  NAND2_X1 U13185 ( .A1(n10628), .A2(n10142), .ZN(n11045) );
  NAND3_X1 U13186 ( .A1(n11045), .A2(n10138), .A3(n9627), .ZN(n10148) );
  NAND3_X1 U13187 ( .A1(n10143), .A2(n11055), .A3(n13800), .ZN(n10147) );
  MUX2_X1 U13188 ( .A(n11056), .B(n10339), .S(n10144), .Z(n10146) );
  OAI211_X1 U13189 ( .C1(n10147), .C2(n10146), .A(n10121), .B(n10145), .ZN(
        n11065) );
  NAND2_X1 U13190 ( .A1(n10150), .A2(n10149), .ZN(n10160) );
  OAI21_X1 U13191 ( .B1(n19687), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n18626), 
        .ZN(n10151) );
  NAND2_X1 U13192 ( .A1(n10153), .A2(n10152), .ZN(n10175) );
  AND2_X2 U13193 ( .A1(n10154), .A2(n10175), .ZN(n10194) );
  INV_X1 U13194 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10156) );
  NOR2_X1 U13195 ( .A1(n10644), .A2(n10127), .ZN(n10159) );
  OAI22_X1 U13196 ( .A1(n10160), .A2(n10159), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10158), .ZN(n10162) );
  NAND2_X1 U13197 ( .A1(n11071), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10163) );
  NAND2_X1 U13198 ( .A1(n10164), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10167) );
  AOI22_X1 U13200 ( .A1(n13450), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n11071), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10166) );
  AND2_X2 U13201 ( .A1(n10167), .A2(n10166), .ZN(n10190) );
  INV_X1 U13202 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10171) );
  INV_X1 U13203 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10168) );
  NAND2_X1 U13204 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10169) );
  OAI211_X1 U13205 ( .C1(n10155), .C2(n10171), .A(n10170), .B(n10169), .ZN(
        n10172) );
  AOI21_X2 U13206 ( .B1(n10739), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10172), .ZN(n10191) );
  NAND2_X1 U13207 ( .A1(n10184), .A2(n10190), .ZN(n10173) );
  NAND2_X1 U13208 ( .A1(n10174), .A2(n10173), .ZN(n10195) );
  NAND2_X1 U13209 ( .A1(n10194), .A2(n10195), .ZN(n10176) );
  NAND2_X1 U13210 ( .A1(n10176), .A2(n10175), .ZN(n10732) );
  NAND2_X1 U13211 ( .A1(n11071), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10177) );
  INV_X1 U13212 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10180) );
  OAI22_X1 U13213 ( .A1(n10835), .A2(n10180), .B1(n18626), .B2(n13763), .ZN(
        n10181) );
  AOI21_X1 U13214 ( .B1(n10848), .B2(P2_EBX_REG_3__SCAN_IN), .A(n10181), .ZN(
        n10182) );
  INV_X1 U13215 ( .A(n10185), .ZN(n10188) );
  INV_X1 U13216 ( .A(n10186), .ZN(n10187) );
  NAND2_X1 U13217 ( .A1(n10188), .A2(n10187), .ZN(n10189) );
  NOR2_X1 U13218 ( .A1(n15399), .A2(n10201), .ZN(n10215) );
  INV_X1 U13219 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12772) );
  INV_X1 U13220 ( .A(n10196), .ZN(n10197) );
  OAI22_X1 U13221 ( .A1(n10384), .A2(n12772), .B1(n10200), .B2(n10392), .ZN(
        n10206) );
  INV_X1 U13222 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10204) );
  INV_X1 U13223 ( .A(n15399), .ZN(n18869) );
  NAND2_X1 U13224 ( .A1(n12618), .A2(n10214), .ZN(n10202) );
  OR2_X2 U13225 ( .A1(n10202), .A2(n13533), .ZN(n10383) );
  OR2_X2 U13226 ( .A1(n10202), .A2(n14217), .ZN(n10379) );
  INV_X1 U13227 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10203) );
  OAI22_X1 U13228 ( .A1(n10204), .A2(n10383), .B1(n10379), .B2(n10203), .ZN(
        n10205) );
  OR2_X2 U13229 ( .A1(n12618), .A2(n14217), .ZN(n10223) );
  NAND2_X1 U13230 ( .A1(n9587), .A2(n15399), .ZN(n10225) );
  INV_X1 U13231 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12765) );
  OAI211_X1 U13232 ( .C1(n19232), .C2(n12765), .A(n10209), .B(n10208), .ZN(
        n10210) );
  NOR2_X1 U13233 ( .A1(n10211), .A2(n10210), .ZN(n10234) );
  NAND2_X1 U13234 ( .A1(n9579), .A2(n9587), .ZN(n10388) );
  INV_X1 U13235 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12773) );
  OAI22_X1 U13236 ( .A1(n12775), .A2(n9670), .B1(n9631), .B2(n12773), .ZN(
        n10213) );
  INV_X1 U13237 ( .A(n10213), .ZN(n10233) );
  INV_X1 U13238 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10217) );
  NOR2_X2 U13239 ( .A1(n10223), .A2(n10221), .ZN(n19203) );
  INV_X1 U13240 ( .A(n10215), .ZN(n10218) );
  OAI22_X1 U13241 ( .A1(n10217), .A2(n10444), .B1(n19132), .B2(n10216), .ZN(
        n10220) );
  OR2_X1 U13242 ( .A1(n9587), .A2(n18869), .ZN(n10222) );
  OR2_X2 U13243 ( .A1(n10226), .A2(n10222), .ZN(n10398) );
  OR2_X2 U13244 ( .A1(n10223), .A2(n10218), .ZN(n10446) );
  INV_X1 U13245 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12764) );
  OAI22_X1 U13246 ( .A1(n19064), .A2(n10398), .B1(n10446), .B2(n12764), .ZN(
        n10219) );
  NOR2_X1 U13247 ( .A1(n10220), .A2(n10219), .ZN(n10232) );
  INV_X1 U13248 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10224) );
  OR2_X2 U13249 ( .A1(n10226), .A2(n10221), .ZN(n19079) );
  OAI22_X1 U13250 ( .A1(n10224), .A2(n19079), .B1(n19170), .B2(n12766), .ZN(
        n10230) );
  OAI22_X1 U13251 ( .A1(n10449), .A2(n10228), .B1(n12774), .B2(n19280), .ZN(
        n10229) );
  NOR2_X1 U13252 ( .A1(n10230), .A2(n10229), .ZN(n10231) );
  NAND4_X1 U13253 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n10270) );
  CLKBUF_X3 U13254 ( .A(n10235), .Z(n12778) );
  AND2_X2 U13255 ( .A1(n12778), .A2(n10023), .ZN(n12747) );
  AOI22_X1 U13256 ( .A1(n12747), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10301), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10244) );
  INV_X1 U13257 ( .A(n10236), .ZN(n12732) );
  AND2_X2 U13258 ( .A1(n9592), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10295) );
  AOI22_X1 U13259 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U13260 ( .A1(n12749), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13261 ( .A1(n10250), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10237) );
  AND2_X1 U13262 ( .A1(n12938), .A2(n10023), .ZN(n10903) );
  AOI22_X1 U13263 ( .A1(n10294), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10903), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10243) );
  AND2_X2 U13264 ( .A1(n12929), .A2(n10023), .ZN(n10292) );
  AOI22_X1 U13265 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13266 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10241) );
  AND2_X1 U13267 ( .A1(n12939), .A2(n10023), .ZN(n10302) );
  AOI22_X1 U13268 ( .A1(n10249), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10302), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10240) );
  NAND3_X1 U13269 ( .A1(n10244), .A2(n10012), .A3(n10006), .ZN(n10860) );
  INV_X1 U13270 ( .A(n10860), .ZN(n10689) );
  OR2_X1 U13271 ( .A1(n10689), .A2(n10208), .ZN(n13233) );
  INV_X1 U13272 ( .A(n13233), .ZN(n10257) );
  AOI22_X1 U13273 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10292), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U13274 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10293), .B1(
        n9590), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13275 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12749), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13276 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10295), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10245) );
  NAND4_X1 U13277 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10256) );
  AOI22_X1 U13278 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10302), .B1(
        n10301), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13279 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U13280 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10903), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U13281 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10917), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10251) );
  NAND4_X1 U13282 ( .A1(n10254), .A2(n10253), .A3(n10252), .A4(n10251), .ZN(
        n10255) );
  NAND2_X1 U13283 ( .A1(n10257), .A2(n10687), .ZN(n10693) );
  AOI22_X1 U13284 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10292), .B1(
        n10294), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13285 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12747), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13286 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U13287 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12749), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10258) );
  NAND4_X1 U13288 ( .A1(n10261), .A2(n10260), .A3(n10259), .A4(n10258), .ZN(
        n10268) );
  AOI22_X1 U13289 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10302), .B1(
        n10301), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13290 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U13291 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10903), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13292 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10262), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10263) );
  NAND4_X1 U13293 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10267) );
  NAND2_X1 U13294 ( .A1(n10693), .A2(n10872), .ZN(n10269) );
  INV_X1 U13295 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10271) );
  INV_X1 U13296 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12825) );
  OAI22_X1 U13297 ( .A1(n10271), .A2(n10380), .B1(n10384), .B2(n12825), .ZN(
        n10275) );
  INV_X1 U13298 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10273) );
  INV_X1 U13299 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10272) );
  OAI22_X1 U13300 ( .A1(n10273), .A2(n10383), .B1(n10379), .B2(n10272), .ZN(
        n10274) );
  OR2_X1 U13301 ( .A1(n10275), .A2(n10274), .ZN(n10277) );
  INV_X1 U13302 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12826) );
  NOR2_X1 U13303 ( .A1(n10388), .A2(n12826), .ZN(n10276) );
  NOR2_X1 U13304 ( .A1(n10277), .A2(n10276), .ZN(n10291) );
  INV_X1 U13305 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U13306 ( .A1(n19203), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10278) );
  OAI211_X1 U13307 ( .C1(n9670), .C2(n12828), .A(n10279), .B(n10278), .ZN(
        n10280) );
  INV_X1 U13308 ( .A(n10280), .ZN(n10290) );
  INV_X1 U13309 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12818) );
  INV_X1 U13310 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12816) );
  OAI22_X1 U13311 ( .A1(n12818), .A2(n10398), .B1(n10446), .B2(n12816), .ZN(
        n10283) );
  INV_X1 U13312 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12827) );
  INV_X1 U13313 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10281) );
  NOR2_X1 U13314 ( .A1(n10283), .A2(n10282), .ZN(n10289) );
  INV_X1 U13315 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10284) );
  INV_X1 U13316 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12817) );
  OAI22_X1 U13317 ( .A1(n10284), .A2(n10449), .B1(n19232), .B2(n12817), .ZN(
        n10287) );
  INV_X1 U13318 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10285) );
  INV_X1 U13319 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12819) );
  OAI22_X1 U13320 ( .A1(n10285), .A2(n19079), .B1(n19170), .B2(n12819), .ZN(
        n10286) );
  NOR2_X1 U13321 ( .A1(n10286), .A2(n10287), .ZN(n10288) );
  NAND4_X1 U13322 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10310) );
  AOI22_X1 U13323 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13324 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12747), .B1(
        n10294), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13325 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10298) );
  AOI22_X1 U13326 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12749), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10297) );
  NAND4_X1 U13327 ( .A1(n10300), .A2(n10299), .A3(n10298), .A4(n10297), .ZN(
        n10308) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13329 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13330 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12697), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13331 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10303) );
  NAND4_X1 U13332 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10307) );
  INV_X1 U13333 ( .A(n10345), .ZN(n10882) );
  NAND2_X1 U13334 ( .A1(n10882), .A2(n9584), .ZN(n10309) );
  NAND2_X1 U13335 ( .A1(n10310), .A2(n10309), .ZN(n10311) );
  NAND2_X1 U13336 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10315) );
  NAND2_X1 U13337 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10314) );
  NAND2_X1 U13338 ( .A1(n10294), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U13339 ( .A1(n12747), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10312) );
  NAND2_X1 U13340 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10319) );
  NAND2_X1 U13341 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10318) );
  NAND2_X1 U13342 ( .A1(n10250), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10317) );
  NAND2_X1 U13343 ( .A1(n10917), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10316) );
  NAND2_X1 U13344 ( .A1(n10249), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10323) );
  NAND2_X1 U13345 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10322) );
  NAND2_X1 U13346 ( .A1(n10903), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10321) );
  NAND2_X1 U13347 ( .A1(n10262), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10320) );
  NAND2_X1 U13348 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10327) );
  NAND2_X1 U13349 ( .A1(n10295), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10326) );
  NAND2_X1 U13350 ( .A1(n12749), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10325) );
  NAND2_X1 U13351 ( .A1(n10296), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10324) );
  MUX2_X1 U13352 ( .A(n19696), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10654) );
  NAND2_X1 U13353 ( .A1(n19703), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10353) );
  NAND2_X1 U13354 ( .A1(n16054), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10343) );
  OAI21_X1 U13355 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16054), .A(
        n10343), .ZN(n10334) );
  XNOR2_X1 U13356 ( .A(n10342), .B(n10334), .ZN(n10660) );
  INV_X1 U13357 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13430) );
  NAND3_X1 U13358 ( .A1(n9656), .A2(n10171), .A3(n13430), .ZN(n10340) );
  NAND2_X1 U13359 ( .A1(n10687), .A2(n10339), .ZN(n10867) );
  NAND2_X1 U13360 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19687), .ZN(
        n10341) );
  NAND2_X1 U13361 ( .A1(n10342), .A2(n10341), .ZN(n10344) );
  NAND2_X1 U13362 ( .A1(n10344), .A2(n10343), .ZN(n10369) );
  XNOR2_X1 U13363 ( .A(n10369), .B(n10368), .ZN(n10617) );
  INV_X1 U13364 ( .A(n10617), .ZN(n10664) );
  MUX2_X1 U13365 ( .A(n10345), .B(n10664), .S(n10127), .Z(n10633) );
  INV_X1 U13366 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10346) );
  MUX2_X1 U13367 ( .A(n10633), .B(n10346), .S(n9656), .Z(n10347) );
  OAI21_X1 U13368 ( .B1(n10349), .B2(n10347), .A(n10376), .ZN(n13619) );
  INV_X1 U13369 ( .A(n10349), .ZN(n10352) );
  NAND2_X1 U13370 ( .A1(n10350), .A2(n10355), .ZN(n10351) );
  NAND2_X1 U13371 ( .A1(n10352), .A2(n10351), .ZN(n13529) );
  INV_X1 U13372 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11051) );
  OAI21_X1 U13373 ( .B1(n19703), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10353), .ZN(n10655) );
  MUX2_X1 U13374 ( .A(n10689), .B(n10655), .S(n10127), .Z(n10632) );
  MUX2_X1 U13375 ( .A(n10632), .B(n13430), .S(n9656), .Z(n18866) );
  NOR2_X1 U13376 ( .A1(n18866), .A2(n13714), .ZN(n13231) );
  INV_X1 U13377 ( .A(n13231), .ZN(n13240) );
  NAND3_X1 U13378 ( .A1(n9656), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U13379 ( .A1(n10355), .A2(n10354), .ZN(n13637) );
  NOR2_X1 U13380 ( .A1(n13240), .A2(n13637), .ZN(n10356) );
  NAND2_X1 U13381 ( .A1(n13240), .A2(n13637), .ZN(n13239) );
  OAI21_X1 U13382 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10356), .A(
        n13239), .ZN(n14194) );
  XNOR2_X1 U13383 ( .A(n13529), .B(n11051), .ZN(n14193) );
  OR2_X1 U13384 ( .A1(n14194), .A2(n14193), .ZN(n14191) );
  OAI21_X1 U13385 ( .B1(n13529), .B2(n11051), .A(n14191), .ZN(n13760) );
  AOI22_X1 U13386 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10292), .B1(
        n9590), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13387 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12747), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10359) );
  AOI22_X1 U13388 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10295), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13389 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12749), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10357) );
  NAND4_X1 U13390 ( .A1(n10360), .A2(n10359), .A3(n10358), .A4(n10357), .ZN(
        n10367) );
  AOI22_X1 U13391 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10903), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13392 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13393 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10301), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13394 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12697), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10362) );
  NAND4_X1 U13395 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10366) );
  NAND2_X1 U13396 ( .A1(n19680), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10370) );
  INV_X1 U13397 ( .A(n10668), .ZN(n10372) );
  MUX2_X1 U13398 ( .A(n10699), .B(n10372), .S(n10127), .Z(n10634) );
  INV_X1 U13399 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10373) );
  MUX2_X1 U13400 ( .A(n10634), .B(n10373), .S(n9930), .Z(n10374) );
  AND2_X1 U13401 ( .A1(n10376), .A2(n10375), .ZN(n10377) );
  OR2_X1 U13402 ( .A1(n10377), .A2(n10423), .ZN(n10378) );
  XNOR2_X1 U13403 ( .A(n10378), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13907) );
  INV_X1 U13404 ( .A(n10378), .ZN(n18848) );
  INV_X1 U13405 ( .A(n10699), .ZN(n10883) );
  INV_X1 U13406 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10382) );
  INV_X1 U13407 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10381) );
  OAI22_X1 U13408 ( .A1(n10382), .A2(n10379), .B1(n10380), .B2(n10381), .ZN(
        n10387) );
  INV_X1 U13409 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10385) );
  INV_X1 U13410 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12878) );
  OAI22_X1 U13411 ( .A1(n10385), .A2(n10383), .B1(n10384), .B2(n12878), .ZN(
        n10386) );
  OR2_X1 U13412 ( .A1(n10387), .A2(n10386), .ZN(n10390) );
  INV_X1 U13413 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12879) );
  NOR2_X1 U13414 ( .A1(n10388), .A2(n12879), .ZN(n10389) );
  NOR2_X1 U13415 ( .A1(n10390), .A2(n10389), .ZN(n10409) );
  INV_X1 U13416 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10391) );
  INV_X1 U13417 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12872) );
  OAI22_X1 U13418 ( .A1(n10391), .A2(n10449), .B1(n19170), .B2(n12872), .ZN(
        n10395) );
  INV_X1 U13419 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10393) );
  INV_X1 U13420 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12880) );
  OAI22_X1 U13421 ( .A1(n10393), .A2(n10392), .B1(n19280), .B2(n12880), .ZN(
        n10394) );
  NOR2_X1 U13422 ( .A1(n10395), .A2(n10394), .ZN(n10408) );
  INV_X1 U13423 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10397) );
  INV_X1 U13424 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10396) );
  OAI22_X1 U13425 ( .A1(n10397), .A2(n19079), .B1(n19132), .B2(n10396), .ZN(
        n10401) );
  INV_X1 U13426 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10399) );
  INV_X1 U13427 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13647) );
  OAI22_X1 U13428 ( .A1(n10399), .A2(n10444), .B1(n10398), .B2(n13647), .ZN(
        n10400) );
  NOR2_X1 U13429 ( .A1(n10401), .A2(n10400), .ZN(n10407) );
  INV_X1 U13430 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12881) );
  INV_X1 U13431 ( .A(n10446), .ZN(n13735) );
  NAND2_X1 U13432 ( .A1(n13735), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13433 ( .A1(n19230), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10403) );
  INV_X1 U13434 ( .A(n10405), .ZN(n10406) );
  NAND4_X1 U13435 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10421) );
  AOI22_X1 U13436 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10292), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13437 ( .A1(n10294), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U13438 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13439 ( .A1(n12749), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10410) );
  NAND4_X1 U13440 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10419) );
  AOI22_X1 U13441 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13442 ( .A1(n10249), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13443 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13444 ( .A1(n10903), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10414) );
  NAND4_X1 U13445 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10418) );
  INV_X1 U13446 ( .A(n10422), .ZN(n10889) );
  NAND2_X1 U13447 ( .A1(n10889), .A2(n9584), .ZN(n10420) );
  INV_X1 U13448 ( .A(n10706), .ZN(n10710) );
  INV_X1 U13449 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10705) );
  NAND3_X1 U13450 ( .A1(n10710), .A2(n10894), .A3(n10705), .ZN(n10428) );
  INV_X1 U13451 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13633) );
  MUX2_X1 U13452 ( .A(n13633), .B(n10422), .S(n10339), .Z(n10424) );
  NOR2_X1 U13453 ( .A1(n10423), .A2(n10424), .ZN(n10425) );
  OR2_X1 U13454 ( .A1(n10472), .A2(n10425), .ZN(n18831) );
  NAND2_X1 U13455 ( .A1(n18831), .A2(n10705), .ZN(n10426) );
  OAI21_X1 U13456 ( .B1(n18831), .B2(n10705), .A(n10426), .ZN(n10427) );
  NAND2_X1 U13457 ( .A1(n10428), .A2(n10427), .ZN(n13989) );
  NAND2_X1 U13458 ( .A1(n13988), .A2(n13989), .ZN(n10431) );
  OAI21_X1 U13459 ( .B1(n10706), .B2(n10478), .A(n18831), .ZN(n10429) );
  NAND2_X1 U13460 ( .A1(n10429), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10430) );
  NAND2_X1 U13461 ( .A1(n10431), .A2(n10430), .ZN(n14051) );
  INV_X1 U13462 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10433) );
  INV_X1 U13463 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10432) );
  OAI22_X1 U13464 ( .A1(n10433), .A2(n10383), .B1(n10380), .B2(n10432), .ZN(
        n10436) );
  INV_X1 U13465 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10434) );
  INV_X1 U13466 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12901) );
  OAI22_X1 U13467 ( .A1(n10434), .A2(n10379), .B1(n10384), .B2(n12901), .ZN(
        n10435) );
  OR2_X1 U13468 ( .A1(n10436), .A2(n10435), .ZN(n10438) );
  INV_X1 U13469 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12903) );
  NOR2_X1 U13470 ( .A1(n10388), .A2(n12903), .ZN(n10437) );
  NOR2_X1 U13471 ( .A1(n10438), .A2(n10437), .ZN(n10456) );
  INV_X1 U13472 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10439) );
  INV_X1 U13473 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12892) );
  OAI22_X1 U13474 ( .A1(n10439), .A2(n19079), .B1(n19170), .B2(n12892), .ZN(
        n10442) );
  INV_X1 U13475 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10440) );
  INV_X1 U13476 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12904) );
  OAI22_X1 U13477 ( .A1(n10440), .A2(n10392), .B1(n19280), .B2(n12904), .ZN(
        n10441) );
  NOR2_X1 U13478 ( .A1(n10442), .A2(n10441), .ZN(n10455) );
  INV_X1 U13479 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10445) );
  INV_X1 U13480 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10443) );
  OAI22_X1 U13481 ( .A1(n10445), .A2(n10444), .B1(n19132), .B2(n10443), .ZN(
        n10448) );
  INV_X1 U13482 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12895) );
  INV_X1 U13483 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12894) );
  OAI22_X1 U13484 ( .A1(n12895), .A2(n10446), .B1(n10398), .B2(n12894), .ZN(
        n10447) );
  NOR2_X1 U13485 ( .A1(n10448), .A2(n10447), .ZN(n10454) );
  INV_X1 U13486 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U13487 ( .A1(n14044), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10451) );
  NAND2_X1 U13488 ( .A1(n19230), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10450) );
  OAI211_X1 U13489 ( .C1(n10402), .C2(n12906), .A(n10451), .B(n10450), .ZN(
        n10452) );
  INV_X1 U13490 ( .A(n10452), .ZN(n10453) );
  NAND4_X1 U13491 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .ZN(
        n10468) );
  AOI22_X1 U13492 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10293), .B1(
        n10292), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13493 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12747), .B1(
        n10294), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13494 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13495 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12749), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10457) );
  NAND4_X1 U13496 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n10466) );
  AOI22_X1 U13497 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13498 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13499 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12697), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13500 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10461) );
  NAND4_X1 U13501 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10465) );
  INV_X1 U13502 ( .A(n10471), .ZN(n10890) );
  NAND2_X1 U13503 ( .A1(n10890), .A2(n9583), .ZN(n10467) );
  INV_X1 U13504 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13657) );
  MUX2_X1 U13505 ( .A(n13657), .B(n10471), .S(n10339), .Z(n10473) );
  NOR2_X1 U13506 ( .A1(n10472), .A2(n10473), .ZN(n10474) );
  OR2_X1 U13507 ( .A1(n10482), .A2(n10474), .ZN(n18820) );
  NAND2_X1 U13508 ( .A1(n10475), .A2(n18820), .ZN(n10476) );
  INV_X1 U13509 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14060) );
  XNOR2_X1 U13510 ( .A(n10476), .B(n14060), .ZN(n14052) );
  NAND2_X1 U13511 ( .A1(n10476), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10477) );
  INV_X1 U13512 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10479) );
  MUX2_X1 U13513 ( .A(n10479), .B(n10478), .S(n10339), .Z(n10481) );
  INV_X1 U13514 ( .A(n10481), .ZN(n10480) );
  XNOR2_X1 U13515 ( .A(n10482), .B(n10480), .ZN(n18813) );
  INV_X1 U13516 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10756) );
  NOR2_X1 U13517 ( .A1(n10339), .A2(n10756), .ZN(n10483) );
  NAND2_X1 U13518 ( .A1(n10485), .A2(n10483), .ZN(n10484) );
  NAND2_X1 U13519 ( .A1(n9704), .A2(n10484), .ZN(n18798) );
  NAND2_X1 U13520 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10716) );
  NOR2_X1 U13521 ( .A1(n18798), .A2(n10716), .ZN(n15991) );
  INV_X1 U13522 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10761) );
  NAND3_X1 U13523 ( .A1(n10493), .A2(P2_EBX_REG_10__SCAN_IN), .A3(n9930), .ZN(
        n10486) );
  OAI211_X1 U13524 ( .C1(n10493), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10486), .B(
        n10591), .ZN(n18776) );
  OR2_X1 U13525 ( .A1(n18776), .A2(n10894), .ZN(n10487) );
  INV_X1 U13526 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16012) );
  NAND2_X1 U13527 ( .A1(n10487), .A2(n16012), .ZN(n15979) );
  NAND2_X1 U13528 ( .A1(n9930), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10488) );
  XNOR2_X1 U13529 ( .A(n9704), .B(n10488), .ZN(n18791) );
  NAND2_X1 U13530 ( .A1(n18791), .A2(n10478), .ZN(n10491) );
  NAND2_X1 U13531 ( .A1(n10491), .A2(n9792), .ZN(n15976) );
  INV_X1 U13532 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16022) );
  OAI21_X1 U13533 ( .B1(n18798), .B2(n10894), .A(n16022), .ZN(n15142) );
  AND4_X1 U13534 ( .A1(n15979), .A2(n15976), .A3(n15140), .A4(n15142), .ZN(
        n10489) );
  NAND2_X1 U13535 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10490) );
  OR2_X1 U13536 ( .A1(n18776), .A2(n10490), .ZN(n15978) );
  INV_X1 U13537 ( .A(n10491), .ZN(n10492) );
  NAND2_X1 U13538 ( .A1(n10492), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15974) );
  AND2_X1 U13539 ( .A1(n15978), .A2(n15974), .ZN(n15134) );
  INV_X1 U13540 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18763) );
  NAND2_X1 U13541 ( .A1(n10494), .A2(n18763), .ZN(n10499) );
  INV_X1 U13542 ( .A(n10494), .ZN(n10495) );
  NAND2_X1 U13543 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10495), .ZN(n10496) );
  NOR2_X1 U13544 ( .A1(n10339), .A2(n10496), .ZN(n10497) );
  NOR2_X1 U13545 ( .A1(n10498), .A2(n10497), .ZN(n18765) );
  NAND2_X1 U13546 ( .A1(n18765), .A2(n10478), .ZN(n15135) );
  INV_X1 U13547 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15371) );
  AND2_X1 U13548 ( .A1(n15134), .A2(n10004), .ZN(n15119) );
  NAND2_X1 U13549 ( .A1(n9930), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10501) );
  INV_X1 U13550 ( .A(n10499), .ZN(n10500) );
  OR2_X1 U13551 ( .A1(n10501), .A2(n10500), .ZN(n10502) );
  NAND2_X1 U13552 ( .A1(n10509), .A2(n10502), .ZN(n18752) );
  NAND2_X1 U13553 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10503) );
  OR2_X1 U13554 ( .A1(n18752), .A2(n10503), .ZN(n15123) );
  AND2_X1 U13555 ( .A1(n15119), .A2(n15123), .ZN(n10504) );
  INV_X1 U13556 ( .A(n15123), .ZN(n10505) );
  NAND2_X1 U13557 ( .A1(n15135), .A2(n15371), .ZN(n15120) );
  OR2_X1 U13558 ( .A1(n10505), .A2(n15120), .ZN(n10506) );
  INV_X1 U13559 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10507) );
  NOR2_X1 U13560 ( .A1(n10339), .A2(n10507), .ZN(n10508) );
  AND2_X1 U13561 ( .A1(n10509), .A2(n10508), .ZN(n10510) );
  OR2_X1 U13562 ( .A1(n10510), .A2(n10537), .ZN(n18741) );
  INV_X1 U13563 ( .A(n18741), .ZN(n10557) );
  AOI21_X1 U13564 ( .B1(n10557), .B2(n10478), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15111) );
  INV_X1 U13565 ( .A(n15111), .ZN(n10513) );
  OR2_X1 U13566 ( .A1(n18752), .A2(n10894), .ZN(n10511) );
  INV_X1 U13567 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15126) );
  NAND2_X1 U13568 ( .A1(n9930), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10535) );
  INV_X1 U13569 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10515) );
  NOR2_X1 U13570 ( .A1(n10339), .A2(n10515), .ZN(n10526) );
  INV_X1 U13571 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10790) );
  INV_X1 U13572 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10516) );
  NOR2_X1 U13573 ( .A1(n10339), .A2(n10516), .ZN(n10530) );
  NAND2_X1 U13574 ( .A1(n9656), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10523) );
  NAND2_X1 U13575 ( .A1(n9930), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10517) );
  NOR2_X1 U13576 ( .A1(n10525), .A2(n10517), .ZN(n10518) );
  OR2_X1 U13577 ( .A1(n10542), .A2(n10518), .ZN(n18684) );
  INV_X1 U13578 ( .A(n18684), .ZN(n10549) );
  AOI21_X1 U13579 ( .B1(n10549), .B2(n10478), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15026) );
  MUX2_X1 U13580 ( .A(P2_EBX_REG_16__SCAN_IN), .B(n9996), .S(n10520), .Z(
        n10521) );
  AND2_X1 U13581 ( .A1(n10521), .A2(n10591), .ZN(n18713) );
  NAND2_X1 U13582 ( .A1(n18713), .A2(n10478), .ZN(n10552) );
  INV_X1 U13583 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15311) );
  XNOR2_X1 U13584 ( .A(n10552), .B(n15311), .ZN(n15080) );
  NOR2_X1 U13585 ( .A1(n10522), .A2(n10523), .ZN(n10524) );
  OR2_X1 U13586 ( .A1(n10525), .A2(n10524), .ZN(n18694) );
  INV_X1 U13587 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15065) );
  INV_X1 U13588 ( .A(n10526), .ZN(n10527) );
  XNOR2_X1 U13589 ( .A(n10528), .B(n10527), .ZN(n18723) );
  NAND2_X1 U13590 ( .A1(n18723), .A2(n10478), .ZN(n10529) );
  INV_X1 U13591 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U13592 ( .A1(n10529), .A2(n15090), .ZN(n15092) );
  INV_X1 U13593 ( .A(n10522), .ZN(n10533) );
  NAND2_X1 U13594 ( .A1(n10531), .A2(n10530), .ZN(n10532) );
  NAND2_X1 U13595 ( .A1(n10533), .A2(n10532), .ZN(n18700) );
  OR2_X1 U13596 ( .A1(n18700), .A2(n10894), .ZN(n10534) );
  INV_X1 U13597 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10554) );
  NAND2_X1 U13598 ( .A1(n10534), .A2(n10554), .ZN(n15023) );
  INV_X1 U13599 ( .A(n10535), .ZN(n10536) );
  XNOR2_X1 U13600 ( .A(n10537), .B(n10536), .ZN(n18730) );
  NAND2_X1 U13601 ( .A1(n18730), .A2(n10478), .ZN(n10538) );
  INV_X1 U13602 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15335) );
  NAND2_X1 U13603 ( .A1(n10538), .A2(n15335), .ZN(n15101) );
  NAND4_X1 U13604 ( .A1(n15061), .A2(n15092), .A3(n15023), .A4(n15101), .ZN(
        n10539) );
  NOR3_X1 U13605 ( .A1(n15026), .A2(n15080), .A3(n10539), .ZN(n10546) );
  NAND2_X1 U13606 ( .A1(n9656), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10540) );
  XNOR2_X1 U13607 ( .A(n10542), .B(n10540), .ZN(n18673) );
  INV_X1 U13608 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15261) );
  NAND2_X1 U13609 ( .A1(n10561), .A2(n15261), .ZN(n15037) );
  INV_X1 U13610 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10541) );
  INV_X1 U13611 ( .A(n10568), .ZN(n10545) );
  NAND3_X1 U13612 ( .A1(n10543), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n9656), .ZN(
        n10544) );
  NAND2_X1 U13613 ( .A1(n10545), .A2(n10544), .ZN(n18658) );
  INV_X1 U13614 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15245) );
  OAI21_X1 U13615 ( .B1(n18658), .B2(n10894), .A(n15245), .ZN(n15022) );
  NAND2_X1 U13616 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10547) );
  OR2_X1 U13617 ( .A1(n18658), .A2(n10547), .ZN(n15021) );
  AND2_X1 U13618 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10548) );
  NAND2_X1 U13619 ( .A1(n10549), .A2(n10548), .ZN(n15048) );
  INV_X1 U13620 ( .A(n18694), .ZN(n10551) );
  AND2_X1 U13621 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10550) );
  NAND2_X1 U13622 ( .A1(n10551), .A2(n10550), .ZN(n15060) );
  NAND2_X1 U13623 ( .A1(n15048), .A2(n15060), .ZN(n15027) );
  INV_X1 U13624 ( .A(n10552), .ZN(n10553) );
  NAND2_X1 U13625 ( .A1(n10553), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12491) );
  OR3_X1 U13626 ( .A1(n18700), .A2(n10894), .A3(n10554), .ZN(n12486) );
  AND2_X1 U13627 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10555) );
  NAND2_X1 U13628 ( .A1(n18730), .A2(n10555), .ZN(n15100) );
  AND2_X1 U13629 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10556) );
  NAND2_X1 U13630 ( .A1(n10557), .A2(n10556), .ZN(n12487) );
  AND2_X1 U13631 ( .A1(n15100), .A2(n12487), .ZN(n10559) );
  AND2_X1 U13632 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13633 ( .A1(n18723), .A2(n10558), .ZN(n15091) );
  NAND4_X1 U13634 ( .A1(n12491), .A2(n12486), .A3(n10559), .A4(n15091), .ZN(
        n10560) );
  NOR2_X1 U13635 ( .A1(n15027), .A2(n10560), .ZN(n10563) );
  INV_X1 U13636 ( .A(n10561), .ZN(n10562) );
  NAND2_X1 U13637 ( .A1(n10562), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15038) );
  INV_X1 U13638 ( .A(n10567), .ZN(n10570) );
  NAND2_X1 U13639 ( .A1(n9656), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10569) );
  OAI21_X1 U13640 ( .B1(n10570), .B2(n10569), .A(n10572), .ZN(n15543) );
  INV_X1 U13641 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15234) );
  OAI21_X1 U13642 ( .B1(n15543), .B2(n10894), .A(n15234), .ZN(n15014) );
  INV_X1 U13643 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10571) );
  NOR2_X1 U13644 ( .A1(n10339), .A2(n10571), .ZN(n10573) );
  NAND2_X1 U13645 ( .A1(n10572), .A2(n10573), .ZN(n10574) );
  NAND2_X1 U13646 ( .A1(n10585), .A2(n10574), .ZN(n13193) );
  NOR2_X1 U13647 ( .A1(n13193), .A2(n10894), .ZN(n10575) );
  XNOR2_X1 U13648 ( .A(n10575), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15002) );
  NAND2_X1 U13649 ( .A1(n10478), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10576) );
  NAND2_X1 U13650 ( .A1(n9656), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10579) );
  INV_X1 U13651 ( .A(n10585), .ZN(n10578) );
  MUX2_X1 U13652 ( .A(n10579), .B(P2_EBX_REG_24__SCAN_IN), .S(n10578), .Z(
        n10580) );
  NAND2_X1 U13653 ( .A1(n10580), .A2(n10591), .ZN(n15948) );
  NOR2_X1 U13654 ( .A1(n15948), .A2(n10894), .ZN(n14992) );
  NAND2_X1 U13655 ( .A1(n10582), .A2(n10581), .ZN(n10584) );
  INV_X1 U13656 ( .A(n14994), .ZN(n10583) );
  INV_X1 U13657 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11090) );
  INV_X1 U13658 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15189) );
  INV_X1 U13659 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14838) );
  AND3_X1 U13660 ( .A1(n9930), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10593), .ZN(
        n10586) );
  NOR2_X1 U13661 ( .A1(n10587), .A2(n15189), .ZN(n10604) );
  NOR2_X1 U13662 ( .A1(n10588), .A2(n14838), .ZN(n10589) );
  NAND2_X1 U13663 ( .A1(n9930), .A2(n10589), .ZN(n10590) );
  AND2_X1 U13664 ( .A1(n10591), .A2(n10590), .ZN(n10592) );
  NAND2_X1 U13665 ( .A1(n10593), .A2(n10592), .ZN(n15933) );
  INV_X1 U13666 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15199) );
  NAND2_X1 U13667 ( .A1(n10602), .A2(n15199), .ZN(n14981) );
  NAND2_X1 U13668 ( .A1(n9930), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10595) );
  OR2_X1 U13669 ( .A1(n10595), .A2(n10594), .ZN(n10596) );
  NAND2_X1 U13670 ( .A1(n10599), .A2(n10596), .ZN(n13208) );
  INV_X1 U13671 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15164) );
  INV_X1 U13672 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10597) );
  NOR2_X1 U13673 ( .A1(n10339), .A2(n10597), .ZN(n10598) );
  NAND2_X1 U13674 ( .A1(n10601), .A2(n10478), .ZN(n14953) );
  INV_X1 U13675 ( .A(n10602), .ZN(n10603) );
  NOR2_X1 U13676 ( .A1(n14983), .A2(n10604), .ZN(n14947) );
  NAND2_X1 U13677 ( .A1(n10605), .A2(n14947), .ZN(n14939) );
  NAND2_X1 U13678 ( .A1(n9930), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10607) );
  XOR2_X1 U13679 ( .A(n10607), .B(n10608), .Z(n15903) );
  INV_X1 U13680 ( .A(n15903), .ZN(n10606) );
  INV_X1 U13681 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15156) );
  OAI21_X1 U13682 ( .B1(n10606), .B2(n10894), .A(n15156), .ZN(n14938) );
  NAND2_X1 U13683 ( .A1(n10608), .A2(n10607), .ZN(n10612) );
  INV_X1 U13684 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10841) );
  NOR2_X1 U13685 ( .A1(n10339), .A2(n10841), .ZN(n10609) );
  XNOR2_X1 U13686 ( .A(n10612), .B(n10609), .ZN(n13160) );
  INV_X1 U13687 ( .A(n13160), .ZN(n10610) );
  AOI21_X1 U13688 ( .B1(n10610), .B2(n10478), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12980) );
  INV_X1 U13689 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11070) );
  OR3_X1 U13690 ( .A1(n13160), .A2(n10894), .A3(n11070), .ZN(n12981) );
  NAND3_X1 U13691 ( .A1(n15903), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10478), .ZN(n14937) );
  INV_X1 U13692 ( .A(n10611), .ZN(n10614) );
  NOR2_X1 U13693 ( .A1(n10612), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10613) );
  MUX2_X1 U13694 ( .A(n10614), .B(n10613), .S(n9930), .Z(n15891) );
  NAND2_X1 U13695 ( .A1(n15891), .A2(n10478), .ZN(n10615) );
  XOR2_X1 U13696 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n10615), .Z(
        n10616) );
  INV_X1 U13697 ( .A(n10655), .ZN(n10657) );
  NOR3_X1 U13698 ( .A1(n10668), .A2(n10660), .A3(n10617), .ZN(n10623) );
  XNOR2_X1 U13699 ( .A(n10654), .B(n10353), .ZN(n10656) );
  NAND2_X1 U13700 ( .A1(n10656), .A2(n10623), .ZN(n10622) );
  NAND2_X1 U13701 ( .A1(n10673), .A2(n10622), .ZN(n16056) );
  AOI211_X1 U13702 ( .C1(n10657), .C2(n10623), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n16056), .ZN(n10627) );
  NAND2_X1 U13703 ( .A1(n10624), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13704 ( .A1(n10625), .A2(n16073), .ZN(n16066) );
  INV_X1 U13705 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18634) );
  OAI21_X1 U13706 ( .B1(n9590), .B2(n16066), .A(n18634), .ZN(n10626) );
  AND2_X1 U13707 ( .A1(n10626), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19700) );
  NOR2_X1 U13708 ( .A1(n16070), .A2(n9584), .ZN(n10629) );
  NAND2_X1 U13709 ( .A1(n19712), .A2(n10629), .ZN(n10639) );
  INV_X1 U13710 ( .A(n10654), .ZN(n10631) );
  OAI21_X1 U13711 ( .B1(n10632), .B2(n10631), .A(n10630), .ZN(n10637) );
  NAND2_X1 U13712 ( .A1(n10634), .A2(n10633), .ZN(n10652) );
  INV_X1 U13713 ( .A(n10652), .ZN(n10636) );
  INV_X1 U13714 ( .A(n10673), .ZN(n10635) );
  AOI21_X1 U13715 ( .B1(n10637), .B2(n10636), .A(n10635), .ZN(n19710) );
  NOR2_X1 U13716 ( .A1(n10208), .A2(n10121), .ZN(n13151) );
  INV_X1 U13717 ( .A(n13151), .ZN(n19728) );
  NAND2_X1 U13718 ( .A1(n19710), .A2(n19708), .ZN(n10638) );
  NAND2_X1 U13719 ( .A1(n10639), .A2(n10638), .ZN(n12978) );
  INV_X1 U13720 ( .A(n12978), .ZN(n10681) );
  OAI21_X1 U13721 ( .B1(n12954), .B2(n11056), .A(n11055), .ZN(n10641) );
  NAND2_X1 U13722 ( .A1(n10640), .A2(n10641), .ZN(n10650) );
  NAND2_X1 U13723 ( .A1(n13754), .A2(n9584), .ZN(n11048) );
  NAND2_X1 U13724 ( .A1(n11048), .A2(n10121), .ZN(n10642) );
  NAND2_X1 U13725 ( .A1(n10642), .A2(n13800), .ZN(n10643) );
  NAND2_X1 U13726 ( .A1(n10643), .A2(n11055), .ZN(n10645) );
  AND2_X1 U13727 ( .A1(n10645), .A2(n10644), .ZN(n10649) );
  NAND2_X1 U13728 ( .A1(n10646), .A2(n13800), .ZN(n10647) );
  NAND2_X1 U13729 ( .A1(n10647), .A2(n13151), .ZN(n11053) );
  NAND4_X1 U13730 ( .A1(n10650), .A2(n10649), .A3(n11053), .A4(n10648), .ZN(
        n11049) );
  NAND2_X1 U13731 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19586) );
  NOR2_X1 U13732 ( .A1(n19587), .A2(n19608), .ZN(n19597) );
  NOR2_X1 U13733 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19600) );
  NAND2_X1 U13734 ( .A1(n19586), .A2(n19730), .ZN(n10678) );
  NOR3_X1 U13735 ( .A1(n10138), .A2(n16056), .A3(n10678), .ZN(n10651) );
  NOR2_X1 U13736 ( .A1(n11049), .A2(n10651), .ZN(n13461) );
  NAND2_X1 U13737 ( .A1(n10652), .A2(n10127), .ZN(n10667) );
  NAND2_X1 U13738 ( .A1(n9627), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18946) );
  NAND2_X1 U13739 ( .A1(n18946), .A2(n10208), .ZN(n10653) );
  MUX2_X1 U13740 ( .A(n10127), .B(n10653), .S(n10660), .Z(n10663) );
  OAI21_X1 U13741 ( .B1(n10655), .B2(n10631), .A(n10332), .ZN(n10659) );
  OAI211_X1 U13742 ( .C1(n10208), .C2(n10657), .A(n10121), .B(n10656), .ZN(
        n10658) );
  OAI211_X1 U13743 ( .C1(n10661), .C2(n10660), .A(n10659), .B(n10658), .ZN(
        n10662) );
  NAND2_X1 U13744 ( .A1(n10663), .A2(n10662), .ZN(n10665) );
  NAND2_X1 U13745 ( .A1(n10665), .A2(n10664), .ZN(n10666) );
  NAND2_X1 U13746 ( .A1(n10667), .A2(n10666), .ZN(n10671) );
  NAND2_X1 U13747 ( .A1(n10668), .A2(n10332), .ZN(n10669) );
  NAND2_X1 U13748 ( .A1(n10671), .A2(n10670), .ZN(n10672) );
  MUX2_X1 U13749 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10672), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n10675) );
  INV_X1 U13750 ( .A(n18942), .ZN(n10677) );
  AOI21_X1 U13751 ( .B1(n10675), .B2(n10121), .A(n11056), .ZN(n10676) );
  NAND2_X1 U13752 ( .A1(n10677), .A2(n10676), .ZN(n10680) );
  NAND3_X1 U13753 ( .A1(n18942), .A2(n13738), .A3(n16063), .ZN(n10679) );
  NAND4_X1 U13754 ( .A1(n10681), .A2(n13461), .A3(n10680), .A4(n10679), .ZN(
        n10682) );
  NAND2_X1 U13755 ( .A1(n18626), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U13756 ( .A1(n10682), .A2(n19720), .ZN(n10686) );
  MUX2_X1 U13757 ( .A(n9865), .B(n13738), .S(n9583), .Z(n10684) );
  NAND2_X1 U13758 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19586), .ZN(n19727) );
  NOR2_X1 U13759 ( .A1(n13152), .A2(n19727), .ZN(n10683) );
  NAND3_X1 U13760 ( .A1(n10684), .A2(n13221), .A3(n10683), .ZN(n10685) );
  NOR2_X1 U13761 ( .A1(n16070), .A2(n10127), .ZN(n19707) );
  NAND2_X1 U13762 ( .A1(n13233), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13232) );
  INV_X1 U13763 ( .A(n13232), .ZN(n10690) );
  INV_X1 U13764 ( .A(n10687), .ZN(n10688) );
  XOR2_X1 U13765 ( .A(n10689), .B(n10688), .Z(n10691) );
  NAND2_X1 U13766 ( .A1(n10690), .A2(n10691), .ZN(n10692) );
  XOR2_X1 U13767 ( .A(n10691), .B(n10690), .Z(n13243) );
  NAND2_X1 U13768 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13243), .ZN(
        n13242) );
  NAND2_X1 U13769 ( .A1(n10692), .A2(n13242), .ZN(n10694) );
  XNOR2_X1 U13770 ( .A(n11051), .B(n10694), .ZN(n14190) );
  XNOR2_X1 U13771 ( .A(n10872), .B(n10693), .ZN(n14189) );
  NAND2_X1 U13772 ( .A1(n14190), .A2(n14189), .ZN(n14188) );
  NAND2_X1 U13773 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10694), .ZN(
        n10695) );
  NAND2_X1 U13774 ( .A1(n14188), .A2(n10695), .ZN(n10696) );
  XNOR2_X1 U13775 ( .A(n10696), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13758) );
  INV_X1 U13776 ( .A(n10696), .ZN(n10697) );
  NAND2_X1 U13777 ( .A1(n10700), .A2(n10701), .ZN(n13897) );
  INV_X1 U13778 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13900) );
  NAND2_X1 U13779 ( .A1(n13897), .A2(n13900), .ZN(n10704) );
  INV_X1 U13780 ( .A(n10700), .ZN(n10703) );
  AND2_X2 U13781 ( .A1(n10704), .A2(n13898), .ZN(n13990) );
  NAND2_X1 U13782 ( .A1(n10706), .A2(n10705), .ZN(n13991) );
  OR2_X1 U13783 ( .A1(n10708), .A2(n10711), .ZN(n10709) );
  NAND2_X1 U13784 ( .A1(n10710), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13992) );
  OR2_X1 U13785 ( .A1(n13992), .A2(n10711), .ZN(n10712) );
  NAND2_X1 U13786 ( .A1(n10713), .A2(n13992), .ZN(n10714) );
  NAND2_X1 U13787 ( .A1(n10714), .A2(n10000), .ZN(n10715) );
  XNOR2_X1 U13788 ( .A(n10707), .B(n10894), .ZN(n10718) );
  OAI21_X1 U13789 ( .B1(n10707), .B2(n10894), .A(n16022), .ZN(n10717) );
  INV_X1 U13790 ( .A(n10718), .ZN(n10719) );
  INV_X1 U13791 ( .A(n15989), .ZN(n10721) );
  NOR2_X1 U13792 ( .A1(n15986), .A2(n10721), .ZN(n10722) );
  AOI21_X1 U13793 ( .B1(n14222), .B2(n10723), .A(n10722), .ZN(n15988) );
  NAND2_X2 U13794 ( .A1(n15988), .A2(n10724), .ZN(n12470) );
  AND3_X1 U13795 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15296) );
  AND2_X1 U13796 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12471) );
  AND2_X1 U13797 ( .A1(n15296), .A2(n12471), .ZN(n12476) );
  NAND2_X1 U13798 ( .A1(n12476), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15284) );
  AND2_X1 U13799 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15376) );
  NAND3_X1 U13800 ( .A1(n15376), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10725) );
  NOR2_X1 U13801 ( .A1(n15284), .A2(n10725), .ZN(n15056) );
  AND2_X1 U13802 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15056), .ZN(
        n10726) );
  OR2_X1 U13803 ( .A1(n15245), .A2(n15261), .ZN(n15011) );
  INV_X1 U13804 ( .A(n15011), .ZN(n10727) );
  NAND2_X1 U13805 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11092) );
  NOR2_X2 U13806 ( .A1(n14972), .A2(n15173), .ZN(n14964) );
  INV_X1 U13807 ( .A(n16040), .ZN(n10731) );
  NAND2_X1 U13808 ( .A1(n14273), .A2(n10731), .ZN(n11102) );
  NAND2_X1 U13809 ( .A1(n10732), .A2(n10733), .ZN(n10738) );
  INV_X1 U13810 ( .A(n10734), .ZN(n10736) );
  NAND2_X1 U13811 ( .A1(n10736), .A2(n10735), .ZN(n10737) );
  NAND2_X1 U13812 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10741) );
  NAND2_X1 U13813 ( .A1(n10847), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10740) );
  OAI211_X1 U13814 ( .C1(n10842), .C2(n10373), .A(n10741), .B(n10740), .ZN(
        n10742) );
  AOI21_X1 U13815 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n10742), .ZN(n13584) );
  NAND2_X1 U13816 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10745) );
  NAND2_X1 U13817 ( .A1(n10847), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10744) );
  OAI211_X1 U13818 ( .C1(n10842), .C2(n13633), .A(n10745), .B(n10744), .ZN(
        n10746) );
  AOI21_X1 U13819 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10746), .ZN(n13632) );
  NAND2_X1 U13820 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10748) );
  NAND2_X1 U13821 ( .A1(n10847), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10747) );
  OAI211_X1 U13822 ( .C1(n10842), .C2(n13657), .A(n10748), .B(n10747), .ZN(
        n10749) );
  AOI21_X1 U13823 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10749), .ZN(n13652) );
  INV_X1 U13824 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16021) );
  OR2_X1 U13825 ( .A1(n9651), .A2(n16021), .ZN(n10753) );
  INV_X1 U13826 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10750) );
  OAI22_X1 U13827 ( .A1(n10835), .A2(n10750), .B1(n18626), .B2(n9802), .ZN(
        n10751) );
  AOI21_X1 U13828 ( .B1(n10848), .B2(P2_EBX_REG_7__SCAN_IN), .A(n10751), .ZN(
        n10752) );
  NAND2_X1 U13829 ( .A1(n10753), .A2(n10752), .ZN(n14224) );
  NAND2_X1 U13830 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10755) );
  NAND2_X1 U13831 ( .A1(n10847), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10754) );
  OAI211_X1 U13832 ( .C1(n10842), .C2(n10756), .A(n10755), .B(n10754), .ZN(
        n10757) );
  AOI21_X1 U13833 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10757), .ZN(n13510) );
  NAND2_X1 U13834 ( .A1(n10758), .A2(n13512), .ZN(n13511) );
  NAND2_X1 U13835 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10760) );
  NAND2_X1 U13836 ( .A1(n10847), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10759) );
  OAI211_X1 U13837 ( .C1(n10842), .C2(n10761), .A(n10760), .B(n10759), .ZN(
        n10762) );
  AOI21_X1 U13838 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10762), .ZN(n13549) );
  OR2_X2 U13839 ( .A1(n13511), .A2(n13549), .ZN(n13564) );
  NAND2_X1 U13840 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10764) );
  NAND2_X1 U13841 ( .A1(n10847), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10763) );
  OAI211_X1 U13842 ( .C1(n10842), .C2(n9925), .A(n10764), .B(n10763), .ZN(
        n10765) );
  AOI21_X1 U13843 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10765), .ZN(n13565) );
  OR2_X1 U13844 ( .A1(n9651), .A2(n15371), .ZN(n10770) );
  INV_X1 U13845 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10767) );
  INV_X1 U13846 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10766) );
  OAI22_X1 U13847 ( .A1(n10835), .A2(n10767), .B1(n18626), .B2(n10766), .ZN(
        n10768) );
  AOI21_X1 U13848 ( .B1(n10848), .B2(P2_EBX_REG_11__SCAN_IN), .A(n10768), .ZN(
        n10769) );
  NAND2_X1 U13849 ( .A1(n10770), .A2(n10769), .ZN(n13658) );
  INV_X1 U13850 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10773) );
  NAND2_X1 U13851 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10772) );
  NAND2_X1 U13852 ( .A1(n10847), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10771) );
  OAI211_X1 U13853 ( .C1(n10842), .C2(n10773), .A(n10772), .B(n10771), .ZN(
        n10774) );
  AOI21_X1 U13854 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10774), .ZN(n13608) );
  INV_X1 U13855 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15346) );
  OR2_X1 U13856 ( .A1(n9651), .A2(n15346), .ZN(n10779) );
  INV_X1 U13857 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10776) );
  INV_X1 U13858 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18742) );
  OAI22_X1 U13859 ( .A1(n10835), .A2(n10776), .B1(n18626), .B2(n18742), .ZN(
        n10777) );
  AOI21_X1 U13860 ( .B1(n10848), .B2(P2_EBX_REG_13__SCAN_IN), .A(n10777), .ZN(
        n10778) );
  OR2_X1 U13861 ( .A1(n9651), .A2(n15090), .ZN(n10782) );
  INV_X1 U13862 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19630) );
  OAI22_X1 U13863 ( .A1(n10835), .A2(n19630), .B1(n18626), .B2(n9816), .ZN(
        n10780) );
  AOI21_X1 U13864 ( .B1(n10848), .B2(P2_EBX_REG_15__SCAN_IN), .A(n10780), .ZN(
        n10781) );
  NAND2_X1 U13865 ( .A1(n10782), .A2(n10781), .ZN(n13887) );
  OR2_X1 U13866 ( .A1(n9651), .A2(n15335), .ZN(n10786) );
  INV_X1 U13867 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19628) );
  INV_X1 U13868 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10783) );
  OAI22_X1 U13869 ( .A1(n10835), .A2(n19628), .B1(n18626), .B2(n10783), .ZN(
        n10784) );
  AOI21_X1 U13870 ( .B1(n10848), .B2(P2_EBX_REG_14__SCAN_IN), .A(n10784), .ZN(
        n10785) );
  NAND2_X1 U13871 ( .A1(n10786), .A2(n10785), .ZN(n13809) );
  AND2_X1 U13872 ( .A1(n13887), .A2(n13809), .ZN(n10787) );
  NAND2_X1 U13873 ( .A1(n13808), .A2(n10787), .ZN(n13886) );
  INV_X1 U13874 ( .A(n13886), .ZN(n10793) );
  NAND2_X1 U13875 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10789) );
  NAND2_X1 U13876 ( .A1(n10847), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10788) );
  OAI211_X1 U13877 ( .C1(n10842), .C2(n10790), .A(n10789), .B(n10788), .ZN(
        n10791) );
  AOI21_X1 U13878 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10791), .ZN(n13935) );
  NAND2_X1 U13879 ( .A1(n10844), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10797) );
  INV_X1 U13880 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19634) );
  INV_X1 U13881 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10794) );
  OAI22_X1 U13882 ( .A1(n10835), .A2(n19634), .B1(n18626), .B2(n10794), .ZN(
        n10795) );
  AOI21_X1 U13883 ( .B1(n10848), .B2(P2_EBX_REG_17__SCAN_IN), .A(n10795), .ZN(
        n10796) );
  OR2_X1 U13884 ( .A1(n9651), .A2(n15065), .ZN(n10800) );
  INV_X1 U13885 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15066) );
  INV_X1 U13886 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13144) );
  OAI22_X1 U13887 ( .A1(n10835), .A2(n15066), .B1(n18626), .B2(n13144), .ZN(
        n10798) );
  AOI21_X1 U13888 ( .B1(n10848), .B2(P2_EBX_REG_18__SCAN_IN), .A(n10798), .ZN(
        n10799) );
  NAND2_X1 U13889 ( .A1(n10800), .A2(n10799), .ZN(n14016) );
  INV_X1 U13890 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15273) );
  OR2_X1 U13891 ( .A1(n9651), .A2(n15273), .ZN(n10803) );
  INV_X1 U13892 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19637) );
  OAI22_X1 U13893 ( .A1(n10835), .A2(n19637), .B1(n18626), .B2(n13123), .ZN(
        n10801) );
  AOI21_X1 U13894 ( .B1(n10848), .B2(P2_EBX_REG_19__SCAN_IN), .A(n10801), .ZN(
        n10802) );
  NAND2_X1 U13895 ( .A1(n10803), .A2(n10802), .ZN(n14088) );
  NAND2_X1 U13896 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U13897 ( .A1(n10847), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10804) );
  OAI211_X1 U13898 ( .C1(n10842), .C2(n10541), .A(n10805), .B(n10804), .ZN(
        n10806) );
  AOI21_X1 U13899 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10806), .ZN(n14875) );
  NAND2_X1 U13900 ( .A1(n10844), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10809) );
  INV_X1 U13901 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19641) );
  INV_X1 U13902 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18659) );
  OAI22_X1 U13903 ( .A1(n10835), .A2(n19641), .B1(n18626), .B2(n18659), .ZN(
        n10807) );
  AOI21_X1 U13904 ( .B1(n10848), .B2(P2_EBX_REG_21__SCAN_IN), .A(n10807), .ZN(
        n10808) );
  OR2_X1 U13905 ( .A1(n9651), .A2(n15234), .ZN(n10814) );
  INV_X1 U13906 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10811) );
  INV_X1 U13907 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10810) );
  OAI22_X1 U13908 ( .A1(n10835), .A2(n10811), .B1(n18626), .B2(n10810), .ZN(
        n10812) );
  AOI21_X1 U13909 ( .B1(n10848), .B2(P2_EBX_REG_22__SCAN_IN), .A(n10812), .ZN(
        n10813) );
  NAND2_X1 U13910 ( .A1(n10814), .A2(n10813), .ZN(n14858) );
  INV_X1 U13911 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15219) );
  OR2_X1 U13912 ( .A1(n9651), .A2(n15219), .ZN(n10817) );
  INV_X1 U13913 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19644) );
  OAI22_X1 U13914 ( .A1(n10835), .A2(n19644), .B1(n18626), .B2(n15004), .ZN(
        n10815) );
  AOI21_X1 U13915 ( .B1(n10848), .B2(P2_EBX_REG_23__SCAN_IN), .A(n10815), .ZN(
        n10816) );
  NAND2_X1 U13916 ( .A1(n10817), .A2(n10816), .ZN(n13196) );
  NAND2_X1 U13917 ( .A1(n13195), .A2(n13196), .ZN(n13194) );
  NAND2_X1 U13918 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U13919 ( .A1(n10847), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10818) );
  OAI211_X1 U13920 ( .C1(n10842), .C2(n9914), .A(n10819), .B(n10818), .ZN(
        n10820) );
  AOI21_X1 U13921 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10820), .ZN(n14847) );
  NOR2_X2 U13922 ( .A1(n13194), .A2(n14847), .ZN(n14834) );
  INV_X1 U13923 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19647) );
  INV_X1 U13924 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14986) );
  OAI22_X1 U13925 ( .A1(n10835), .A2(n19647), .B1(n18626), .B2(n14986), .ZN(
        n10821) );
  INV_X1 U13926 ( .A(n10821), .ZN(n10822) );
  OAI21_X1 U13927 ( .B1(n10842), .B2(n14838), .A(n10822), .ZN(n10823) );
  AOI21_X1 U13928 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10823), .ZN(n14837) );
  NAND2_X1 U13929 ( .A1(n10844), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10827) );
  INV_X1 U13930 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19649) );
  INV_X1 U13931 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13111) );
  OAI22_X1 U13932 ( .A1(n10835), .A2(n19649), .B1(n18626), .B2(n13111), .ZN(
        n10825) );
  AOI21_X1 U13933 ( .B1(n10848), .B2(P2_EBX_REG_26__SCAN_IN), .A(n10825), .ZN(
        n10826) );
  OR2_X1 U13934 ( .A1(n9651), .A2(n15173), .ZN(n10830) );
  INV_X1 U13935 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19651) );
  INV_X1 U13936 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14965) );
  OAI22_X1 U13937 ( .A1(n10835), .A2(n19651), .B1(n18626), .B2(n14965), .ZN(
        n10828) );
  AOI21_X1 U13938 ( .B1(n10848), .B2(P2_EBX_REG_27__SCAN_IN), .A(n10828), .ZN(
        n10829) );
  NAND2_X1 U13939 ( .A1(n10830), .A2(n10829), .ZN(n13211) );
  OR2_X1 U13940 ( .A1(n9651), .A2(n15164), .ZN(n10834) );
  INV_X1 U13941 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n14956) );
  INV_X1 U13942 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10831) );
  OAI22_X1 U13943 ( .A1(n10835), .A2(n14956), .B1(n18626), .B2(n10831), .ZN(
        n10832) );
  AOI21_X1 U13944 ( .B1(n10848), .B2(P2_EBX_REG_28__SCAN_IN), .A(n10832), .ZN(
        n10833) );
  NAND2_X1 U13945 ( .A1(n10834), .A2(n10833), .ZN(n14815) );
  OR2_X1 U13946 ( .A1(n9651), .A2(n15156), .ZN(n10838) );
  INV_X1 U13947 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19653) );
  INV_X1 U13948 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14942) );
  OAI22_X1 U13949 ( .A1(n10835), .A2(n19653), .B1(n18626), .B2(n14942), .ZN(
        n10836) );
  AOI21_X1 U13950 ( .B1(n10848), .B2(P2_EBX_REG_29__SCAN_IN), .A(n10836), .ZN(
        n10837) );
  NAND2_X1 U13951 ( .A1(n10838), .A2(n10837), .ZN(n12921) );
  NAND2_X1 U13952 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10840) );
  NAND2_X1 U13953 ( .A1(n10847), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10839) );
  OAI211_X1 U13954 ( .C1(n10842), .C2(n10841), .A(n10840), .B(n10839), .ZN(
        n10843) );
  AOI21_X1 U13955 ( .B1(n10844), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10843), .ZN(n12984) );
  INV_X1 U13956 ( .A(n12984), .ZN(n10845) );
  NAND2_X1 U13957 ( .A1(n10846), .A2(n10845), .ZN(n12987) );
  INV_X1 U13958 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U13959 ( .A1(n10847), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10850) );
  NAND2_X1 U13960 ( .A1(n10848), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n10849) );
  OAI211_X1 U13961 ( .C1(n9651), .C2(n13103), .A(n10850), .B(n10849), .ZN(
        n10851) );
  INV_X1 U13962 ( .A(n10851), .ZN(n10852) );
  OAI21_X1 U13963 ( .B1(n9583), .B2(n13714), .A(n19697), .ZN(n10857) );
  NOR2_X1 U13964 ( .A1(n10855), .A2(n10863), .ZN(n10862) );
  AOI211_X1 U13965 ( .C1(n12957), .C2(P2_EAX_REG_0__SCAN_IN), .A(n10857), .B(
        n10856), .ZN(n13282) );
  INV_X1 U13966 ( .A(n10863), .ZN(n10858) );
  MUX2_X1 U13967 ( .A(n12957), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        P2_STATE2_REG_3__SCAN_IN), .Z(n10859) );
  NOR2_X1 U13968 ( .A1(n13282), .A2(n13281), .ZN(n13280) );
  INV_X1 U13969 ( .A(n10876), .ZN(n11037) );
  INV_X1 U13970 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13713) );
  NOR2_X1 U13971 ( .A1(n13800), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10861) );
  INV_X1 U13972 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19007) );
  INV_X1 U13973 ( .A(n10862), .ZN(n10990) );
  OAI222_X1 U13974 ( .A1(n11037), .A2(n13713), .B1(n11024), .B2(n19007), .C1(
        n10990), .C2(n10168), .ZN(n10868) );
  XNOR2_X1 U13975 ( .A(n13280), .B(n10868), .ZN(n13309) );
  NAND2_X1 U13976 ( .A1(n10864), .A2(n13800), .ZN(n10865) );
  MUX2_X1 U13977 ( .A(n10865), .B(n19696), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10866) );
  OAI21_X1 U13978 ( .B1(n10867), .B2(n10863), .A(n10866), .ZN(n13308) );
  OAI21_X1 U13979 ( .B1(n13309), .B2(n13308), .A(n9680), .ZN(n10869) );
  INV_X1 U13980 ( .A(n10869), .ZN(n10874) );
  AOI21_X1 U13981 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n10870), .ZN(n10871) );
  OAI21_X1 U13982 ( .B1(n10872), .B2(n11005), .A(n10871), .ZN(n10873) );
  XNOR2_X1 U13983 ( .A(n10874), .B(n10873), .ZN(n13519) );
  INV_X1 U13984 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19005) );
  OAI222_X1 U13985 ( .A1(n11037), .A2(n11051), .B1(n11024), .B2(n19005), .C1(
        n10990), .C2(n10128), .ZN(n13518) );
  NOR2_X1 U13986 ( .A1(n13519), .A2(n13518), .ZN(n13517) );
  NOR2_X1 U13987 ( .A1(n10874), .A2(n10873), .ZN(n10875) );
  NAND2_X1 U13988 ( .A1(n11030), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10878) );
  NAND2_X1 U13989 ( .A1(n11041), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10877) );
  OAI211_X1 U13990 ( .C1(n19680), .C2(n19697), .A(n10878), .B(n10877), .ZN(
        n10879) );
  INV_X1 U13991 ( .A(n10879), .ZN(n10881) );
  NAND2_X1 U13992 ( .A1(n11027), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10880) );
  OAI211_X1 U13993 ( .C1(n10882), .C2(n11005), .A(n10881), .B(n10880), .ZN(
        n13620) );
  NAND2_X1 U13994 ( .A1(n13621), .A2(n13620), .ZN(n13622) );
  AOI22_X1 U13995 ( .A1(n11030), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11041), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10886) );
  NAND2_X1 U13996 ( .A1(n11027), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10885) );
  OR2_X1 U13997 ( .A1(n11005), .A2(n10883), .ZN(n10884) );
  AOI22_X1 U13998 ( .A1(n11030), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11041), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10888) );
  NAND2_X1 U13999 ( .A1(n11027), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10887) );
  OAI211_X1 U14000 ( .C1(n10889), .C2(n11005), .A(n10888), .B(n10887), .ZN(
        n13996) );
  OR2_X1 U14001 ( .A1(n11005), .A2(n10890), .ZN(n10891) );
  NAND2_X1 U14002 ( .A1(n11027), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U14003 ( .A1(n11030), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n10892) );
  OAI211_X1 U14004 ( .C1(n11037), .C2(n14060), .A(n10893), .B(n10892), .ZN(
        n14053) );
  OR2_X1 U14005 ( .A1(n11005), .A2(n10894), .ZN(n10895) );
  AOI22_X1 U14006 ( .A1(n11030), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11041), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U14007 ( .A1(n11027), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10897) );
  NAND2_X1 U14008 ( .A1(n10898), .A2(n10897), .ZN(n14226) );
  AOI22_X1 U14009 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10294), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U14010 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U14011 ( .A1(n12749), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U14012 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10899) );
  NAND4_X1 U14013 ( .A1(n10902), .A2(n10901), .A3(n10900), .A4(n10899), .ZN(
        n10909) );
  AOI22_X1 U14014 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10302), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U14015 ( .A1(n10249), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U14016 ( .A1(n10250), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10903), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10905) );
  AOI22_X1 U14017 ( .A1(n10917), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10904) );
  NAND4_X1 U14018 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n10908) );
  NAND2_X1 U14019 ( .A1(n10962), .A2(n13514), .ZN(n10912) );
  AOI22_X1 U14020 ( .A1(n11030), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11041), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10911) );
  NAND2_X1 U14021 ( .A1(n11027), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14022 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U14023 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12747), .B1(
        n10294), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U14024 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U14025 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10913) );
  NAND4_X1 U14026 ( .A1(n10916), .A2(n10915), .A3(n10914), .A4(n10913), .ZN(
        n10923) );
  AOI22_X1 U14027 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U14028 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U14029 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12697), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U14030 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10918) );
  NAND4_X1 U14031 ( .A1(n10921), .A2(n10920), .A3(n10919), .A4(n10918), .ZN(
        n10922) );
  NOR2_X1 U14032 ( .A1(n10923), .A2(n10922), .ZN(n13546) );
  AOI22_X1 U14033 ( .A1(n11030), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11041), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10925) );
  NAND2_X1 U14034 ( .A1(n11027), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10924) );
  OAI211_X1 U14035 ( .C1(n13546), .C2(n11005), .A(n10925), .B(n10924), .ZN(
        n15387) );
  AOI22_X1 U14036 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10292), .B1(
        n9590), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U14037 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12747), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U14038 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U14039 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U14040 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10935) );
  AOI22_X1 U14041 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12697), .B1(
        n10903), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U14042 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U14043 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U14044 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10917), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10930) );
  NAND4_X1 U14045 ( .A1(n10933), .A2(n10932), .A3(n10931), .A4(n10930), .ZN(
        n10934) );
  NOR2_X1 U14046 ( .A1(n10935), .A2(n10934), .ZN(n13560) );
  AOI22_X1 U14047 ( .A1(n11030), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10936) );
  OAI21_X1 U14048 ( .B1(n13560), .B2(n11005), .A(n10936), .ZN(n10937) );
  AOI21_X1 U14049 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n11027), .A(n10937), 
        .ZN(n16007) );
  AOI22_X1 U14050 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14051 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12747), .B1(
        n10294), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14052 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14053 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10938) );
  NAND4_X1 U14054 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10947) );
  AOI22_X1 U14055 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U14056 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U14057 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12697), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14058 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10942) );
  NAND4_X1 U14059 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n10946) );
  NOR2_X1 U14060 ( .A1(n10947), .A2(n10946), .ZN(n13663) );
  NAND2_X1 U14061 ( .A1(n11030), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n10949) );
  NAND2_X1 U14062 ( .A1(n11041), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10948) );
  AND2_X1 U14063 ( .A1(n10949), .A2(n10948), .ZN(n10951) );
  NAND2_X1 U14064 ( .A1(n11027), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10950) );
  OAI211_X1 U14065 ( .C1(n11005), .C2(n13663), .A(n10951), .B(n10950), .ZN(
        n15373) );
  NAND2_X1 U14066 ( .A1(n15372), .A2(n15373), .ZN(n15359) );
  AOI22_X1 U14067 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10293), .B1(
        n10294), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U14068 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10292), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U14069 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12748), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14070 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10295), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10952) );
  NAND4_X1 U14071 ( .A1(n10955), .A2(n10954), .A3(n10953), .A4(n10952), .ZN(
        n10961) );
  AOI22_X1 U14072 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12697), .B1(
        n10903), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U14073 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U14074 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10301), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U14075 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10262), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10956) );
  NAND4_X1 U14076 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n10960) );
  OR2_X1 U14077 ( .A1(n10961), .A2(n10960), .ZN(n13614) );
  NAND2_X1 U14078 ( .A1(n10962), .A2(n13614), .ZN(n10965) );
  AOI22_X1 U14079 ( .A1(n11030), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U14080 ( .A1(n10862), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U14081 ( .A1(n11030), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U14082 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10292), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U14083 ( .A1(n10294), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U14084 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U14085 ( .A1(n12749), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10967) );
  NAND4_X1 U14086 ( .A1(n10970), .A2(n10969), .A3(n10968), .A4(n10967), .ZN(
        n10976) );
  AOI22_X1 U14087 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U14088 ( .A1(n10249), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U14089 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U14090 ( .A1(n10903), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10971) );
  NAND4_X1 U14091 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10975) );
  NOR2_X1 U14092 ( .A1(n10976), .A2(n10975), .ZN(n12668) );
  OR2_X1 U14093 ( .A1(n11005), .A2(n12668), .ZN(n10978) );
  NAND2_X1 U14094 ( .A1(n11027), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U14095 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10292), .B1(
        n9590), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U14096 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12747), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U14097 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U14098 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10980) );
  NAND4_X1 U14099 ( .A1(n10983), .A2(n10982), .A3(n10981), .A4(n10980), .ZN(
        n10989) );
  AOI22_X1 U14100 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U14101 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U14102 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10917), .B1(
        n10903), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U14103 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12697), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10984) );
  NAND4_X1 U14104 ( .A1(n10987), .A2(n10986), .A3(n10985), .A4(n10984), .ZN(
        n10988) );
  NOR2_X1 U14105 ( .A1(n10989), .A2(n10988), .ZN(n12667) );
  AOI22_X1 U14106 ( .A1(n11030), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U14107 ( .A1(n11027), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10991) );
  OAI211_X1 U14108 ( .C1(n12667), .C2(n11005), .A(n10992), .B(n10991), .ZN(
        n15328) );
  AOI22_X1 U14109 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U14110 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12747), .B1(
        n10294), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U14111 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14112 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10993) );
  NAND4_X1 U14113 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n11002) );
  AOI22_X1 U14114 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14115 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14116 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10302), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14117 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10997) );
  NAND4_X1 U14118 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11001) );
  NOR2_X1 U14119 ( .A1(n11002), .A2(n11001), .ZN(n13892) );
  AOI22_X1 U14120 ( .A1(n11030), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11004) );
  NAND2_X1 U14121 ( .A1(n11027), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11003) );
  OAI211_X1 U14122 ( .C1(n13892), .C2(n11005), .A(n11004), .B(n11003), .ZN(
        n15314) );
  NAND2_X1 U14123 ( .A1(n15313), .A2(n15314), .ZN(n15315) );
  INV_X1 U14124 ( .A(n15315), .ZN(n15300) );
  NAND2_X1 U14125 ( .A1(n11030), .A2(P2_EAX_REG_16__SCAN_IN), .ZN(n11007) );
  NAND2_X1 U14126 ( .A1(n11041), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11006) );
  AND2_X1 U14127 ( .A1(n11007), .A2(n11006), .ZN(n11009) );
  NAND2_X1 U14128 ( .A1(n11027), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U14129 ( .A1(n11009), .A2(n11008), .ZN(n15301) );
  NAND2_X1 U14130 ( .A1(n15300), .A2(n15301), .ZN(n15303) );
  AOI22_X1 U14131 ( .A1(n11030), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U14132 ( .A1(n11027), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U14133 ( .A1(n11030), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11013) );
  NAND2_X1 U14134 ( .A1(n11027), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11012) );
  AOI22_X1 U14135 ( .A1(n11030), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11015) );
  NAND2_X1 U14136 ( .A1(n11027), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11014) );
  NAND2_X1 U14137 ( .A1(n11027), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11017) );
  NAND2_X1 U14138 ( .A1(n11030), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n11016) );
  OAI211_X1 U14139 ( .C1(n11037), .C2(n15261), .A(n11017), .B(n11016), .ZN(
        n15254) );
  AOI22_X1 U14140 ( .A1(n11030), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11019) );
  NAND2_X1 U14141 ( .A1(n11027), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14142 ( .A1(n11030), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11021) );
  NAND2_X1 U14143 ( .A1(n11027), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11020) );
  INV_X1 U14144 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n18962) );
  NAND2_X1 U14145 ( .A1(n11027), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U14146 ( .A1(n11041), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11022) );
  OAI211_X1 U14147 ( .C1(n18962), .C2(n11024), .A(n11023), .B(n11022), .ZN(
        n13200) );
  NAND2_X1 U14148 ( .A1(n13199), .A2(n13200), .ZN(n13198) );
  AOI22_X1 U14149 ( .A1(n11030), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11026) );
  NAND2_X1 U14150 ( .A1(n11027), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11025) );
  AND2_X1 U14151 ( .A1(n11026), .A2(n11025), .ZN(n14912) );
  AOI22_X1 U14152 ( .A1(n11030), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11029) );
  NAND2_X1 U14153 ( .A1(n11027), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U14154 ( .A1(n11027), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11032) );
  NAND2_X1 U14155 ( .A1(n11030), .A2(P2_EAX_REG_26__SCAN_IN), .ZN(n11031) );
  OAI211_X1 U14156 ( .C1(n11037), .C2(n15189), .A(n11032), .B(n11031), .ZN(
        n14897) );
  NAND2_X1 U14157 ( .A1(n11027), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11034) );
  NAND2_X1 U14158 ( .A1(n10861), .A2(P2_EAX_REG_27__SCAN_IN), .ZN(n11033) );
  OAI211_X1 U14159 ( .C1(n11037), .C2(n15173), .A(n11034), .B(n11033), .ZN(
        n13215) );
  NAND2_X1 U14160 ( .A1(n11027), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U14161 ( .A1(n10861), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n11035) );
  OAI211_X1 U14162 ( .C1(n11037), .C2(n15156), .A(n11036), .B(n11035), .ZN(
        n14282) );
  INV_X1 U14163 ( .A(n14282), .ZN(n11040) );
  AOI22_X1 U14164 ( .A1(n11030), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11039) );
  NAND2_X1 U14165 ( .A1(n10862), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11038) );
  AND2_X1 U14166 ( .A1(n11039), .A2(n11038), .ZN(n14882) );
  NAND2_X1 U14167 ( .A1(n9896), .A2(n10002), .ZN(n14284) );
  AOI22_X1 U14168 ( .A1(n10861), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11041), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11043) );
  NAND2_X1 U14169 ( .A1(n10862), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11042) );
  AND2_X1 U14170 ( .A1(n11043), .A2(n11042), .ZN(n12956) );
  AOI222_X1 U14171 ( .A1(n10862), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10861), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11041), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11044) );
  XNOR2_X1 U14172 ( .A(n12955), .B(n11044), .ZN(n15890) );
  INV_X1 U14173 ( .A(n11045), .ZN(n11046) );
  AND2_X1 U14174 ( .A1(n13717), .A2(n11046), .ZN(n16058) );
  INV_X1 U14175 ( .A(n16058), .ZN(n13447) );
  OAI21_X1 U14176 ( .B1(n9584), .B2(n9721), .A(n13447), .ZN(n11047) );
  INV_X1 U14177 ( .A(n15056), .ZN(n11085) );
  NOR2_X1 U14178 ( .A1(n16022), .A2(n16021), .ZN(n16020) );
  INV_X1 U14179 ( .A(n16060), .ZN(n11050) );
  NAND2_X1 U14180 ( .A1(n11075), .A2(n11050), .ZN(n12473) );
  INV_X1 U14181 ( .A(n12473), .ZN(n14207) );
  NOR2_X1 U14182 ( .A1(n13714), .A2(n13713), .ZN(n14202) );
  INV_X1 U14183 ( .A(n14202), .ZN(n13306) );
  NOR2_X1 U14184 ( .A1(n11051), .A2(n13306), .ZN(n14209) );
  NOR2_X1 U14185 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14202), .ZN(
        n14208) );
  INV_X1 U14186 ( .A(n14208), .ZN(n11077) );
  NAND2_X1 U14187 ( .A1(n11052), .A2(n10208), .ZN(n13718) );
  NAND2_X1 U14188 ( .A1(n13718), .A2(n11053), .ZN(n11067) );
  OAI22_X1 U14189 ( .A1(n11054), .A2(n11056), .B1(n10121), .B2(n11055), .ZN(
        n11057) );
  INV_X1 U14190 ( .A(n11057), .ZN(n11064) );
  NAND2_X1 U14191 ( .A1(n11059), .A2(n11058), .ZN(n11060) );
  NAND2_X1 U14192 ( .A1(n11060), .A2(n11054), .ZN(n11062) );
  NAND2_X1 U14193 ( .A1(n11062), .A2(n11061), .ZN(n11063) );
  NAND3_X1 U14194 ( .A1(n11065), .A2(n11064), .A3(n11063), .ZN(n11066) );
  AOI21_X1 U14195 ( .B1(n11067), .B2(n13778), .A(n11066), .ZN(n15398) );
  INV_X1 U14196 ( .A(n10158), .ZN(n13454) );
  NAND2_X1 U14197 ( .A1(n15398), .A2(n13454), .ZN(n11068) );
  NAND2_X1 U14198 ( .A1(n11075), .A2(n11068), .ZN(n12468) );
  NAND2_X1 U14199 ( .A1(n12473), .A2(n12468), .ZN(n13307) );
  OAI211_X1 U14200 ( .C1(n14207), .C2(n14209), .A(n11077), .B(n13307), .ZN(
        n16046) );
  NOR2_X1 U14201 ( .A1(n16047), .A2(n16046), .ZN(n13994) );
  NAND3_X1 U14202 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n13994), .ZN(n14055) );
  NOR2_X1 U14203 ( .A1(n14060), .A2(n14055), .ZN(n16024) );
  NAND2_X1 U14204 ( .A1(n16020), .A2(n16024), .ZN(n15385) );
  NOR2_X1 U14205 ( .A1(n11085), .A2(n15385), .ZN(n15271) );
  AND2_X1 U14206 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U14207 ( .A1(n15271), .A2(n11087), .ZN(n15244) );
  NAND2_X1 U14208 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15220) );
  NOR2_X1 U14209 ( .A1(n15233), .A2(n15220), .ZN(n15208) );
  NAND2_X1 U14210 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15208), .ZN(
        n15196) );
  INV_X1 U14211 ( .A(n15196), .ZN(n11069) );
  NAND2_X1 U14212 ( .A1(n10728), .A2(n11069), .ZN(n15153) );
  NOR2_X1 U14213 ( .A1(n15153), .A2(n15173), .ZN(n15161) );
  NAND3_X1 U14214 ( .A1(n15161), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13072) );
  NOR3_X1 U14215 ( .A1(n13072), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n11070), .ZN(n11073) );
  INV_X1 U14216 ( .A(n15127), .ZN(n14056) );
  NAND2_X1 U14217 ( .A1(n15392), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14268) );
  INV_X1 U14218 ( .A(n14268), .ZN(n11072) );
  OR2_X1 U14219 ( .A1(n12468), .A2(n14202), .ZN(n11076) );
  OR2_X1 U14220 ( .A1(n11075), .A2(n15392), .ZN(n13343) );
  INV_X1 U14221 ( .A(n13307), .ZN(n13344) );
  NOR2_X1 U14222 ( .A1(n12468), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14201) );
  OAI211_X1 U14223 ( .C1(n12473), .C2(n11077), .A(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n14204), .ZN(n11078) );
  NOR2_X1 U14224 ( .A1(n14201), .A2(n11078), .ZN(n16048) );
  NOR2_X1 U14225 ( .A1(n16014), .A2(n16048), .ZN(n13905) );
  AND2_X1 U14226 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11079) );
  NOR2_X1 U14227 ( .A1(n16014), .A2(n11079), .ZN(n11080) );
  NOR2_X1 U14228 ( .A1(n13905), .A2(n11080), .ZN(n14061) );
  NAND2_X1 U14229 ( .A1(n13307), .A2(n14060), .ZN(n11081) );
  NAND2_X1 U14230 ( .A1(n14061), .A2(n11081), .ZN(n16025) );
  INV_X1 U14231 ( .A(n16025), .ZN(n11084) );
  INV_X1 U14232 ( .A(n16020), .ZN(n11082) );
  NAND2_X1 U14233 ( .A1(n13307), .A2(n11082), .ZN(n11083) );
  NAND2_X1 U14234 ( .A1(n11084), .A2(n11083), .ZN(n12469) );
  OR2_X1 U14235 ( .A1(n12469), .A2(n11085), .ZN(n11086) );
  NAND2_X1 U14236 ( .A1(n11086), .A2(n11094), .ZN(n15274) );
  OR2_X1 U14237 ( .A1(n16014), .A2(n11087), .ZN(n11088) );
  AND2_X1 U14238 ( .A1(n15274), .A2(n11088), .ZN(n15246) );
  NAND2_X1 U14239 ( .A1(n15246), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11089) );
  NAND2_X1 U14240 ( .A1(n11094), .A2(n11089), .ZN(n15235) );
  AOI21_X1 U14241 ( .B1(n13307), .B2(n15220), .A(n11090), .ZN(n11091) );
  NAND2_X1 U14242 ( .A1(n15235), .A2(n11091), .ZN(n15207) );
  NAND2_X1 U14243 ( .A1(n15207), .A2(n11094), .ZN(n15200) );
  NAND2_X1 U14244 ( .A1(n11094), .A2(n11092), .ZN(n11093) );
  NAND2_X1 U14245 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11095) );
  OAI21_X1 U14246 ( .B1(n11095), .B2(n15156), .A(n11094), .ZN(n11096) );
  NAND2_X1 U14247 ( .A1(n15174), .A2(n11096), .ZN(n13073) );
  NOR2_X1 U14248 ( .A1(n13344), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11097) );
  OAI21_X1 U14249 ( .B1(n13073), .B2(n11097), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11098) );
  OAI211_X1 U14250 ( .C1(n14271), .C2(n16008), .A(n11099), .B(n11098), .ZN(
        n11100) );
  NAND3_X1 U14251 ( .A1(n11103), .A2(n11102), .A3(n11101), .ZN(P2_U3015) );
  AND2_X2 U14252 ( .A1(n11113), .A2(n13682), .ZN(n12064) );
  AOI22_X1 U14253 ( .A1(n12064), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11325), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11108) );
  AND2_X2 U14254 ( .A1(n13682), .A2(n11111), .ZN(n11298) );
  AOI22_X1 U14255 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U14256 ( .A1(n9653), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11292), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11106) );
  AND2_X4 U14257 ( .A1(n11109), .A2(n11113), .ZN(n11409) );
  AOI22_X1 U14258 ( .A1(n11277), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11117) );
  AND2_X2 U14259 ( .A1(n13682), .A2(n13669), .ZN(n11300) );
  AOI22_X1 U14260 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11115) );
  NAND2_X1 U14261 ( .A1(n12064), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14262 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11122) );
  NAND2_X1 U14263 ( .A1(n11325), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11121) );
  NAND2_X1 U14264 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U14265 ( .A1(n11276), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U14266 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11126) );
  NAND2_X1 U14267 ( .A1(n11277), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U14268 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14269 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11131) );
  NAND2_X1 U14270 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11130) );
  NAND2_X1 U14271 ( .A1(n9653), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11129) );
  NAND2_X1 U14272 ( .A1(n11292), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11128) );
  NAND2_X1 U14273 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11135) );
  NAND2_X1 U14274 ( .A1(n11326), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14275 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U14276 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14277 ( .A1(n11612), .A2(n11249), .ZN(n11266) );
  NAND2_X1 U14278 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11143) );
  NAND2_X1 U14279 ( .A1(n11276), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U14280 ( .A1(n11277), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11141) );
  NAND2_X1 U14281 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11140) );
  NAND2_X1 U14282 ( .A1(n12064), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U14283 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11146) );
  NAND2_X1 U14284 ( .A1(n11325), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11145) );
  NAND2_X1 U14285 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11144) );
  NAND2_X1 U14286 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11151) );
  NAND2_X1 U14287 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11150) );
  NAND2_X1 U14288 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11149) );
  NAND2_X1 U14289 ( .A1(n11292), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11148) );
  NAND2_X1 U14290 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11155) );
  NAND2_X1 U14291 ( .A1(n11326), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11154) );
  NAND2_X1 U14292 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11153) );
  NAND2_X1 U14293 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11152) );
  AOI22_X1 U14294 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n9653), .ZN(n11163) );
  AOI22_X1 U14295 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11325), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14296 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11292), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11161) );
  AOI22_X1 U14297 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11160) );
  AOI22_X1 U14298 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14299 ( .A1(n11277), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11276), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14300 ( .A1(n11326), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14301 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14302 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11326), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11173) );
  AOI22_X1 U14303 ( .A1(n11276), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11223), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14304 ( .A1(n11277), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14305 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11170) );
  NAND4_X1 U14306 ( .A1(n11173), .A2(n11172), .A3(n11171), .A4(n11170), .ZN(
        n11179) );
  AOI22_X1 U14307 ( .A1(n12064), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11325), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14308 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11332), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14309 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11175) );
  AOI22_X1 U14310 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11292), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11174) );
  NAND4_X1 U14311 ( .A1(n11177), .A2(n11176), .A3(n11175), .A4(n11174), .ZN(
        n11178) );
  NAND2_X1 U14312 ( .A1(n11248), .A2(n11254), .ZN(n11181) );
  AOI22_X1 U14313 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14314 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14315 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11326), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11182) );
  NAND3_X1 U14316 ( .A1(n11184), .A2(n11183), .A3(n11182), .ZN(n11187) );
  AOI22_X1 U14317 ( .A1(n11277), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14318 ( .A1(n12064), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11325), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14319 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11989), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14320 ( .A1(n11276), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11278), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14321 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11292), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11188) );
  NAND2_X2 U14322 ( .A1(n11193), .A2(n11192), .ZN(n19983) );
  NAND2_X1 U14323 ( .A1(n9993), .A2(n9599), .ZN(n11195) );
  NAND2_X2 U14324 ( .A1(n11242), .A2(n11249), .ZN(n11244) );
  NAND2_X1 U14325 ( .A1(n11244), .A2(n19983), .ZN(n11194) );
  NAND2_X1 U14326 ( .A1(n12064), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11201) );
  NAND2_X1 U14327 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11200) );
  NAND2_X1 U14328 ( .A1(n11325), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11199) );
  NAND2_X1 U14329 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11198) );
  NAND2_X1 U14330 ( .A1(n11277), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11204) );
  NAND2_X1 U14331 ( .A1(n11276), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11203) );
  NAND2_X1 U14332 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11202) );
  NAND3_X1 U14333 ( .A1(n11204), .A2(n11203), .A3(n11202), .ZN(n11205) );
  NAND2_X1 U14334 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11209) );
  NAND2_X1 U14335 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11208) );
  NAND2_X1 U14336 ( .A1(n11292), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11207) );
  NAND2_X1 U14337 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11214) );
  NAND2_X1 U14338 ( .A1(n11275), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11213) );
  NAND2_X1 U14339 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11212) );
  NAND2_X1 U14340 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11211) );
  AND4_X2 U14341 ( .A1(n11214), .A2(n11213), .A3(n11212), .A4(n11211), .ZN(
        n11215) );
  NAND4_X4 U14342 ( .A1(n11218), .A2(n11217), .A3(n11216), .A4(n11215), .ZN(
        n12501) );
  NAND2_X1 U14343 ( .A1(n12064), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11222) );
  NAND2_X1 U14344 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11221) );
  NAND2_X1 U14345 ( .A1(n11325), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11220) );
  NAND2_X1 U14346 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11219) );
  NAND2_X1 U14347 ( .A1(n11276), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11227) );
  NAND2_X1 U14348 ( .A1(n11223), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11226) );
  NAND2_X1 U14349 ( .A1(n11277), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11225) );
  NAND2_X1 U14350 ( .A1(n11278), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11224) );
  NAND2_X1 U14351 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11231) );
  NAND2_X1 U14352 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11230) );
  NAND2_X1 U14353 ( .A1(n11989), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11229) );
  NAND2_X1 U14354 ( .A1(n11292), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11228) );
  NAND2_X1 U14355 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11235) );
  NAND2_X1 U14356 ( .A1(n11326), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11234) );
  NAND2_X1 U14357 ( .A1(n11300), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11233) );
  NAND2_X1 U14358 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11232) );
  NAND2_X1 U14359 ( .A1(n9640), .A2(n14302), .ZN(n11241) );
  NAND2_X1 U14360 ( .A1(n19983), .A2(n12501), .ZN(n11240) );
  NAND2_X1 U14361 ( .A1(n11241), .A2(n11240), .ZN(n13021) );
  NAND2_X1 U14362 ( .A1(n12997), .A2(n19979), .ZN(n13398) );
  OAI211_X1 U14363 ( .C1(n11243), .C2(n13251), .A(n13385), .B(n13398), .ZN(
        n11246) );
  NAND2_X1 U14364 ( .A1(n11255), .A2(n11270), .ZN(n11247) );
  NAND2_X1 U14365 ( .A1(n11256), .A2(n19994), .ZN(n11250) );
  NAND2_X1 U14366 ( .A1(n11267), .A2(n11250), .ZN(n13023) );
  XNOR2_X1 U14367 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12596) );
  INV_X1 U14368 ( .A(n13386), .ZN(n11260) );
  NAND2_X1 U14369 ( .A1(n11254), .A2(n11270), .ZN(n13004) );
  OAI21_X1 U14370 ( .B1(n14300), .B2(n12596), .A(n13019), .ZN(n11261) );
  NOR2_X1 U14371 ( .A1(n13013), .A2(n11261), .ZN(n11317) );
  NAND2_X1 U14372 ( .A1(n13038), .A2(n11317), .ZN(n11262) );
  NAND2_X2 U14373 ( .A1(n11262), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11357) );
  MUX2_X1 U14374 ( .A(n12104), .B(n15583), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11264) );
  OAI21_X2 U14375 ( .B1(n11357), .B2(n11263), .A(n11264), .ZN(n11321) );
  NAND3_X1 U14376 ( .A1(n12998), .A2(n14796), .A3(n19979), .ZN(n11273) );
  INV_X1 U14377 ( .A(n14800), .ZN(n20625) );
  NOR2_X1 U14378 ( .A1(n20625), .A2(n20790), .ZN(n11272) );
  INV_X1 U14379 ( .A(n14302), .ZN(n14305) );
  NAND2_X1 U14380 ( .A1(n11266), .A2(n19987), .ZN(n11269) );
  INV_X1 U14381 ( .A(n11267), .ZN(n11268) );
  INV_X1 U14382 ( .A(n13251), .ZN(n20642) );
  AOI22_X1 U14383 ( .A1(n13249), .A2(n11269), .B1(n11268), .B2(n20642), .ZN(
        n11271) );
  INV_X1 U14384 ( .A(n11258), .ZN(n13671) );
  OR2_X1 U14385 ( .A1(n13671), .A2(n11270), .ZN(n13034) );
  NAND2_X1 U14386 ( .A1(n11265), .A2(n10015), .ZN(n11320) );
  AOI22_X1 U14387 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11275), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14388 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14389 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14390 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11279) );
  NAND4_X1 U14391 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11291) );
  AOI22_X1 U14392 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11289) );
  BUF_X1 U14394 ( .A(n11332), .Z(n11283) );
  AOI22_X1 U14395 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11288) );
  BUF_X1 U14396 ( .A(n11297), .Z(n11285) );
  AOI22_X1 U14397 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14398 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11286) );
  NAND4_X1 U14399 ( .A1(n11289), .A2(n11288), .A3(n11287), .A4(n11286), .ZN(
        n11290) );
  NAND2_X1 U14400 ( .A1(n11243), .A2(n11515), .ZN(n11309) );
  NOR2_X1 U14401 ( .A1(n11408), .A2(n11515), .ZN(n11381) );
  AOI22_X1 U14402 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14403 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14404 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14405 ( .A1(n11363), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11293) );
  NAND4_X1 U14406 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n11306) );
  AOI22_X1 U14407 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14408 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14410 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14411 ( .A1(n11327), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11300), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11301) );
  NAND4_X1 U14412 ( .A1(n11304), .A2(n11303), .A3(n11302), .A4(n11301), .ZN(
        n11305) );
  MUX2_X1 U14413 ( .A(n11512), .B(n11381), .S(n11395), .Z(n11307) );
  INV_X1 U14414 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11311) );
  AOI21_X1 U14415 ( .B1(n12997), .B2(n11395), .A(n20790), .ZN(n11310) );
  NAND2_X1 U14416 ( .A1(n12997), .A2(n19987), .ZN(n11396) );
  OAI21_X1 U14417 ( .B1(n13251), .B2(n11395), .A(n11396), .ZN(n11312) );
  INV_X1 U14418 ( .A(n11312), .ZN(n11313) );
  OAI21_X1 U14419 ( .B1(n11611), .B2(n11541), .A(n11313), .ZN(n13432) );
  NAND2_X1 U14420 ( .A1(n13432), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13433) );
  INV_X1 U14421 ( .A(n15583), .ZN(n15576) );
  NAND2_X1 U14422 ( .A1(n15576), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11349) );
  NAND2_X1 U14423 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11355) );
  OAI21_X1 U14424 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11355), .ZN(n20287) );
  OR2_X1 U14425 ( .A1(n12104), .A2(n20287), .ZN(n11315) );
  AND2_X1 U14426 ( .A1(n11349), .A2(n11315), .ZN(n11316) );
  OAI21_X2 U14427 ( .B1(n11357), .B2(n11314), .A(n11316), .ZN(n11319) );
  INV_X1 U14428 ( .A(n11317), .ZN(n11318) );
  XNOR2_X2 U14429 ( .A(n11319), .B(n11348), .ZN(n20071) );
  INV_X1 U14430 ( .A(n20071), .ZN(n11323) );
  INV_X1 U14431 ( .A(n11408), .ZN(n11339) );
  AOI22_X1 U14432 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14433 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14434 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14435 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11328) );
  NAND4_X1 U14436 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11338) );
  AOI22_X1 U14437 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14438 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14439 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14440 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11333) );
  NAND4_X1 U14441 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n11337) );
  NAND2_X1 U14442 ( .A1(n11386), .A2(n19979), .ZN(n11344) );
  XNOR2_X1 U14443 ( .A(n11395), .B(n11394), .ZN(n11341) );
  OAI211_X1 U14444 ( .C1(n11341), .C2(n13251), .A(n11340), .B(n19994), .ZN(
        n11342) );
  INV_X1 U14445 ( .A(n11342), .ZN(n11343) );
  NAND2_X1 U14446 ( .A1(n11344), .A2(n11343), .ZN(n11345) );
  NAND2_X1 U14447 ( .A1(n13489), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13490) );
  INV_X1 U14448 ( .A(n11345), .ZN(n11346) );
  OR2_X1 U14449 ( .A1(n13433), .A2(n11346), .ZN(n11347) );
  INV_X1 U14450 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19954) );
  INV_X1 U14451 ( .A(n11348), .ZN(n11351) );
  NAND2_X1 U14452 ( .A1(n11349), .A2(n11314), .ZN(n11350) );
  NAND2_X1 U14453 ( .A1(n11351), .A2(n11350), .ZN(n11352) );
  INV_X1 U14454 ( .A(n11355), .ZN(n11354) );
  NAND2_X1 U14455 ( .A1(n11354), .A2(n15558), .ZN(n20328) );
  NAND2_X1 U14456 ( .A1(n11355), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11356) );
  NAND2_X1 U14457 ( .A1(n15576), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11359) );
  AOI22_X1 U14458 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14459 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14460 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14461 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11364) );
  NAND4_X1 U14462 ( .A1(n11367), .A2(n11366), .A3(n11365), .A4(n11364), .ZN(
        n11375) );
  AOI22_X1 U14463 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14464 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14465 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14466 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11370) );
  NAND4_X1 U14467 ( .A1(n11373), .A2(n11372), .A3(n11371), .A4(n11370), .ZN(
        n11374) );
  INV_X1 U14468 ( .A(n11407), .ZN(n11382) );
  AOI22_X1 U14469 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11382), .B2(n11376), .ZN(n11377) );
  INV_X1 U14470 ( .A(n11512), .ZN(n11380) );
  INV_X1 U14471 ( .A(n11381), .ZN(n11385) );
  NAND2_X1 U14472 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U14473 ( .A1(n11382), .A2(n11394), .ZN(n11383) );
  INV_X1 U14474 ( .A(n11387), .ZN(n11388) );
  NOR2_X1 U14475 ( .A1(n11389), .A2(n11388), .ZN(n11390) );
  NAND2_X1 U14476 ( .A1(n11395), .A2(n11394), .ZN(n11427) );
  XNOR2_X1 U14477 ( .A(n11427), .B(n11426), .ZN(n11398) );
  INV_X1 U14478 ( .A(n11396), .ZN(n11397) );
  AOI21_X1 U14479 ( .B1(n11398), .B2(n20642), .A(n11397), .ZN(n11399) );
  NAND2_X1 U14480 ( .A1(n11400), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11401) );
  INV_X1 U14481 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19933) );
  NAND3_X1 U14482 ( .A1(n20363), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20203) );
  INV_X1 U14483 ( .A(n20203), .ZN(n11402) );
  NAND2_X1 U14484 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11402), .ZN(
        n20201) );
  NAND2_X1 U14485 ( .A1(n20363), .A2(n20201), .ZN(n11403) );
  NOR3_X1 U14486 ( .A1(n20363), .A2(n15558), .A3(n11542), .ZN(n20500) );
  NAND2_X1 U14487 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20500), .ZN(
        n20494) );
  NAND2_X1 U14488 ( .A1(n11403), .A2(n20494), .ZN(n20234) );
  OAI22_X1 U14489 ( .A1(n12104), .A2(n20234), .B1(n15583), .B2(n20363), .ZN(
        n11404) );
  INV_X1 U14490 ( .A(n11404), .ZN(n11405) );
  NAND2_X1 U14491 ( .A1(n20233), .A2(n20790), .ZN(n11421) );
  AOI22_X1 U14492 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14493 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14494 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14495 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11410) );
  NAND4_X1 U14496 ( .A1(n11413), .A2(n11412), .A3(n11411), .A4(n11410), .ZN(
        n11419) );
  AOI22_X1 U14497 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14498 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14499 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14500 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11414) );
  NAND4_X1 U14501 ( .A1(n11417), .A2(n11416), .A3(n11415), .A4(n11414), .ZN(
        n11418) );
  AOI22_X1 U14502 ( .A1(n11555), .A2(n11467), .B1(n11581), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11420) );
  NAND2_X1 U14503 ( .A1(n11424), .A2(n19961), .ZN(n11425) );
  OR2_X1 U14504 ( .A1(n11624), .A2(n11541), .ZN(n11431) );
  NAND2_X1 U14505 ( .A1(n11427), .A2(n11426), .ZN(n11470) );
  INV_X1 U14506 ( .A(n11467), .ZN(n11428) );
  XNOR2_X1 U14507 ( .A(n11470), .B(n11428), .ZN(n11429) );
  NAND2_X1 U14508 ( .A1(n11429), .A2(n20642), .ZN(n11430) );
  NAND2_X1 U14509 ( .A1(n11431), .A2(n11430), .ZN(n13602) );
  NAND2_X1 U14510 ( .A1(n11432), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11433) );
  AOI22_X1 U14511 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14512 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12076), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14513 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14514 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12075), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11434) );
  NAND4_X1 U14515 ( .A1(n11437), .A2(n11436), .A3(n11435), .A4(n11434), .ZN(
        n11443) );
  AOI22_X1 U14516 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12043), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14517 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11284), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14518 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14519 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11438) );
  NAND4_X1 U14520 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n11442) );
  NAND2_X1 U14521 ( .A1(n11555), .A2(n11468), .ZN(n11445) );
  NAND2_X1 U14522 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11444) );
  NAND2_X1 U14523 ( .A1(n11445), .A2(n11444), .ZN(n11453) );
  INV_X1 U14524 ( .A(n11541), .ZN(n11511) );
  NAND2_X1 U14525 ( .A1(n11599), .A2(n11511), .ZN(n11449) );
  NAND2_X1 U14526 ( .A1(n11470), .A2(n11467), .ZN(n11446) );
  XNOR2_X1 U14527 ( .A(n11446), .B(n11468), .ZN(n11447) );
  NAND2_X1 U14528 ( .A1(n11447), .A2(n20642), .ZN(n11448) );
  NAND2_X1 U14529 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  INV_X1 U14530 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19922) );
  NAND2_X1 U14531 ( .A1(n11450), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11451) );
  AOI22_X1 U14532 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14533 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14534 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14535 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11455) );
  NAND4_X1 U14536 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(
        n11464) );
  AOI22_X1 U14537 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14538 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14539 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14540 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11459) );
  NAND4_X1 U14541 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n11463) );
  NAND2_X1 U14542 ( .A1(n11555), .A2(n11494), .ZN(n11466) );
  NAND2_X1 U14543 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11465) );
  NAND2_X1 U14544 ( .A1(n11466), .A2(n11465), .ZN(n11487) );
  AND2_X1 U14545 ( .A1(n11468), .A2(n11467), .ZN(n11469) );
  NAND2_X1 U14546 ( .A1(n11470), .A2(n11469), .ZN(n11496) );
  XNOR2_X1 U14547 ( .A(n11496), .B(n11494), .ZN(n11471) );
  NAND2_X1 U14548 ( .A1(n11471), .A2(n20642), .ZN(n11472) );
  INV_X1 U14549 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20699) );
  NAND2_X1 U14550 ( .A1(n11473), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11474) );
  AOI22_X1 U14551 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14552 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14553 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14554 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11475) );
  NAND4_X1 U14555 ( .A1(n11478), .A2(n11477), .A3(n11476), .A4(n11475), .ZN(
        n11484) );
  AOI22_X1 U14556 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14557 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14558 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14559 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14560 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11483) );
  NAND2_X1 U14561 ( .A1(n11555), .A2(n11505), .ZN(n11486) );
  NAND2_X1 U14562 ( .A1(n11581), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11485) );
  OR2_X1 U14563 ( .A1(n11491), .A2(n11490), .ZN(n11493) );
  NAND3_X1 U14564 ( .A1(n9668), .A2(n11511), .A3(n11653), .ZN(n11499) );
  INV_X1 U14565 ( .A(n11494), .ZN(n11495) );
  OR2_X1 U14566 ( .A1(n11496), .A2(n11495), .ZN(n11504) );
  XNOR2_X1 U14567 ( .A(n11504), .B(n11505), .ZN(n11497) );
  NAND2_X1 U14568 ( .A1(n11497), .A2(n20642), .ZN(n11498) );
  INV_X1 U14569 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15855) );
  NAND2_X1 U14570 ( .A1(n15751), .A2(n15855), .ZN(n11500) );
  INV_X1 U14571 ( .A(n15751), .ZN(n11501) );
  NAND2_X1 U14572 ( .A1(n11501), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11502) );
  AOI22_X1 U14573 ( .A1(n11555), .A2(n11515), .B1(n11581), .B2(
        P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11503) );
  OR2_X1 U14574 ( .A1(n11654), .A2(n11541), .ZN(n11509) );
  INV_X1 U14575 ( .A(n11504), .ZN(n11506) );
  NAND2_X1 U14576 ( .A1(n11506), .A2(n11505), .ZN(n11514) );
  XNOR2_X1 U14577 ( .A(n11514), .B(n11515), .ZN(n11507) );
  NAND2_X1 U14578 ( .A1(n11507), .A2(n20642), .ZN(n11508) );
  NAND2_X1 U14579 ( .A1(n11509), .A2(n11508), .ZN(n11510) );
  OR2_X1 U14580 ( .A1(n11510), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15746) );
  NAND2_X1 U14581 ( .A1(n11510), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15745) );
  AND2_X1 U14582 ( .A1(n11512), .A2(n11511), .ZN(n11513) );
  INV_X1 U14583 ( .A(n11514), .ZN(n11516) );
  NAND3_X1 U14584 ( .A1(n11516), .A2(n20642), .A3(n11515), .ZN(n11517) );
  NAND2_X1 U14585 ( .A1(n11528), .A2(n11517), .ZN(n14003) );
  OR2_X1 U14586 ( .A1(n14003), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11518) );
  NAND2_X1 U14587 ( .A1(n14003), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11519) );
  INV_X1 U14588 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14025) );
  NAND2_X1 U14589 ( .A1(n9597), .A2(n14025), .ZN(n11520) );
  INV_X1 U14590 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15797) );
  INV_X1 U14591 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11521) );
  INV_X1 U14592 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12552) );
  INV_X1 U14593 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15814) );
  NAND2_X1 U14594 ( .A1(n11528), .A2(n15814), .ZN(n11523) );
  NAND2_X1 U14595 ( .A1(n14625), .A2(n11523), .ZN(n14641) );
  NAND2_X1 U14596 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11524) );
  AND2_X1 U14597 ( .A1(n11528), .A2(n11524), .ZN(n14632) );
  NOR2_X1 U14598 ( .A1(n14641), .A2(n14632), .ZN(n14624) );
  INV_X1 U14599 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U14600 ( .A1(n11528), .A2(n14782), .ZN(n14639) );
  INV_X1 U14601 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15809) );
  NAND2_X1 U14602 ( .A1(n11528), .A2(n15809), .ZN(n11525) );
  AND2_X1 U14603 ( .A1(n14639), .A2(n11525), .ZN(n11526) );
  NAND2_X1 U14604 ( .A1(n14624), .A2(n11526), .ZN(n14609) );
  OR2_X1 U14605 ( .A1(n11528), .A2(n15809), .ZN(n11527) );
  NAND2_X1 U14606 ( .A1(n14625), .A2(n11527), .ZN(n11531) );
  NOR2_X1 U14607 ( .A1(n11528), .A2(n15797), .ZN(n14613) );
  NOR2_X1 U14608 ( .A1(n11531), .A2(n14613), .ZN(n15710) );
  XNOR2_X1 U14609 ( .A(n11528), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14615) );
  NAND2_X1 U14610 ( .A1(n11528), .A2(n15797), .ZN(n14614) );
  NAND2_X1 U14611 ( .A1(n14615), .A2(n14614), .ZN(n11529) );
  INV_X1 U14612 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14634) );
  INV_X1 U14613 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15738) );
  AND3_X1 U14614 ( .A1(n14634), .A2(n15738), .A3(n14782), .ZN(n11530) );
  NOR2_X1 U14615 ( .A1(n9597), .A2(n11530), .ZN(n14623) );
  XNOR2_X1 U14616 ( .A(n15735), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14603) );
  INV_X1 U14617 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20747) );
  INV_X1 U14618 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14751) );
  INV_X1 U14619 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14743) );
  NAND2_X1 U14620 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11533) );
  INV_X1 U14621 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14703) );
  INV_X1 U14622 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14723) );
  NAND2_X1 U14623 ( .A1(n14703), .A2(n14723), .ZN(n14254) );
  NAND3_X1 U14624 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14698) );
  INV_X1 U14625 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13064) );
  NAND2_X1 U14626 ( .A1(n11536), .A2(n15735), .ZN(n14551) );
  NAND2_X1 U14627 ( .A1(n14533), .A2(n14551), .ZN(n11537) );
  INV_X1 U14628 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14682) );
  INV_X1 U14629 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14690) );
  NAND2_X1 U14630 ( .A1(n14682), .A2(n14690), .ZN(n14678) );
  NOR2_X2 U14631 ( .A1(n14535), .A2(n9998), .ZN(n14525) );
  NAND2_X1 U14632 ( .A1(n14525), .A2(n9649), .ZN(n14514) );
  AND2_X1 U14633 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13066) );
  AND2_X1 U14634 ( .A1(n15735), .A2(n13066), .ZN(n11538) );
  INV_X1 U14635 ( .A(n13023), .ZN(n11540) );
  NAND2_X1 U14636 ( .A1(n14796), .A2(n12997), .ZN(n11539) );
  MUX2_X1 U14637 ( .A(n11542), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11553) );
  NAND2_X1 U14638 ( .A1(n20416), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11556) );
  NAND2_X1 U14639 ( .A1(n11553), .A2(n11552), .ZN(n11544) );
  NAND2_X1 U14640 ( .A1(n11542), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11543) );
  NAND2_X1 U14641 ( .A1(n11544), .A2(n11543), .ZN(n11566) );
  MUX2_X1 U14642 ( .A(n15558), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11565) );
  NAND2_X1 U14643 ( .A1(n11566), .A2(n11565), .ZN(n11546) );
  NAND2_X1 U14644 ( .A1(n15558), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11545) );
  NOR2_X1 U14645 ( .A1(n11104), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14646 ( .A1(n11548), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11549) );
  NAND2_X1 U14647 ( .A1(n11577), .A2(n12443), .ZN(n11590) );
  NAND2_X1 U14648 ( .A1(n12443), .A2(n11555), .ZN(n11588) );
  XNOR2_X1 U14649 ( .A(n11551), .B(n11550), .ZN(n12440) );
  XNOR2_X1 U14650 ( .A(n11553), .B(n11552), .ZN(n12438) );
  AOI22_X1 U14651 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11255), .B1(n11555), 
        .B2(n19979), .ZN(n11564) );
  INV_X1 U14652 ( .A(n11564), .ZN(n11554) );
  NOR2_X1 U14653 ( .A1(n12438), .A2(n11554), .ZN(n11562) );
  INV_X1 U14654 ( .A(n11555), .ZN(n11572) );
  OAI21_X1 U14655 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20416), .A(
        n11556), .ZN(n11558) );
  NOR2_X1 U14656 ( .A1(n11572), .A2(n11558), .ZN(n11561) );
  NAND2_X1 U14657 ( .A1(n11255), .A2(n12501), .ZN(n11557) );
  NAND2_X1 U14658 ( .A1(n11557), .A2(n11253), .ZN(n11571) );
  INV_X1 U14659 ( .A(n11558), .ZN(n11559) );
  OAI211_X1 U14660 ( .C1(n12997), .C2(n11244), .A(n11571), .B(n11559), .ZN(
        n11560) );
  OAI21_X1 U14661 ( .B1(n11577), .B2(n11561), .A(n11560), .ZN(n11563) );
  NAND2_X1 U14662 ( .A1(n11562), .A2(n11563), .ZN(n11570) );
  NAND2_X1 U14663 ( .A1(n11564), .A2(n19979), .ZN(n11583) );
  OAI211_X1 U14664 ( .C1(n11564), .C2(n11563), .A(n12438), .B(n11583), .ZN(
        n11569) );
  XNOR2_X1 U14665 ( .A(n11566), .B(n11565), .ZN(n12439) );
  NAND2_X1 U14666 ( .A1(n11581), .A2(n12439), .ZN(n11567) );
  OAI211_X1 U14667 ( .C1(n11572), .C2(n12439), .A(n11567), .B(n11571), .ZN(
        n11568) );
  NAND3_X1 U14668 ( .A1(n11570), .A2(n11569), .A3(n11568), .ZN(n11574) );
  AOI22_X1 U14669 ( .A1(n11575), .A2(n12440), .B1(n11574), .B2(n11573), .ZN(
        n11576) );
  AOI21_X1 U14670 ( .B1(n11577), .B2(n12440), .A(n11576), .ZN(n11585) );
  INV_X1 U14671 ( .A(n12441), .ZN(n11580) );
  NOR2_X1 U14672 ( .A1(n11581), .A2(n11580), .ZN(n11584) );
  NAND2_X1 U14673 ( .A1(n11581), .A2(n12441), .ZN(n11582) );
  OAI22_X1 U14674 ( .A1(n11585), .A2(n11584), .B1(n11583), .B2(n11582), .ZN(
        n11586) );
  AOI21_X1 U14675 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20790), .A(
        n11586), .ZN(n11587) );
  NAND2_X1 U14676 ( .A1(n11588), .A2(n11587), .ZN(n11589) );
  NAND3_X1 U14677 ( .A1(n13015), .A2(n11245), .A3(n14301), .ZN(n15564) );
  NAND2_X1 U14678 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11626) );
  INV_X1 U14679 ( .A(n11626), .ZN(n11591) );
  INV_X1 U14680 ( .A(n11637), .ZN(n11639) );
  INV_X1 U14681 ( .A(n11592), .ZN(n11629) );
  INV_X1 U14682 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11593) );
  NAND2_X1 U14683 ( .A1(n11629), .A2(n11593), .ZN(n11594) );
  NAND2_X1 U14684 ( .A1(n11639), .A2(n11594), .ZN(n19915) );
  INV_X1 U14685 ( .A(n11633), .ZN(n11617) );
  INV_X1 U14686 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13683) );
  NAND2_X1 U14687 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11596) );
  NAND2_X1 U14688 ( .A1(n12096), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11595) );
  OAI211_X1 U14689 ( .C1(n11617), .C2(n13683), .A(n11596), .B(n11595), .ZN(
        n11597) );
  NOR2_X4 U14690 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12496) );
  MUX2_X1 U14691 ( .A(n19915), .B(n11597), .S(n12087), .Z(n11598) );
  AOI21_X1 U14692 ( .B1(n11599), .B2(n11783), .A(n11598), .ZN(n13543) );
  INV_X1 U14693 ( .A(n13543), .ZN(n11636) );
  INV_X1 U14694 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11601) );
  XNOR2_X1 U14695 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13950) );
  AOI21_X1 U14696 ( .B1(n12496), .B2(n13950), .A(n12095), .ZN(n11600) );
  OAI21_X1 U14697 ( .B1(n12090), .B2(n11601), .A(n11600), .ZN(n11602) );
  AOI21_X1 U14698 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n11633), .A(
        n11602), .ZN(n11603) );
  NAND2_X1 U14699 ( .A1(n12095), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11623) );
  XNOR2_X2 U14700 ( .A(n11606), .B(n11605), .ZN(n13691) );
  NAND2_X1 U14701 ( .A1(n13691), .A2(n11783), .ZN(n11610) );
  INV_X1 U14702 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11607) );
  INV_X1 U14703 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13488) );
  OAI22_X1 U14704 ( .A1(n12090), .A2(n11607), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13488), .ZN(n11608) );
  AOI21_X1 U14705 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11633), .A(
        n11608), .ZN(n11609) );
  NAND2_X1 U14706 ( .A1(n11610), .A2(n11609), .ZN(n13361) );
  NAND2_X1 U14707 ( .A1(n11611), .A2(n11612), .ZN(n11613) );
  NAND2_X1 U14708 ( .A1(n11613), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13353) );
  NAND2_X1 U14709 ( .A1(n12096), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U14710 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11615) );
  OAI211_X1 U14711 ( .C1(n11617), .C2(n11263), .A(n11616), .B(n11615), .ZN(
        n11618) );
  AOI21_X1 U14712 ( .B1(n11614), .B2(n11783), .A(n11618), .ZN(n11619) );
  OR2_X1 U14713 ( .A1(n13353), .A2(n11619), .ZN(n13354) );
  INV_X1 U14714 ( .A(n11619), .ZN(n13355) );
  OR2_X1 U14715 ( .A1(n13355), .A2(n12087), .ZN(n11620) );
  NAND2_X1 U14716 ( .A1(n13354), .A2(n11620), .ZN(n13360) );
  NAND2_X1 U14717 ( .A1(n13361), .A2(n13360), .ZN(n13502) );
  NAND2_X2 U14718 ( .A1(n13500), .A2(n11623), .ZN(n13542) );
  INV_X1 U14719 ( .A(n11624), .ZN(n11625) );
  NAND2_X1 U14720 ( .A1(n11625), .A2(n11783), .ZN(n11635) );
  INV_X1 U14721 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11631) );
  INV_X1 U14722 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11627) );
  NAND2_X1 U14723 ( .A1(n11627), .A2(n11626), .ZN(n11628) );
  NAND2_X1 U14724 ( .A1(n11629), .A2(n11628), .ZN(n13870) );
  AOI22_X1 U14725 ( .A1(n13870), .A2(n12496), .B1(n12095), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11630) );
  OAI21_X1 U14726 ( .B1(n12090), .B2(n11631), .A(n11630), .ZN(n11632) );
  AOI21_X1 U14727 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11633), .A(
        n11632), .ZN(n11634) );
  NAND2_X1 U14728 ( .A1(n11635), .A2(n11634), .ZN(n13541) );
  NAND3_X1 U14729 ( .A1(n11636), .A2(n13542), .A3(n13541), .ZN(n13539) );
  INV_X1 U14730 ( .A(n13539), .ZN(n11645) );
  INV_X1 U14731 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13598) );
  INV_X1 U14732 ( .A(n11646), .ZN(n11648) );
  INV_X1 U14733 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11638) );
  NAND2_X1 U14734 ( .A1(n11639), .A2(n11638), .ZN(n11640) );
  NAND2_X1 U14735 ( .A1(n11648), .A2(n11640), .ZN(n19812) );
  AOI22_X1 U14736 ( .A1(n19812), .A2(n12496), .B1(n12095), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11641) );
  OAI21_X1 U14737 ( .B1(n12090), .B2(n13598), .A(n11641), .ZN(n11642) );
  AOI21_X1 U14738 ( .B1(n11643), .B2(n11783), .A(n11642), .ZN(n13596) );
  INV_X1 U14739 ( .A(n13596), .ZN(n11644) );
  INV_X1 U14740 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11651) );
  INV_X1 U14741 ( .A(n11656), .ZN(n11658) );
  INV_X1 U14742 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14743 ( .A1(n11648), .A2(n11647), .ZN(n11649) );
  NAND2_X1 U14744 ( .A1(n11658), .A2(n11649), .ZN(n19805) );
  AOI22_X1 U14745 ( .A1(n19805), .A2(n12496), .B1(n12095), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11650) );
  OAI21_X1 U14746 ( .B1(n12090), .B2(n11651), .A(n11650), .ZN(n11652) );
  INV_X1 U14747 ( .A(n11654), .ZN(n11655) );
  NAND2_X1 U14748 ( .A1(n11655), .A2(n11783), .ZN(n11665) );
  INV_X1 U14749 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11662) );
  INV_X1 U14750 ( .A(n11681), .ZN(n11660) );
  INV_X1 U14751 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11657) );
  NAND2_X1 U14752 ( .A1(n11658), .A2(n11657), .ZN(n11659) );
  NAND2_X1 U14753 ( .A1(n11660), .A2(n11659), .ZN(n19791) );
  AOI22_X1 U14754 ( .A1(n19791), .A2(n12496), .B1(n12095), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14755 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14756 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14757 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14758 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11666) );
  NAND4_X1 U14759 ( .A1(n11669), .A2(n11668), .A3(n11667), .A4(n11666), .ZN(
        n11675) );
  AOI22_X1 U14760 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14761 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14762 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14763 ( .A1(n12073), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11670) );
  NAND4_X1 U14764 ( .A1(n11673), .A2(n11672), .A3(n11671), .A4(n11670), .ZN(
        n11674) );
  OAI21_X1 U14765 ( .B1(n11675), .B2(n11674), .A(n11783), .ZN(n11679) );
  NAND2_X1 U14766 ( .A1(n12096), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11678) );
  XNOR2_X1 U14767 ( .A(n11681), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n19777) );
  NAND2_X1 U14768 ( .A1(n19777), .A2(n12496), .ZN(n11677) );
  NAND2_X1 U14769 ( .A1(n12095), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11676) );
  XOR2_X1 U14770 ( .A(n19768), .B(n11696), .Z(n19765) );
  INV_X1 U14771 ( .A(n19765), .ZN(n14028) );
  AOI22_X1 U14772 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14773 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14774 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14775 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11682) );
  NAND4_X1 U14776 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11691) );
  AOI22_X1 U14777 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14778 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14779 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14780 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11686) );
  NAND4_X1 U14781 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11690) );
  OAI21_X1 U14782 ( .B1(n11691), .B2(n11690), .A(n11783), .ZN(n11694) );
  NAND2_X1 U14783 ( .A1(n12096), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11693) );
  NAND2_X1 U14784 ( .A1(n12095), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11692) );
  NAND3_X1 U14785 ( .A1(n11694), .A2(n11693), .A3(n11692), .ZN(n11695) );
  AOI21_X1 U14786 ( .B1(n14028), .B2(n12496), .A(n11695), .ZN(n13943) );
  XNOR2_X1 U14787 ( .A(n11712), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13978) );
  NAND2_X1 U14788 ( .A1(n13978), .A2(n12496), .ZN(n11711) );
  INV_X1 U14789 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13986) );
  INV_X1 U14790 ( .A(n12095), .ZN(n11823) );
  INV_X1 U14791 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14652) );
  OAI22_X1 U14792 ( .A1(n12090), .A2(n13986), .B1(n11823), .B2(n14652), .ZN(
        n11709) );
  AOI22_X1 U14793 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14794 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14795 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14796 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11697) );
  NAND4_X1 U14797 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11706) );
  AOI22_X1 U14798 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14799 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14800 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U14801 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11701) );
  NAND4_X1 U14802 ( .A1(n11704), .A2(n11703), .A3(n11702), .A4(n11701), .ZN(
        n11705) );
  NOR2_X1 U14803 ( .A1(n11706), .A2(n11705), .ZN(n11707) );
  NOR2_X1 U14804 ( .A1(n11752), .A2(n11707), .ZN(n11708) );
  NOR2_X1 U14805 ( .A1(n11709), .A2(n11708), .ZN(n11710) );
  NAND2_X1 U14806 ( .A1(n11711), .A2(n11710), .ZN(n13970) );
  INV_X1 U14807 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14068) );
  OAI21_X1 U14808 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11713), .A(
        n11740), .ZN(n15743) );
  AOI22_X1 U14809 ( .A1(n12496), .A2(n15743), .B1(n12095), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11714) );
  OAI21_X1 U14810 ( .B1(n12090), .B2(n14068), .A(n11714), .ZN(n14065) );
  AOI22_X1 U14811 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14812 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14813 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14814 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11715) );
  NAND4_X1 U14815 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(
        n11724) );
  AOI22_X1 U14816 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14817 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14818 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14819 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11719) );
  NAND4_X1 U14820 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11723) );
  NOR2_X1 U14821 ( .A1(n11724), .A2(n11723), .ZN(n11725) );
  NOR2_X1 U14822 ( .A1(n11752), .A2(n11725), .ZN(n14092) );
  XOR2_X1 U14823 ( .A(n14108), .B(n11757), .Z(n14644) );
  AOI22_X1 U14824 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14825 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U14826 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14827 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11726) );
  NAND4_X1 U14828 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11735) );
  AOI22_X1 U14829 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14830 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14831 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14832 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11730) );
  NAND4_X1 U14833 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11734) );
  NOR2_X1 U14834 ( .A1(n11735), .A2(n11734), .ZN(n11736) );
  OAI22_X1 U14835 ( .A1(n11752), .A2(n11736), .B1(n11823), .B2(n14108), .ZN(
        n11738) );
  INV_X1 U14836 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14135) );
  NOR2_X1 U14837 ( .A1(n12090), .A2(n14135), .ZN(n11737) );
  NOR2_X1 U14838 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  OAI21_X1 U14839 ( .B1(n14644), .B2(n12087), .A(n11739), .ZN(n14103) );
  XOR2_X1 U14840 ( .A(n15686), .B(n11740), .Z(n15730) );
  AOI22_X1 U14841 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11368), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14842 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11284), .B1(
        n11285), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14843 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14844 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11741) );
  NAND4_X1 U14845 ( .A1(n11744), .A2(n11743), .A3(n11742), .A4(n11741), .ZN(
        n11750) );
  AOI22_X1 U14846 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U14847 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11283), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U14848 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U14849 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11745) );
  NAND4_X1 U14850 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n11749) );
  NOR2_X1 U14851 ( .A1(n11750), .A2(n11749), .ZN(n11751) );
  OAI22_X1 U14852 ( .A1(n11752), .A2(n11751), .B1(n11823), .B2(n15686), .ZN(
        n11754) );
  INV_X1 U14853 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14101) );
  NOR2_X1 U14854 ( .A1(n12090), .A2(n14101), .ZN(n11753) );
  NOR2_X1 U14855 ( .A1(n11754), .A2(n11753), .ZN(n11755) );
  OAI21_X1 U14856 ( .B1(n15730), .B2(n12087), .A(n11755), .ZN(n14095) );
  XNOR2_X1 U14857 ( .A(n11774), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15672) );
  AOI22_X1 U14858 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U14859 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14860 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14861 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11758) );
  NAND4_X1 U14862 ( .A1(n11761), .A2(n11760), .A3(n11759), .A4(n11758), .ZN(
        n11767) );
  AOI22_X1 U14863 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U14864 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14865 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14866 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11762) );
  NAND4_X1 U14867 ( .A1(n11765), .A2(n11764), .A3(n11763), .A4(n11762), .ZN(
        n11766) );
  OAI21_X1 U14868 ( .B1(n11767), .B2(n11766), .A(n11783), .ZN(n11770) );
  NAND2_X1 U14869 ( .A1(n12096), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U14870 ( .A1(n12095), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11768) );
  NAND3_X1 U14871 ( .A1(n11770), .A2(n11769), .A3(n11768), .ZN(n11771) );
  AOI21_X1 U14872 ( .B1(n15672), .B2(n12496), .A(n11771), .ZN(n14073) );
  NAND2_X1 U14873 ( .A1(n11773), .A2(n11772), .ZN(n14070) );
  XOR2_X1 U14874 ( .A(n15664), .B(n11792), .Z(n15725) );
  INV_X1 U14875 ( .A(n15725), .ZN(n11790) );
  AOI22_X1 U14876 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14877 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11409), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14878 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14879 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11775) );
  NAND4_X1 U14880 ( .A1(n11778), .A2(n11777), .A3(n11776), .A4(n11775), .ZN(
        n11785) );
  AOI22_X1 U14881 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14882 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14883 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14884 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11779) );
  NAND4_X1 U14885 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11784) );
  OAI21_X1 U14886 ( .B1(n11785), .B2(n11784), .A(n11783), .ZN(n11788) );
  NAND2_X1 U14887 ( .A1(n12096), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11787) );
  NAND2_X1 U14888 ( .A1(n12095), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11786) );
  NAND3_X1 U14889 ( .A1(n11788), .A2(n11787), .A3(n11786), .ZN(n11789) );
  AOI21_X1 U14890 ( .B1(n11790), .B2(n12496), .A(n11789), .ZN(n14118) );
  INV_X1 U14891 ( .A(n14118), .ZN(n11791) );
  INV_X1 U14892 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14617) );
  XNOR2_X1 U14893 ( .A(n11811), .B(n14617), .ZN(n14619) );
  NAND2_X1 U14894 ( .A1(n14619), .A2(n12496), .ZN(n11810) );
  AOI22_X1 U14895 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14896 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U14897 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14898 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11793) );
  NAND4_X1 U14899 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11805) );
  AOI22_X1 U14900 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14901 ( .A1(n11275), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11332), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11801) );
  AOI21_X1 U14902 ( .B1(n12065), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n12496), .ZN(n11798) );
  NAND2_X1 U14903 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11797) );
  AND2_X1 U14904 ( .A1(n11798), .A2(n11797), .ZN(n11800) );
  AOI22_X1 U14905 ( .A1(n12073), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11799) );
  NAND4_X1 U14906 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11804) );
  INV_X1 U14907 ( .A(n14796), .ZN(n11803) );
  NAND2_X1 U14908 ( .A1(n12059), .A2(n12087), .ZN(n11899) );
  OAI21_X1 U14909 ( .B1(n11805), .B2(n11804), .A(n11899), .ZN(n11808) );
  NAND2_X1 U14910 ( .A1(n12096), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n11807) );
  NAND2_X1 U14911 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11806) );
  NAND3_X1 U14912 ( .A1(n11808), .A2(n11807), .A3(n11806), .ZN(n11809) );
  NAND2_X1 U14913 ( .A1(n11810), .A2(n11809), .ZN(n14149) );
  XOR2_X1 U14914 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11828), .Z(
        n15715) );
  AOI22_X1 U14915 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14916 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14917 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14918 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11812) );
  NAND4_X1 U14919 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11821) );
  AOI22_X1 U14920 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14921 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11332), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U14922 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U14923 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11816) );
  NAND4_X1 U14924 ( .A1(n11819), .A2(n11818), .A3(n11817), .A4(n11816), .ZN(
        n11820) );
  OR2_X1 U14925 ( .A1(n11821), .A2(n11820), .ZN(n11826) );
  INV_X1 U14926 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n11824) );
  INV_X1 U14927 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11822) );
  OAI22_X1 U14928 ( .A1(n12090), .A2(n11824), .B1(n11823), .B2(n11822), .ZN(
        n11825) );
  AOI21_X1 U14929 ( .B1(n12085), .B2(n11826), .A(n11825), .ZN(n11827) );
  OAI21_X1 U14930 ( .B1(n15715), .B2(n12087), .A(n11827), .ZN(n14461) );
  XNOR2_X1 U14931 ( .A(n11861), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15649) );
  AOI22_X1 U14932 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U14933 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11332), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11833) );
  NAND2_X1 U14934 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11830) );
  NAND2_X1 U14935 ( .A1(n12065), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11829) );
  AND3_X1 U14936 ( .A1(n11830), .A2(n12087), .A3(n11829), .ZN(n11832) );
  AOI22_X1 U14937 ( .A1(n12073), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11831) );
  NAND4_X1 U14938 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11840) );
  AOI22_X1 U14939 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11275), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14940 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14941 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14942 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11835) );
  NAND4_X1 U14943 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11839) );
  OR2_X1 U14944 ( .A1(n11840), .A2(n11839), .ZN(n11843) );
  INV_X1 U14945 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n11841) );
  OAI22_X1 U14946 ( .A1(n12090), .A2(n11841), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14601), .ZN(n11842) );
  AOI21_X1 U14947 ( .B1(n11899), .B2(n11843), .A(n11842), .ZN(n11844) );
  AOI21_X1 U14948 ( .B1(n15649), .B2(n12496), .A(n11844), .ZN(n14451) );
  NOR2_X2 U14949 ( .A1(n14448), .A2(n11845), .ZN(n14442) );
  AOI22_X1 U14950 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14951 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14952 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14953 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11846) );
  NAND4_X1 U14954 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n11855) );
  AOI22_X1 U14955 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14956 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14957 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U14958 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11850) );
  NAND4_X1 U14959 ( .A1(n11853), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n11854) );
  NOR2_X1 U14960 ( .A1(n11855), .A2(n11854), .ZN(n11860) );
  INV_X1 U14961 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U14962 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11856) );
  OAI211_X1 U14963 ( .C1(n12090), .C2(n11857), .A(n12087), .B(n11856), .ZN(
        n11858) );
  INV_X1 U14964 ( .A(n11858), .ZN(n11859) );
  OAI21_X1 U14965 ( .B1(n12059), .B2(n11860), .A(n11859), .ZN(n11864) );
  OAI21_X1 U14966 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11862), .A(
        n11904), .ZN(n15707) );
  OR2_X1 U14967 ( .A1(n15707), .A2(n12087), .ZN(n11863) );
  AOI22_X1 U14968 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14969 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14970 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14971 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11865) );
  NAND4_X1 U14972 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(
        n11874) );
  AOI22_X1 U14973 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14974 ( .A1(n11275), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14975 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14976 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11869) );
  NAND4_X1 U14977 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11873) );
  NOR2_X1 U14978 ( .A1(n11874), .A2(n11873), .ZN(n11879) );
  INV_X1 U14979 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n11876) );
  NAND2_X1 U14980 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11875) );
  OAI211_X1 U14981 ( .C1(n12090), .C2(n11876), .A(n12087), .B(n11875), .ZN(
        n11877) );
  INV_X1 U14982 ( .A(n11877), .ZN(n11878) );
  OAI21_X1 U14983 ( .B1(n12059), .B2(n11879), .A(n11878), .ZN(n11885) );
  INV_X1 U14984 ( .A(n11881), .ZN(n11882) );
  INV_X1 U14985 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14590) );
  NAND2_X1 U14986 ( .A1(n11882), .A2(n14590), .ZN(n11883) );
  AND2_X1 U14987 ( .A1(n11921), .A2(n11883), .ZN(n15611) );
  NAND2_X1 U14988 ( .A1(n15611), .A2(n12496), .ZN(n11884) );
  NAND2_X1 U14989 ( .A1(n11885), .A2(n11884), .ZN(n14435) );
  AOI22_X1 U14990 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12043), .B1(
        n11332), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14991 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11890) );
  NAND2_X1 U14992 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11887) );
  NAND2_X1 U14993 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11886) );
  AND3_X1 U14994 ( .A1(n11887), .A2(n11886), .A3(n12087), .ZN(n11889) );
  AOI22_X1 U14995 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11888) );
  NAND4_X1 U14996 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11897) );
  AOI22_X1 U14997 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14998 ( .A1(n11275), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14999 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U15000 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11892) );
  NAND4_X1 U15001 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11896) );
  OR2_X1 U15002 ( .A1(n11897), .A2(n11896), .ZN(n11898) );
  NAND2_X1 U15003 ( .A1(n11899), .A2(n11898), .ZN(n11903) );
  INV_X1 U15004 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n11900) );
  INV_X1 U15005 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15624) );
  OAI22_X1 U15006 ( .A1(n12090), .A2(n11900), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15624), .ZN(n11901) );
  INV_X1 U15007 ( .A(n11901), .ZN(n11902) );
  NAND2_X1 U15008 ( .A1(n11903), .A2(n11902), .ZN(n11906) );
  XNOR2_X1 U15009 ( .A(n11904), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15630) );
  NAND2_X1 U15010 ( .A1(n15630), .A2(n12496), .ZN(n11905) );
  NAND2_X1 U15011 ( .A1(n11906), .A2(n11905), .ZN(n14439) );
  AOI22_X1 U15012 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11275), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15013 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15014 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U15015 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U15016 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11917) );
  AOI22_X1 U15017 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15018 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15019 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U15020 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U15021 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  OAI21_X1 U15022 ( .B1(n11917), .B2(n11916), .A(n12085), .ZN(n11920) );
  INV_X1 U15023 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14578) );
  AOI21_X1 U15024 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14578), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11918) );
  AOI21_X1 U15025 ( .B1(n12096), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11918), .ZN(
        n11919) );
  XNOR2_X1 U15026 ( .A(n11921), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14580) );
  AOI22_X1 U15027 ( .A1(n11920), .A2(n11919), .B1(n12496), .B2(n14580), .ZN(
        n14400) );
  NAND2_X1 U15028 ( .A1(n11923), .A2(n14392), .ZN(n11924) );
  NAND2_X1 U15029 ( .A1(n11963), .A2(n11924), .ZN(n14574) );
  AOI22_X1 U15030 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15031 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U15032 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15033 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11925) );
  NAND4_X1 U15034 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(
        n11934) );
  AOI22_X1 U15035 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U15036 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U15037 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15038 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11929) );
  NAND4_X1 U15039 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n11933) );
  NOR2_X1 U15040 ( .A1(n11934), .A2(n11933), .ZN(n11960) );
  AOI22_X1 U15041 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15042 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15043 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U15044 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11935) );
  NAND4_X1 U15045 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11944) );
  AOI22_X1 U15046 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11942) );
  AOI22_X1 U15047 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15048 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15049 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11939) );
  NAND4_X1 U15050 ( .A1(n11942), .A2(n11941), .A3(n11940), .A4(n11939), .ZN(
        n11943) );
  NOR2_X1 U15051 ( .A1(n11944), .A2(n11943), .ZN(n11959) );
  XNOR2_X1 U15052 ( .A(n11960), .B(n11959), .ZN(n11947) );
  OAI21_X1 U15053 ( .B1(n20641), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n20640), .ZN(n11946) );
  NAND2_X1 U15054 ( .A1(n12096), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n11945) );
  OAI211_X1 U15055 ( .C1(n12059), .C2(n11947), .A(n11946), .B(n11945), .ZN(
        n11948) );
  OAI21_X1 U15056 ( .B1(n12087), .B2(n14574), .A(n11948), .ZN(n14390) );
  AOI22_X1 U15057 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U15058 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U15059 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15060 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11949) );
  NAND4_X1 U15061 ( .A1(n11952), .A2(n11951), .A3(n11950), .A4(n11949), .ZN(
        n11958) );
  AOI22_X1 U15062 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U15063 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15064 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15065 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11953) );
  NAND4_X1 U15066 ( .A1(n11956), .A2(n11955), .A3(n11954), .A4(n11953), .ZN(
        n11957) );
  OR2_X1 U15067 ( .A1(n11958), .A2(n11957), .ZN(n11979) );
  NOR2_X1 U15068 ( .A1(n11960), .A2(n11959), .ZN(n11980) );
  XOR2_X1 U15069 ( .A(n11979), .B(n11980), .Z(n11961) );
  NAND2_X1 U15070 ( .A1(n11961), .A2(n12085), .ZN(n11965) );
  INV_X1 U15071 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14565) );
  NOR2_X1 U15072 ( .A1(n14565), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11962) );
  AOI211_X1 U15073 ( .C1(n12096), .C2(P1_EAX_REG_24__SCAN_IN), .A(n12496), .B(
        n11962), .ZN(n11964) );
  XOR2_X1 U15074 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n11966), .Z(
        n14569) );
  AOI22_X1 U15075 ( .A1(n11965), .A2(n11964), .B1(n12496), .B2(n14569), .ZN(
        n14378) );
  NAND2_X1 U15076 ( .A1(n14376), .A2(n14378), .ZN(n14360) );
  INV_X1 U15077 ( .A(n11967), .ZN(n11968) );
  INV_X1 U15078 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14366) );
  OAI21_X1 U15079 ( .B1(n11968), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n12000), .ZN(n14557) );
  AOI22_X1 U15080 ( .A1(n11332), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15081 ( .A1(n11368), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15082 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U15083 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U15084 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11978) );
  AOI22_X1 U15085 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15086 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11284), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15087 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15088 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11973) );
  NAND4_X1 U15089 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11977) );
  NOR2_X1 U15090 ( .A1(n11978), .A2(n11977), .ZN(n11997) );
  NAND2_X1 U15091 ( .A1(n11980), .A2(n11979), .ZN(n11996) );
  XNOR2_X1 U15092 ( .A(n11997), .B(n11996), .ZN(n11983) );
  AOI21_X1 U15093 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20640), .A(
        n12496), .ZN(n11982) );
  NAND2_X1 U15094 ( .A1(n12096), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n11981) );
  OAI211_X1 U15095 ( .C1(n11983), .C2(n12059), .A(n11982), .B(n11981), .ZN(
        n11984) );
  OAI21_X1 U15096 ( .B1(n12087), .B2(n14557), .A(n11984), .ZN(n14361) );
  NOR2_X2 U15097 ( .A1(n14360), .A2(n14361), .ZN(n14348) );
  AOI22_X1 U15098 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15099 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15100 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15101 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11985) );
  NAND4_X1 U15102 ( .A1(n11988), .A2(n11987), .A3(n11986), .A4(n11985), .ZN(
        n11995) );
  AOI22_X1 U15103 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15104 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15105 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15106 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11990) );
  NAND4_X1 U15107 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11994) );
  NOR2_X1 U15108 ( .A1(n11997), .A2(n11996), .ZN(n12017) );
  XOR2_X1 U15109 ( .A(n12016), .B(n12017), .Z(n11998) );
  NAND2_X1 U15110 ( .A1(n11998), .A2(n12085), .ZN(n12002) );
  INV_X1 U15111 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14545) );
  NOR2_X1 U15112 ( .A1(n14545), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11999) );
  AOI211_X1 U15113 ( .C1(n12096), .C2(P1_EAX_REG_26__SCAN_IN), .A(n12496), .B(
        n11999), .ZN(n12001) );
  XOR2_X1 U15114 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(n12003), .Z(
        n14549) );
  AOI22_X1 U15115 ( .A1(n12002), .A2(n12001), .B1(n12496), .B2(n14549), .ZN(
        n14350) );
  NAND2_X1 U15116 ( .A1(n14348), .A2(n14350), .ZN(n14335) );
  INV_X1 U15117 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14341) );
  NAND2_X1 U15118 ( .A1(n12004), .A2(n14341), .ZN(n12005) );
  NAND2_X1 U15119 ( .A1(n12039), .A2(n12005), .ZN(n14538) );
  AOI22_X1 U15120 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11369), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U15121 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15122 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U15123 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12006) );
  NAND4_X1 U15124 ( .A1(n12009), .A2(n12008), .A3(n12007), .A4(n12006), .ZN(
        n12015) );
  AOI22_X1 U15125 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12043), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15126 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11284), .B1(
        n11299), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15127 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15128 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12010) );
  NAND4_X1 U15129 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12010), .ZN(
        n12014) );
  NOR2_X1 U15130 ( .A1(n12015), .A2(n12014), .ZN(n12033) );
  NAND2_X1 U15131 ( .A1(n12017), .A2(n12016), .ZN(n12032) );
  XNOR2_X1 U15132 ( .A(n12033), .B(n12032), .ZN(n12020) );
  AOI21_X1 U15133 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20640), .A(
        n12496), .ZN(n12019) );
  NAND2_X1 U15134 ( .A1(n12096), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12018) );
  OAI211_X1 U15135 ( .C1(n12020), .C2(n12059), .A(n12019), .B(n12018), .ZN(
        n12021) );
  OAI21_X1 U15136 ( .B1(n12087), .B2(n14538), .A(n12021), .ZN(n14337) );
  AOI22_X1 U15137 ( .A1(n12043), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15138 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11332), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15139 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15140 ( .A1(n11369), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12022) );
  NAND4_X1 U15141 ( .A1(n12025), .A2(n12024), .A3(n12023), .A4(n12022), .ZN(
        n12031) );
  AOI22_X1 U15142 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11275), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15143 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15144 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15145 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U15146 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12030) );
  OR2_X1 U15147 ( .A1(n12031), .A2(n12030), .ZN(n12055) );
  NOR2_X1 U15148 ( .A1(n12033), .A2(n12032), .ZN(n12056) );
  XOR2_X1 U15149 ( .A(n12055), .B(n12056), .Z(n12034) );
  NAND2_X1 U15150 ( .A1(n12034), .A2(n12085), .ZN(n12038) );
  INV_X1 U15151 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14260) );
  NOR2_X1 U15152 ( .A1(n14260), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12035) );
  AOI211_X1 U15153 ( .C1(n12096), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12496), .B(
        n12035), .ZN(n12037) );
  INV_X1 U15154 ( .A(n12039), .ZN(n12036) );
  XOR2_X1 U15155 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n12036), .Z(
        n14326) );
  AOI22_X1 U15156 ( .A1(n12038), .A2(n12037), .B1(n12496), .B2(n14326), .ZN(
        n14261) );
  NAND2_X1 U15157 ( .A1(n12040), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12102) );
  INV_X1 U15158 ( .A(n12040), .ZN(n12041) );
  INV_X1 U15159 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U15160 ( .A1(n12041), .A2(n14312), .ZN(n12042) );
  NAND2_X1 U15161 ( .A1(n12102), .A2(n12042), .ZN(n14528) );
  AOI22_X1 U15162 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12043), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15163 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15164 ( .A1(n11284), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15165 ( .A1(n12075), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12045) );
  NAND4_X1 U15166 ( .A1(n12048), .A2(n12047), .A3(n12046), .A4(n12045), .ZN(
        n12054) );
  AOI22_X1 U15167 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15168 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15169 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15170 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11363), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12049) );
  NAND4_X1 U15171 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(
        n12053) );
  NOR2_X1 U15172 ( .A1(n12054), .A2(n12053), .ZN(n12063) );
  NAND2_X1 U15173 ( .A1(n12056), .A2(n12055), .ZN(n12062) );
  XNOR2_X1 U15174 ( .A(n12063), .B(n12062), .ZN(n12060) );
  AOI21_X1 U15175 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20640), .A(
        n12496), .ZN(n12058) );
  NAND2_X1 U15176 ( .A1(n12096), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12057) );
  OAI211_X1 U15177 ( .C1(n12060), .C2(n12059), .A(n12058), .B(n12057), .ZN(
        n12061) );
  OAI21_X1 U15178 ( .B1(n12087), .B2(n14528), .A(n12061), .ZN(n14310) );
  NOR2_X1 U15179 ( .A1(n12063), .A2(n12062), .ZN(n12084) );
  AOI22_X1 U15180 ( .A1(n11285), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12064), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15181 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11369), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15182 ( .A1(n11409), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12065), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15183 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12044), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15184 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12082) );
  AOI22_X1 U15185 ( .A1(n11275), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11368), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15186 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12071), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15187 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15188 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12075), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U15189 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12081) );
  NOR2_X1 U15190 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  XNOR2_X1 U15191 ( .A(n12084), .B(n12083), .ZN(n12086) );
  NAND2_X1 U15192 ( .A1(n12086), .A2(n12085), .ZN(n12094) );
  INV_X1 U15193 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12089) );
  NAND2_X1 U15194 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12088) );
  OAI211_X1 U15195 ( .C1(n12090), .C2(n12089), .A(n12088), .B(n12087), .ZN(
        n12091) );
  INV_X1 U15196 ( .A(n12091), .ZN(n12093) );
  XNOR2_X1 U15197 ( .A(n12102), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14517) );
  AND2_X1 U15198 ( .A1(n14517), .A2(n12496), .ZN(n12092) );
  AOI21_X1 U15199 ( .B1(n12094), .B2(n12093), .A(n12092), .ZN(n13086) );
  AOI22_X1 U15200 ( .A1(n12096), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12095), .ZN(n12097) );
  NAND3_X1 U15201 ( .A1(n20790), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15883) );
  INV_X1 U15202 ( .A(n15883), .ZN(n12099) );
  NAND2_X1 U15203 ( .A1(n12500), .A2(n19911), .ZN(n12109) );
  NAND2_X1 U15204 ( .A1(n20493), .A2(n12104), .ZN(n20646) );
  NAND2_X1 U15205 ( .A1(n20646), .A2(n20790), .ZN(n12100) );
  NAND2_X1 U15206 ( .A1(n20790), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15577) );
  NAND2_X1 U15207 ( .A1(n20641), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12101) );
  INV_X1 U15208 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14519) );
  INV_X1 U15209 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12607) );
  NAND2_X1 U15210 ( .A1(n12105), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n13057) );
  NAND2_X1 U15211 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12106) );
  OAI211_X1 U15212 ( .C1(n19916), .C2(n13866), .A(n13057), .B(n12106), .ZN(
        n12107) );
  OAI211_X1 U15213 ( .C1(n13018), .C2(n19746), .A(n12109), .B(n12108), .ZN(
        P1_U2968) );
  NOR2_X2 U15214 ( .A1(n12118), .A2(n16651), .ZN(n16872) );
  AOI22_X1 U15215 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15216 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9586), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12113) );
  NOR2_X1 U15217 ( .A1(n16651), .A2(n12120), .ZN(n12162) );
  AOI22_X1 U15218 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12112) );
  NOR2_X2 U15219 ( .A1(n12118), .A2(n12115), .ZN(n12172) );
  AOI22_X1 U15220 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12111) );
  NAND4_X1 U15221 ( .A1(n12114), .A2(n12113), .A3(n12112), .A4(n12111), .ZN(
        n12126) );
  NOR2_X2 U15222 ( .A1(n12116), .A2(n12119), .ZN(n12206) );
  CLKBUF_X3 U15223 ( .A(n12206), .Z(n16941) );
  AOI22_X1 U15224 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15225 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15226 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15227 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12121) );
  NAND4_X1 U15228 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  AOI22_X1 U15229 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15230 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15231 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15232 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U15233 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12137) );
  AOI22_X1 U15234 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15235 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15236 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15237 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U15238 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12136) );
  AOI22_X1 U15239 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15240 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15241 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15242 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12138) );
  NAND4_X1 U15243 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12148) );
  AOI22_X1 U15244 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15245 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12163), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15246 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15247 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12143) );
  NAND4_X1 U15248 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12147) );
  AOI22_X1 U15249 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16942), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15250 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n16916), .ZN(n12152) );
  AOI22_X1 U15251 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12110), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15252 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12245), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12177), .ZN(n12150) );
  NAND4_X1 U15253 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12161) );
  AOI22_X1 U15254 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n12163), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n15473), .ZN(n12159) );
  AOI22_X1 U15255 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9594), .B1(
        n16683), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15256 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9585), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n12206), .ZN(n12157) );
  AOI22_X1 U15257 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n9601), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n16922), .ZN(n12156) );
  NAND4_X1 U15258 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12160) );
  OR2_X2 U15259 ( .A1(n12161), .A2(n12160), .ZN(n12394) );
  AOI22_X1 U15260 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15261 ( .A1(n12162), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12207), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15262 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12163), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15263 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12245), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12164) );
  INV_X1 U15264 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U15265 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12168) );
  OAI21_X1 U15266 ( .B1(n12258), .B2(n16982), .A(n12168), .ZN(n12171) );
  AOI22_X1 U15267 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15268 ( .A1(n12206), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12174) );
  NAND4_X1 U15269 ( .A1(n9997), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n17129) );
  NAND2_X1 U15270 ( .A1(n12394), .A2(n17129), .ZN(n12201) );
  NOR2_X1 U15271 ( .A1(n17123), .A2(n12201), .ZN(n12199) );
  AOI22_X1 U15272 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15273 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12185) );
  INV_X1 U15274 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20786) );
  INV_X2 U15275 ( .A(n16840), .ZN(n16933) );
  AOI22_X1 U15276 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12176) );
  OAI21_X1 U15277 ( .B1(n15453), .B2(n20786), .A(n12176), .ZN(n12183) );
  AOI22_X1 U15278 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15279 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15280 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15281 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12178) );
  NAND4_X1 U15282 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12182) );
  AOI211_X1 U15283 ( .C1(n16877), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n12183), .B(n12182), .ZN(n12184) );
  NAND3_X1 U15284 ( .A1(n12186), .A2(n12185), .A3(n12184), .ZN(n17119) );
  NAND2_X1 U15285 ( .A1(n12199), .A2(n17119), .ZN(n12198) );
  AOI22_X1 U15286 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9585), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15287 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15288 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12187) );
  OAI21_X1 U15289 ( .B1(n15453), .B2(n20774), .A(n12187), .ZN(n12193) );
  AOI22_X1 U15290 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15291 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15292 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15293 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12188) );
  NAND4_X1 U15294 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12192) );
  AOI211_X1 U15295 ( .C1(n16945), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n12193), .B(n12192), .ZN(n12194) );
  NAND3_X1 U15296 ( .A1(n12196), .A2(n12195), .A3(n12194), .ZN(n17111) );
  INV_X1 U15297 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17654) );
  INV_X1 U15298 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17747) );
  INV_X1 U15299 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17836) );
  NOR2_X1 U15300 ( .A1(n17836), .A2(n17822), .ZN(n17814) );
  NAND2_X1 U15301 ( .A1(n17814), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17783) );
  NOR2_X1 U15302 ( .A1(n17783), .A2(n17794), .ZN(n17442) );
  NAND2_X1 U15303 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17442), .ZN(
        n17754) );
  NOR2_X1 U15304 ( .A1(n17771), .A2(n17754), .ZN(n17435) );
  NAND2_X1 U15305 ( .A1(n17435), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17733) );
  XOR2_X1 U15306 ( .A(n17111), .B(n12197), .Z(n12224) );
  XOR2_X1 U15307 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12224), .Z(
        n17541) );
  XOR2_X1 U15308 ( .A(n17115), .B(n12198), .Z(n12222) );
  XOR2_X1 U15309 ( .A(n17119), .B(n12199), .Z(n12200) );
  NAND2_X1 U15310 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12200), .ZN(
        n12221) );
  XOR2_X1 U15311 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12200), .Z(
        n17570) );
  XOR2_X1 U15312 ( .A(n17123), .B(n12201), .Z(n12217) );
  INV_X1 U15313 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17914) );
  XNOR2_X1 U15314 ( .A(n12215), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17591) );
  NAND2_X1 U15315 ( .A1(n17141), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12214) );
  AOI22_X1 U15316 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12110), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15317 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15318 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12163), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15319 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12202) );
  NAND4_X1 U15320 ( .A1(n12205), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        n12213) );
  AOI22_X1 U15321 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15322 ( .A1(n12206), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15323 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15324 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12208) );
  NAND4_X1 U15325 ( .A1(n12211), .A2(n12210), .A3(n12209), .A4(n12208), .ZN(
        n12212) );
  NOR2_X1 U15326 ( .A1(n12213), .A2(n12212), .ZN(n17608) );
  NOR2_X1 U15327 ( .A1(n17608), .A2(n18583), .ZN(n17607) );
  NAND2_X1 U15328 ( .A1(n17599), .A2(n17607), .ZN(n17598) );
  NAND2_X1 U15329 ( .A1(n12214), .A2(n17598), .ZN(n17590) );
  NAND2_X1 U15330 ( .A1(n17591), .A2(n17590), .ZN(n17589) );
  OR2_X1 U15331 ( .A1(n17914), .A2(n12215), .ZN(n12216) );
  NAND2_X1 U15332 ( .A1(n17589), .A2(n12216), .ZN(n12219) );
  NAND2_X1 U15333 ( .A1(n12217), .A2(n12219), .ZN(n12220) );
  XNOR2_X1 U15334 ( .A(n12219), .B(n12218), .ZN(n17580) );
  NAND2_X1 U15335 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17580), .ZN(
        n17579) );
  NAND2_X1 U15336 ( .A1(n12222), .A2(n12223), .ZN(n17557) );
  NAND2_X1 U15337 ( .A1(n17558), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17555) );
  NAND2_X1 U15338 ( .A1(n17557), .A2(n17555), .ZN(n17540) );
  NAND2_X1 U15339 ( .A1(n17541), .A2(n17540), .ZN(n17539) );
  NAND2_X1 U15340 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12224), .ZN(
        n12225) );
  NAND2_X1 U15341 ( .A1(n17539), .A2(n12225), .ZN(n12227) );
  AOI21_X1 U15342 ( .B1(n17108), .B2(n16158), .A(n17518), .ZN(n12228) );
  XNOR2_X1 U15343 ( .A(n12227), .B(n12226), .ZN(n17529) );
  NAND2_X1 U15344 ( .A1(n12228), .A2(n12227), .ZN(n12229) );
  NOR2_X2 U15345 ( .A1(n12382), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12230) );
  INV_X1 U15346 ( .A(n12230), .ZN(n12231) );
  AND2_X1 U15347 ( .A1(n12382), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17400) );
  NAND2_X1 U15348 ( .A1(n17771), .A2(n17794), .ZN(n17422) );
  NOR4_X1 U15349 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n17422), .ZN(n12232) );
  AOI21_X1 U15350 ( .B1(n17419), .B2(n12232), .A(n17518), .ZN(n12235) );
  INV_X1 U15351 ( .A(n12235), .ZN(n12233) );
  OAI221_X1 U15352 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n9847), .C1(
        n17747), .C2(n12234), .A(n12233), .ZN(n17388) );
  NOR2_X1 U15353 ( .A1(n12235), .A2(n12234), .ZN(n17402) );
  NAND2_X1 U15354 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17384) );
  INV_X1 U15355 ( .A(n17384), .ZN(n17729) );
  INV_X1 U15356 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17694) );
  NAND2_X1 U15357 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17695) );
  NOR3_X1 U15358 ( .A1(n17693), .A2(n17694), .A3(n17695), .ZN(n17331) );
  NAND2_X1 U15359 ( .A1(n17331), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17640) );
  NOR2_X1 U15360 ( .A1(n17668), .A2(n17640), .ZN(n17639) );
  NAND2_X1 U15361 ( .A1(n17729), .A2(n17639), .ZN(n17294) );
  NAND2_X1 U15362 ( .A1(n17693), .A2(n9847), .ZN(n17381) );
  NOR2_X1 U15363 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17381), .ZN(
        n12236) );
  INV_X1 U15364 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n20755) );
  NAND2_X1 U15365 ( .A1(n12236), .A2(n20755), .ZN(n17338) );
  INV_X1 U15366 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17691) );
  NAND3_X1 U15367 ( .A1(n17332), .A2(n17691), .A3(n17668), .ZN(n12237) );
  INV_X1 U15368 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17663) );
  NAND2_X1 U15369 ( .A1(n17300), .A2(n17663), .ZN(n17299) );
  NOR2_X1 U15370 ( .A1(n17384), .A2(n17402), .ZN(n17337) );
  NAND3_X1 U15371 ( .A1(n17299), .A2(n17639), .A3(n17383), .ZN(n12241) );
  NAND2_X1 U15372 ( .A1(n9847), .A2(n17299), .ZN(n17284) );
  NAND2_X1 U15373 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17614) );
  OR2_X1 U15374 ( .A1(n12241), .A2(n17614), .ZN(n12242) );
  NOR2_X2 U15375 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n12244), .ZN(
        n16166) );
  INV_X1 U15376 ( .A(n16166), .ZN(n12418) );
  NAND2_X1 U15377 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n12244), .ZN(
        n16157) );
  NAND2_X1 U15378 ( .A1(n12418), .A2(n16157), .ZN(n17258) );
  NAND2_X1 U15379 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17518), .ZN(
        n15529) );
  OAI21_X1 U15380 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17518), .A(
        n15529), .ZN(n16165) );
  AOI22_X1 U15381 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15382 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15383 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12207), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12247) );
  CLKBUF_X3 U15384 ( .A(n12245), .Z(n16936) );
  AOI22_X1 U15385 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12246) );
  NAND4_X1 U15386 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12257) );
  AOI22_X1 U15387 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n9594), .ZN(n12255) );
  AOI22_X1 U15388 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16917), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15389 ( .A1(n16877), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15390 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12252) );
  NAND4_X1 U15391 ( .A1(n12255), .A2(n12254), .A3(n12253), .A4(n12252), .ZN(
        n12256) );
  AOI22_X1 U15392 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15393 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15394 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12259) );
  OAI21_X1 U15395 ( .B1(n12280), .B2(n16813), .A(n12259), .ZN(n12265) );
  AOI22_X1 U15396 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15397 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15398 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15399 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12260) );
  NAND4_X1 U15400 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12264) );
  NAND2_X1 U15401 ( .A1(n16612), .A2(n18605), .ZN(n12342) );
  NAND2_X1 U15402 ( .A1(n17960), .A2(n17955), .ZN(n12336) );
  NAND2_X1 U15403 ( .A1(n12342), .A2(n12336), .ZN(n18619) );
  AOI22_X1 U15404 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15405 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15406 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12269) );
  OAI21_X1 U15407 ( .B1(n12280), .B2(n20785), .A(n12269), .ZN(n12275) );
  AOI22_X1 U15408 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15409 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9585), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15410 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15411 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12270) );
  NAND4_X1 U15412 ( .A1(n12273), .A2(n12272), .A3(n12271), .A4(n12270), .ZN(
        n12274) );
  AOI22_X1 U15413 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15414 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12288) );
  INV_X1 U15415 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U15416 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12279) );
  OAI21_X1 U15417 ( .B1(n12280), .B2(n16971), .A(n12279), .ZN(n12286) );
  AOI22_X1 U15418 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15419 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15420 ( .A1(n16877), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15421 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12163), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12281) );
  NAND4_X1 U15422 ( .A1(n12284), .A2(n12283), .A3(n12282), .A4(n12281), .ZN(
        n12285) );
  AOI211_X1 U15423 ( .C1(n16944), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n12286), .B(n12285), .ZN(n12287) );
  NAND3_X1 U15424 ( .A1(n12289), .A2(n12288), .A3(n12287), .ZN(n15510) );
  AOI22_X1 U15425 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15426 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15427 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15428 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12290) );
  NAND4_X1 U15429 ( .A1(n12293), .A2(n12292), .A3(n12291), .A4(n12290), .ZN(
        n12299) );
  AOI22_X1 U15430 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15431 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16922), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15432 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15433 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9586), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12294) );
  NAND4_X1 U15434 ( .A1(n12297), .A2(n12296), .A3(n12295), .A4(n12294), .ZN(
        n12298) );
  AOI22_X1 U15435 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15436 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15437 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15438 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12300) );
  NAND4_X1 U15439 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12309) );
  AOI22_X1 U15440 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15441 ( .A1(n16877), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15442 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15443 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12304) );
  NAND4_X1 U15444 ( .A1(n12307), .A2(n12306), .A3(n12305), .A4(n12304), .ZN(
        n12308) );
  AOI22_X1 U15445 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15446 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15447 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12163), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15448 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12310) );
  NAND4_X1 U15449 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12319) );
  AOI22_X1 U15450 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15451 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16922), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15452 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15453 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12314) );
  NAND4_X1 U15454 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n12318) );
  AOI22_X1 U15455 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15456 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15457 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15458 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12320) );
  NAND4_X1 U15459 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12320), .ZN(
        n12329) );
  AOI22_X1 U15460 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15461 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15462 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15463 ( .A1(n12110), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12324) );
  NAND4_X1 U15464 ( .A1(n12327), .A2(n12326), .A3(n12325), .A4(n12324), .ZN(
        n12328) );
  NOR2_X1 U15465 ( .A1(n17989), .A2(n17969), .ZN(n12334) );
  NAND2_X1 U15466 ( .A1(n15510), .A2(n17983), .ZN(n18400) );
  NAND2_X1 U15467 ( .A1(n17965), .A2(n17969), .ZN(n18399) );
  AND2_X1 U15468 ( .A1(n17960), .A2(n14173), .ZN(n12332) );
  NAND2_X1 U15469 ( .A1(n17969), .A2(n12340), .ZN(n12330) );
  INV_X1 U15470 ( .A(n17983), .ZN(n15513) );
  NAND2_X1 U15471 ( .A1(n15509), .A2(n15513), .ZN(n12341) );
  INV_X1 U15472 ( .A(n12341), .ZN(n15511) );
  NAND2_X1 U15473 ( .A1(n17973), .A2(n15511), .ZN(n12343) );
  INV_X1 U15474 ( .A(n15491), .ZN(n12331) );
  NOR3_X1 U15475 ( .A1(n17960), .A2(n12334), .A3(n12333), .ZN(n12350) );
  INV_X1 U15476 ( .A(n17969), .ZN(n12339) );
  INV_X1 U15477 ( .A(n12335), .ZN(n12337) );
  NAND2_X1 U15478 ( .A1(n17983), .A2(n15509), .ZN(n18423) );
  AOI21_X1 U15479 ( .B1(n17077), .B2(n18423), .A(n12336), .ZN(n15490) );
  OAI21_X1 U15480 ( .B1(n12337), .B2(n15490), .A(n12339), .ZN(n12338) );
  OAI21_X1 U15481 ( .B1(n12340), .B2(n12339), .A(n12338), .ZN(n12349) );
  NAND3_X1 U15482 ( .A1(n17965), .A2(n12342), .A3(n12341), .ZN(n12345) );
  OAI22_X1 U15483 ( .A1(n17989), .A2(n12345), .B1(n12344), .B2(n12343), .ZN(
        n12346) );
  OAI22_X1 U15484 ( .A1(n18573), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18433), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12359) );
  OAI22_X1 U15485 ( .A1(n18580), .A2(n18428), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12365) );
  OAI21_X1 U15486 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18573), .A(
        n12352), .ZN(n12353) );
  NAND2_X1 U15487 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12353), .ZN(
        n12355) );
  OAI22_X1 U15488 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18437), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12353), .ZN(n12357) );
  AOI21_X1 U15489 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12355), .A(
        n12357), .ZN(n12354) );
  NOR2_X1 U15490 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18437), .ZN(
        n12356) );
  AOI22_X1 U15491 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12357), .B1(
        n12356), .B2(n12355), .ZN(n12361) );
  NAND2_X1 U15492 ( .A1(n12360), .A2(n12359), .ZN(n12358) );
  AOI21_X1 U15493 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18586), .A(
        n12364), .ZN(n12369) );
  NAND3_X1 U15494 ( .A1(n12365), .A2(n12361), .A3(n12369), .ZN(n12362) );
  NAND3_X1 U15495 ( .A1(n12366), .A2(n12367), .A3(n12362), .ZN(n15517) );
  INV_X1 U15496 ( .A(n15517), .ZN(n18386) );
  XNOR2_X1 U15497 ( .A(n18605), .B(n17965), .ZN(n15507) );
  INV_X1 U15498 ( .A(n12367), .ZN(n12370) );
  XNOR2_X1 U15499 ( .A(n12365), .B(n12364), .ZN(n12368) );
  AOI21_X1 U15500 ( .B1(n12370), .B2(n12369), .A(n15508), .ZN(n18390) );
  AOI211_X1 U15501 ( .C1(n12371), .C2(n16165), .A(n16154), .B(n17498), .ZN(
        n12372) );
  INV_X1 U15502 ( .A(n12372), .ZN(n12416) );
  OAI21_X1 U15503 ( .B1(n18617), .B2(n18566), .A(n18555), .ZN(n18602) );
  INV_X1 U15504 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16275) );
  NOR2_X1 U15505 ( .A1(n18566), .A2(n16275), .ZN(n17512) );
  INV_X1 U15506 ( .A(n17512), .ZN(n17566) );
  INV_X1 U15507 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12375) );
  NAND2_X1 U15508 ( .A1(n16598), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17476) );
  NAND4_X1 U15509 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16527) );
  AND2_X2 U15510 ( .A1(n16526), .A2(n12374), .ZN(n17479) );
  NAND2_X1 U15511 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U15512 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17290) );
  INV_X1 U15513 ( .A(n16298), .ZN(n16308) );
  INV_X1 U15514 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16309) );
  NAND2_X1 U15515 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16307), .ZN(
        n16297) );
  NOR2_X2 U15516 ( .A1(n16297), .A2(n12375), .ZN(n12427) );
  AOI21_X1 U15517 ( .B1(n12375), .B2(n16297), .A(n12427), .ZN(n16349) );
  INV_X1 U15518 ( .A(n16349), .ZN(n12380) );
  NOR2_X1 U15519 ( .A1(n17288), .A2(n17290), .ZN(n17271) );
  NAND2_X1 U15520 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17271), .ZN(
        n12377) );
  INV_X1 U15521 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16360) );
  NOR2_X1 U15522 ( .A1(n12377), .A2(n16360), .ZN(n12425) );
  INV_X1 U15523 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18608) );
  NAND2_X1 U15524 ( .A1(n18608), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18464) );
  NAND2_X1 U15525 ( .A1(n18617), .A2(n18555), .ZN(n16272) );
  INV_X1 U15526 ( .A(n18191), .ZN(n18287) );
  AOI22_X1 U15527 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .B1(n18566), .B2(n18617), .ZN(n18461) );
  AOI21_X1 U15528 ( .B1(n17353), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18329), .ZN(n17289) );
  NAND3_X1 U15529 ( .A1(n12425), .A2(n12375), .A3(n17446), .ZN(n12379) );
  NOR3_X1 U15530 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17289), .A3(
        n12377), .ZN(n17261) );
  OAI21_X1 U15531 ( .B1(n16298), .B2(n18464), .A(n17609), .ZN(n12376) );
  AOI21_X1 U15532 ( .B1(n17512), .B2(n12377), .A(n12376), .ZN(n17275) );
  OAI21_X1 U15533 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17354), .A(
        n17275), .ZN(n17262) );
  OAI21_X1 U15534 ( .B1(n17261), .B2(n17262), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12378) );
  OAI211_X1 U15535 ( .C1(n17450), .C2(n12380), .A(n12379), .B(n12378), .ZN(
        n12413) );
  INV_X1 U15536 ( .A(n17108), .ZN(n12381) );
  NOR2_X2 U15537 ( .A1(n12381), .A2(n17612), .ZN(n17520) );
  INV_X1 U15538 ( .A(n17331), .ZN(n17675) );
  NOR2_X1 U15539 ( .A1(n17384), .A2(n17675), .ZN(n17679) );
  AND2_X1 U15540 ( .A1(n17679), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17618) );
  NOR2_X1 U15541 ( .A1(n17668), .A2(n17663), .ZN(n17642) );
  INV_X1 U15542 ( .A(n17642), .ZN(n17619) );
  NOR2_X1 U15543 ( .A1(n17619), .A2(n17614), .ZN(n15524) );
  INV_X1 U15544 ( .A(n17733), .ZN(n17401) );
  NOR2_X1 U15545 ( .A1(n17518), .A2(n12382), .ZN(n17487) );
  INV_X1 U15546 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17846) );
  NAND2_X1 U15547 ( .A1(n17401), .A2(n17808), .ZN(n17681) );
  NAND2_X1 U15548 ( .A1(n15506), .A2(n17752), .ZN(n17615) );
  NOR2_X1 U15549 ( .A1(n17608), .A2(n17141), .ZN(n12390) );
  NOR2_X1 U15550 ( .A1(n12390), .A2(n17129), .ZN(n12388) );
  NOR2_X1 U15551 ( .A1(n12388), .A2(n17123), .ZN(n12387) );
  NAND2_X1 U15552 ( .A1(n12387), .A2(n17119), .ZN(n12385) );
  NOR2_X1 U15553 ( .A1(n17115), .A2(n12385), .ZN(n12384) );
  NAND2_X1 U15554 ( .A1(n12384), .A2(n17111), .ZN(n12383) );
  NOR2_X1 U15555 ( .A1(n17108), .A2(n12383), .ZN(n12408) );
  XOR2_X1 U15556 ( .A(n12383), .B(n17108), .Z(n17531) );
  XOR2_X1 U15557 ( .A(n12384), .B(n17111), .Z(n12401) );
  XOR2_X1 U15558 ( .A(n12385), .B(n17115), .Z(n12386) );
  NAND2_X1 U15559 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12386), .ZN(
        n12400) );
  XOR2_X1 U15560 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12386), .Z(
        n17551) );
  XOR2_X1 U15561 ( .A(n12387), .B(n17119), .Z(n12398) );
  XOR2_X1 U15562 ( .A(n17123), .B(n12388), .Z(n12389) );
  NAND2_X1 U15563 ( .A1(n12389), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12396) );
  XOR2_X1 U15564 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12389), .Z(
        n17577) );
  XOR2_X1 U15565 ( .A(n17129), .B(n12390), .Z(n12391) );
  OR2_X1 U15566 ( .A1(n17914), .A2(n12391), .ZN(n12395) );
  XOR2_X1 U15567 ( .A(n17914), .B(n12391), .Z(n17588) );
  INV_X1 U15568 ( .A(n17608), .ZN(n15607) );
  AOI21_X1 U15569 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12394), .A(
        n15607), .ZN(n12393) );
  NOR2_X1 U15570 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12394), .ZN(
        n12392) );
  AOI221_X1 U15571 ( .B1(n15607), .B2(n12394), .C1(n12393), .C2(n18583), .A(
        n12392), .ZN(n17587) );
  NAND2_X1 U15572 ( .A1(n17588), .A2(n17587), .ZN(n17586) );
  NAND2_X1 U15573 ( .A1(n12395), .A2(n17586), .ZN(n17576) );
  NAND2_X1 U15574 ( .A1(n17577), .A2(n17576), .ZN(n17575) );
  NAND2_X1 U15575 ( .A1(n12396), .A2(n17575), .ZN(n12397) );
  NAND2_X1 U15576 ( .A1(n12398), .A2(n12397), .ZN(n12399) );
  XOR2_X1 U15577 ( .A(n12398), .B(n12397), .Z(n17564) );
  NAND2_X1 U15578 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17564), .ZN(
        n17563) );
  NAND2_X1 U15579 ( .A1(n12399), .A2(n17563), .ZN(n17550) );
  NAND2_X1 U15580 ( .A1(n17551), .A2(n17550), .ZN(n17549) );
  NAND2_X1 U15581 ( .A1(n12400), .A2(n17549), .ZN(n12402) );
  NAND2_X1 U15582 ( .A1(n12401), .A2(n12402), .ZN(n12403) );
  XOR2_X1 U15583 ( .A(n12402), .B(n12401), .Z(n17544) );
  NAND2_X1 U15584 ( .A1(n17544), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17543) );
  NAND2_X1 U15585 ( .A1(n12403), .A2(n17543), .ZN(n17532) );
  NAND2_X1 U15586 ( .A1(n12404), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12407) );
  INV_X1 U15587 ( .A(n12407), .ZN(n12405) );
  NAND2_X1 U15588 ( .A1(n12408), .A2(n12405), .ZN(n12409) );
  NAND2_X1 U15589 ( .A1(n17531), .A2(n17532), .ZN(n17530) );
  NAND2_X1 U15590 ( .A1(n12408), .A2(n12407), .ZN(n12406) );
  OAI211_X1 U15591 ( .C1(n12408), .C2(n12407), .A(n17530), .B(n12406), .ZN(
        n17852) );
  NAND2_X1 U15592 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17852), .ZN(
        n17851) );
  NAND2_X1 U15593 ( .A1(n17805), .A2(n17401), .ZN(n17682) );
  NAND2_X1 U15594 ( .A1(n17760), .A2(n15506), .ZN(n17616) );
  AOI22_X1 U15595 ( .A1(n17520), .A2(n17615), .B1(n17601), .B2(n17616), .ZN(
        n17270) );
  NAND2_X1 U15596 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17270), .ZN(
        n17263) );
  NAND2_X1 U15597 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17263), .ZN(
        n12411) );
  NOR2_X1 U15598 ( .A1(n17520), .A2(n17601), .ZN(n17359) );
  NOR2_X1 U15599 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18618) );
  NAND3_X2 U15600 ( .A1(n18608), .A2(n18617), .A3(n18618), .ZN(n17930) );
  OAI21_X1 U15601 ( .B1(n12411), .B2(n17359), .A(n12410), .ZN(n12412) );
  NAND2_X1 U15602 ( .A1(n15506), .A2(n17391), .ZN(n16115) );
  INV_X1 U15603 ( .A(n16115), .ZN(n17264) );
  INV_X1 U15604 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16153) );
  NAND2_X1 U15605 ( .A1(n17518), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12417) );
  INV_X1 U15606 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16135) );
  OAI22_X1 U15607 ( .A1(n17518), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n12417), .B2(n16135), .ZN(n12424) );
  INV_X1 U15608 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18567) );
  INV_X1 U15609 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15536) );
  NOR3_X1 U15610 ( .A1(n15529), .A2(n16157), .A3(n15536), .ZN(n15589) );
  AOI21_X1 U15611 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18567), .A(
        n15589), .ZN(n12419) );
  NAND2_X1 U15612 ( .A1(n15530), .A2(n15536), .ZN(n15590) );
  NAND2_X1 U15613 ( .A1(n9847), .A2(n15590), .ZN(n12421) );
  NAND2_X1 U15614 ( .A1(n12419), .A2(n12421), .ZN(n12423) );
  NOR2_X1 U15615 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18567), .ZN(
        n16142) );
  AOI22_X1 U15616 ( .A1(n17518), .A2(n18567), .B1(n16142), .B2(n9847), .ZN(
        n12420) );
  AOI21_X1 U15617 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15589), .A(
        n12420), .ZN(n12422) );
  AOI22_X1 U15618 ( .A1(n12424), .A2(n12423), .B1(n12422), .B2(n12421), .ZN(
        n16144) );
  NAND2_X1 U15619 ( .A1(n16144), .A2(n17519), .ZN(n12436) );
  INV_X1 U15620 ( .A(n12427), .ZN(n16120) );
  INV_X1 U15621 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16321) );
  NAND2_X1 U15622 ( .A1(n17932), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n16145) );
  INV_X1 U15623 ( .A(n16145), .ZN(n12430) );
  NAND2_X1 U15624 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n12425), .ZN(
        n16124) );
  NOR2_X1 U15625 ( .A1(n16337), .A2(n16124), .ZN(n12426) );
  NAND2_X1 U15626 ( .A1(n12426), .A2(n17446), .ZN(n16108) );
  XNOR2_X1 U15627 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12428) );
  NOR2_X1 U15628 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17354), .ZN(
        n16121) );
  OR2_X1 U15629 ( .A1(n17980), .A2(n12426), .ZN(n16125) );
  OAI211_X1 U15630 ( .C1(n12427), .C2(n18464), .A(n16125), .B(n17609), .ZN(
        n16118) );
  NOR2_X1 U15631 ( .A1(n16121), .A2(n16118), .ZN(n16107) );
  OAI22_X1 U15632 ( .A1(n16108), .A2(n12428), .B1(n16107), .B2(n16321), .ZN(
        n12429) );
  AOI211_X1 U15633 ( .C1(n17465), .C2(n9589), .A(n12430), .B(n12429), .ZN(
        n12435) );
  INV_X1 U15634 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n20690) );
  NOR2_X1 U15635 ( .A1(n16153), .A2(n20690), .ZN(n16116) );
  NAND2_X1 U15636 ( .A1(n16116), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16134) );
  NOR2_X1 U15637 ( .A1(n17615), .A2(n16134), .ZN(n16129) );
  NAND2_X1 U15638 ( .A1(n16129), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12431) );
  XOR2_X1 U15639 ( .A(n12431), .B(n18567), .Z(n16138) );
  NAND2_X1 U15640 ( .A1(n16138), .A2(n17520), .ZN(n12434) );
  NOR3_X1 U15641 ( .A1(n16134), .A2(n17616), .A3(n16135), .ZN(n12432) );
  XOR2_X1 U15642 ( .A(n18567), .B(n12432), .Z(n16140) );
  OR2_X1 U15643 ( .A1(n16140), .A2(n17613), .ZN(n12433) );
  NAND2_X1 U15644 ( .A1(n12436), .A2(n10013), .ZN(P3_U2799) );
  NOR4_X1 U15645 ( .A1(n12441), .A2(n12440), .A3(n12439), .A4(n12438), .ZN(
        n12442) );
  OR2_X1 U15646 ( .A1(n12443), .A2(n12442), .ZN(n14297) );
  OR2_X1 U15647 ( .A1(n14297), .A2(n13250), .ZN(n12447) );
  NAND2_X1 U15648 ( .A1(n13015), .A2(n14302), .ZN(n13421) );
  OAI21_X1 U15649 ( .B1(n12444), .B2(n13250), .A(n13421), .ZN(n12445) );
  NAND2_X1 U15650 ( .A1(n12445), .A2(n14301), .ZN(n12446) );
  INV_X1 U15651 ( .A(n11254), .ZN(n13095) );
  NAND4_X1 U15652 ( .A1(n13095), .A2(n11243), .A3(n14307), .A4(n11270), .ZN(
        n13087) );
  AND2_X1 U15653 ( .A1(n14482), .A2(n13095), .ZN(n12450) );
  NAND2_X1 U15654 ( .A1(n12500), .A2(n12450), .ZN(n12467) );
  NOR4_X1 U15655 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12454) );
  NOR4_X1 U15656 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12453) );
  NOR4_X1 U15657 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12452) );
  NOR4_X1 U15658 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12451) );
  AND4_X1 U15659 ( .A1(n12454), .A2(n12453), .A3(n12452), .A4(n12451), .ZN(
        n12459) );
  NOR4_X1 U15660 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12457) );
  NOR4_X1 U15661 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12456) );
  NOR4_X1 U15662 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12455) );
  INV_X1 U15663 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20576) );
  AND4_X1 U15664 ( .A1(n12457), .A2(n12456), .A3(n12455), .A4(n20576), .ZN(
        n12458) );
  NAND2_X1 U15665 ( .A1(n12459), .A2(n12458), .ZN(n12460) );
  NOR3_X1 U15666 ( .A1(n14506), .A2(n19957), .A3(n13004), .ZN(n12461) );
  AOI22_X1 U15667 ( .A1(n14510), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14506), .ZN(n12462) );
  INV_X1 U15668 ( .A(n12462), .ZN(n12465) );
  INV_X1 U15669 ( .A(n19957), .ZN(n19959) );
  NOR2_X1 U15670 ( .A1(n13004), .A2(n19959), .ZN(n12463) );
  NAND2_X1 U15671 ( .A1(n14482), .A2(n12463), .ZN(n14484) );
  INV_X1 U15672 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16173) );
  NOR2_X1 U15673 ( .A1(n14484), .A2(n16173), .ZN(n12464) );
  NOR2_X1 U15674 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  NAND2_X1 U15675 ( .A1(n12467), .A2(n12466), .ZN(P1_U2873) );
  INV_X1 U15676 ( .A(n12468), .ZN(n12475) );
  NOR2_X1 U15677 ( .A1(n9792), .A2(n12469), .ZN(n16013) );
  AND2_X1 U15678 ( .A1(n15376), .A2(n16013), .ZN(n15287) );
  AOI21_X1 U15679 ( .B1(n15296), .B2(n15287), .A(n16014), .ZN(n15321) );
  INV_X1 U15680 ( .A(n12471), .ZN(n12472) );
  AOI21_X1 U15681 ( .B1(n16040), .B2(n12473), .A(n15084), .ZN(n12474) );
  NOR2_X1 U15682 ( .A1(n9792), .A2(n15385), .ZN(n16011) );
  NAND2_X1 U15683 ( .A1(n15376), .A2(n16011), .ZN(n15344) );
  INV_X1 U15684 ( .A(n15344), .ZN(n15297) );
  AOI22_X1 U15685 ( .A1(n15084), .A2(n10731), .B1(n12476), .B2(n15297), .ZN(
        n12484) );
  AND2_X1 U15686 ( .A1(n13933), .A2(n12477), .ZN(n12479) );
  OR2_X1 U15687 ( .A1(n12479), .A2(n12478), .ZN(n13966) );
  INV_X1 U15688 ( .A(n13966), .ZN(n18703) );
  NAND2_X1 U15689 ( .A1(n15303), .A2(n12480), .ZN(n12481) );
  NAND2_X1 U15690 ( .A1(n15281), .A2(n12481), .ZN(n18709) );
  NAND2_X1 U15691 ( .A1(n15127), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15073) );
  OAI21_X1 U15692 ( .B1(n16036), .B2(n18709), .A(n15073), .ZN(n12482) );
  AOI21_X1 U15693 ( .B1(n18703), .B2(n16038), .A(n12482), .ZN(n12483) );
  OAI21_X1 U15694 ( .B1(n12484), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12483), .ZN(n12485) );
  NAND2_X1 U15695 ( .A1(n15023), .A2(n12486), .ZN(n15024) );
  INV_X1 U15696 ( .A(n12487), .ZN(n15110) );
  INV_X1 U15697 ( .A(n15101), .ZN(n12489) );
  INV_X1 U15698 ( .A(n15091), .ZN(n12490) );
  XOR2_X1 U15699 ( .A(n15024), .B(n15025), .Z(n15078) );
  INV_X1 U15700 ( .A(n14297), .ZN(n12493) );
  NAND2_X1 U15701 ( .A1(n14303), .A2(n14307), .ZN(n14292) );
  NAND2_X1 U15702 ( .A1(n20640), .A2(n20553), .ZN(n20643) );
  NAND2_X1 U15703 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13688), .ZN(n15581) );
  AND2_X1 U15704 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20790), .ZN(n12495) );
  NAND2_X1 U15705 ( .A1(n12496), .A2(n12495), .ZN(n12497) );
  OAI211_X1 U15706 ( .C1(n15581), .C2(n20790), .A(n19942), .B(n12497), .ZN(
        n12498) );
  NAND2_X1 U15707 ( .A1(n12500), .A2(n19809), .ZN(n12617) );
  BUF_X2 U15708 ( .A(n13022), .Z(n12565) );
  INV_X1 U15709 ( .A(n19987), .ZN(n12502) );
  NAND2_X1 U15710 ( .A1(n12583), .A2(n19941), .ZN(n12504) );
  INV_X1 U15711 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13882) );
  NAND2_X1 U15712 ( .A1(n13410), .A2(n13882), .ZN(n12503) );
  NAND3_X1 U15713 ( .A1(n12504), .A2(n12565), .A3(n12503), .ZN(n12505) );
  NAND2_X1 U15714 ( .A1(n12583), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12508) );
  INV_X1 U15715 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12506) );
  NAND2_X1 U15716 ( .A1(n12565), .A2(n12506), .ZN(n12507) );
  NAND2_X1 U15717 ( .A1(n12508), .A2(n12507), .ZN(n13414) );
  XNOR2_X1 U15718 ( .A(n12509), .B(n13414), .ZN(n13411) );
  NAND2_X1 U15719 ( .A1(n13411), .A2(n13410), .ZN(n13409) );
  NAND2_X1 U15720 ( .A1(n13409), .A2(n12509), .ZN(n13505) );
  INV_X1 U15721 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13953) );
  NAND2_X1 U15722 ( .A1(n12577), .A2(n13953), .ZN(n12513) );
  NAND2_X1 U15723 ( .A1(n12583), .A2(n19954), .ZN(n12511) );
  NAND2_X1 U15724 ( .A1(n13410), .A2(n13953), .ZN(n12510) );
  NAND3_X1 U15725 ( .A1(n12511), .A2(n12565), .A3(n12510), .ZN(n12512) );
  AND2_X1 U15726 ( .A1(n12513), .A2(n12512), .ZN(n13504) );
  MUX2_X1 U15727 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12516) );
  OAI21_X1 U15728 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13413), .A(
        n12516), .ZN(n13555) );
  INV_X1 U15729 ( .A(n12583), .ZN(n12576) );
  MUX2_X1 U15730 ( .A(n12577), .B(n12576), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12518) );
  NAND2_X1 U15731 ( .A1(n12576), .A2(n12520), .ZN(n12541) );
  OAI21_X1 U15732 ( .B1(n13410), .B2(n19922), .A(n12541), .ZN(n12517) );
  NOR2_X1 U15733 ( .A1(n12518), .A2(n12517), .ZN(n13568) );
  INV_X1 U15734 ( .A(n12580), .ZN(n12519) );
  INV_X1 U15735 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19850) );
  NAND2_X1 U15736 ( .A1(n12519), .A2(n19850), .ZN(n12523) );
  NAND2_X1 U15737 ( .A1(n12565), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12521) );
  OAI211_X1 U15738 ( .C1(n12520), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12583), .B(
        n12521), .ZN(n12522) );
  AND2_X1 U15739 ( .A1(n12523), .A2(n12522), .ZN(n15873) );
  NAND2_X1 U15740 ( .A1(n15874), .A2(n15873), .ZN(n15876) );
  MUX2_X1 U15741 ( .A(n12577), .B(n12576), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12526) );
  NAND2_X1 U15742 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12520), .ZN(
        n12524) );
  NAND2_X1 U15743 ( .A1(n12541), .A2(n12524), .ZN(n12525) );
  NAND2_X1 U15744 ( .A1(n12565), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12528) );
  OAI211_X1 U15745 ( .C1(n12520), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12583), .B(
        n12528), .ZN(n12529) );
  OAI21_X1 U15746 ( .B1(n12580), .B2(P1_EBX_REG_7__SCAN_IN), .A(n12529), .ZN(
        n13703) );
  MUX2_X1 U15747 ( .A(n12586), .B(n12583), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12532) );
  NAND2_X1 U15748 ( .A1(n12520), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12530) );
  AND2_X1 U15749 ( .A1(n12541), .A2(n12530), .ZN(n12531) );
  NAND2_X1 U15750 ( .A1(n12532), .A2(n12531), .ZN(n13827) );
  NAND2_X1 U15751 ( .A1(n12565), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12533) );
  OAI211_X1 U15752 ( .C1(n12520), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12583), .B(
        n12533), .ZN(n12534) );
  OAI21_X1 U15753 ( .B1(n12580), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12534), .ZN(
        n15837) );
  MUX2_X1 U15754 ( .A(n12577), .B(n12576), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12537) );
  NAND2_X1 U15755 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n12520), .ZN(
        n12535) );
  NAND2_X1 U15756 ( .A1(n12541), .A2(n12535), .ZN(n12536) );
  NOR2_X1 U15757 ( .A1(n12537), .A2(n12536), .ZN(n13976) );
  NOR2_X2 U15758 ( .A1(n15840), .A2(n13976), .ZN(n14081) );
  MUX2_X1 U15759 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12539) );
  OR2_X1 U15760 ( .A1(n13413), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12538) );
  MUX2_X1 U15761 ( .A(n12586), .B(n12583), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12543) );
  NAND2_X1 U15762 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n12520), .ZN(
        n12540) );
  AND2_X1 U15763 ( .A1(n12541), .A2(n12540), .ZN(n12542) );
  NAND2_X1 U15764 ( .A1(n12543), .A2(n12542), .ZN(n14124) );
  MUX2_X1 U15765 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12544) );
  OAI21_X1 U15766 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13413), .A(
        n12544), .ZN(n14106) );
  MUX2_X1 U15767 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12545) );
  OAI21_X1 U15768 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n13413), .A(
        n12545), .ZN(n12546) );
  INV_X1 U15769 ( .A(n12546), .ZN(n14119) );
  NAND2_X1 U15770 ( .A1(n12583), .A2(n15809), .ZN(n12549) );
  INV_X1 U15771 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U15772 ( .A1(n13410), .A2(n12547), .ZN(n12548) );
  NAND3_X1 U15773 ( .A1(n12549), .A2(n12565), .A3(n12548), .ZN(n12550) );
  OAI21_X1 U15774 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(n12586), .A(n12550), .ZN(
        n14120) );
  NAND2_X1 U15775 ( .A1(n14119), .A2(n14120), .ZN(n12551) );
  NAND2_X1 U15776 ( .A1(n12583), .A2(n12552), .ZN(n12554) );
  INV_X1 U15777 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14161) );
  NAND2_X1 U15778 ( .A1(n13410), .A2(n14161), .ZN(n12553) );
  NAND3_X1 U15779 ( .A1(n12554), .A2(n12565), .A3(n12553), .ZN(n12555) );
  OAI21_X1 U15780 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(n12586), .A(n12555), .ZN(
        n14153) );
  MUX2_X1 U15781 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12557) );
  OR2_X1 U15782 ( .A1(n13413), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12556) );
  INV_X1 U15783 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14455) );
  NAND2_X1 U15784 ( .A1(n12577), .A2(n14455), .ZN(n12561) );
  INV_X1 U15785 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15700) );
  NAND2_X1 U15786 ( .A1(n12583), .A2(n15700), .ZN(n12559) );
  NAND2_X1 U15787 ( .A1(n13410), .A2(n14455), .ZN(n12558) );
  NAND3_X1 U15788 ( .A1(n12559), .A2(n12565), .A3(n12558), .ZN(n12560) );
  MUX2_X1 U15789 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12562) );
  OAI21_X1 U15790 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13413), .A(
        n12562), .ZN(n14445) );
  MUX2_X1 U15791 ( .A(n12586), .B(n12583), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12564) );
  NAND2_X1 U15792 ( .A1(n12520), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12563) );
  NAND2_X1 U15793 ( .A1(n12564), .A2(n12563), .ZN(n14441) );
  MUX2_X1 U15794 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12566) );
  OAI21_X1 U15795 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13413), .A(
        n12566), .ZN(n14431) );
  NOR2_X2 U15796 ( .A1(n14440), .A2(n14431), .ZN(n14401) );
  INV_X1 U15797 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U15798 ( .A1(n12577), .A2(n14428), .ZN(n12570) );
  INV_X1 U15799 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15763) );
  NAND2_X1 U15800 ( .A1(n12583), .A2(n15763), .ZN(n12568) );
  NAND2_X1 U15801 ( .A1(n13410), .A2(n14428), .ZN(n12567) );
  NAND3_X1 U15802 ( .A1(n12568), .A2(n12565), .A3(n12567), .ZN(n12569) );
  AND2_X1 U15803 ( .A1(n12570), .A2(n12569), .ZN(n14402) );
  INV_X1 U15804 ( .A(n14402), .ZN(n12571) );
  NAND2_X1 U15805 ( .A1(n14401), .A2(n12571), .ZN(n14404) );
  MUX2_X1 U15806 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12572) );
  OAI21_X1 U15807 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n13413), .A(
        n12572), .ZN(n14387) );
  NAND2_X1 U15808 ( .A1(n12583), .A2(n14723), .ZN(n12573) );
  OAI211_X1 U15809 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n12520), .A(n12573), .B(
        n12565), .ZN(n12574) );
  OAI21_X1 U15810 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n12586), .A(n12574), .ZN(
        n14375) );
  MUX2_X1 U15811 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12575) );
  OAI21_X1 U15812 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n13413), .A(
        n12575), .ZN(n14362) );
  MUX2_X1 U15813 ( .A(n12577), .B(n12576), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12579) );
  AND2_X1 U15814 ( .A1(n12520), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12578) );
  NOR2_X1 U15815 ( .A1(n12579), .A2(n12578), .ZN(n14351) );
  MUX2_X1 U15816 ( .A(n12580), .B(n12565), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12582) );
  OR2_X1 U15817 ( .A1(n13413), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12581) );
  AND2_X1 U15818 ( .A1(n12582), .A2(n12581), .ZN(n14332) );
  AND2_X2 U15819 ( .A1(n14331), .A2(n14332), .ZN(n14334) );
  NAND2_X1 U15820 ( .A1(n12583), .A2(n14682), .ZN(n12584) );
  OAI211_X1 U15821 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n12520), .A(n12584), .B(
        n12565), .ZN(n12585) );
  OAI21_X1 U15822 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(n12586), .A(n12585), .ZN(
        n14323) );
  INV_X1 U15823 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14420) );
  NAND2_X1 U15824 ( .A1(n13410), .A2(n14420), .ZN(n12588) );
  OR2_X1 U15825 ( .A1(n13413), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12587) );
  NAND2_X1 U15826 ( .A1(n12587), .A2(n12588), .ZN(n13092) );
  MUX2_X1 U15827 ( .A(n12588), .B(n13092), .S(n12565), .Z(n14316) );
  NOR2_X2 U15828 ( .A1(n14322), .A2(n14316), .ZN(n14318) );
  AND2_X1 U15829 ( .A1(n12520), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12590) );
  AOI21_X1 U15830 ( .B1(n13413), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12590), .ZN(
        n13094) );
  AOI22_X1 U15831 ( .A1(n13413), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12520), .ZN(n12593) );
  XNOR2_X2 U15832 ( .A(n12594), .B(n12593), .ZN(n14419) );
  NAND2_X1 U15833 ( .A1(n19979), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12602) );
  AND2_X1 U15834 ( .A1(n20647), .A2(n20641), .ZN(n15575) );
  NOR2_X1 U15835 ( .A1(n12602), .A2(n15575), .ZN(n12595) );
  NOR2_X1 U15836 ( .A1(n12596), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15599) );
  OAI21_X1 U15837 ( .B1(n19979), .B2(n15599), .A(n20647), .ZN(n13005) );
  NOR2_X1 U15838 ( .A1(n13005), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12604) );
  NAND2_X1 U15839 ( .A1(n15677), .A2(n14405), .ZN(n19789) );
  INV_X1 U15840 ( .A(n19789), .ZN(n13975) );
  AND2_X1 U15841 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n12610) );
  INV_X1 U15842 ( .A(n14405), .ZN(n14365) );
  INV_X1 U15843 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20722) );
  INV_X1 U15844 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15675) );
  NAND2_X1 U15845 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .ZN(n13973) );
  INV_X1 U15846 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n19786) );
  INV_X1 U15847 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19804) );
  NAND2_X1 U15848 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19799) );
  OR3_X1 U15849 ( .A1(n19786), .A2(n19804), .A3(n19799), .ZN(n19764) );
  INV_X1 U15850 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n19774) );
  NOR3_X1 U15851 ( .A1(n19764), .A2(n14651), .A3(n19774), .ZN(n13974) );
  INV_X1 U15852 ( .A(n13974), .ZN(n12597) );
  NAND2_X1 U15853 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14109) );
  NOR3_X1 U15854 ( .A1(n13973), .A2(n12597), .A3(n14109), .ZN(n12598) );
  NAND4_X1 U15855 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .A4(n12598), .ZN(n15676) );
  NOR2_X1 U15856 ( .A1(n15675), .A2(n15676), .ZN(n14167) );
  NAND3_X1 U15857 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n15640) );
  INV_X1 U15858 ( .A(n15640), .ZN(n15641) );
  NAND3_X1 U15859 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14167), .A3(n15641), 
        .ZN(n15636) );
  NOR2_X1 U15860 ( .A1(n20722), .A2(n15636), .ZN(n15622) );
  INV_X1 U15861 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15609) );
  INV_X1 U15862 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15633) );
  NOR2_X1 U15863 ( .A1(n15609), .A2(n15633), .ZN(n14409) );
  AND2_X1 U15864 ( .A1(n14409), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n12599) );
  NAND2_X1 U15865 ( .A1(n15622), .A2(n12599), .ZN(n14391) );
  INV_X1 U15866 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14572) );
  OR2_X1 U15867 ( .A1(n14391), .A2(n14572), .ZN(n14382) );
  NAND2_X1 U15868 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n12600) );
  NOR2_X1 U15869 ( .A1(n14382), .A2(n12600), .ZN(n14353) );
  NAND2_X1 U15870 ( .A1(n14353), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14340) );
  NAND2_X1 U15871 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n12601) );
  OR2_X1 U15872 ( .A1(n14340), .A2(n12601), .ZN(n12608) );
  OAI21_X1 U15873 ( .B1(n14365), .B2(n12608), .A(n19789), .ZN(n14311) );
  OAI21_X1 U15874 ( .B1(n13975), .B2(n12610), .A(n14311), .ZN(n14249) );
  INV_X1 U15875 ( .A(n12602), .ZN(n12603) );
  NOR2_X1 U15876 ( .A1(n12604), .A2(n12603), .ZN(n12605) );
  INV_X1 U15877 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14418) );
  OAI22_X1 U15878 ( .A1(n19825), .A2(n14418), .B1(n12607), .B2(n19769), .ZN(
        n12613) );
  INV_X1 U15879 ( .A(n12608), .ZN(n12609) );
  NAND2_X1 U15880 ( .A1(n15623), .A2(n12609), .ZN(n14315) );
  INV_X1 U15881 ( .A(n12610), .ZN(n12611) );
  NOR3_X1 U15882 ( .A1(n14315), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n12611), 
        .ZN(n12612) );
  AOI211_X1 U15883 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14249), .A(n12613), 
        .B(n12612), .ZN(n12614) );
  NAND2_X1 U15884 ( .A1(n12617), .A2(n12616), .ZN(P1_U2809) );
  NAND2_X1 U15885 ( .A1(n13444), .A2(n12635), .ZN(n12623) );
  NAND2_X1 U15886 ( .A1(n13785), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12619) );
  NOR2_X1 U15887 ( .A1(n19687), .A2(n19696), .ZN(n19450) );
  OAI21_X1 U15888 ( .B1(n12626), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19681), .ZN(n12620) );
  NOR2_X1 U15889 ( .A1(n12620), .A2(n19517), .ZN(n12621) );
  AOI21_X1 U15890 ( .B1(n12636), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12621), .ZN(n12622) );
  NOR2_X1 U15891 ( .A1(n12863), .A2(n12818), .ZN(n12624) );
  NAND2_X1 U15892 ( .A1(n12645), .A2(n12624), .ZN(n13575) );
  NAND2_X1 U15893 ( .A1(n13533), .A2(n12635), .ZN(n12630) );
  NAND2_X1 U15894 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19347) );
  NAND2_X1 U15895 ( .A1(n19347), .A2(n19687), .ZN(n12628) );
  INV_X1 U15896 ( .A(n12626), .ZN(n12627) );
  AND2_X1 U15897 ( .A1(n19390), .A2(n19681), .ZN(n19164) );
  AOI21_X1 U15898 ( .B1(n12636), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n19164), .ZN(n12629) );
  INV_X1 U15899 ( .A(n13383), .ZN(n12642) );
  NAND2_X1 U15900 ( .A1(n12636), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12633) );
  NAND2_X1 U15901 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19696), .ZN(
        n19200) );
  NAND2_X1 U15902 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19703), .ZN(
        n19317) );
  NAND2_X1 U15903 ( .A1(n19200), .A2(n19317), .ZN(n19163) );
  NAND2_X1 U15904 ( .A1(n19681), .A2(n19163), .ZN(n19322) );
  NAND2_X1 U15905 ( .A1(n12633), .A2(n19322), .ZN(n12634) );
  INV_X1 U15906 ( .A(n12635), .ZN(n12990) );
  AOI22_X1 U15907 ( .A1(n12636), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19681), .B2(n19703), .ZN(n12637) );
  NAND2_X1 U15908 ( .A1(n13286), .A2(n13287), .ZN(n12641) );
  INV_X1 U15909 ( .A(n15405), .ZN(n12639) );
  NAND2_X1 U15910 ( .A1(n12639), .A2(n12638), .ZN(n12640) );
  NAND2_X1 U15911 ( .A1(n12642), .A2(n9702), .ZN(n12644) );
  NAND2_X1 U15912 ( .A1(n12645), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13577) );
  NAND4_X1 U15913 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .A4(P2_INSTQUEUE_REG_0__5__SCAN_IN), 
        .ZN(n12646) );
  AOI22_X1 U15914 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15915 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10294), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15916 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15917 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12647) );
  NAND4_X1 U15918 ( .A1(n12650), .A2(n12649), .A3(n12648), .A4(n12647), .ZN(
        n12656) );
  AOI22_X1 U15919 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U15920 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15921 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10302), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U15922 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12651) );
  NAND4_X1 U15923 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        n12655) );
  NOR2_X1 U15924 ( .A1(n12656), .A2(n12655), .ZN(n13963) );
  INV_X1 U15925 ( .A(n13963), .ZN(n12671) );
  AOI22_X1 U15926 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10292), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15927 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U15928 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12658) );
  AOI22_X1 U15929 ( .A1(n12749), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12657) );
  NAND4_X1 U15930 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n12666) );
  AOI22_X1 U15931 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15932 ( .A1(n10249), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15933 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U15934 ( .A1(n10903), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12661) );
  NAND4_X1 U15935 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12665) );
  OR2_X1 U15936 ( .A1(n12666), .A2(n12665), .ZN(n13936) );
  INV_X1 U15937 ( .A(n12667), .ZN(n13813) );
  INV_X1 U15938 ( .A(n12668), .ZN(n13819) );
  INV_X1 U15939 ( .A(n13663), .ZN(n12669) );
  NOR2_X1 U15940 ( .A1(n13546), .A2(n13560), .ZN(n13561) );
  AND2_X1 U15941 ( .A1(n12669), .A2(n13561), .ZN(n13612) );
  AND2_X1 U15942 ( .A1(n13614), .A2(n13612), .ZN(n13613) );
  INV_X1 U15943 ( .A(n13892), .ZN(n12670) );
  AOI22_X1 U15944 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U15945 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10294), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U15946 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U15947 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12673) );
  NAND4_X1 U15948 ( .A1(n12676), .A2(n12675), .A3(n12674), .A4(n12673), .ZN(
        n12682) );
  AOI22_X1 U15949 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U15950 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12679) );
  AOI22_X1 U15951 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12697), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U15952 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12677) );
  NAND4_X1 U15953 ( .A1(n12680), .A2(n12679), .A3(n12678), .A4(n12677), .ZN(
        n12681) );
  NOR2_X1 U15954 ( .A1(n12682), .A2(n12681), .ZN(n14019) );
  AOI22_X1 U15955 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15956 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n9590), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U15957 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12748), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15958 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12683) );
  NAND4_X1 U15959 ( .A1(n12686), .A2(n12685), .A3(n12684), .A4(n12683), .ZN(
        n12692) );
  AOI22_X1 U15960 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12690) );
  AOI22_X1 U15961 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U15962 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12697), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U15963 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12687) );
  NAND4_X1 U15964 ( .A1(n12690), .A2(n12689), .A3(n12688), .A4(n12687), .ZN(
        n12691) );
  AND2_X2 U15965 ( .A1(n14018), .A2(n14086), .ZN(n14084) );
  AOI22_X1 U15966 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15967 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9590), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U15968 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U15969 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12693) );
  NAND4_X1 U15970 ( .A1(n12696), .A2(n12695), .A3(n12694), .A4(n12693), .ZN(
        n12703) );
  AOI22_X1 U15971 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15972 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U15973 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12697), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U15974 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12698) );
  NAND4_X1 U15975 ( .A1(n12701), .A2(n12700), .A3(n12699), .A4(n12698), .ZN(
        n12702) );
  AOI22_X1 U15976 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10292), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15977 ( .A1(n10294), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U15978 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15979 ( .A1(n12749), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10296), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12704) );
  NAND4_X1 U15980 ( .A1(n12707), .A2(n12706), .A3(n12705), .A4(n12704), .ZN(
        n12713) );
  AOI22_X1 U15981 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15982 ( .A1(n10249), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15983 ( .A1(n10302), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15984 ( .A1(n10903), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12708) );
  NAND4_X1 U15985 ( .A1(n12711), .A2(n12710), .A3(n12709), .A4(n12708), .ZN(
        n12712) );
  NOR2_X1 U15986 ( .A1(n12713), .A2(n12712), .ZN(n14869) );
  AOI22_X1 U15987 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15988 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n9590), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15989 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12748), .B1(
        n10295), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U15990 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12714) );
  NAND4_X1 U15991 ( .A1(n12717), .A2(n12716), .A3(n12715), .A4(n12714), .ZN(
        n12723) );
  AOI22_X1 U15992 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15993 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15994 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12697), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U15995 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12718) );
  NAND4_X1 U15996 ( .A1(n12721), .A2(n12720), .A3(n12719), .A4(n12718), .ZN(
        n12722) );
  NOR2_X1 U15997 ( .A1(n12723), .A2(n12722), .ZN(n14860) );
  INV_X1 U15998 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12727) );
  INV_X1 U15999 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12726) );
  OAI22_X1 U16000 ( .A1(n12724), .A2(n12727), .B1(n12907), .B2(n12726), .ZN(
        n12731) );
  INV_X1 U16001 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19260) );
  INV_X1 U16002 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13848) );
  OAI22_X1 U16003 ( .A1(n12902), .A2(n19260), .B1(n12905), .B2(n13848), .ZN(
        n12730) );
  NOR2_X1 U16004 ( .A1(n12731), .A2(n12730), .ZN(n12735) );
  AOI22_X1 U16005 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U16006 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9592), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12733) );
  XNOR2_X1 U16007 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12932) );
  NAND4_X1 U16008 ( .A1(n12735), .A2(n12734), .A3(n12733), .A4(n12932), .ZN(
        n12746) );
  INV_X1 U16009 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12737) );
  INV_X1 U16010 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12736) );
  OAI22_X1 U16011 ( .A1(n12724), .A2(n12737), .B1(n12902), .B2(n12736), .ZN(
        n12741) );
  INV_X1 U16012 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12739) );
  INV_X1 U16013 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12738) );
  OAI22_X1 U16014 ( .A1(n12907), .A2(n12739), .B1(n12905), .B2(n12738), .ZN(
        n12740) );
  NOR2_X1 U16015 ( .A1(n12741), .A2(n12740), .ZN(n12744) );
  AOI22_X1 U16016 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U16017 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9591), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12742) );
  NAND4_X1 U16018 ( .A1(n12744), .A2(n12743), .A3(n12942), .A4(n12742), .ZN(
        n12745) );
  AND2_X1 U16019 ( .A1(n12746), .A2(n12745), .ZN(n12786) );
  NAND2_X1 U16020 ( .A1(n10208), .A2(n12786), .ZN(n12760) );
  AOI22_X1 U16021 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10292), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12753) );
  AOI22_X1 U16022 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9590), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U16023 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10295), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16024 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10296), .B1(
        n12749), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12750) );
  NAND4_X1 U16025 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12759) );
  AOI22_X1 U16026 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10301), .B1(
        n10250), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U16027 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10361), .B1(
        n10249), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U16028 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10302), .B1(
        n10917), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U16029 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10903), .B1(
        n10262), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12754) );
  NAND4_X1 U16030 ( .A1(n12757), .A2(n12756), .A3(n12755), .A4(n12754), .ZN(
        n12758) );
  NOR2_X1 U16031 ( .A1(n12759), .A2(n12758), .ZN(n12762) );
  XOR2_X1 U16032 ( .A(n12760), .B(n12762), .Z(n12785) );
  NAND2_X1 U16033 ( .A1(n9584), .A2(n12786), .ZN(n14854) );
  NOR2_X1 U16034 ( .A1(n14852), .A2(n14854), .ZN(n14853) );
  INV_X1 U16035 ( .A(n12762), .ZN(n12763) );
  AND2_X1 U16036 ( .A1(n12763), .A2(n12786), .ZN(n12784) );
  OAI22_X1 U16037 ( .A1(n12724), .A2(n12765), .B1(n12902), .B2(n12764), .ZN(
        n12768) );
  OAI22_X1 U16038 ( .A1(n12907), .A2(n12766), .B1(n12905), .B2(n19064), .ZN(
        n12767) );
  NOR2_X1 U16039 ( .A1(n12768), .A2(n12767), .ZN(n12771) );
  AOI22_X1 U16040 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U16041 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12769) );
  NAND4_X1 U16042 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12932), .ZN(
        n12783) );
  OAI22_X1 U16043 ( .A1(n12724), .A2(n12773), .B1(n12902), .B2(n12772), .ZN(
        n12777) );
  OAI22_X1 U16044 ( .A1(n12907), .A2(n12775), .B1(n12905), .B2(n12774), .ZN(
        n12776) );
  NOR2_X1 U16045 ( .A1(n12777), .A2(n12776), .ZN(n12781) );
  AOI22_X1 U16046 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12780) );
  AOI22_X1 U16047 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12779) );
  NAND4_X1 U16048 ( .A1(n12781), .A2(n12780), .A3(n12942), .A4(n12779), .ZN(
        n12782) );
  AND2_X1 U16049 ( .A1(n12783), .A2(n12782), .ZN(n12787) );
  NAND2_X1 U16050 ( .A1(n12784), .A2(n12787), .ZN(n12790) );
  OAI211_X1 U16051 ( .C1(n12784), .C2(n12787), .A(n13574), .B(n12790), .ZN(
        n14844) );
  INV_X1 U16052 ( .A(n12786), .ZN(n12788) );
  NAND2_X1 U16053 ( .A1(n9583), .A2(n12787), .ZN(n14846) );
  NOR3_X1 U16054 ( .A1(n9978), .A2(n12788), .A3(n14846), .ZN(n12789) );
  INV_X1 U16055 ( .A(n12790), .ZN(n12809) );
  INV_X1 U16056 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12791) );
  INV_X1 U16057 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13741) );
  OAI22_X1 U16058 ( .A1(n12724), .A2(n12791), .B1(n12902), .B2(n13741), .ZN(
        n12794) );
  INV_X1 U16059 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12792) );
  OAI22_X1 U16060 ( .A1(n12907), .A2(n12792), .B1(n12905), .B2(n13853), .ZN(
        n12793) );
  NOR2_X1 U16061 ( .A1(n12794), .A2(n12793), .ZN(n12797) );
  AOI22_X1 U16062 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U16063 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12795) );
  NAND4_X1 U16064 ( .A1(n12797), .A2(n12796), .A3(n12795), .A4(n12932), .ZN(
        n12808) );
  INV_X1 U16065 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12799) );
  INV_X1 U16066 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12798) );
  OAI22_X1 U16067 ( .A1(n12724), .A2(n12799), .B1(n12902), .B2(n12798), .ZN(
        n12803) );
  INV_X1 U16068 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12801) );
  INV_X1 U16069 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12800) );
  OAI22_X1 U16070 ( .A1(n12907), .A2(n12801), .B1(n12905), .B2(n12800), .ZN(
        n12802) );
  NOR2_X1 U16071 ( .A1(n12803), .A2(n12802), .ZN(n12806) );
  AOI22_X1 U16072 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U16073 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12804) );
  NAND4_X1 U16074 ( .A1(n12806), .A2(n12805), .A3(n12942), .A4(n12804), .ZN(
        n12807) );
  AND2_X1 U16075 ( .A1(n12808), .A2(n12807), .ZN(n12811) );
  NAND2_X1 U16076 ( .A1(n12809), .A2(n12811), .ZN(n12836) );
  OAI211_X1 U16077 ( .C1(n12809), .C2(n12811), .A(n13574), .B(n12836), .ZN(
        n12814) );
  XNOR2_X1 U16078 ( .A(n12813), .B(n12810), .ZN(n14833) );
  INV_X1 U16079 ( .A(n12811), .ZN(n12812) );
  NOR2_X1 U16080 ( .A1(n10208), .A2(n12812), .ZN(n14832) );
  NAND2_X1 U16081 ( .A1(n14833), .A2(n14832), .ZN(n14831) );
  OAI22_X1 U16082 ( .A1(n12724), .A2(n12817), .B1(n12902), .B2(n12816), .ZN(
        n12821) );
  OAI22_X1 U16083 ( .A1(n12907), .A2(n12819), .B1(n12905), .B2(n12818), .ZN(
        n12820) );
  NOR2_X1 U16084 ( .A1(n12821), .A2(n12820), .ZN(n12824) );
  AOI22_X1 U16085 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U16086 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12822) );
  NAND4_X1 U16087 ( .A1(n12824), .A2(n12823), .A3(n12822), .A4(n12932), .ZN(
        n12835) );
  OAI22_X1 U16088 ( .A1(n12724), .A2(n12826), .B1(n12902), .B2(n12825), .ZN(
        n12830) );
  OAI22_X1 U16089 ( .A1(n12907), .A2(n12828), .B1(n12905), .B2(n12827), .ZN(
        n12829) );
  NOR2_X1 U16090 ( .A1(n12830), .A2(n12829), .ZN(n12833) );
  AOI22_X1 U16091 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U16092 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12831) );
  NAND4_X1 U16093 ( .A1(n12833), .A2(n12832), .A3(n12942), .A4(n12831), .ZN(
        n12834) );
  NAND2_X1 U16094 ( .A1(n12835), .A2(n12834), .ZN(n12838) );
  AOI21_X1 U16095 ( .B1(n12836), .B2(n12838), .A(n12863), .ZN(n12837) );
  NAND2_X1 U16096 ( .A1(n12837), .A2(n12864), .ZN(n12840) );
  NOR2_X1 U16097 ( .A1(n10208), .A2(n12838), .ZN(n14824) );
  INV_X1 U16098 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12844) );
  INV_X1 U16099 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12843) );
  OAI22_X1 U16100 ( .A1(n12724), .A2(n12844), .B1(n12902), .B2(n12843), .ZN(
        n12848) );
  INV_X1 U16101 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12846) );
  INV_X1 U16102 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12845) );
  OAI22_X1 U16103 ( .A1(n12907), .A2(n12846), .B1(n12905), .B2(n12845), .ZN(
        n12847) );
  NOR2_X1 U16104 ( .A1(n12848), .A2(n12847), .ZN(n12851) );
  AOI22_X1 U16105 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U16106 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12849) );
  NAND4_X1 U16107 ( .A1(n12851), .A2(n12850), .A3(n12849), .A4(n12932), .ZN(
        n12862) );
  INV_X1 U16108 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12853) );
  INV_X1 U16109 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12852) );
  OAI22_X1 U16110 ( .A1(n12724), .A2(n12853), .B1(n12902), .B2(n12852), .ZN(
        n12857) );
  INV_X1 U16111 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12855) );
  INV_X1 U16112 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12854) );
  OAI22_X1 U16113 ( .A1(n12907), .A2(n12855), .B1(n12905), .B2(n12854), .ZN(
        n12856) );
  NOR2_X1 U16114 ( .A1(n12857), .A2(n12856), .ZN(n12860) );
  AOI22_X1 U16115 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U16116 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12858) );
  NAND4_X1 U16117 ( .A1(n12860), .A2(n12859), .A3(n12942), .A4(n12858), .ZN(
        n12861) );
  NAND2_X1 U16118 ( .A1(n12862), .A2(n12861), .ZN(n12867) );
  NOR2_X1 U16119 ( .A1(n12864), .A2(n12867), .ZN(n12890) );
  AOI211_X1 U16120 ( .C1(n12867), .C2(n12864), .A(n12863), .B(n12890), .ZN(
        n12865) );
  INV_X1 U16121 ( .A(n12867), .ZN(n12868) );
  NAND2_X1 U16122 ( .A1(n9584), .A2(n12868), .ZN(n14819) );
  INV_X1 U16123 ( .A(n12869), .ZN(n12889) );
  INV_X1 U16124 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12871) );
  INV_X1 U16125 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12870) );
  OAI22_X1 U16126 ( .A1(n12724), .A2(n12871), .B1(n12902), .B2(n12870), .ZN(
        n12874) );
  OAI22_X1 U16127 ( .A1(n12907), .A2(n12872), .B1(n12905), .B2(n13647), .ZN(
        n12873) );
  NOR2_X1 U16128 ( .A1(n12874), .A2(n12873), .ZN(n12877) );
  AOI22_X1 U16129 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U16130 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12875) );
  NAND4_X1 U16131 ( .A1(n12877), .A2(n12876), .A3(n12875), .A4(n12932), .ZN(
        n12888) );
  OAI22_X1 U16132 ( .A1(n12724), .A2(n12879), .B1(n12902), .B2(n12878), .ZN(
        n12883) );
  OAI22_X1 U16133 ( .A1(n12907), .A2(n12881), .B1(n12905), .B2(n12880), .ZN(
        n12882) );
  NOR2_X1 U16134 ( .A1(n12883), .A2(n12882), .ZN(n12886) );
  AOI22_X1 U16135 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12885) );
  AOI22_X1 U16136 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12884) );
  NAND4_X1 U16137 ( .A1(n12886), .A2(n12885), .A3(n12942), .A4(n12884), .ZN(
        n12887) );
  AND2_X1 U16138 ( .A1(n12888), .A2(n12887), .ZN(n14811) );
  INV_X1 U16139 ( .A(n12890), .ZN(n14810) );
  NAND2_X1 U16140 ( .A1(n10208), .A2(n14811), .ZN(n12891) );
  NOR2_X1 U16141 ( .A1(n14810), .A2(n12891), .ZN(n12916) );
  INV_X1 U16142 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12893) );
  OAI22_X1 U16143 ( .A1(n12724), .A2(n12893), .B1(n12907), .B2(n12892), .ZN(
        n12897) );
  OAI22_X1 U16144 ( .A1(n12902), .A2(n12895), .B1(n12905), .B2(n12894), .ZN(
        n12896) );
  NOR2_X1 U16145 ( .A1(n12897), .A2(n12896), .ZN(n12900) );
  AOI22_X1 U16146 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12899) );
  INV_X1 U16147 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n19123) );
  AOI22_X1 U16148 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12898) );
  NAND4_X1 U16149 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12932), .ZN(
        n12914) );
  OAI22_X1 U16150 ( .A1(n12724), .A2(n12903), .B1(n12902), .B2(n12901), .ZN(
        n12909) );
  OAI22_X1 U16151 ( .A1(n12907), .A2(n12906), .B1(n12905), .B2(n12904), .ZN(
        n12908) );
  NOR2_X1 U16152 ( .A1(n12909), .A2(n12908), .ZN(n12912) );
  AOI22_X1 U16153 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U16154 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12910) );
  NAND4_X1 U16155 ( .A1(n12912), .A2(n12911), .A3(n12942), .A4(n12910), .ZN(
        n12913) );
  AND2_X1 U16156 ( .A1(n12914), .A2(n12913), .ZN(n12915) );
  NAND2_X1 U16157 ( .A1(n12916), .A2(n12915), .ZN(n12926) );
  OAI21_X1 U16158 ( .B1(n12916), .B2(n12915), .A(n12926), .ZN(n12917) );
  INV_X1 U16159 ( .A(n12928), .ZN(n12920) );
  NAND2_X1 U16160 ( .A1(n12918), .A2(n12917), .ZN(n14281) );
  NAND2_X1 U16161 ( .A1(n16055), .A2(n16058), .ZN(n13462) );
  XNOR2_X1 U16162 ( .A(n14813), .B(n12921), .ZN(n15906) );
  NAND2_X1 U16163 ( .A1(n14873), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12922) );
  INV_X1 U16164 ( .A(n12926), .ZN(n12927) );
  NOR2_X1 U16165 ( .A1(n12928), .A2(n12927), .ZN(n12950) );
  AOI22_X1 U16166 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16167 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12930) );
  NAND2_X1 U16168 ( .A1(n12931), .A2(n12930), .ZN(n12948) );
  AOI22_X1 U16169 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12939), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U16170 ( .A1(n12938), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12933) );
  NAND3_X1 U16171 ( .A1(n12934), .A2(n12933), .A3(n12932), .ZN(n12947) );
  AOI22_X1 U16172 ( .A1(n12778), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12935), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U16173 ( .A1(n10033), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10236), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12936) );
  NAND2_X1 U16174 ( .A1(n12937), .A2(n12936), .ZN(n12946) );
  AOI22_X1 U16175 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12938), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U16176 ( .A1(n12941), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12940), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12943) );
  NAND3_X1 U16177 ( .A1(n12944), .A2(n12943), .A3(n12942), .ZN(n12945) );
  OAI22_X1 U16178 ( .A1(n12948), .A2(n12947), .B1(n12946), .B2(n12945), .ZN(
        n12949) );
  XNOR2_X1 U16179 ( .A(n12950), .B(n12949), .ZN(n14280) );
  INV_X1 U16180 ( .A(n9721), .ZN(n16057) );
  NAND2_X1 U16181 ( .A1(n16057), .A2(n13221), .ZN(n16065) );
  NAND2_X1 U16182 ( .A1(n11054), .A2(n19586), .ZN(n16062) );
  OAI22_X1 U16183 ( .A1(n16055), .A2(n16060), .B1(n16065), .B2(n16062), .ZN(
        n13464) );
  AND2_X1 U16184 ( .A1(n12951), .A2(n16067), .ZN(n12952) );
  AOI21_X1 U16185 ( .B1(n12956), .B2(n14284), .A(n12955), .ZN(n13164) );
  NOR4_X1 U16186 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12962) );
  NOR4_X1 U16187 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12961) );
  NOR4_X1 U16188 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12960) );
  NOR4_X1 U16189 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12959) );
  NAND4_X1 U16190 ( .A1(n12962), .A2(n12961), .A3(n12960), .A4(n12959), .ZN(
        n12967) );
  NOR4_X1 U16191 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12965) );
  NOR4_X1 U16192 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12964) );
  NOR4_X1 U16193 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12963) );
  NAND4_X1 U16194 ( .A1(n12965), .A2(n12964), .A3(n12963), .A4(n19611), .ZN(
        n12966) );
  NAND2_X1 U16195 ( .A1(n18891), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12971) );
  INV_X1 U16196 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12969) );
  OR2_X1 U16197 ( .A1(n18891), .A2(n12969), .ZN(n12970) );
  NAND2_X1 U16198 ( .A1(n12971), .A2(n12970), .ZN(n18894) );
  INV_X1 U16199 ( .A(n18894), .ZN(n12973) );
  INV_X1 U16200 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12972) );
  OAI22_X1 U16201 ( .A1(n14928), .A2(n12973), .B1(n18922), .B2(n12972), .ZN(
        n12974) );
  AOI21_X1 U16202 ( .B1(n13164), .B2(n18932), .A(n12974), .ZN(n12977) );
  AOI22_X1 U16203 ( .A1(n18884), .A2(BUF2_REG_30__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12976) );
  OAI21_X1 U16204 ( .B1(n14280), .B2(n18936), .A(n10003), .ZN(P2_U2889) );
  XNOR2_X1 U16205 ( .A(n14941), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13081) );
  NAND2_X1 U16206 ( .A1(n12979), .A2(n14937), .ZN(n12983) );
  NAND2_X1 U16207 ( .A1(n9764), .A2(n12981), .ZN(n12982) );
  NAND2_X1 U16208 ( .A1(n12985), .A2(n12984), .ZN(n12986) );
  NAND2_X1 U16209 ( .A1(n12987), .A2(n12986), .ZN(n14277) );
  NOR2_X1 U16210 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19669) );
  OR2_X1 U16211 ( .A1(n19681), .A2(n19669), .ZN(n19671) );
  NAND2_X1 U16212 ( .A1(n19671), .A2(n19729), .ZN(n12988) );
  AND2_X1 U16213 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19688) );
  NOR2_X1 U16214 ( .A1(n14277), .A2(n19057), .ZN(n12993) );
  NAND2_X1 U16215 ( .A1(n19668), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12989) );
  NAND2_X1 U16216 ( .A1(n12990), .A2(n12989), .ZN(n13236) );
  NAND2_X1 U16217 ( .A1(n13139), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13137) );
  NAND2_X1 U16218 ( .A1(n13138), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13135) );
  NAND2_X1 U16219 ( .A1(n13134), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13131) );
  NAND2_X1 U16220 ( .A1(n13121), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13120) );
  NAND2_X1 U16221 ( .A1(n13119), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13118) );
  OR2_X1 U16222 ( .A1(n13111), .A2(n14986), .ZN(n13109) );
  OR2_X1 U16223 ( .A1(n13109), .A2(n14965), .ZN(n13106) );
  NOR2_X1 U16224 ( .A1(n14942), .A2(n13105), .ZN(n13099) );
  AND2_X1 U16225 ( .A1(n13101), .A2(n13099), .ZN(n13149) );
  NAND2_X1 U16226 ( .A1(n15392), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U16227 ( .A1(n15105), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12991) );
  OAI211_X1 U16228 ( .C1(n15144), .C2(n15897), .A(n13074), .B(n12991), .ZN(
        n12992) );
  NOR2_X1 U16229 ( .A1(n12993), .A2(n12992), .ZN(n12994) );
  NAND3_X1 U16230 ( .A1(n12996), .A2(n12995), .A3(n12994), .ZN(P2_U2984) );
  INV_X1 U16231 ( .A(n12492), .ZN(n13001) );
  INV_X1 U16232 ( .A(n13015), .ZN(n13000) );
  NOR2_X1 U16233 ( .A1(n11266), .A2(n11253), .ZN(n13037) );
  NOR2_X1 U16234 ( .A1(n13037), .A2(n12997), .ZN(n12999) );
  AND2_X1 U16235 ( .A1(n12999), .A2(n12998), .ZN(n13031) );
  AOI21_X1 U16236 ( .B1(n13001), .B2(n13000), .A(n13031), .ZN(n13397) );
  INV_X1 U16237 ( .A(n15599), .ZN(n14304) );
  NAND2_X1 U16238 ( .A1(n19979), .A2(n14304), .ZN(n13002) );
  NAND2_X1 U16239 ( .A1(n13002), .A2(n20647), .ZN(n13003) );
  OR2_X1 U16240 ( .A1(n14297), .A2(n13003), .ZN(n13008) );
  OAI211_X1 U16241 ( .C1(n9621), .C2(n13005), .A(n12501), .B(n13004), .ZN(
        n13006) );
  NAND2_X1 U16242 ( .A1(n13006), .A2(n14301), .ZN(n13007) );
  MUX2_X1 U16243 ( .A(n13008), .B(n13007), .S(n9599), .Z(n13011) );
  INV_X1 U16244 ( .A(n13037), .ZN(n13009) );
  OR2_X1 U16245 ( .A1(n14301), .A2(n13009), .ZN(n13010) );
  NAND3_X1 U16246 ( .A1(n13397), .A2(n13011), .A3(n13010), .ZN(n13012) );
  INV_X1 U16247 ( .A(n13013), .ZN(n13016) );
  OR2_X1 U16248 ( .A1(n11245), .A2(n14302), .ZN(n13014) );
  NAND2_X1 U16249 ( .A1(n13015), .A2(n13014), .ZN(n14296) );
  OAI211_X1 U16250 ( .C1(n11243), .C2(n13019), .A(n13016), .B(n14296), .ZN(
        n13017) );
  OR2_X1 U16251 ( .A1(n9621), .A2(n13251), .ZN(n15580) );
  OAI21_X1 U16252 ( .B1(n13019), .B2(n11180), .A(n15580), .ZN(n13020) );
  NOR2_X1 U16253 ( .A1(n14419), .A2(n19945), .ZN(n13070) );
  INV_X1 U16254 ( .A(n20820), .ZN(n13033) );
  NAND2_X1 U16255 ( .A1(n13023), .A2(n12589), .ZN(n13029) );
  INV_X1 U16256 ( .A(n13398), .ZN(n13864) );
  NAND2_X1 U16257 ( .A1(n11244), .A2(n13864), .ZN(n13028) );
  INV_X1 U16258 ( .A(n11340), .ZN(n13024) );
  NAND2_X1 U16259 ( .A1(n13024), .A2(n13413), .ZN(n13027) );
  OAI21_X1 U16260 ( .B1(n9599), .B2(n11270), .A(n11254), .ZN(n13025) );
  OAI21_X1 U16261 ( .B1(n13025), .B2(n11258), .A(n19979), .ZN(n13026) );
  NAND4_X1 U16262 ( .A1(n13029), .A2(n13028), .A3(n13027), .A4(n13026), .ZN(
        n13030) );
  NOR2_X1 U16263 ( .A1(n13031), .A2(n13030), .ZN(n13032) );
  NAND2_X1 U16264 ( .A1(n13033), .A2(n13032), .ZN(n13388) );
  OAI21_X1 U16265 ( .B1(n13385), .B2(n12501), .A(n13034), .ZN(n13035) );
  OR2_X1 U16266 ( .A1(n13388), .A2(n13035), .ZN(n13036) );
  INV_X1 U16267 ( .A(n14763), .ZN(n14737) );
  NAND2_X1 U16268 ( .A1(n13038), .A2(n13037), .ZN(n14295) );
  INV_X1 U16269 ( .A(n14295), .ZN(n13039) );
  AND2_X1 U16270 ( .A1(n13864), .A2(n11245), .ZN(n13041) );
  INV_X1 U16271 ( .A(n15854), .ZN(n15790) );
  NOR2_X1 U16272 ( .A1(n19954), .A2(n19941), .ZN(n15849) );
  NAND2_X1 U16273 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19919) );
  NOR2_X1 U16274 ( .A1(n20699), .A2(n19919), .ZN(n13060) );
  NAND2_X1 U16275 ( .A1(n15849), .A2(n13060), .ZN(n14779) );
  INV_X1 U16276 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15862) );
  INV_X1 U16277 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15866) );
  NOR3_X1 U16278 ( .A1(n15862), .A2(n15866), .A3(n15855), .ZN(n15830) );
  NAND3_X1 U16279 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15830), .ZN(n14778) );
  NOR2_X1 U16280 ( .A1(n15738), .A2(n14778), .ZN(n14785) );
  NAND2_X1 U16281 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14785), .ZN(
        n14760) );
  NOR2_X1 U16282 ( .A1(n14779), .A2(n14760), .ZN(n15812) );
  AND4_X1 U16283 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14767) );
  AND3_X1 U16284 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n14767), .ZN(n14738) );
  NAND2_X1 U16285 ( .A1(n15812), .A2(n14738), .ZN(n14739) );
  NAND2_X1 U16286 ( .A1(n19940), .A2(n14739), .ZN(n13046) );
  INV_X1 U16287 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19937) );
  NAND2_X1 U16288 ( .A1(n14763), .A2(n19937), .ZN(n13043) );
  NOR2_X1 U16289 ( .A1(n13042), .A2(n12105), .ZN(n13434) );
  INV_X1 U16290 ( .A(n13434), .ZN(n14764) );
  OAI21_X1 U16291 ( .B1(n19937), .B2(n19941), .A(n19954), .ZN(n13058) );
  NAND2_X1 U16292 ( .A1(n13060), .A2(n13058), .ZN(n15847) );
  NOR2_X1 U16293 ( .A1(n14760), .A2(n15847), .ZN(n14766) );
  AND2_X1 U16294 ( .A1(n14766), .A2(n14738), .ZN(n13044) );
  OR2_X1 U16295 ( .A1(n19936), .A2(n13044), .ZN(n13045) );
  AND3_X1 U16296 ( .A1(n13046), .A2(n15848), .A3(n13045), .ZN(n14749) );
  AND2_X1 U16297 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U16298 ( .A1(n14749), .A2(n14740), .ZN(n13048) );
  OR2_X1 U16299 ( .A1(n15854), .A2(n19938), .ZN(n13047) );
  NAND2_X1 U16300 ( .A1(n13048), .A2(n13047), .ZN(n15762) );
  NAND2_X1 U16301 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15767) );
  NAND2_X1 U16302 ( .A1(n15854), .A2(n15767), .ZN(n13049) );
  NAND2_X1 U16303 ( .A1(n15762), .A2(n13049), .ZN(n14728) );
  NOR2_X1 U16304 ( .A1(n19936), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13050) );
  OR2_X1 U16305 ( .A1(n14728), .A2(n13050), .ZN(n14718) );
  AOI22_X1 U16306 ( .A1(n13059), .A2(n14698), .B1(n14763), .B2(n11535), .ZN(
        n13051) );
  OAI21_X1 U16307 ( .B1(n13436), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n13051), .ZN(n13052) );
  INV_X1 U16308 ( .A(n14711), .ZN(n13056) );
  INV_X1 U16309 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13424) );
  INV_X1 U16310 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14662) );
  NAND2_X1 U16311 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13053) );
  AND2_X1 U16312 ( .A1(n15854), .A2(n13053), .ZN(n13054) );
  NOR2_X1 U16313 ( .A1(n14711), .A2(n13054), .ZN(n14687) );
  INV_X1 U16314 ( .A(n13066), .ZN(n14679) );
  NAND2_X1 U16315 ( .A1(n15854), .A2(n14679), .ZN(n13055) );
  NAND2_X1 U16316 ( .A1(n14687), .A2(n13055), .ZN(n14670) );
  AOI211_X1 U16317 ( .C1(n9649), .C2(n15854), .A(n14662), .B(n14670), .ZN(
        n14661) );
  AOI211_X1 U16318 ( .C1(n15790), .C2(n13056), .A(n13424), .B(n14661), .ZN(
        n13069) );
  INV_X1 U16319 ( .A(n13057), .ZN(n13068) );
  INV_X1 U16320 ( .A(n13058), .ZN(n19950) );
  NAND2_X1 U16321 ( .A1(n15849), .A2(n19935), .ZN(n15853) );
  INV_X1 U16322 ( .A(n14760), .ZN(n13062) );
  AND4_X1 U16323 ( .A1(n14738), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n14740), .ZN(n13061) );
  NAND2_X1 U16324 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  NOR2_X1 U16325 ( .A1(n14698), .A2(n13064), .ZN(n13065) );
  AND2_X1 U16326 ( .A1(n14734), .A2(n13065), .ZN(n14691) );
  AND2_X1 U16327 ( .A1(n14691), .A2(n13066), .ZN(n14671) );
  NAND2_X1 U16328 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n14671), .ZN(
        n14663) );
  NOR3_X1 U16329 ( .A1(n14662), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14663), .ZN(n13067) );
  NOR4_X2 U16330 ( .A1(n13070), .A2(n13069), .A3(n13068), .A4(n13067), .ZN(
        n13071) );
  NAND2_X1 U16331 ( .A1(n13164), .A2(n15354), .ZN(n13079) );
  NOR2_X1 U16332 ( .A1(n13072), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13077) );
  INV_X1 U16333 ( .A(n13073), .ZN(n13075) );
  NOR2_X1 U16334 ( .A1(n13077), .A2(n13076), .ZN(n13078) );
  OAI21_X1 U16335 ( .B1(n14277), .B2(n16008), .A(n9992), .ZN(n13080) );
  OR2_X1 U16336 ( .A1(n13081), .A2(n16040), .ZN(n13084) );
  NAND2_X1 U16337 ( .A1(n13082), .A2(n16044), .ZN(n13083) );
  NAND3_X1 U16338 ( .A1(n13085), .A2(n13084), .A3(n13083), .ZN(P2_U3016) );
  INV_X1 U16339 ( .A(n13087), .ZN(n13088) );
  NAND3_X1 U16340 ( .A1(n13089), .A2(n13410), .A3(n13088), .ZN(n13090) );
  NAND2_X1 U16341 ( .A1(n14521), .A2(n19847), .ZN(n13098) );
  INV_X1 U16342 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14246) );
  INV_X1 U16343 ( .A(n13096), .ZN(n13097) );
  AND2_X1 U16344 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n13099), .ZN(
        n13100) );
  INV_X1 U16345 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13102) );
  NOR2_X1 U16346 ( .A1(n13104), .A2(n13105), .ZN(n13147) );
  NOR2_X1 U16347 ( .A1(n13104), .A2(n13106), .ZN(n13110) );
  NOR2_X1 U16348 ( .A1(n13110), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13107) );
  OR2_X1 U16349 ( .A1(n13147), .A2(n13107), .ZN(n14958) );
  INV_X1 U16350 ( .A(n14958), .ZN(n15915) );
  OR2_X1 U16351 ( .A1(n13104), .A2(n13109), .ZN(n13113) );
  AOI21_X1 U16352 ( .B1(n14965), .B2(n13113), .A(n13110), .ZN(n14967) );
  OR2_X1 U16353 ( .A1(n13104), .A2(n14986), .ZN(n13114) );
  NAND2_X1 U16354 ( .A1(n13114), .A2(n13111), .ZN(n13112) );
  NAND2_X1 U16355 ( .A1(n13113), .A2(n13112), .ZN(n14976) );
  INV_X1 U16356 ( .A(n14976), .ZN(n15924) );
  INV_X1 U16357 ( .A(n13114), .ZN(n13115) );
  AOI21_X1 U16358 ( .B1(n14986), .B2(n13104), .A(n13115), .ZN(n15938) );
  OR2_X1 U16359 ( .A1(n13116), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13117) );
  NAND2_X1 U16360 ( .A1(n13104), .A2(n13117), .ZN(n14996) );
  INV_X1 U16361 ( .A(n14996), .ZN(n15946) );
  AOI21_X1 U16362 ( .B1(n15004), .B2(n13118), .A(n13116), .ZN(n15006) );
  OAI21_X1 U16363 ( .B1(n13119), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n13118), .ZN(n15017) );
  INV_X1 U16364 ( .A(n15017), .ZN(n15541) );
  AOI21_X1 U16365 ( .B1(n13120), .B2(n18659), .A(n13119), .ZN(n18656) );
  OAI21_X1 U16366 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13121), .A(
        n13120), .ZN(n15044) );
  INV_X1 U16367 ( .A(n15044), .ZN(n18670) );
  AND2_X1 U16368 ( .A1(n13122), .A2(n13123), .ZN(n13124) );
  OR2_X1 U16369 ( .A1(n13121), .A2(n13124), .ZN(n15055) );
  INV_X1 U16370 ( .A(n15055), .ZN(n18681) );
  AOI21_X1 U16371 ( .B1(n13126), .B2(n13125), .A(n9703), .ZN(n18712) );
  NOR2_X1 U16372 ( .A1(n13128), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13129) );
  OR2_X1 U16373 ( .A1(n13127), .A2(n13129), .ZN(n18735) );
  INV_X1 U16374 ( .A(n18735), .ZN(n13142) );
  AOI21_X1 U16375 ( .B1(n18753), .B2(n9658), .A(n13130), .ZN(n18757) );
  AOI21_X1 U16376 ( .B1(n18787), .B2(n13131), .A(n13132), .ZN(n18781) );
  AOI21_X1 U16377 ( .B1(n18799), .B2(n13133), .A(n13134), .ZN(n18804) );
  AOI21_X1 U16378 ( .B1(n18821), .B2(n13135), .A(n13136), .ZN(n18826) );
  AOI21_X1 U16379 ( .B1(n20762), .B2(n13137), .A(n13138), .ZN(n19048) );
  AOI21_X1 U16380 ( .B1(n13638), .B2(n13530), .A(n13139), .ZN(n14195) );
  AOI22_X1 U16381 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13638), .B2(n19729), .ZN(
        n13643) );
  NAND2_X1 U16382 ( .A1(n18878), .A2(n13643), .ZN(n13642) );
  NOR2_X1 U16383 ( .A1(n14195), .A2(n13642), .ZN(n13617) );
  OAI21_X1 U16384 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13139), .A(
        n13137), .ZN(n13764) );
  NAND2_X1 U16385 ( .A1(n13617), .A2(n13764), .ZN(n18853) );
  NOR2_X1 U16386 ( .A1(n19048), .A2(n18853), .ZN(n18833) );
  OAI21_X1 U16387 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13138), .A(
        n13135), .ZN(n18834) );
  NAND2_X1 U16388 ( .A1(n18833), .A2(n18834), .ZN(n18824) );
  OAI21_X1 U16389 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13136), .A(
        n13133), .ZN(n18812) );
  NAND2_X1 U16390 ( .A1(n18809), .A2(n18812), .ZN(n18802) );
  NOR2_X1 U16391 ( .A1(n18804), .A2(n18802), .ZN(n18788) );
  OAI21_X1 U16392 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n13134), .A(
        n13131), .ZN(n18790) );
  NAND2_X1 U16393 ( .A1(n18788), .A2(n18790), .ZN(n18779) );
  OAI21_X1 U16394 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13132), .A(
        n9658), .ZN(n18775) );
  NAND2_X1 U16395 ( .A1(n18772), .A2(n18775), .ZN(n18770) );
  NOR2_X1 U16396 ( .A1(n18757), .A2(n18770), .ZN(n18744) );
  INV_X1 U16397 ( .A(n13130), .ZN(n13140) );
  AOI21_X1 U16398 ( .B1(n18742), .B2(n13140), .A(n13128), .ZN(n18746) );
  INV_X1 U16399 ( .A(n18746), .ZN(n13141) );
  NAND2_X1 U16400 ( .A1(n18744), .A2(n13141), .ZN(n18733) );
  OR2_X1 U16401 ( .A1(n13127), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13143) );
  NAND2_X1 U16402 ( .A1(n13143), .A2(n13125), .ZN(n18722) );
  NAND2_X1 U16403 ( .A1(n18720), .A2(n18722), .ZN(n18710) );
  NOR2_X1 U16404 ( .A1(n18712), .A2(n18710), .ZN(n18706) );
  XNOR2_X1 U16405 ( .A(n9703), .B(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18705) );
  NAND2_X1 U16406 ( .A1(n9703), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13145) );
  NAND2_X1 U16407 ( .A1(n13145), .A2(n13144), .ZN(n13146) );
  NAND2_X1 U16408 ( .A1(n13146), .A2(n13122), .ZN(n15067) );
  INV_X1 U16409 ( .A(n15067), .ZN(n18691) );
  NOR2_X1 U16410 ( .A1(n18681), .A2(n18680), .ZN(n18679) );
  NOR2_X1 U16411 ( .A1(n15541), .A2(n15540), .ZN(n15539) );
  NOR2_X1 U16412 ( .A1(n18810), .A2(n15539), .ZN(n13191) );
  NOR2_X1 U16413 ( .A1(n15006), .A2(n13191), .ZN(n13190) );
  NOR2_X1 U16414 ( .A1(n15924), .A2(n15923), .ZN(n15922) );
  NOR2_X1 U16415 ( .A1(n18810), .A2(n15922), .ZN(n13207) );
  NOR2_X1 U16416 ( .A1(n14967), .A2(n13207), .ZN(n13206) );
  NOR2_X1 U16417 ( .A1(n18810), .A2(n13206), .ZN(n15916) );
  NOR2_X1 U16418 ( .A1(n15915), .A2(n15916), .ZN(n15914) );
  NOR2_X1 U16419 ( .A1(n13147), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13148) );
  NOR2_X1 U16420 ( .A1(n13149), .A2(n13148), .ZN(n15901) );
  NOR2_X1 U16421 ( .A1(n15902), .A2(n15901), .ZN(n15900) );
  NAND4_X1 U16422 ( .A1(n19729), .A2(n19504), .A3(n19668), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19582) );
  NAND2_X1 U16423 ( .A1(n19668), .A2(n16063), .ZN(n13156) );
  INV_X1 U16424 ( .A(n13156), .ZN(n13150) );
  AND2_X1 U16425 ( .A1(n13151), .A2(n13150), .ZN(n16050) );
  NOR3_X1 U16426 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13152), .A3(n19697), 
        .ZN(n16100) );
  OR2_X1 U16427 ( .A1(n15392), .A2(n16100), .ZN(n13153) );
  NAND3_X1 U16428 ( .A1(n9865), .A2(n13221), .A3(n13154), .ZN(n13222) );
  INV_X1 U16429 ( .A(n19586), .ZN(n19722) );
  OAI21_X1 U16430 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19722), .A(
        P2_EBX_REG_31__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U16431 ( .A1(n19043), .A2(n13156), .ZN(n15893) );
  INV_X1 U16432 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15894) );
  OR2_X1 U16433 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19722), .ZN(n13165) );
  NAND2_X1 U16434 ( .A1(n15894), .A2(n13165), .ZN(n13157) );
  OR2_X1 U16435 ( .A1(n13222), .A2(n13157), .ZN(n13158) );
  NAND2_X2 U16436 ( .A1(n15893), .A2(n13158), .ZN(n18861) );
  AOI22_X1 U16437 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18861), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18862), .ZN(n13159) );
  OAI21_X1 U16438 ( .B1(n13160), .B2(n18865), .A(n13159), .ZN(n13161) );
  AOI21_X1 U16439 ( .B1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18842), .A(
        n13161), .ZN(n13162) );
  AOI21_X1 U16440 ( .B1(n18859), .B2(n13164), .A(n13163), .ZN(n13167) );
  NOR2_X2 U16441 ( .A1(n13255), .A2(n13165), .ZN(n18868) );
  INV_X1 U16442 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20636) );
  NOR3_X1 U16443 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20636), .ZN(n13170) );
  NOR4_X1 U16444 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13169) );
  NAND4_X1 U16445 ( .A1(n19957), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13170), .A4(
        n13169), .ZN(U214) );
  INV_X1 U16446 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19705) );
  NOR2_X1 U16447 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n19705), .ZN(n13172) );
  NOR4_X1 U16448 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13171) );
  INV_X1 U16449 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19660) );
  NAND4_X1 U16450 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13172), .A3(n13171), .A4(
        n19660), .ZN(n13173) );
  NOR2_X1 U16451 ( .A1(n18891), .A2(n13173), .ZN(n16172) );
  NAND2_X1 U16452 ( .A1(n16172), .A2(U214), .ZN(U212) );
  INV_X1 U16453 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17377) );
  NAND2_X1 U16454 ( .A1(n13174), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17404) );
  NOR2_X1 U16455 ( .A1(n13175), .A2(n17404), .ZN(n16464) );
  NAND2_X1 U16456 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16464), .ZN(
        n17365) );
  NOR2_X1 U16457 ( .A1(n17377), .A2(n17365), .ZN(n16447) );
  NAND2_X1 U16458 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16447), .ZN(
        n17323) );
  AOI22_X1 U16459 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17325), .B1(
        n17350), .B2(n17323), .ZN(n17352) );
  INV_X1 U16460 ( .A(n17323), .ZN(n13176) );
  INV_X1 U16461 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16658) );
  INV_X1 U16462 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17415) );
  NOR2_X1 U16463 ( .A1(n17415), .A2(n17404), .ZN(n16477) );
  AND2_X1 U16464 ( .A1(n16658), .A2(n16477), .ZN(n16466) );
  AOI211_X1 U16465 ( .C1(n17352), .C2(n13177), .A(n16302), .B(n18460), .ZN(
        n13189) );
  NOR3_X1 U16466 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16638) );
  NAND2_X1 U16467 ( .A1(n16638), .A2(n16968), .ZN(n16631) );
  NOR2_X1 U16468 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16631), .ZN(n16611) );
  INV_X1 U16469 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16955) );
  NAND2_X1 U16470 ( .A1(n16611), .A2(n16955), .ZN(n16603) );
  NAND2_X1 U16471 ( .A1(n16588), .A2(n16581), .ZN(n16579) );
  INV_X1 U16472 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16851) );
  NAND2_X1 U16473 ( .A1(n16560), .A2(n16851), .ZN(n16539) );
  NAND2_X1 U16474 ( .A1(n16538), .A2(n16534), .ZN(n16533) );
  INV_X1 U16475 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16505) );
  NAND2_X1 U16476 ( .A1(n16515), .A2(n16505), .ZN(n16504) );
  NAND2_X1 U16477 ( .A1(n16489), .A2(n16483), .ZN(n16481) );
  INV_X1 U16478 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16797) );
  NAND2_X1 U16479 ( .A1(n16469), .A2(n16797), .ZN(n16460) );
  INV_X1 U16480 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16770) );
  NAND2_X1 U16481 ( .A1(n16445), .A2(n16770), .ZN(n16436) );
  NAND2_X1 U16482 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18599) );
  INV_X1 U16483 ( .A(n18599), .ZN(n18606) );
  INV_X1 U16484 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n13181) );
  NOR2_X1 U16485 ( .A1(n13181), .A2(n17960), .ZN(n13179) );
  OAI211_X2 U16486 ( .C1(n18606), .C2(P3_STATEBS16_REG_SCAN_IN), .A(n13182), 
        .B(n13179), .ZN(n16665) );
  AOI211_X1 U16487 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16436), .A(n16431), .B(
        n16665), .ZN(n13188) );
  NAND2_X1 U16488 ( .A1(n18617), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18323) );
  OR2_X1 U16489 ( .A1(n18455), .A2(n18323), .ZN(n18450) );
  INV_X2 U16490 ( .A(n18615), .ZN(n18543) );
  NAND2_X2 U16491 ( .A1(n18543), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18541) );
  NOR2_X1 U16492 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16274) );
  INV_X1 U16493 ( .A(n16274), .ZN(n18466) );
  NAND3_X1 U16494 ( .A1(n18480), .A2(n18541), .A3(n18466), .ZN(n18472) );
  OAI211_X1 U16495 ( .C1(n18605), .C2(n18604), .A(n18599), .B(n16275), .ZN(
        n18445) );
  OAI211_X2 U16496 ( .C1(n13181), .C2(n17960), .A(n18445), .B(n13182), .ZN(
        n16666) );
  INV_X1 U16497 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n15409) );
  OAI22_X1 U16498 ( .A1(n17350), .A2(n16656), .B1(n16666), .B2(n15409), .ZN(
        n13187) );
  INV_X1 U16499 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18514) );
  NAND2_X1 U16500 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16473) );
  NOR2_X1 U16501 ( .A1(n18514), .A2(n16473), .ZN(n16440) );
  NAND3_X1 U16502 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16440), .ZN(n13184) );
  INV_X1 U16503 ( .A(n18445), .ZN(n13183) );
  INV_X1 U16504 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18491) );
  INV_X1 U16505 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18488) );
  NAND3_X1 U16506 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16624) );
  NOR3_X1 U16507 ( .A1(n18491), .A2(n18488), .A3(n16624), .ZN(n16574) );
  NAND4_X1 U16508 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16574), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n16500) );
  NAND3_X1 U16509 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_9__SCAN_IN), .ZN(n16501) );
  NOR2_X1 U16510 ( .A1(n16500), .A2(n16501), .ZN(n16516) );
  NAND2_X1 U16511 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16516), .ZN(n16508) );
  NOR2_X1 U16512 ( .A1(n18506), .A2(n16508), .ZN(n16491) );
  NAND3_X1 U16513 ( .A1(n16648), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n16491), 
        .ZN(n16487) );
  NOR2_X1 U16514 ( .A1(n13184), .A2(n16487), .ZN(n13185) );
  INV_X1 U16515 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18521) );
  NAND2_X1 U16516 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16491), .ZN(n16490) );
  NOR3_X1 U16517 ( .A1(n18521), .A2(n16490), .A3(n13184), .ZN(n16426) );
  OAI21_X1 U16518 ( .B1(n16426), .B2(n16659), .A(n16669), .ZN(n16422) );
  MUX2_X1 U16519 ( .A(n13185), .B(n16422), .S(P3_REIP_REG_20__SCAN_IN), .Z(
        n13186) );
  AOI211_X1 U16520 ( .C1(n15006), .C2(n13191), .A(n13190), .B(n19582), .ZN(
        n13205) );
  AOI22_X1 U16521 ( .A1(n18861), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18862), .ZN(n13192) );
  INV_X1 U16522 ( .A(n13192), .ZN(n13204) );
  OAI22_X1 U16523 ( .A1(n15004), .A2(n18871), .B1(n13193), .B2(n18865), .ZN(
        n13203) );
  OR2_X1 U16524 ( .A1(n13195), .A2(n13196), .ZN(n13197) );
  NAND2_X1 U16525 ( .A1(n13194), .A2(n13197), .ZN(n15218) );
  OR2_X1 U16526 ( .A1(n13199), .A2(n13200), .ZN(n13201) );
  NAND2_X1 U16527 ( .A1(n13198), .A2(n13201), .ZN(n15224) );
  OAI22_X1 U16528 ( .A1(n15218), .A2(n18858), .B1(n15224), .B2(n18841), .ZN(
        n13202) );
  AOI211_X1 U16529 ( .C1(n14967), .C2(n13207), .A(n13206), .B(n19582), .ZN(
        n13220) );
  OAI22_X1 U16530 ( .A1(n19651), .A2(n18845), .B1(n13208), .B2(n18865), .ZN(
        n13219) );
  AOI22_X1 U16531 ( .A1(n18861), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18842), .ZN(n13209) );
  INV_X1 U16532 ( .A(n13209), .ZN(n13218) );
  NOR2_X1 U16533 ( .A1(n14827), .A2(n13211), .ZN(n13212) );
  OR2_X1 U16534 ( .A1(n13214), .A2(n13215), .ZN(n13216) );
  NAND2_X1 U16535 ( .A1(n13213), .A2(n13216), .ZN(n15177) );
  OAI22_X1 U16536 ( .A1(n15172), .A2(n18858), .B1(n15177), .B2(n18841), .ZN(
        n13217) );
  OR4_X1 U16537 ( .A1(n13220), .A2(n13219), .A3(n13218), .A4(n13217), .ZN(
        P2_U2828) );
  INV_X1 U16538 ( .A(n10640), .ZN(n18941) );
  NAND3_X1 U16539 ( .A1(n18941), .A2(n19720), .A3(n13221), .ZN(n18851) );
  INV_X1 U16540 ( .A(n18851), .ZN(n18872) );
  INV_X1 U16541 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13224) );
  INV_X1 U16542 ( .A(n19681), .ZN(n19454) );
  NOR2_X1 U16543 ( .A1(n19454), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13225) );
  INV_X1 U16544 ( .A(n13225), .ZN(n13223) );
  OAI211_X1 U16545 ( .C1(n18872), .C2(n13224), .A(n13223), .B(n13222), .ZN(
        P2_U2814) );
  INV_X1 U16546 ( .A(n11054), .ZN(n13228) );
  INV_X1 U16547 ( .A(n19724), .ZN(n13227) );
  OAI21_X1 U16548 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n13225), .A(n13227), 
        .ZN(n13226) );
  OAI21_X1 U16549 ( .B1(n13228), .B2(n13227), .A(n13226), .ZN(P2_U3612) );
  INV_X1 U16550 ( .A(n18866), .ZN(n13229) );
  NOR2_X1 U16551 ( .A1(n13229), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13230) );
  NOR2_X1 U16552 ( .A1(n13231), .A2(n13230), .ZN(n13342) );
  NAND2_X1 U16553 ( .A1(n15127), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13337) );
  INV_X1 U16554 ( .A(n13337), .ZN(n13235) );
  OAI21_X1 U16555 ( .B1(n13233), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13232), .ZN(n13338) );
  NOR2_X1 U16556 ( .A1(n15996), .A2(n13338), .ZN(n13234) );
  AOI211_X1 U16557 ( .C1(n13342), .C2(n19050), .A(n13235), .B(n13234), .ZN(
        n13238) );
  OAI21_X1 U16558 ( .B1(n15105), .B2(n13236), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13237) );
  OAI211_X1 U16559 ( .C1(n19057), .C2(n15399), .A(n13238), .B(n13237), .ZN(
        P2_U3014) );
  OAI21_X1 U16560 ( .B1(n13637), .B2(n13240), .A(n13239), .ZN(n13241) );
  XOR2_X1 U16561 ( .A(n13241), .B(n13713), .Z(n13315) );
  OAI21_X1 U16562 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13243), .A(
        n13242), .ZN(n13312) );
  NAND2_X1 U16563 ( .A1(n15127), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13305) );
  OAI21_X1 U16564 ( .B1(n15996), .B2(n13312), .A(n13305), .ZN(n13245) );
  MUX2_X1 U16565 ( .A(n19049), .B(n15105), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13244) );
  AOI211_X1 U16566 ( .C1(n19050), .C2(n13315), .A(n13245), .B(n13244), .ZN(
        n13246) );
  OAI21_X1 U16567 ( .B1(n10212), .B2(n19057), .A(n13246), .ZN(P2_U3013) );
  INV_X1 U16568 ( .A(n20645), .ZN(n13248) );
  NAND2_X1 U16569 ( .A1(n20418), .A2(n20553), .ZN(n19743) );
  INV_X1 U16570 ( .A(n19743), .ZN(n13980) );
  OAI21_X1 U16571 ( .B1(n13980), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13248), 
        .ZN(n13247) );
  OAI21_X1 U16572 ( .B1(n13249), .B2(n13248), .A(n13247), .ZN(P1_U3487) );
  AND2_X1 U16573 ( .A1(n13251), .A2(n13250), .ZN(n13252) );
  NAND2_X1 U16574 ( .A1(n13317), .A2(n11253), .ZN(n13364) );
  INV_X1 U16575 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14130) );
  NAND2_X1 U16576 ( .A1(n13317), .A2(n19979), .ZN(n13318) );
  INV_X1 U16577 ( .A(DATAI_15_), .ZN(n13254) );
  INV_X1 U16578 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13253) );
  MUX2_X1 U16579 ( .A(n13254), .B(n13253), .S(n19957), .Z(n14131) );
  INV_X1 U16580 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20791) );
  OAI222_X1 U16581 ( .A1(n13364), .A2(n14130), .B1(n13318), .B2(n14131), .C1(
        n13317), .C2(n20791), .ZN(P1_U2967) );
  INV_X1 U16582 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20697) );
  INV_X1 U16583 ( .A(n13255), .ZN(n13256) );
  NOR2_X2 U16584 ( .A1(n13271), .A2(n19043), .ZN(n19016) );
  NAND2_X1 U16585 ( .A1(n19016), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13259) );
  NAND2_X1 U16586 ( .A1(n18891), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13258) );
  INV_X1 U16587 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16210) );
  OR2_X1 U16588 ( .A1(n18891), .A2(n16210), .ZN(n13257) );
  NAND2_X1 U16589 ( .A1(n13258), .A2(n13257), .ZN(n18902) );
  NAND2_X1 U16590 ( .A1(n13271), .A2(n18902), .ZN(n13349) );
  OAI211_X1 U16591 ( .C1(n20697), .C2(n18943), .A(n13259), .B(n13349), .ZN(
        P2_U2977) );
  INV_X1 U16592 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n18993) );
  NAND2_X1 U16593 ( .A1(n19016), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13262) );
  NAND2_X1 U16594 ( .A1(n18891), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13261) );
  INV_X1 U16595 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16214) );
  OR2_X1 U16596 ( .A1(n18891), .A2(n16214), .ZN(n13260) );
  NAND2_X1 U16597 ( .A1(n13261), .A2(n13260), .ZN(n18908) );
  NAND2_X1 U16598 ( .A1(n13271), .A2(n18908), .ZN(n13347) );
  OAI211_X1 U16599 ( .C1(n18993), .C2(n18943), .A(n13262), .B(n13347), .ZN(
        P2_U2975) );
  INV_X1 U16600 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18982) );
  NAND2_X1 U16601 ( .A1(n19016), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13263) );
  NAND2_X1 U16602 ( .A1(n13271), .A2(n18894), .ZN(n13267) );
  OAI211_X1 U16603 ( .C1(n18982), .C2(n18943), .A(n13263), .B(n13267), .ZN(
        P2_U2981) );
  INV_X1 U16604 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18991) );
  NAND2_X1 U16605 ( .A1(n19016), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13266) );
  NAND2_X1 U16606 ( .A1(n18891), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13265) );
  INV_X1 U16607 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16212) );
  OR2_X1 U16608 ( .A1(n18891), .A2(n16212), .ZN(n13264) );
  NAND2_X1 U16609 ( .A1(n13265), .A2(n13264), .ZN(n18905) );
  NAND2_X1 U16610 ( .A1(n13271), .A2(n18905), .ZN(n13351) );
  OAI211_X1 U16611 ( .C1(n18991), .C2(n18943), .A(n13266), .B(n13351), .ZN(
        P2_U2976) );
  NAND2_X1 U16612 ( .A1(n19016), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13268) );
  OAI211_X1 U16613 ( .C1(n12972), .C2(n18943), .A(n13268), .B(n13267), .ZN(
        P2_U2966) );
  INV_X1 U16614 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18985) );
  NAND2_X1 U16615 ( .A1(n19016), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U16616 ( .A1(n18891), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13270) );
  INV_X1 U16617 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16207) );
  OR2_X1 U16618 ( .A1(n18891), .A2(n16207), .ZN(n13269) );
  NAND2_X1 U16619 ( .A1(n13270), .A2(n13269), .ZN(n18898) );
  NAND2_X1 U16620 ( .A1(n13271), .A2(n18898), .ZN(n13273) );
  OAI211_X1 U16621 ( .C1(n18985), .C2(n18943), .A(n13272), .B(n13273), .ZN(
        P2_U2979) );
  INV_X1 U16622 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n18952) );
  NAND2_X1 U16623 ( .A1(n19016), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13274) );
  OAI211_X1 U16624 ( .C1(n18952), .C2(n18943), .A(n13274), .B(n13273), .ZN(
        P2_U2964) );
  INV_X1 U16625 ( .A(n13275), .ZN(n13276) );
  OAI22_X1 U16626 ( .A1(n18891), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n18892), .ZN(n19024) );
  OAI21_X1 U16627 ( .B1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B2(
        P2_STATE2_REG_3__SCAN_IN), .A(n10863), .ZN(n13277) );
  AOI21_X1 U16628 ( .B1(n13282), .B2(n13281), .A(n13280), .ZN(n18860) );
  INV_X1 U16629 ( .A(n18860), .ZN(n13339) );
  NOR2_X1 U16630 ( .A1(n19698), .A2(n13339), .ZN(n18935) );
  INV_X1 U16631 ( .A(n18935), .ZN(n13283) );
  OAI211_X1 U16632 ( .C1(n18873), .C2(n18860), .A(n13283), .B(n18890), .ZN(
        n13285) );
  AOI22_X1 U16633 ( .A1(n18932), .A2(n18860), .B1(n18931), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13284) );
  OAI211_X1 U16634 ( .C1(n18940), .C2(n19024), .A(n13285), .B(n13284), .ZN(
        P2_U2919) );
  XNOR2_X1 U16635 ( .A(n13286), .B(n13287), .ZN(n19692) );
  MUX2_X1 U16636 ( .A(n10171), .B(n10212), .S(n14840), .Z(n13288) );
  OAI21_X1 U16637 ( .B1(n19689), .B2(n14880), .A(n13288), .ZN(P2_U2886) );
  INV_X1 U16638 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13293) );
  INV_X1 U16639 ( .A(n15550), .ZN(n13289) );
  NAND2_X1 U16640 ( .A1(n13289), .A2(n15580), .ZN(n13291) );
  NAND2_X1 U16641 ( .A1(n14301), .A2(n15599), .ZN(n13394) );
  NOR2_X1 U16642 ( .A1(n19740), .A2(n13394), .ZN(n13290) );
  NAND2_X1 U16643 ( .A1(n19854), .A2(n12501), .ZN(n13486) );
  NAND2_X1 U16644 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15884) );
  NAND2_X1 U16645 ( .A1(n20790), .A2(n14789), .ZN(n19853) );
  NOR2_X4 U16646 ( .A1(n19854), .A2(n19873), .ZN(n19872) );
  AOI22_X1 U16647 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13292) );
  OAI21_X1 U16648 ( .B1(n13293), .B2(n13486), .A(n13292), .ZN(P1_U2909) );
  INV_X1 U16649 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U16650 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13294) );
  OAI21_X1 U16651 ( .B1(n13295), .B2(n13486), .A(n13294), .ZN(P1_U2908) );
  INV_X1 U16652 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U16653 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13296) );
  OAI21_X1 U16654 ( .B1(n13297), .B2(n13486), .A(n13296), .ZN(P1_U2907) );
  AOI22_X1 U16655 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13298) );
  OAI21_X1 U16656 ( .B1(n12089), .B2(n13486), .A(n13298), .ZN(P1_U2906) );
  INV_X1 U16657 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16658 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13299) );
  OAI21_X1 U16659 ( .B1(n13300), .B2(n13486), .A(n13299), .ZN(P1_U2912) );
  INV_X1 U16660 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13302) );
  AOI22_X1 U16661 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13301) );
  OAI21_X1 U16662 ( .B1(n13302), .B2(n13486), .A(n13301), .ZN(P1_U2911) );
  INV_X1 U16663 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13304) );
  AOI22_X1 U16664 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13303) );
  OAI21_X1 U16665 ( .B1(n13304), .B2(n13486), .A(n13303), .ZN(P1_U2910) );
  OAI21_X1 U16666 ( .B1(n13343), .B2(n13713), .A(n13305), .ZN(n13314) );
  OAI211_X1 U16667 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n13307), .B(n13306), .ZN(n13311) );
  XNOR2_X1 U16668 ( .A(n13309), .B(n13308), .ZN(n19694) );
  NAND2_X1 U16669 ( .A1(n15354), .A2(n19694), .ZN(n13310) );
  OAI211_X1 U16670 ( .C1(n13312), .C2(n16040), .A(n13311), .B(n13310), .ZN(
        n13313) );
  AOI211_X1 U16671 ( .C1(n16044), .C2(n13315), .A(n13314), .B(n13313), .ZN(
        n13316) );
  OAI21_X1 U16672 ( .B1(n10212), .B2(n16008), .A(n13316), .ZN(P2_U3045) );
  INV_X2 U16673 ( .A(n13317), .ZN(n19904) );
  AOI22_X1 U16674 ( .A1(n19905), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13321) );
  INV_X1 U16675 ( .A(DATAI_7_), .ZN(n13320) );
  NAND2_X1 U16676 ( .A1(n19957), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13319) );
  OAI21_X1 U16677 ( .B1(n19957), .B2(n13320), .A(n13319), .ZN(n14486) );
  NAND2_X1 U16678 ( .A1(n19890), .A2(n14486), .ZN(n13375) );
  NAND2_X1 U16679 ( .A1(n13321), .A2(n13375), .ZN(P1_U2959) );
  AOI22_X1 U16680 ( .A1(n19905), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U16681 ( .A1(n19959), .A2(DATAI_5_), .ZN(n13323) );
  NAND2_X1 U16682 ( .A1(n19957), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13322) );
  AND2_X1 U16683 ( .A1(n13323), .A2(n13322), .ZN(n19995) );
  INV_X1 U16684 ( .A(n19995), .ZN(n14494) );
  NAND2_X1 U16685 ( .A1(n19890), .A2(n14494), .ZN(n13370) );
  NAND2_X1 U16686 ( .A1(n13324), .A2(n13370), .ZN(P1_U2957) );
  AOI22_X1 U16687 ( .A1(n19905), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13327) );
  NAND2_X1 U16688 ( .A1(n19959), .A2(DATAI_4_), .ZN(n13326) );
  NAND2_X1 U16689 ( .A1(n19957), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13325) );
  AND2_X1 U16690 ( .A1(n13326), .A2(n13325), .ZN(n19991) );
  INV_X1 U16691 ( .A(n19991), .ZN(n14497) );
  NAND2_X1 U16692 ( .A1(n19890), .A2(n14497), .ZN(n13365) );
  NAND2_X1 U16693 ( .A1(n13327), .A2(n13365), .ZN(P1_U2956) );
  AOI22_X1 U16694 ( .A1(n19905), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U16695 ( .A1(n19959), .A2(DATAI_2_), .ZN(n13329) );
  NAND2_X1 U16696 ( .A1(n19957), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13328) );
  AND2_X1 U16697 ( .A1(n13329), .A2(n13328), .ZN(n19984) );
  INV_X1 U16698 ( .A(n19984), .ZN(n14503) );
  NAND2_X1 U16699 ( .A1(n19890), .A2(n14503), .ZN(n13373) );
  NAND2_X1 U16700 ( .A1(n13330), .A2(n13373), .ZN(P1_U2954) );
  AOI22_X1 U16701 ( .A1(n19905), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13333) );
  NAND2_X1 U16702 ( .A1(n19959), .A2(DATAI_6_), .ZN(n13332) );
  NAND2_X1 U16703 ( .A1(n19957), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13331) );
  INV_X1 U16704 ( .A(n19998), .ZN(n14490) );
  NAND2_X1 U16705 ( .A1(n19890), .A2(n14490), .ZN(n13377) );
  NAND2_X1 U16706 ( .A1(n13333), .A2(n13377), .ZN(P1_U2958) );
  AOI22_X1 U16707 ( .A1(n19905), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13336) );
  NAND2_X1 U16708 ( .A1(n19959), .A2(DATAI_3_), .ZN(n13335) );
  NAND2_X1 U16709 ( .A1(n19957), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13334) );
  AND2_X1 U16710 ( .A1(n13335), .A2(n13334), .ZN(n19988) );
  INV_X1 U16711 ( .A(n19988), .ZN(n14500) );
  NAND2_X1 U16712 ( .A1(n19890), .A2(n14500), .ZN(n13367) );
  NAND2_X1 U16713 ( .A1(n13336), .A2(n13367), .ZN(P1_U2955) );
  OAI21_X1 U16714 ( .B1(n16008), .B2(n15399), .A(n13337), .ZN(n13341) );
  OAI22_X1 U16715 ( .A1(n16036), .A2(n13339), .B1(n16040), .B2(n13338), .ZN(
        n13340) );
  AOI211_X1 U16716 ( .C1(n16044), .C2(n13342), .A(n13341), .B(n13340), .ZN(
        n13346) );
  MUX2_X1 U16717 ( .A(n13344), .B(n13343), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13345) );
  NAND2_X1 U16718 ( .A1(n13346), .A2(n13345), .ZN(P2_U3046) );
  INV_X1 U16719 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n18960) );
  NAND2_X1 U16720 ( .A1(n19044), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13348) );
  OAI211_X1 U16721 ( .C1(n18960), .C2(n18943), .A(n13348), .B(n13347), .ZN(
        P2_U2960) );
  INV_X1 U16722 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n18956) );
  NAND2_X1 U16723 ( .A1(n19044), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13350) );
  OAI211_X1 U16724 ( .C1(n18956), .C2(n18943), .A(n13350), .B(n13349), .ZN(
        P2_U2962) );
  INV_X1 U16725 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n18958) );
  NAND2_X1 U16726 ( .A1(n19044), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13352) );
  OAI211_X1 U16727 ( .C1(n18943), .C2(n18958), .A(n13352), .B(n13351), .ZN(
        P2_U2961) );
  INV_X1 U16728 ( .A(n13353), .ZN(n13356) );
  OAI21_X1 U16729 ( .B1(n13356), .B2(n13355), .A(n13354), .ZN(n13929) );
  NAND2_X1 U16730 ( .A1(n11266), .A2(n11254), .ZN(n13357) );
  NAND2_X1 U16731 ( .A1(n19959), .A2(DATAI_0_), .ZN(n13359) );
  NAND2_X1 U16732 ( .A1(n19957), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13358) );
  AND2_X1 U16733 ( .A1(n13359), .A2(n13358), .ZN(n19971) );
  INV_X1 U16734 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19876) );
  OAI222_X1 U16735 ( .A1(n13929), .A2(n14493), .B1(n14137), .B2(n19971), .C1(
        n14482), .C2(n19876), .ZN(P1_U2904) );
  OAI21_X1 U16736 ( .B1(n13361), .B2(n13360), .A(n13502), .ZN(n13885) );
  NAND2_X1 U16737 ( .A1(n19959), .A2(DATAI_1_), .ZN(n13363) );
  NAND2_X1 U16738 ( .A1(n19957), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13362) );
  AND2_X1 U16739 ( .A1(n13363), .A2(n13362), .ZN(n19980) );
  OAI222_X1 U16740 ( .A1(n13885), .A2(n14493), .B1(n14137), .B2(n19980), .C1(
        n14482), .C2(n11607), .ZN(P1_U2903) );
  INV_X2 U16741 ( .A(n13364), .ZN(n19905) );
  AOI22_X1 U16742 ( .A1(n19905), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13366) );
  NAND2_X1 U16743 ( .A1(n13366), .A2(n13365), .ZN(P1_U2941) );
  AOI22_X1 U16744 ( .A1(n19905), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13368) );
  NAND2_X1 U16745 ( .A1(n13368), .A2(n13367), .ZN(P1_U2940) );
  AOI22_X1 U16746 ( .A1(n19905), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13369) );
  INV_X1 U16747 ( .A(n19971), .ZN(n14157) );
  NAND2_X1 U16748 ( .A1(n19890), .A2(n14157), .ZN(n13379) );
  NAND2_X1 U16749 ( .A1(n13369), .A2(n13379), .ZN(P1_U2952) );
  AOI22_X1 U16750 ( .A1(n19905), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13371) );
  NAND2_X1 U16751 ( .A1(n13371), .A2(n13370), .ZN(P1_U2942) );
  AOI22_X1 U16752 ( .A1(n19905), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13372) );
  INV_X1 U16753 ( .A(n19980), .ZN(n14508) );
  NAND2_X1 U16754 ( .A1(n19890), .A2(n14508), .ZN(n13381) );
  NAND2_X1 U16755 ( .A1(n13372), .A2(n13381), .ZN(P1_U2938) );
  AOI22_X1 U16756 ( .A1(n19905), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13374) );
  NAND2_X1 U16757 ( .A1(n13374), .A2(n13373), .ZN(P1_U2939) );
  AOI22_X1 U16758 ( .A1(n19905), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13376) );
  NAND2_X1 U16759 ( .A1(n13376), .A2(n13375), .ZN(P1_U2944) );
  AOI22_X1 U16760 ( .A1(n19905), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U16761 ( .A1(n13378), .A2(n13377), .ZN(P1_U2943) );
  AOI22_X1 U16762 ( .A1(n19905), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13380) );
  NAND2_X1 U16763 ( .A1(n13380), .A2(n13379), .ZN(P1_U2937) );
  AOI22_X1 U16764 ( .A1(n19905), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13382) );
  NAND2_X1 U16765 ( .A1(n13382), .A2(n13381), .ZN(P1_U2953) );
  INV_X1 U16766 ( .A(n19171), .ZN(n19682) );
  MUX2_X1 U16767 ( .A(n10131), .B(n14217), .S(n14840), .Z(n13384) );
  OAI21_X1 U16768 ( .B1(n19682), .B2(n14880), .A(n13384), .ZN(P2_U2885) );
  AND3_X1 U16769 ( .A1(n13386), .A2(n13385), .A3(n9621), .ZN(n13387) );
  NAND2_X1 U16770 ( .A1(n12437), .A2(n13387), .ZN(n13389) );
  NOR2_X1 U16771 ( .A1(n13389), .A2(n13388), .ZN(n14794) );
  INV_X1 U16772 ( .A(n14794), .ZN(n13672) );
  NOR2_X1 U16773 ( .A1(n14796), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13390) );
  AOI21_X1 U16774 ( .B1(n11614), .B2(n13672), .A(n13390), .ZN(n15552) );
  INV_X1 U16775 ( .A(n15552), .ZN(n13392) );
  OAI22_X1 U16776 ( .A1(n20553), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20623), .ZN(n13391) );
  AOI21_X1 U16777 ( .B1(n13392), .B2(n14800), .A(n13391), .ZN(n13404) );
  INV_X1 U16778 ( .A(n9621), .ZN(n13395) );
  INV_X1 U16779 ( .A(n13394), .ZN(n15574) );
  OAI211_X1 U16780 ( .C1(n15550), .C2(n13395), .A(n15574), .B(n20647), .ZN(
        n13396) );
  OAI211_X1 U16781 ( .C1(n13398), .C2(n19983), .A(n13397), .B(n13396), .ZN(
        n13400) );
  NOR2_X1 U16782 ( .A1(n13400), .A2(n13399), .ZN(n13402) );
  INV_X1 U16783 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19747) );
  NAND2_X1 U16784 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14789), .ZN(n15888) );
  OAI22_X1 U16785 ( .A1(n13684), .A2(n19740), .B1(n19747), .B2(n15888), .ZN(
        n13406) );
  AOI21_X1 U16786 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20790), .A(n13406), 
        .ZN(n14808) );
  AOI21_X1 U16787 ( .B1(n15550), .B2(n14800), .A(n14808), .ZN(n13403) );
  OAI22_X1 U16788 ( .A1(n13404), .A2(n14808), .B1(n13403), .B2(n11263), .ZN(
        P1_U3474) );
  INV_X1 U16789 ( .A(n20113), .ZN(n20360) );
  XNOR2_X1 U16790 ( .A(n13405), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19831) );
  INV_X1 U16791 ( .A(n12437), .ZN(n13407) );
  NAND3_X1 U16792 ( .A1(n13407), .A2(n14800), .A3(n13406), .ZN(n13408) );
  INV_X1 U16793 ( .A(n14808), .ZN(n20627) );
  OAI22_X1 U16794 ( .A1(n19831), .A2(n13408), .B1(n13683), .B2(n20627), .ZN(
        P1_U3468) );
  OAI21_X1 U16795 ( .B1(n13411), .B2(n13410), .A(n13409), .ZN(n13877) );
  AOI22_X1 U16796 ( .A1(n19846), .A2(n13877), .B1(n14446), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13412) );
  OAI21_X1 U16797 ( .B1(n13885), .B2(n14463), .A(n13412), .ZN(P1_U2871) );
  OR2_X1 U16798 ( .A1(n13413), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13415) );
  AND2_X1 U16799 ( .A1(n13415), .A2(n13414), .ZN(n13925) );
  AOI22_X1 U16800 ( .A1(n19846), .A2(n13925), .B1(P1_EBX_REG_0__SCAN_IN), .B2(
        n14446), .ZN(n13416) );
  OAI21_X1 U16801 ( .B1(n13929), .B2(n14463), .A(n13416), .ZN(P1_U2872) );
  INV_X1 U16802 ( .A(n13418), .ZN(n14802) );
  NAND2_X1 U16803 ( .A1(n14802), .A2(n11358), .ZN(n13675) );
  NAND2_X1 U16804 ( .A1(n13418), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13670) );
  NAND2_X1 U16805 ( .A1(n13675), .A2(n13670), .ZN(n13425) );
  NOR2_X1 U16806 ( .A1(n13671), .A2(n13425), .ZN(n13420) );
  XNOR2_X1 U16807 ( .A(n11358), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13419) );
  AOI22_X1 U16808 ( .A1(n14794), .A2(n13420), .B1(n15550), .B2(n13419), .ZN(
        n13423) );
  NAND2_X1 U16809 ( .A1(n14295), .A2(n13421), .ZN(n13677) );
  NAND2_X1 U16810 ( .A1(n13677), .A2(n13425), .ZN(n13422) );
  OAI211_X1 U16811 ( .C1(n13417), .C2(n14794), .A(n13423), .B(n13422), .ZN(
        n13667) );
  AOI22_X1 U16812 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19941), .B2(n13424), .ZN(
        n14807) );
  NAND2_X1 U16813 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14806) );
  INV_X1 U16814 ( .A(n14806), .ZN(n13427) );
  INV_X1 U16815 ( .A(n20623), .ZN(n14801) );
  INV_X1 U16816 ( .A(n13425), .ZN(n13426) );
  AOI222_X1 U16817 ( .A1(n13667), .A2(n14800), .B1(n14807), .B2(n13427), .C1(
        n14801), .C2(n13426), .ZN(n13428) );
  MUX2_X1 U16818 ( .A(n13428), .B(n11358), .S(n14808), .Z(n13429) );
  INV_X1 U16819 ( .A(n13429), .ZN(P1_U3472) );
  MUX2_X1 U16820 ( .A(n15399), .B(n13430), .S(n14873), .Z(n13431) );
  OAI21_X1 U16821 ( .B1(n19698), .B2(n14880), .A(n13431), .ZN(P2_U2887) );
  OAI21_X1 U16822 ( .B1(n13432), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13433), .ZN(n13470) );
  INV_X1 U16823 ( .A(n13436), .ZN(n13435) );
  AOI21_X1 U16824 ( .B1(n19937), .B2(n13435), .A(n13434), .ZN(n13499) );
  AOI22_X1 U16825 ( .A1(n13499), .A2(n14761), .B1(n19937), .B2(n13436), .ZN(
        n13437) );
  INV_X1 U16826 ( .A(n13437), .ZN(n13439) );
  AND2_X1 U16827 ( .A1(n12105), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13473) );
  AOI21_X1 U16828 ( .B1(n19925), .B2(n13925), .A(n13473), .ZN(n13438) );
  OAI211_X1 U16829 ( .C1(n19946), .C2(n13470), .A(n13439), .B(n13438), .ZN(
        P1_U3031) );
  MUX2_X1 U16830 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n13444), .S(n14840), .Z(
        n13445) );
  AOI21_X1 U16831 ( .B1(n19678), .B2(n14870), .A(n13445), .ZN(n13446) );
  INV_X1 U16832 ( .A(n13446), .ZN(P2_U2884) );
  INV_X1 U16833 ( .A(n15398), .ZN(n13715) );
  NAND2_X1 U16834 ( .A1(n13444), .A2(n13715), .ZN(n13460) );
  NAND2_X1 U16835 ( .A1(n16060), .A2(n13447), .ZN(n13913) );
  INV_X1 U16836 ( .A(n13448), .ZN(n13449) );
  NAND2_X1 U16837 ( .A1(n13449), .A2(n16054), .ZN(n13914) );
  NAND2_X1 U16838 ( .A1(n13450), .A2(n10624), .ZN(n13451) );
  NAND2_X1 U16839 ( .A1(n13451), .A2(n12732), .ZN(n13452) );
  AOI21_X1 U16840 ( .B1(n13913), .B2(n13914), .A(n13452), .ZN(n13458) );
  INV_X1 U16841 ( .A(n10624), .ZN(n13453) );
  NAND2_X1 U16842 ( .A1(n13450), .A2(n13453), .ZN(n13919) );
  NAND2_X1 U16843 ( .A1(n13919), .A2(n13914), .ZN(n13456) );
  NAND2_X1 U16844 ( .A1(n13454), .A2(n10161), .ZN(n13455) );
  AND2_X1 U16845 ( .A1(n13455), .A2(n12732), .ZN(n13915) );
  NOR2_X1 U16846 ( .A1(n13456), .A2(n13915), .ZN(n13457) );
  MUX2_X1 U16847 ( .A(n13458), .B(n13457), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13459) );
  NAND2_X1 U16848 ( .A1(n13460), .A2(n13459), .ZN(n16051) );
  AOI22_X1 U16849 ( .A1(n19678), .A2(n16049), .B1(n19669), .B2(n16051), .ZN(
        n13469) );
  NAND2_X1 U16850 ( .A1(n13462), .A2(n13461), .ZN(n13463) );
  NOR2_X1 U16851 ( .A1(n13464), .A2(n13463), .ZN(n13466) );
  NAND3_X1 U16852 ( .A1(n18942), .A2(n18941), .A3(n16063), .ZN(n13465) );
  NAND2_X1 U16853 ( .A1(n13466), .A2(n13465), .ZN(n16077) );
  NAND2_X1 U16854 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n16095) );
  NOR2_X1 U16855 ( .A1(n19729), .A2(n16095), .ZN(n16103) );
  INV_X1 U16856 ( .A(n16103), .ZN(n16097) );
  OAI22_X1 U16857 ( .A1(n16097), .A2(n18634), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19697), .ZN(n13467) );
  AOI21_X1 U16858 ( .B1(n16077), .B2(n19720), .A(n13467), .ZN(n15502) );
  NAND2_X1 U16859 ( .A1(n15502), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13468) );
  OAI21_X1 U16860 ( .B1(n13469), .B2(n15502), .A(n13468), .ZN(P2_U3596) );
  INV_X1 U16861 ( .A(n13470), .ZN(n13474) );
  INV_X1 U16862 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13923) );
  AOI21_X1 U16863 ( .B1(n14653), .B2(n13471), .A(n13923), .ZN(n13472) );
  AOI211_X1 U16864 ( .C1(n13474), .C2(n19912), .A(n13473), .B(n13472), .ZN(
        n13475) );
  OAI21_X1 U16865 ( .B1(n19960), .B2(n13929), .A(n13475), .ZN(P1_U2999) );
  INV_X1 U16866 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U16867 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13476) );
  OAI21_X1 U16868 ( .B1(n13477), .B2(n13486), .A(n13476), .ZN(P1_U2920) );
  AOI22_X1 U16869 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13478) );
  OAI21_X1 U16870 ( .B1(n11824), .B2(n13486), .A(n13478), .ZN(P1_U2919) );
  AOI22_X1 U16871 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13479) );
  OAI21_X1 U16872 ( .B1(n11841), .B2(n13486), .A(n13479), .ZN(P1_U2918) );
  AOI22_X1 U16873 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13480) );
  OAI21_X1 U16874 ( .B1(n11900), .B2(n13486), .A(n13480), .ZN(P1_U2916) );
  AOI22_X1 U16875 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13481) );
  OAI21_X1 U16876 ( .B1(n11876), .B2(n13486), .A(n13481), .ZN(P1_U2915) );
  INV_X1 U16877 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U16878 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13482) );
  OAI21_X1 U16879 ( .B1(n13483), .B2(n13486), .A(n13482), .ZN(P1_U2914) );
  INV_X1 U16880 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14483) );
  AOI22_X1 U16881 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13484) );
  OAI21_X1 U16882 ( .B1(n14483), .B2(n13486), .A(n13484), .ZN(P1_U2913) );
  AOI22_X1 U16883 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13485) );
  OAI21_X1 U16884 ( .B1(n11857), .B2(n13486), .A(n13485), .ZN(P1_U2917) );
  INV_X1 U16885 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13878) );
  NOR2_X1 U16886 ( .A1(n19942), .A2(n13878), .ZN(n13495) );
  NOR2_X1 U16887 ( .A1(n14653), .A2(n13488), .ZN(n13487) );
  AOI211_X1 U16888 ( .C1(n15731), .C2(n13488), .A(n13495), .B(n13487), .ZN(
        n13492) );
  OR2_X1 U16889 ( .A1(n13489), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13496) );
  NAND3_X1 U16890 ( .A1(n13496), .A2(n13490), .A3(n19912), .ZN(n13491) );
  OAI211_X1 U16891 ( .C1(n13885), .C2(n19960), .A(n13492), .B(n13491), .ZN(
        P1_U2998) );
  NOR3_X1 U16892 ( .A1(n15790), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13493), .ZN(n13494) );
  AOI211_X1 U16893 ( .C1(n19925), .C2(n13877), .A(n13495), .B(n13494), .ZN(
        n13498) );
  NAND3_X1 U16894 ( .A1(n13496), .A2(n13490), .A3(n19929), .ZN(n13497) );
  OAI211_X1 U16895 ( .C1(n13499), .C2(n19941), .A(n13498), .B(n13497), .ZN(
        P1_U3030) );
  INV_X1 U16896 ( .A(n13500), .ZN(n13501) );
  AOI21_X1 U16897 ( .B1(n13503), .B2(n13502), .A(n13501), .ZN(n13593) );
  INV_X1 U16898 ( .A(n13593), .ZN(n13960) );
  INV_X2 U16899 ( .A(n19847), .ZN(n14463) );
  NAND2_X1 U16900 ( .A1(n13505), .A2(n13504), .ZN(n13506) );
  NAND2_X1 U16901 ( .A1(n13556), .A2(n13506), .ZN(n19944) );
  INV_X1 U16902 ( .A(n19944), .ZN(n13507) );
  AOI22_X1 U16903 ( .A1(n19846), .A2(n13507), .B1(n14446), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13508) );
  OAI21_X1 U16904 ( .B1(n13960), .B2(n14463), .A(n13508), .ZN(P1_U2870) );
  OAI222_X1 U16905 ( .A1(n13960), .A2(n14493), .B1(n14137), .B2(n19984), .C1(
        n14482), .C2(n11601), .ZN(P1_U2902) );
  INV_X1 U16906 ( .A(n13510), .ZN(n13512) );
  OAI21_X1 U16907 ( .B1(n10758), .B2(n13512), .A(n13511), .ZN(n16026) );
  INV_X1 U16908 ( .A(n13611), .ZN(n13547) );
  OAI211_X1 U16909 ( .C1(n13513), .C2(n13514), .A(n13547), .B(n14870), .ZN(
        n13516) );
  NAND2_X1 U16910 ( .A1(n14873), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13515) );
  OAI211_X1 U16911 ( .C1(n16026), .C2(n14873), .A(n13516), .B(n13515), .ZN(
        P2_U2879) );
  AOI21_X1 U16912 ( .B1(n13519), .B2(n13518), .A(n13517), .ZN(n14211) );
  XNOR2_X1 U16913 ( .A(n19682), .B(n14211), .ZN(n13524) );
  INV_X1 U16914 ( .A(n19694), .ZN(n13520) );
  NAND2_X1 U16915 ( .A1(n19689), .A2(n13520), .ZN(n13521) );
  OAI21_X1 U16916 ( .B1(n19689), .B2(n13520), .A(n13521), .ZN(n18934) );
  NOR2_X1 U16917 ( .A1(n18934), .A2(n18935), .ZN(n18933) );
  INV_X1 U16918 ( .A(n13521), .ZN(n13522) );
  NOR2_X1 U16919 ( .A1(n18933), .A2(n13522), .ZN(n13523) );
  NOR2_X1 U16920 ( .A1(n13523), .A2(n13524), .ZN(n13854) );
  AOI21_X1 U16921 ( .B1(n13524), .B2(n13523), .A(n13854), .ZN(n13527) );
  OAI22_X1 U16922 ( .A1(n18891), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n18892), .ZN(n19028) );
  INV_X1 U16923 ( .A(n19028), .ZN(n15969) );
  AOI22_X1 U16924 ( .A1(n18913), .A2(n15969), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n18931), .ZN(n13526) );
  INV_X1 U16925 ( .A(n14211), .ZN(n19685) );
  NAND2_X1 U16926 ( .A1(n19685), .A2(n18932), .ZN(n13525) );
  OAI211_X1 U16927 ( .C1(n13527), .C2(n18936), .A(n13526), .B(n13525), .ZN(
        P2_U2917) );
  XOR2_X1 U16928 ( .A(n13542), .B(n13541), .Z(n13605) );
  INV_X1 U16929 ( .A(n13605), .ZN(n13876) );
  OAI222_X1 U16930 ( .A1(n13876), .A2(n14493), .B1(n14137), .B2(n19988), .C1(
        n14482), .C2(n11631), .ZN(P1_U2901) );
  NAND2_X1 U16931 ( .A1(n13108), .A2(n13642), .ZN(n13528) );
  XNOR2_X1 U16932 ( .A(n14195), .B(n13528), .ZN(n13537) );
  OAI22_X1 U16933 ( .A1(n10128), .A2(n18845), .B1(n13529), .B2(n18865), .ZN(
        n13532) );
  OAI22_X1 U16934 ( .A1(n14211), .A2(n18841), .B1(n13530), .B2(n18871), .ZN(
        n13531) );
  AOI211_X1 U16935 ( .C1(P2_EBX_REG_2__SCAN_IN), .C2(n18861), .A(n13532), .B(
        n13531), .ZN(n13535) );
  NAND2_X1 U16936 ( .A1(n13533), .A2(n18868), .ZN(n13534) );
  OAI211_X1 U16937 ( .C1(n18851), .C2(n19682), .A(n13535), .B(n13534), .ZN(
        n13536) );
  AOI21_X1 U16938 ( .B1(n13537), .B2(n18838), .A(n13536), .ZN(n13538) );
  INV_X1 U16939 ( .A(n13538), .ZN(P2_U2853) );
  NAND2_X1 U16940 ( .A1(n13542), .A2(n13541), .ZN(n13544) );
  NAND2_X1 U16941 ( .A1(n13544), .A2(n13543), .ZN(n13545) );
  AND2_X1 U16942 ( .A1(n13540), .A2(n13545), .ZN(n19910) );
  INV_X1 U16943 ( .A(n19910), .ZN(n13571) );
  INV_X1 U16944 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20749) );
  OAI222_X1 U16945 ( .A1(n13571), .A2(n14493), .B1(n14137), .B2(n19991), .C1(
        n14482), .C2(n20749), .ZN(P1_U2900) );
  INV_X1 U16946 ( .A(n13546), .ZN(n13548) );
  OR2_X1 U16947 ( .A1(n13547), .A2(n13546), .ZN(n13559) );
  OAI211_X1 U16948 ( .C1(n13611), .C2(n13548), .A(n14870), .B(n13559), .ZN(
        n13553) );
  NAND2_X1 U16949 ( .A1(n13511), .A2(n13549), .ZN(n13550) );
  NAND2_X1 U16950 ( .A1(n13564), .A2(n13550), .ZN(n18793) );
  INV_X1 U16951 ( .A(n18793), .ZN(n13551) );
  NAND2_X1 U16952 ( .A1(n13551), .A2(n14840), .ZN(n13552) );
  OAI211_X1 U16953 ( .C1(n14840), .C2(n10761), .A(n13553), .B(n13552), .ZN(
        P2_U2878) );
  INV_X1 U16954 ( .A(n13569), .ZN(n13554) );
  AOI21_X1 U16955 ( .B1(n13556), .B2(n13555), .A(n13554), .ZN(n19926) );
  INV_X1 U16956 ( .A(n19926), .ZN(n13558) );
  INV_X1 U16957 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13557) );
  OAI222_X1 U16958 ( .A1(n13558), .A2(n14465), .B1(n19851), .B2(n13557), .C1(
        n14463), .C2(n13876), .ZN(P1_U2869) );
  INV_X1 U16959 ( .A(n13559), .ZN(n13563) );
  INV_X1 U16960 ( .A(n13560), .ZN(n13562) );
  NAND2_X1 U16961 ( .A1(n13611), .A2(n13561), .ZN(n13662) );
  OAI211_X1 U16962 ( .C1(n13563), .C2(n13562), .A(n14870), .B(n13662), .ZN(
        n13567) );
  AOI21_X1 U16963 ( .B1(n13565), .B2(n13564), .A(n13659), .ZN(n16006) );
  NAND2_X1 U16964 ( .A1(n16006), .A2(n14840), .ZN(n13566) );
  OAI211_X1 U16965 ( .C1(n14840), .C2(n9925), .A(n13567), .B(n13566), .ZN(
        P2_U2877) );
  AND2_X1 U16966 ( .A1(n13569), .A2(n13568), .ZN(n13570) );
  NOR2_X1 U16967 ( .A1(n15874), .A2(n13570), .ZN(n19918) );
  INV_X1 U16968 ( .A(n19918), .ZN(n13572) );
  INV_X1 U16969 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19826) );
  OAI222_X1 U16970 ( .A1(n13572), .A2(n14465), .B1(n19851), .B2(n19826), .C1(
        n14463), .C2(n13571), .ZN(P1_U2868) );
  INV_X1 U16971 ( .A(n13442), .ZN(n13573) );
  AOI21_X1 U16972 ( .B1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13785), .A(
        n13573), .ZN(n13576) );
  NAND2_X1 U16973 ( .A1(n13574), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13578) );
  NAND3_X1 U16974 ( .A1(n13576), .A2(n13575), .A3(n13578), .ZN(n13582) );
  INV_X1 U16975 ( .A(n13576), .ZN(n13581) );
  INV_X1 U16976 ( .A(n13577), .ZN(n13580) );
  INV_X1 U16977 ( .A(n13578), .ZN(n13579) );
  OAI21_X1 U16978 ( .B1(n13581), .B2(n13580), .A(n13579), .ZN(n13648) );
  NAND2_X1 U16979 ( .A1(n13582), .A2(n13648), .ZN(n18915) );
  NAND2_X1 U16980 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  NAND2_X1 U16981 ( .A1(n13583), .A2(n13586), .ZN(n19056) );
  MUX2_X1 U16982 ( .A(n10373), .B(n19056), .S(n14840), .Z(n13587) );
  OAI21_X1 U16983 ( .B1(n18915), .B2(n14880), .A(n13587), .ZN(P2_U2883) );
  OAI21_X1 U16984 ( .B1(n13588), .B2(n13590), .A(n13589), .ZN(n19947) );
  AOI22_X1 U16985 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13591) );
  OAI21_X1 U16986 ( .B1(n19916), .B2(n13950), .A(n13591), .ZN(n13592) );
  AOI21_X1 U16987 ( .B1(n13593), .B2(n19911), .A(n13592), .ZN(n13594) );
  OAI21_X1 U16988 ( .B1(n19746), .B2(n19947), .A(n13594), .ZN(P1_U2997) );
  NAND2_X1 U16989 ( .A1(n13540), .A2(n13596), .ZN(n13597) );
  AND2_X1 U16990 ( .A1(n13595), .A2(n13597), .ZN(n19848) );
  INV_X1 U16991 ( .A(n19848), .ZN(n13599) );
  OAI222_X1 U16992 ( .A1(n13599), .A2(n14493), .B1(n14137), .B2(n19995), .C1(
        n13598), .C2(n14482), .ZN(P1_U2899) );
  OAI21_X1 U16993 ( .B1(n13600), .B2(n13602), .A(n9641), .ZN(n19927) );
  NAND2_X1 U16994 ( .A1(n12105), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n19923) );
  NAND2_X1 U16995 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13603) );
  OAI211_X1 U16996 ( .C1(n19916), .C2(n13870), .A(n19923), .B(n13603), .ZN(
        n13604) );
  AOI21_X1 U16997 ( .B1(n13605), .B2(n19911), .A(n13604), .ZN(n13606) );
  OAI21_X1 U16998 ( .B1(n19927), .B2(n19746), .A(n13606), .ZN(P1_U2996) );
  INV_X1 U16999 ( .A(n13607), .ZN(n13610) );
  OAI21_X1 U17000 ( .B1(n13610), .B2(n10775), .A(n13609), .ZN(n18762) );
  AND2_X1 U17001 ( .A1(n13611), .A2(n13612), .ZN(n13661) );
  NAND2_X1 U17002 ( .A1(n13611), .A2(n13613), .ZN(n13817) );
  OAI211_X1 U17003 ( .C1(n13661), .C2(n13614), .A(n13817), .B(n14870), .ZN(
        n13616) );
  NAND2_X1 U17004 ( .A1(n14873), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13615) );
  OAI211_X1 U17005 ( .C1(n18762), .C2(n14873), .A(n13616), .B(n13615), .ZN(
        P2_U2875) );
  NOR2_X1 U17006 ( .A1(n18810), .A2(n13617), .ZN(n13618) );
  XNOR2_X1 U17007 ( .A(n13618), .B(n13764), .ZN(n13629) );
  OAI22_X1 U17008 ( .A1(n10180), .A2(n18845), .B1(n13619), .B2(n18865), .ZN(
        n13625) );
  INV_X1 U17009 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13763) );
  OR2_X1 U17010 ( .A1(n13621), .A2(n13620), .ZN(n13623) );
  NAND2_X1 U17011 ( .A1(n13623), .A2(n13622), .ZN(n19676) );
  OAI22_X1 U17012 ( .A1(n13763), .A2(n18871), .B1(n18841), .B2(n19676), .ZN(
        n13624) );
  AOI211_X1 U17013 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n18861), .A(n13625), .B(
        n13624), .ZN(n13627) );
  NAND2_X1 U17014 ( .A1(n13444), .A2(n18868), .ZN(n13626) );
  OAI211_X1 U17015 ( .C1(n18851), .C2(n13855), .A(n13627), .B(n13626), .ZN(
        n13628) );
  AOI21_X1 U17016 ( .B1(n13629), .B2(n18838), .A(n13628), .ZN(n13630) );
  INV_X1 U17017 ( .A(n13630), .ZN(P2_U2852) );
  XOR2_X1 U17018 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13648), .Z(n13636)
         );
  INV_X1 U17019 ( .A(n13653), .ZN(n13631) );
  AOI21_X1 U17020 ( .B1(n13632), .B2(n13583), .A(n13631), .ZN(n18836) );
  NOR2_X1 U17021 ( .A1(n14840), .A2(n13633), .ZN(n13634) );
  AOI21_X1 U17022 ( .B1(n18836), .B2(n14840), .A(n13634), .ZN(n13635) );
  OAI21_X1 U17023 ( .B1(n13636), .B2(n14880), .A(n13635), .ZN(P2_U2882) );
  OAI22_X1 U17024 ( .A1(n18845), .A2(n10168), .B1(n13637), .B2(n18865), .ZN(
        n13640) );
  INV_X1 U17025 ( .A(n18861), .ZN(n18777) );
  OAI22_X1 U17026 ( .A1(n18777), .A2(n10171), .B1(n13638), .B2(n18871), .ZN(
        n13639) );
  AOI211_X1 U17027 ( .C1(n18859), .C2(n19694), .A(n13640), .B(n13639), .ZN(
        n13641) );
  OAI21_X1 U17028 ( .B1(n10212), .B2(n18858), .A(n13641), .ZN(n13645) );
  NAND2_X1 U17029 ( .A1(n18838), .A2(n18810), .ZN(n18870) );
  OAI211_X1 U17030 ( .C1(n18878), .C2(n13643), .A(n13108), .B(n13642), .ZN(
        n13712) );
  OAI22_X1 U17031 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18870), .B1(
        n13712), .B2(n19582), .ZN(n13644) );
  AOI211_X1 U17032 ( .C1(n18872), .C2(n19692), .A(n13645), .B(n13644), .ZN(
        n13646) );
  INV_X1 U17033 ( .A(n13646), .ZN(P2_U2854) );
  NOR2_X1 U17034 ( .A1(n13648), .A2(n13647), .ZN(n13651) );
  INV_X1 U17035 ( .A(n13649), .ZN(n13650) );
  OAI211_X1 U17036 ( .C1(n13651), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14870), .B(n13650), .ZN(n13656) );
  AND2_X1 U17037 ( .A1(n13653), .A2(n13652), .ZN(n13654) );
  NAND2_X1 U17038 ( .A1(n9716), .A2(n14840), .ZN(n13655) );
  OAI211_X1 U17039 ( .C1(n14840), .C2(n13657), .A(n13656), .B(n13655), .ZN(
        P2_U2881) );
  OAI21_X1 U17040 ( .B1(n13659), .B2(n13658), .A(n13607), .ZN(n13660) );
  INV_X1 U17041 ( .A(n13660), .ZN(n18769) );
  NOR2_X1 U17042 ( .A1(n14840), .A2(n18763), .ZN(n13665) );
  AOI211_X1 U17043 ( .C1(n13663), .C2(n13662), .A(n14880), .B(n13661), .ZN(
        n13664) );
  AOI211_X1 U17044 ( .C1(n18769), .C2(n14840), .A(n13665), .B(n13664), .ZN(
        n13666) );
  INV_X1 U17045 ( .A(n13666), .ZN(P2_U2876) );
  INV_X1 U17046 ( .A(n20233), .ZN(n13873) );
  MUX2_X1 U17047 ( .A(n13667), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n13684), .Z(n15557) );
  NOR2_X1 U17048 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20553), .ZN(n13685) );
  AOI22_X1 U17049 ( .A1(n15557), .A2(n20553), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13685), .ZN(n13681) );
  NAND2_X1 U17050 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U17051 ( .A1(n13669), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n11104), .B2(n13668), .ZN(n13674) );
  AOI21_X1 U17052 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13670), .A(
        n11369), .ZN(n20624) );
  NOR3_X1 U17053 ( .A1(n13672), .A2(n20624), .A3(n13671), .ZN(n13673) );
  AOI21_X1 U17054 ( .B1(n15550), .B2(n13674), .A(n13673), .ZN(n13679) );
  XNOR2_X1 U17055 ( .A(n13675), .B(n11104), .ZN(n13676) );
  NAND2_X1 U17056 ( .A1(n13677), .A2(n13676), .ZN(n13678) );
  OAI211_X1 U17057 ( .C1(n13873), .C2(n14794), .A(n13679), .B(n13678), .ZN(
        n20622) );
  INV_X1 U17058 ( .A(n13684), .ZN(n15548) );
  MUX2_X1 U17059 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20622), .S(
        n15548), .Z(n15562) );
  AOI22_X1 U17060 ( .A1(n13685), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20553), .B2(n15562), .ZN(n13680) );
  NOR2_X1 U17061 ( .A1(n13681), .A2(n13680), .ZN(n15570) );
  INV_X1 U17062 ( .A(n13682), .ZN(n14803) );
  NAND2_X1 U17063 ( .A1(n15570), .A2(n14803), .ZN(n14790) );
  OAI21_X1 U17064 ( .B1(n19831), .B2(n12437), .A(n15548), .ZN(n13687) );
  AOI21_X1 U17065 ( .B1(n13684), .B2(n13683), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13686) );
  AOI22_X1 U17066 ( .A1(n13687), .A2(n13686), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13685), .ZN(n15572) );
  AND3_X1 U17067 ( .A1(n14790), .A2(n15572), .A3(n19747), .ZN(n13689) );
  INV_X1 U17068 ( .A(n20119), .ZN(n19965) );
  INV_X1 U17069 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20371) );
  NAND2_X1 U17070 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20371), .ZN(n14791) );
  AND2_X1 U17071 ( .A1(n19956), .A2(n14791), .ZN(n13695) );
  INV_X1 U17072 ( .A(n13695), .ZN(n14187) );
  INV_X1 U17073 ( .A(n19956), .ZN(n14183) );
  NOR2_X1 U17074 ( .A1(n14183), .A2(n20493), .ZN(n14185) );
  NAND2_X1 U17075 ( .A1(n13691), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20333) );
  NOR2_X1 U17076 ( .A1(n13690), .A2(n20333), .ZN(n14182) );
  INV_X1 U17077 ( .A(n20333), .ZN(n20497) );
  NAND2_X1 U17078 ( .A1(n20112), .A2(n20497), .ZN(n20205) );
  OAI21_X1 U17079 ( .B1(n14182), .B2(n11624), .A(n20205), .ZN(n13692) );
  AOI22_X1 U17080 ( .A1(n14185), .A2(n13692), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14183), .ZN(n13693) );
  OAI21_X1 U17081 ( .B1(n13873), .B2(n14187), .A(n13693), .ZN(P1_U3475) );
  OAI211_X1 U17082 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n13691), .A(n14185), 
        .B(n20333), .ZN(n13697) );
  NAND2_X1 U17083 ( .A1(n13695), .A2(n9648), .ZN(n13696) );
  OAI211_X1 U17084 ( .C1(n11542), .C2(n19956), .A(n13697), .B(n13696), .ZN(
        P1_U3477) );
  OR2_X1 U17085 ( .A1(n9642), .A2(n13700), .ZN(n13701) );
  AND2_X1 U17086 ( .A1(n13698), .A2(n13701), .ZN(n19801) );
  INV_X1 U17087 ( .A(n19801), .ZN(n13702) );
  INV_X1 U17088 ( .A(n14486), .ZN(n20004) );
  OAI222_X1 U17089 ( .A1(n13702), .A2(n14493), .B1(n14137), .B2(n20004), .C1(
        n14482), .C2(n11662), .ZN(P1_U2897) );
  INV_X1 U17090 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13708) );
  NAND2_X1 U17091 ( .A1(n19801), .A2(n19847), .ZN(n13707) );
  AND2_X1 U17092 ( .A1(n13704), .A2(n13703), .ZN(n13705) );
  NOR2_X1 U17093 ( .A1(n13828), .A2(n13705), .ZN(n19792) );
  NAND2_X1 U17094 ( .A1(n19792), .A2(n19846), .ZN(n13706) );
  OAI211_X1 U17095 ( .C1(n13708), .C2(n19851), .A(n13707), .B(n13706), .ZN(
        P1_U2865) );
  AND2_X1 U17096 ( .A1(n13595), .A2(n13709), .ZN(n13710) );
  NOR2_X1 U17097 ( .A1(n9642), .A2(n13710), .ZN(n19842) );
  INV_X1 U17098 ( .A(n19842), .ZN(n13711) );
  OAI222_X1 U17099 ( .A1(n13711), .A2(n14493), .B1(n14137), .B2(n19998), .C1(
        n14482), .C2(n11651), .ZN(P1_U2898) );
  OAI21_X1 U17100 ( .B1(n13108), .B2(n13713), .A(n13712), .ZN(n13920) );
  INV_X1 U17101 ( .A(n13920), .ZN(n13726) );
  AOI221_X1 U17102 ( .B1(n18878), .B2(n13108), .C1(n13714), .C2(n18810), .A(
        n18626), .ZN(n15407) );
  NAND2_X1 U17103 ( .A1(n9587), .A2(n13715), .ZN(n13725) );
  INV_X1 U17104 ( .A(n13717), .ZN(n13719) );
  NAND2_X1 U17105 ( .A1(n13719), .A2(n13718), .ZN(n15400) );
  INV_X1 U17106 ( .A(n13720), .ZN(n13722) );
  NAND2_X1 U17107 ( .A1(n9634), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13721) );
  NAND2_X1 U17108 ( .A1(n13722), .A2(n13721), .ZN(n13723) );
  AOI22_X1 U17109 ( .A1(n10016), .A2(n13450), .B1(n15400), .B2(n13723), .ZN(
        n13724) );
  NAND2_X1 U17110 ( .A1(n13725), .A2(n13724), .ZN(n16078) );
  AOI222_X1 U17111 ( .A1(n13726), .A2(n15407), .B1(n19692), .B2(n16049), .C1(
        n16078), .C2(n19669), .ZN(n13728) );
  NAND2_X1 U17112 ( .A1(n15502), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13727) );
  OAI21_X1 U17113 ( .B1(n13728), .B2(n15502), .A(n13727), .ZN(P2_U3600) );
  NAND2_X1 U17114 ( .A1(n13855), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19201) );
  NAND2_X1 U17115 ( .A1(n19680), .A2(n19450), .ZN(n13737) );
  OAI21_X1 U17116 ( .B1(n19201), .B2(n19670), .A(n13737), .ZN(n13733) );
  INV_X1 U17117 ( .A(n19347), .ZN(n13729) );
  NAND2_X1 U17118 ( .A1(n19680), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19234) );
  INV_X1 U17119 ( .A(n19234), .ZN(n19165) );
  NAND2_X1 U17120 ( .A1(n13729), .A2(n19165), .ZN(n19282) );
  OAI211_X1 U17121 ( .C1(n10446), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19282), 
        .B(n19454), .ZN(n13731) );
  OAI21_X1 U17122 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n19729), .ZN(n19726) );
  INV_X1 U17123 ( .A(n19726), .ZN(n16093) );
  AND2_X1 U17124 ( .A1(n13731), .A2(n19515), .ZN(n13732) );
  NAND2_X1 U17125 ( .A1(n13733), .A2(n13732), .ZN(n19275) );
  INV_X1 U17126 ( .A(n19275), .ZN(n19261) );
  AOI22_X2 U17127 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n13795), .ZN(n19535) );
  INV_X1 U17128 ( .A(n19535), .ZN(n19145) );
  INV_X1 U17129 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16183) );
  INV_X1 U17130 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17963) );
  OAI22_X2 U17131 ( .A1(n16183), .A2(n13798), .B1(n17963), .B2(n13797), .ZN(
        n19532) );
  AOI22_X1 U17132 ( .A1(n19306), .A2(n19145), .B1(n19274), .B2(n19532), .ZN(
        n13740) );
  INV_X1 U17133 ( .A(n19282), .ZN(n19285) );
  OAI21_X1 U17134 ( .B1(n13735), .B2(n19285), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13736) );
  OAI21_X1 U17135 ( .B1(n13737), .B2(n19454), .A(n13736), .ZN(n19273) );
  NAND2_X1 U17136 ( .A1(n15969), .A2(n19515), .ZN(n19530) );
  NAND2_X1 U17137 ( .A1(n13738), .A2(n13799), .ZN(n19529) );
  AOI22_X1 U17138 ( .A1(n19273), .A2(n19470), .B1(n19469), .B2(n19285), .ZN(
        n13739) );
  OAI211_X1 U17139 ( .C1(n19261), .C2(n13741), .A(n13740), .B(n13739), .ZN(
        P2_U3106) );
  NAND2_X1 U17140 ( .A1(n19687), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19349) );
  NOR2_X1 U17141 ( .A1(n19349), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13748) );
  INV_X1 U17142 ( .A(n13748), .ZN(n19278) );
  NAND2_X1 U17143 ( .A1(n19511), .A2(n19083), .ZN(n13742) );
  NAND2_X1 U17144 ( .A1(n13742), .A2(n19681), .ZN(n13749) );
  NOR2_X1 U17145 ( .A1(n19278), .A2(n13749), .ZN(n13744) );
  NOR2_X1 U17146 ( .A1(n19200), .A2(n19349), .ZN(n19315) );
  INV_X1 U17147 ( .A(n19315), .ZN(n13801) );
  AOI21_X1 U17148 ( .B1(n10383), .B2(n13801), .A(n19504), .ZN(n13743) );
  INV_X1 U17149 ( .A(n19024), .ZN(n18881) );
  NAND2_X1 U17150 ( .A1(n18881), .A2(n19515), .ZN(n19509) );
  OR2_X1 U17151 ( .A1(n10383), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13746) );
  NOR2_X1 U17152 ( .A1(n19681), .A2(n19315), .ZN(n13745) );
  AOI21_X1 U17153 ( .B1(n13746), .B2(n13745), .A(n19392), .ZN(n13747) );
  INV_X1 U17154 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16200) );
  INV_X1 U17155 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n17949) );
  OAI22_X2 U17156 ( .A1(n16200), .A2(n13798), .B1(n17949), .B2(n13797), .ZN(
        n19518) );
  INV_X1 U17157 ( .A(n19518), .ZN(n13839) );
  AOI22_X1 U17158 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n13795), .ZN(n19521) );
  INV_X1 U17159 ( .A(n19521), .ZN(n19323) );
  NOR2_X2 U17160 ( .A1(n10121), .A2(n13750), .ZN(n19451) );
  AOI22_X1 U17161 ( .A1(n19323), .A2(n19299), .B1(n19451), .B2(n19315), .ZN(
        n13751) );
  OAI21_X1 U17162 ( .B1(n13839), .B2(n19336), .A(n13751), .ZN(n13752) );
  AOI21_X1 U17163 ( .B1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B2(n13804), .A(
        n13752), .ZN(n13753) );
  OAI21_X1 U17164 ( .B1(n13807), .B2(n19509), .A(n13753), .ZN(P2_U3120) );
  OAI22_X1 U17165 ( .A1(n18891), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n18892), .ZN(n19032) );
  INV_X1 U17166 ( .A(n19032), .ZN(n15963) );
  NAND2_X1 U17167 ( .A1(n15963), .A2(n19515), .ZN(n19544) );
  AOI22_X1 U17168 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n13795), .ZN(n19549) );
  AOI22_X1 U17169 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n13795), .ZN(n19485) );
  AOI22_X1 U17170 ( .A1(n19546), .A2(n19299), .B1(n19315), .B2(n19479), .ZN(
        n13755) );
  OAI21_X1 U17171 ( .B1(n19549), .B2(n19336), .A(n13755), .ZN(n13756) );
  AOI21_X1 U17172 ( .B1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B2(n13804), .A(
        n13756), .ZN(n13757) );
  OAI21_X1 U17173 ( .B1(n13807), .B2(n19544), .A(n13757), .ZN(P2_U3124) );
  XNOR2_X1 U17174 ( .A(n13759), .B(n13758), .ZN(n16041) );
  XNOR2_X1 U17175 ( .A(n13760), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13761) );
  XNOR2_X1 U17176 ( .A(n13762), .B(n13761), .ZN(n16043) );
  NAND2_X1 U17177 ( .A1(n16043), .A2(n19050), .ZN(n13768) );
  NAND2_X1 U17178 ( .A1(n15392), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16035) );
  OAI21_X1 U17179 ( .B1(n19061), .B2(n13763), .A(n16035), .ZN(n13766) );
  NOR2_X1 U17180 ( .A1(n15144), .A2(n13764), .ZN(n13765) );
  AOI211_X1 U17181 ( .C1(n16001), .C2(n13444), .A(n13766), .B(n13765), .ZN(
        n13767) );
  OAI211_X1 U17182 ( .C1(n16041), .C2(n15996), .A(n13768), .B(n13767), .ZN(
        P2_U3011) );
  NAND2_X1 U17183 ( .A1(n13698), .A2(n13770), .ZN(n13771) );
  AND2_X1 U17184 ( .A1(n13769), .A2(n13771), .ZN(n19784) );
  INV_X1 U17185 ( .A(n19784), .ZN(n13830) );
  INV_X1 U17186 ( .A(n14137), .ZN(n14078) );
  INV_X1 U17187 ( .A(DATAI_8_), .ZN(n13773) );
  NAND2_X1 U17188 ( .A1(n19957), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13772) );
  OAI21_X1 U17189 ( .B1(n19957), .B2(n13773), .A(n13772), .ZN(n19877) );
  AOI22_X1 U17190 ( .A1(n14078), .A2(n19877), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14506), .ZN(n13774) );
  OAI21_X1 U17191 ( .B1(n13830), .B2(n14493), .A(n13774), .ZN(P1_U2896) );
  AOI22_X1 U17192 ( .A1(n18892), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n18891), .ZN(n19034) );
  INV_X1 U17193 ( .A(n19034), .ZN(n18914) );
  NAND2_X1 U17194 ( .A1(n18914), .A2(n19515), .ZN(n19551) );
  AOI22_X1 U17195 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n13795), .ZN(n19491) );
  AOI22_X1 U17196 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n13795), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n13796), .ZN(n19558) );
  NAND2_X1 U17197 ( .A1(n10339), .A2(n13799), .ZN(n19550) );
  OAI22_X1 U17198 ( .A1(n19558), .A2(n19311), .B1(n13801), .B2(n19550), .ZN(
        n13775) );
  AOI21_X1 U17199 ( .B1(n19343), .B2(n19553), .A(n13775), .ZN(n13777) );
  NAND2_X1 U17200 ( .A1(n13804), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n13776) );
  OAI211_X1 U17201 ( .C1(n13807), .C2(n19551), .A(n13777), .B(n13776), .ZN(
        P2_U3125) );
  AOI22_X1 U17202 ( .A1(n18892), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n18891), .ZN(n19030) );
  NOR2_X2 U17203 ( .A1(n19030), .A2(n19392), .ZN(n19475) );
  INV_X1 U17204 ( .A(n19475), .ZN(n19537) );
  AOI22_X1 U17205 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n13795), .ZN(n19542) );
  AOI22_X1 U17206 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n13795), .ZN(n19478) );
  NAND2_X1 U17207 ( .A1(n13778), .A2(n13799), .ZN(n19536) );
  OAI22_X1 U17208 ( .A1(n19478), .A2(n19311), .B1(n13801), .B2(n19536), .ZN(
        n13779) );
  AOI21_X1 U17209 ( .B1(n19343), .B2(n19474), .A(n13779), .ZN(n13781) );
  NAND2_X1 U17210 ( .A1(n13804), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13780) );
  OAI211_X1 U17211 ( .C1(n13807), .C2(n19537), .A(n13781), .B(n13780), .ZN(
        P2_U3123) );
  INV_X1 U17212 ( .A(n19532), .ZN(n13850) );
  OAI22_X1 U17213 ( .A1(n13850), .A2(n19311), .B1(n19529), .B2(n13801), .ZN(
        n13782) );
  AOI21_X1 U17214 ( .B1(n19145), .B2(n19343), .A(n13782), .ZN(n13784) );
  NAND2_X1 U17215 ( .A1(n13804), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13783) );
  OAI211_X1 U17216 ( .C1(n13807), .C2(n19530), .A(n13784), .B(n13783), .ZN(
        P2_U3122) );
  OAI22_X1 U17217 ( .A1(n18891), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n18892), .ZN(n19036) );
  INV_X1 U17218 ( .A(n19036), .ZN(n15957) );
  NAND2_X1 U17219 ( .A1(n15957), .A2(n19515), .ZN(n19560) );
  INV_X1 U17220 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16191) );
  INV_X1 U17221 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17038) );
  NAND2_X1 U17222 ( .A1(n13785), .A2(n13799), .ZN(n19559) );
  AOI22_X1 U17223 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n13795), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n13796), .ZN(n19412) );
  NAND2_X1 U17224 ( .A1(n19562), .A2(n19299), .ZN(n13786) );
  OAI21_X1 U17225 ( .B1(n13801), .B2(n19559), .A(n13786), .ZN(n13787) );
  AOI21_X1 U17226 ( .B1(n19343), .B2(n19408), .A(n13787), .ZN(n13789) );
  NAND2_X1 U17227 ( .A1(n13804), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13788) );
  OAI211_X1 U17228 ( .C1(n13807), .C2(n19560), .A(n13789), .B(n13788), .ZN(
        P2_U3126) );
  AOI22_X1 U17229 ( .A1(n18892), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n18891), .ZN(n19026) );
  NOR2_X2 U17230 ( .A1(n19026), .A2(n19392), .ZN(n19466) );
  INV_X1 U17231 ( .A(n19466), .ZN(n19523) );
  AOI22_X2 U17232 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n13795), .ZN(n19528) );
  INV_X1 U17233 ( .A(n19528), .ZN(n19142) );
  INV_X1 U17234 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16185) );
  INV_X1 U17235 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n13790) );
  OAI22_X2 U17236 ( .A1(n16185), .A2(n13798), .B1(n13790), .B2(n13797), .ZN(
        n19525) );
  INV_X1 U17237 ( .A(n19525), .ZN(n13791) );
  NAND2_X1 U17238 ( .A1(n10208), .A2(n13799), .ZN(n19522) );
  OAI22_X1 U17239 ( .A1(n13791), .A2(n19311), .B1(n13801), .B2(n19522), .ZN(
        n13792) );
  AOI21_X1 U17240 ( .B1(n19343), .B2(n19142), .A(n13792), .ZN(n13794) );
  NAND2_X1 U17241 ( .A1(n13804), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13793) );
  OAI211_X1 U17242 ( .C1(n13807), .C2(n19523), .A(n13794), .B(n13793), .ZN(
        P2_U3121) );
  AOI22_X1 U17243 ( .A1(n18892), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n18891), .ZN(n19038) );
  NOR2_X2 U17244 ( .A1(n19038), .A2(n19392), .ZN(n19500) );
  INV_X1 U17245 ( .A(n19500), .ZN(n19568) );
  AOI22_X2 U17246 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n13796), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n13795), .ZN(n19577) );
  INV_X1 U17247 ( .A(n19577), .ZN(n19158) );
  INV_X1 U17248 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16997) );
  OAI22_X2 U17249 ( .A1(n16173), .A2(n13798), .B1(n16997), .B2(n13797), .ZN(
        n19571) );
  INV_X1 U17250 ( .A(n19571), .ZN(n13802) );
  NAND2_X1 U17251 ( .A1(n13800), .A2(n13799), .ZN(n19566) );
  OAI22_X1 U17252 ( .A1(n13802), .A2(n19311), .B1(n13801), .B2(n19566), .ZN(
        n13803) );
  AOI21_X1 U17253 ( .B1(n19343), .B2(n19158), .A(n13803), .ZN(n13806) );
  NAND2_X1 U17254 ( .A1(n13804), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n13805) );
  OAI211_X1 U17255 ( .C1(n13807), .C2(n19568), .A(n13806), .B(n13805), .ZN(
        P2_U3127) );
  AND2_X1 U17256 ( .A1(n13808), .A2(n13809), .ZN(n13888) );
  NOR2_X1 U17257 ( .A1(n13808), .A2(n13809), .ZN(n13810) );
  NAND2_X1 U17258 ( .A1(n13611), .A2(n13811), .ZN(n13818) );
  INV_X1 U17259 ( .A(n13818), .ZN(n13814) );
  NAND2_X1 U17260 ( .A1(n13611), .A2(n13812), .ZN(n13891) );
  OAI211_X1 U17261 ( .C1(n13814), .C2(n13813), .A(n14870), .B(n13891), .ZN(
        n13816) );
  NAND2_X1 U17262 ( .A1(n14873), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13815) );
  OAI211_X1 U17263 ( .C1(n18740), .C2(n14873), .A(n13816), .B(n13815), .ZN(
        P2_U2873) );
  INV_X1 U17264 ( .A(n13817), .ZN(n13820) );
  OAI211_X1 U17265 ( .C1(n13820), .C2(n13819), .A(n14870), .B(n13818), .ZN(
        n13826) );
  INV_X1 U17266 ( .A(n13808), .ZN(n13823) );
  NAND2_X1 U17267 ( .A1(n13609), .A2(n13821), .ZN(n13822) );
  NAND2_X1 U17268 ( .A1(n13823), .A2(n13822), .ZN(n18747) );
  INV_X1 U17269 ( .A(n18747), .ZN(n13824) );
  NAND2_X1 U17270 ( .A1(n13824), .A2(n14840), .ZN(n13825) );
  OAI211_X1 U17271 ( .C1(n14840), .C2(n10507), .A(n13826), .B(n13825), .ZN(
        P2_U2874) );
  OR2_X1 U17272 ( .A1(n13828), .A2(n13827), .ZN(n13829) );
  NAND2_X1 U17273 ( .A1(n15838), .A2(n13829), .ZN(n19780) );
  INV_X1 U17274 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13831) );
  OAI222_X1 U17275 ( .A1(n19780), .A2(n14465), .B1(n19851), .B2(n13831), .C1(
        n14463), .C2(n13830), .ZN(P1_U2864) );
  NAND2_X1 U17276 ( .A1(n19576), .A2(n19095), .ZN(n13833) );
  NAND2_X1 U17277 ( .A1(n13833), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13834) );
  NAND2_X1 U17278 ( .A1(n13834), .A2(n19681), .ZN(n13845) );
  INV_X1 U17279 ( .A(n19517), .ZN(n19567) );
  NAND2_X1 U17280 ( .A1(n19680), .A2(n19687), .ZN(n19131) );
  NOR3_X2 U17281 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19131), .ZN(n19074) );
  INV_X1 U17282 ( .A(n19074), .ZN(n13838) );
  NAND2_X1 U17283 ( .A1(n19567), .A2(n13838), .ZN(n13841) );
  OR2_X1 U17284 ( .A1(n13845), .A2(n13841), .ZN(n13837) );
  OAI211_X1 U17285 ( .C1(n10398), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n13838), 
        .B(n19454), .ZN(n13835) );
  AND2_X1 U17286 ( .A1(n13835), .A2(n19515), .ZN(n13836) );
  INV_X1 U17287 ( .A(n19076), .ZN(n19065) );
  INV_X1 U17288 ( .A(n19451), .ZN(n19508) );
  OAI22_X1 U17289 ( .A1(n13839), .A2(n19095), .B1(n19508), .B2(n13838), .ZN(
        n13840) );
  AOI21_X1 U17290 ( .B1(n19554), .B2(n19323), .A(n13840), .ZN(n13847) );
  INV_X1 U17291 ( .A(n13841), .ZN(n13844) );
  INV_X1 U17292 ( .A(n10398), .ZN(n13842) );
  OAI21_X1 U17293 ( .B1(n13842), .B2(n19074), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13843) );
  NAND2_X1 U17294 ( .A1(n19075), .A2(n19462), .ZN(n13846) );
  OAI211_X1 U17295 ( .C1(n19065), .C2(n13848), .A(n13847), .B(n13846), .ZN(
        P2_U3048) );
  AOI22_X1 U17296 ( .A1(n19145), .A2(n19104), .B1(n19469), .B2(n19074), .ZN(
        n13849) );
  OAI21_X1 U17297 ( .B1(n13850), .B2(n19576), .A(n13849), .ZN(n13851) );
  AOI21_X1 U17298 ( .B1(n19470), .B2(n19075), .A(n13851), .ZN(n13852) );
  OAI21_X1 U17299 ( .B1(n19065), .B2(n13853), .A(n13852), .ZN(P2_U3050) );
  AOI21_X1 U17300 ( .B1(n14211), .B2(n19682), .A(n13854), .ZN(n18927) );
  XNOR2_X1 U17301 ( .A(n13855), .B(n19676), .ZN(n18926) );
  NOR2_X1 U17302 ( .A1(n18927), .A2(n18926), .ZN(n18925) );
  AOI21_X1 U17303 ( .B1(n19676), .B2(n13855), .A(n18925), .ZN(n13858) );
  INV_X1 U17304 ( .A(n13622), .ZN(n13856) );
  XNOR2_X1 U17305 ( .A(n13857), .B(n13856), .ZN(n18843) );
  NOR2_X1 U17306 ( .A1(n13858), .A2(n18843), .ZN(n18916) );
  XNOR2_X1 U17307 ( .A(n18916), .B(n18915), .ZN(n13861) );
  AOI22_X1 U17308 ( .A1(n18932), .A2(n18843), .B1(n18931), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13860) );
  NAND2_X1 U17309 ( .A1(n18913), .A2(n15963), .ZN(n13859) );
  OAI211_X1 U17310 ( .C1(n13861), .C2(n18936), .A(n13860), .B(n13859), .ZN(
        P2_U2915) );
  OAI21_X1 U17311 ( .B1(n13863), .B2(n14305), .A(n15655), .ZN(n19833) );
  INV_X1 U17312 ( .A(n19833), .ZN(n13959) );
  INV_X1 U17313 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n19943) );
  NOR2_X1 U17314 ( .A1(n13878), .A2(n19943), .ZN(n13862) );
  OAI21_X1 U17315 ( .B1(n13862), .B2(n15677), .A(n14405), .ZN(n13972) );
  INV_X1 U17316 ( .A(n13863), .ZN(n13865) );
  NAND2_X1 U17317 ( .A1(n13865), .A2(n13864), .ZN(n19830) );
  NAND2_X2 U17318 ( .A1(n14405), .A2(n13867), .ZN(n19821) );
  NAND2_X1 U17319 ( .A1(n19797), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n13869) );
  INV_X1 U17320 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20577) );
  NAND3_X1 U17321 ( .A1(n15623), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .ZN(n13971) );
  INV_X1 U17322 ( .A(n13971), .ZN(n19819) );
  AOI22_X1 U17323 ( .A1(n19823), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20577), .B2(n19819), .ZN(n13868) );
  OAI211_X1 U17324 ( .C1(n19821), .C2(n13870), .A(n13869), .B(n13868), .ZN(
        n13871) );
  AOI21_X1 U17325 ( .B1(n19828), .B2(n19926), .A(n13871), .ZN(n13872) );
  OAI21_X1 U17326 ( .B1(n13873), .B2(n19830), .A(n13872), .ZN(n13874) );
  AOI21_X1 U17327 ( .B1(n13972), .B2(P1_REIP_REG_3__SCAN_IN), .A(n13874), .ZN(
        n13875) );
  OAI21_X1 U17328 ( .B1(n13876), .B2(n13959), .A(n13875), .ZN(P1_U2837) );
  INV_X1 U17329 ( .A(n19830), .ZN(n13956) );
  AOI22_X1 U17330 ( .A1(n15623), .A2(n13878), .B1(n19828), .B2(n13877), .ZN(
        n13881) );
  OAI22_X1 U17331 ( .A1(n19821), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13878), .B2(n14405), .ZN(n13879) );
  AOI21_X1 U17332 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19823), .A(
        n13879), .ZN(n13880) );
  OAI211_X1 U17333 ( .C1(n13882), .C2(n19825), .A(n13881), .B(n13880), .ZN(
        n13883) );
  AOI21_X1 U17334 ( .B1(n9648), .B2(n13956), .A(n13883), .ZN(n13884) );
  OAI21_X1 U17335 ( .B1(n13885), .B2(n13959), .A(n13884), .ZN(P1_U2839) );
  OR2_X1 U17336 ( .A1(n13888), .A2(n13887), .ZN(n13889) );
  NAND2_X1 U17337 ( .A1(n13886), .A2(n13889), .ZN(n18725) );
  INV_X1 U17338 ( .A(n18725), .ZN(n13895) );
  NOR2_X1 U17339 ( .A1(n14840), .A2(n10515), .ZN(n13894) );
  AND2_X1 U17340 ( .A1(n13611), .A2(n13890), .ZN(n13937) );
  AOI211_X1 U17341 ( .C1(n13892), .C2(n13891), .A(n14880), .B(n13937), .ZN(
        n13893) );
  AOI211_X1 U17342 ( .C1(n13895), .C2(n14840), .A(n13894), .B(n13893), .ZN(
        n13896) );
  INV_X1 U17343 ( .A(n13896), .ZN(P2_U2872) );
  NAND2_X1 U17344 ( .A1(n13898), .A2(n13897), .ZN(n13899) );
  XNOR2_X1 U17345 ( .A(n13899), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19053) );
  INV_X1 U17346 ( .A(n19053), .ZN(n13911) );
  NAND2_X1 U17347 ( .A1(n13994), .A2(n13900), .ZN(n13903) );
  INV_X1 U17348 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19612) );
  NOR2_X1 U17349 ( .A1(n19612), .A2(n14056), .ZN(n13901) );
  AOI21_X1 U17350 ( .B1(n15354), .B2(n18843), .A(n13901), .ZN(n13902) );
  OAI211_X1 U17351 ( .C1(n19056), .C2(n16008), .A(n13903), .B(n13902), .ZN(
        n13904) );
  AOI21_X1 U17352 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13905), .A(
        n13904), .ZN(n13910) );
  INV_X1 U17353 ( .A(n13907), .ZN(n13908) );
  XNOR2_X1 U17354 ( .A(n13906), .B(n13908), .ZN(n19051) );
  NAND2_X1 U17355 ( .A1(n19051), .A2(n16044), .ZN(n13909) );
  OAI211_X1 U17356 ( .C1(n13911), .C2(n16040), .A(n13910), .B(n13909), .ZN(
        P2_U3042) );
  INV_X1 U17357 ( .A(n13914), .ZN(n13912) );
  NOR3_X1 U17358 ( .A1(n13915), .A2(n10236), .A3(n13912), .ZN(n13917) );
  AOI21_X1 U17359 ( .B1(n13915), .B2(n13914), .A(n13913), .ZN(n13916) );
  OAI222_X1 U17360 ( .A1(n13919), .A2(n13918), .B1(n14217), .B2(n15398), .C1(
        n13917), .C2(n13916), .ZN(n16052) );
  AOI222_X1 U17361 ( .A1(n16052), .A2(n19669), .B1(n15407), .B2(n13920), .C1(
        n19171), .C2(n16049), .ZN(n13921) );
  INV_X1 U17362 ( .A(n15502), .ZN(n15504) );
  MUX2_X1 U17363 ( .A(n16054), .B(n13921), .S(n15504), .Z(n13922) );
  INV_X1 U17364 ( .A(n13922), .ZN(P2_U3599) );
  AOI21_X1 U17365 ( .B1(n19769), .B2(n19821), .A(n13923), .ZN(n13924) );
  AOI21_X1 U17366 ( .B1(n19797), .B2(P1_EBX_REG_0__SCAN_IN), .A(n13924), .ZN(
        n13928) );
  NAND2_X1 U17367 ( .A1(n19789), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13927) );
  NAND2_X1 U17368 ( .A1(n19828), .A2(n13925), .ZN(n13926) );
  NAND3_X1 U17369 ( .A1(n13928), .A2(n13927), .A3(n13926), .ZN(n13931) );
  NOR2_X1 U17370 ( .A1(n13929), .A2(n13959), .ZN(n13930) );
  AOI211_X1 U17371 ( .C1(n13956), .C2(n11614), .A(n13931), .B(n13930), .ZN(
        n13932) );
  INV_X1 U17372 ( .A(n13932), .ZN(P1_U2840) );
  INV_X1 U17373 ( .A(n13933), .ZN(n13934) );
  AOI21_X1 U17374 ( .B1(n13935), .B2(n13886), .A(n13934), .ZN(n18716) );
  INV_X1 U17375 ( .A(n18716), .ZN(n15307) );
  OR2_X1 U17376 ( .A1(n13937), .A2(n13936), .ZN(n13939) );
  NAND2_X1 U17377 ( .A1(n13611), .A2(n13938), .ZN(n13962) );
  AND2_X1 U17378 ( .A1(n13939), .A2(n13962), .ZN(n18886) );
  NAND2_X1 U17379 ( .A1(n18886), .A2(n14870), .ZN(n13941) );
  NAND2_X1 U17380 ( .A1(n14873), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13940) );
  OAI211_X1 U17381 ( .C1(n15307), .C2(n14873), .A(n13941), .B(n13940), .ZN(
        P2_U2871) );
  AND2_X1 U17382 ( .A1(n13769), .A2(n13943), .ZN(n13944) );
  NOR2_X1 U17383 ( .A1(n13942), .A2(n13944), .ZN(n19838) );
  INV_X1 U17384 ( .A(n19838), .ZN(n13948) );
  INV_X1 U17385 ( .A(DATAI_9_), .ZN(n13946) );
  NAND2_X1 U17386 ( .A1(n19957), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13945) );
  OAI21_X1 U17387 ( .B1(n19957), .B2(n13946), .A(n13945), .ZN(n19879) );
  AOI22_X1 U17388 ( .A1(n14078), .A2(n19879), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14506), .ZN(n13947) );
  OAI21_X1 U17389 ( .B1(n13948), .B2(n14493), .A(n13947), .ZN(P1_U2895) );
  NOR2_X1 U17390 ( .A1(n15677), .A2(n13878), .ZN(n13949) );
  OAI21_X1 U17391 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(n13949), .A(n13972), .ZN(
        n13958) );
  INV_X1 U17392 ( .A(n13417), .ZN(n19968) );
  NOR2_X1 U17393 ( .A1(n19793), .A2(n19944), .ZN(n13955) );
  INV_X1 U17394 ( .A(n13950), .ZN(n13951) );
  AOI22_X1 U17395 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19823), .B1(
        n19766), .B2(n13951), .ZN(n13952) );
  OAI21_X1 U17396 ( .B1(n19825), .B2(n13953), .A(n13952), .ZN(n13954) );
  AOI211_X1 U17397 ( .C1(n19968), .C2(n13956), .A(n13955), .B(n13954), .ZN(
        n13957) );
  OAI211_X1 U17398 ( .C1(n13960), .C2(n13959), .A(n13958), .B(n13957), .ZN(
        P1_U2838) );
  INV_X1 U17399 ( .A(n14020), .ZN(n13961) );
  AOI21_X1 U17400 ( .B1(n13963), .B2(n13962), .A(n13961), .ZN(n14031) );
  NAND2_X1 U17401 ( .A1(n14031), .A2(n14870), .ZN(n13965) );
  NAND2_X1 U17402 ( .A1(n14873), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13964) );
  OAI211_X1 U17403 ( .C1(n13966), .C2(n14873), .A(n13965), .B(n13964), .ZN(
        P2_U2870) );
  INV_X1 U17404 ( .A(n13968), .ZN(n13969) );
  OAI21_X1 U17405 ( .B1(n13942), .B2(n13970), .A(n13969), .ZN(n14658) );
  NOR2_X1 U17406 ( .A1(n13973), .A2(n13971), .ZN(n19815) );
  INV_X1 U17407 ( .A(n19815), .ZN(n19798) );
  NOR2_X1 U17408 ( .A1(n19764), .A2(n19798), .ZN(n19771) );
  AOI21_X1 U17409 ( .B1(n15623), .B2(n13973), .A(n13972), .ZN(n19835) );
  OAI21_X1 U17410 ( .B1(n13975), .B2(n13974), .A(n19835), .ZN(n15696) );
  OAI221_X1 U17411 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n19771), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(P1_REIP_REG_9__SCAN_IN), .A(n15696), 
        .ZN(n13983) );
  AND2_X1 U17412 ( .A1(n15840), .A2(n13976), .ZN(n13977) );
  OR2_X1 U17413 ( .A1(n13977), .A2(n14081), .ZN(n15831) );
  INV_X1 U17414 ( .A(n13978), .ZN(n14655) );
  AOI22_X1 U17415 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n19797), .B1(n14655), 
        .B2(n19766), .ZN(n13979) );
  OAI21_X1 U17416 ( .B1(n19793), .B2(n15831), .A(n13979), .ZN(n13981) );
  NAND2_X1 U17417 ( .A1(n14405), .A2(n13980), .ZN(n19820) );
  AOI211_X1 U17418 ( .C1(n19823), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n13981), .B(n19775), .ZN(n13982) );
  OAI211_X1 U17419 ( .C1(n14658), .C2(n15655), .A(n13983), .B(n13982), .ZN(
        P1_U2830) );
  INV_X1 U17420 ( .A(DATAI_10_), .ZN(n13985) );
  NAND2_X1 U17421 ( .A1(n19957), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13984) );
  OAI21_X1 U17422 ( .B1(n19957), .B2(n13985), .A(n13984), .ZN(n19881) );
  INV_X1 U17423 ( .A(n19881), .ZN(n13987) );
  OAI222_X1 U17424 ( .A1(n14658), .A2(n14493), .B1(n14137), .B2(n13987), .C1(
        n13986), .C2(n14482), .ZN(P1_U2894) );
  XNOR2_X1 U17425 ( .A(n13988), .B(n9622), .ZN(n14014) );
  NAND2_X1 U17426 ( .A1(n13992), .A2(n13991), .ZN(n13993) );
  XNOR2_X1 U17427 ( .A(n13990), .B(n13993), .ZN(n14011) );
  AOI21_X1 U17428 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13994), .A(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13999) );
  XNOR2_X1 U17429 ( .A(n13996), .B(n13995), .ZN(n18919) );
  NAND2_X1 U17430 ( .A1(n15127), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n14008) );
  OAI21_X1 U17431 ( .B1(n16036), .B2(n18919), .A(n14008), .ZN(n13997) );
  AOI21_X1 U17432 ( .B1(n18836), .B2(n16038), .A(n13997), .ZN(n13998) );
  OAI21_X1 U17433 ( .B1(n14061), .B2(n13999), .A(n13998), .ZN(n14000) );
  AOI21_X1 U17434 ( .B1(n14011), .B2(n10731), .A(n14000), .ZN(n14001) );
  OAI21_X1 U17435 ( .B1(n14014), .B2(n16034), .A(n14001), .ZN(P2_U3041) );
  XOR2_X1 U17436 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14003), .Z(
        n14004) );
  XNOR2_X1 U17437 ( .A(n14002), .B(n14004), .ZN(n15856) );
  AOI22_X1 U17438 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14005) );
  OAI21_X1 U17439 ( .B1(n19916), .B2(n19777), .A(n14005), .ZN(n14006) );
  AOI21_X1 U17440 ( .B1(n19784), .B2(n19911), .A(n14006), .ZN(n14007) );
  OAI21_X1 U17441 ( .B1(n15856), .B2(n19746), .A(n14007), .ZN(P1_U2991) );
  INV_X1 U17442 ( .A(n14008), .ZN(n14010) );
  INV_X1 U17443 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20756) );
  OAI22_X1 U17444 ( .A1(n19061), .A2(n20756), .B1(n15144), .B2(n18834), .ZN(
        n14009) );
  AOI211_X1 U17445 ( .C1(n18836), .C2(n16001), .A(n14010), .B(n14009), .ZN(
        n14013) );
  NAND2_X1 U17446 ( .A1(n14011), .A2(n19052), .ZN(n14012) );
  OAI211_X1 U17447 ( .C1(n14014), .C2(n15995), .A(n14013), .B(n14012), .ZN(
        P2_U3009) );
  INV_X1 U17448 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14015) );
  OAI222_X1 U17449 ( .A1(n15831), .A2(n14465), .B1(n19851), .B2(n14015), .C1(
        n14463), .C2(n14658), .ZN(P1_U2862) );
  NOR2_X1 U17450 ( .A1(n12478), .A2(n14016), .ZN(n14017) );
  OR2_X1 U17451 ( .A1(n14089), .A2(n14017), .ZN(n18698) );
  AND2_X1 U17452 ( .A1(n14020), .A2(n14019), .ZN(n14021) );
  NOR2_X1 U17453 ( .A1(n14018), .A2(n14021), .ZN(n15970) );
  NAND2_X1 U17454 ( .A1(n15970), .A2(n14870), .ZN(n14023) );
  NAND2_X1 U17455 ( .A1(n14873), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14022) );
  OAI211_X1 U17456 ( .C1(n18698), .C2(n14873), .A(n14023), .B(n14022), .ZN(
        P2_U2869) );
  MUX2_X1 U17457 ( .A(n14025), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n15735), .Z(n14026) );
  XNOR2_X1 U17458 ( .A(n14024), .B(n14026), .ZN(n15836) );
  AOI22_X1 U17459 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14027) );
  OAI21_X1 U17460 ( .B1(n19916), .B2(n14028), .A(n14027), .ZN(n14029) );
  AOI21_X1 U17461 ( .B1(n19838), .B2(n19911), .A(n14029), .ZN(n14030) );
  OAI21_X1 U17462 ( .B1(n15836), .B2(n19746), .A(n14030), .ZN(P1_U2990) );
  INV_X1 U17463 ( .A(n14031), .ZN(n14038) );
  INV_X1 U17464 ( .A(n18709), .ZN(n14036) );
  INV_X1 U17465 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n18974) );
  OAI22_X1 U17466 ( .A1(n14928), .A2(n19026), .B1(n18922), .B2(n18974), .ZN(
        n14035) );
  INV_X1 U17467 ( .A(n18884), .ZN(n14932) );
  INV_X1 U17468 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14033) );
  INV_X1 U17469 ( .A(n18883), .ZN(n14930) );
  INV_X1 U17470 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14032) );
  OAI22_X1 U17471 ( .A1(n14932), .A2(n14033), .B1(n14930), .B2(n14032), .ZN(
        n14034) );
  AOI211_X1 U17472 ( .C1(n18932), .C2(n14036), .A(n14035), .B(n14034), .ZN(
        n14037) );
  OAI21_X1 U17473 ( .B1(n14038), .B2(n18936), .A(n14037), .ZN(P2_U2902) );
  NOR2_X1 U17474 ( .A1(n19317), .A2(n19131), .ZN(n19124) );
  AOI21_X1 U17475 ( .B1(n14044), .B2(n19697), .A(n19124), .ZN(n14042) );
  NOR2_X1 U17476 ( .A1(n19322), .A2(n19131), .ZN(n14040) );
  AOI221_X1 U17477 ( .B1(n19126), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19157), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n14040), .ZN(n14041) );
  MUX2_X1 U17478 ( .A(n14042), .B(n14041), .S(n19681), .Z(n14043) );
  INV_X1 U17479 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14048) );
  AOI22_X1 U17480 ( .A1(n19157), .A2(n19518), .B1(n19126), .B2(n19323), .ZN(
        n14047) );
  OAI21_X1 U17481 ( .B1(n14044), .B2(n19124), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14045) );
  OAI21_X1 U17482 ( .B1(n19131), .B2(n19322), .A(n14045), .ZN(n19125) );
  AOI22_X1 U17483 ( .A1(n19125), .A2(n19462), .B1(n19451), .B2(n19124), .ZN(
        n14046) );
  OAI211_X1 U17484 ( .C1(n19130), .C2(n14048), .A(n14047), .B(n14046), .ZN(
        P2_U3064) );
  OAI21_X1 U17485 ( .B1(n14050), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14049), .ZN(n16000) );
  XOR2_X1 U17486 ( .A(n14052), .B(n14051), .Z(n16002) );
  XNOR2_X1 U17487 ( .A(n14054), .B(n14053), .ZN(n18912) );
  NOR2_X1 U17488 ( .A1(n16036), .A2(n18912), .ZN(n14058) );
  INV_X1 U17489 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19616) );
  OAI22_X1 U17490 ( .A1(n14056), .A2(n19616), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14055), .ZN(n14057) );
  AOI211_X1 U17491 ( .C1(n9716), .C2(n16038), .A(n14058), .B(n14057), .ZN(
        n14059) );
  OAI21_X1 U17492 ( .B1(n14061), .B2(n14060), .A(n14059), .ZN(n14062) );
  AOI21_X1 U17493 ( .B1(n16002), .B2(n16044), .A(n14062), .ZN(n14063) );
  OAI21_X1 U17494 ( .B1(n16040), .B2(n16000), .A(n14063), .ZN(P2_U3040) );
  OAI21_X1 U17495 ( .B1(n13968), .B2(n14065), .A(n14064), .ZN(n14094) );
  XNOR2_X1 U17496 ( .A(n14094), .B(n14092), .ZN(n15740) );
  INV_X1 U17497 ( .A(n15740), .ZN(n14083) );
  INV_X1 U17498 ( .A(DATAI_11_), .ZN(n14067) );
  NAND2_X1 U17499 ( .A1(n19957), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14066) );
  OAI21_X1 U17500 ( .B1(n19957), .B2(n14067), .A(n14066), .ZN(n19883) );
  INV_X1 U17501 ( .A(n19883), .ZN(n14069) );
  OAI222_X1 U17502 ( .A1(n14083), .A2(n14493), .B1(n14137), .B2(n14069), .C1(
        n14068), .C2(n14482), .ZN(P1_U2893) );
  NAND2_X1 U17503 ( .A1(n14072), .A2(n14073), .ZN(n14074) );
  NAND2_X1 U17504 ( .A1(n14070), .A2(n14074), .ZN(n15674) );
  XNOR2_X1 U17505 ( .A(n14105), .B(n14120), .ZN(n15804) );
  AOI22_X1 U17506 ( .A1(n15804), .A2(n19846), .B1(n14446), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14075) );
  OAI21_X1 U17507 ( .B1(n15674), .B2(n14463), .A(n14075), .ZN(P1_U2858) );
  INV_X1 U17508 ( .A(DATAI_14_), .ZN(n14077) );
  NAND2_X1 U17509 ( .A1(n19957), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14076) );
  OAI21_X1 U17510 ( .B1(n19957), .B2(n14077), .A(n14076), .ZN(n19889) );
  AOI22_X1 U17511 ( .A1(n14078), .A2(n19889), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14506), .ZN(n14079) );
  OAI21_X1 U17512 ( .B1(n15674), .B2(n14493), .A(n14079), .ZN(P1_U2890) );
  NOR2_X1 U17513 ( .A1(n14081), .A2(n14080), .ZN(n14082) );
  OR2_X1 U17514 ( .A1(n14125), .A2(n14082), .ZN(n15822) );
  INV_X1 U17515 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15692) );
  OAI222_X1 U17516 ( .A1(n15822), .A2(n14465), .B1(n15692), .B2(n19851), .C1(
        n14463), .C2(n14083), .ZN(P1_U2861) );
  INV_X1 U17517 ( .A(n14084), .ZN(n14085) );
  OAI21_X1 U17518 ( .B1(n14018), .B2(n14086), .A(n14085), .ZN(n14147) );
  OAI21_X1 U17519 ( .B1(n14089), .B2(n14088), .A(n14087), .ZN(n15053) );
  NOR2_X1 U17520 ( .A1(n15053), .A2(n14873), .ZN(n14090) );
  AOI21_X1 U17521 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14873), .A(n14090), .ZN(
        n14091) );
  OAI21_X1 U17522 ( .B1(n14147), .B2(n14880), .A(n14091), .ZN(P2_U2868) );
  INV_X1 U17523 ( .A(n14092), .ZN(n14093) );
  OAI21_X1 U17524 ( .B1(n14094), .B2(n14093), .A(n14064), .ZN(n14096) );
  INV_X1 U17525 ( .A(n14096), .ZN(n14098) );
  INV_X1 U17526 ( .A(n14095), .ZN(n14097) );
  AND2_X1 U17527 ( .A1(n14096), .A2(n14095), .ZN(n14104) );
  AOI21_X1 U17528 ( .B1(n14098), .B2(n14097), .A(n14104), .ZN(n15729) );
  INV_X1 U17529 ( .A(n15729), .ZN(n14128) );
  INV_X1 U17530 ( .A(DATAI_12_), .ZN(n14100) );
  NAND2_X1 U17531 ( .A1(n19957), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14099) );
  OAI21_X1 U17532 ( .B1(n19957), .B2(n14100), .A(n14099), .ZN(n19885) );
  INV_X1 U17533 ( .A(n19885), .ZN(n14102) );
  OAI222_X1 U17534 ( .A1(n14128), .A2(n14493), .B1(n14137), .B2(n14102), .C1(
        n14101), .C2(n14482), .ZN(P1_U2892) );
  OAI21_X1 U17535 ( .B1(n14104), .B2(n14103), .A(n14072), .ZN(n14647) );
  INV_X1 U17536 ( .A(n14105), .ZN(n14121) );
  AOI21_X1 U17537 ( .B1(n14106), .B2(n14127), .A(n14121), .ZN(n15815) );
  AOI22_X1 U17538 ( .A1(n15815), .A2(n19828), .B1(n19797), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14107) );
  OAI211_X1 U17539 ( .C1(n19769), .C2(n14108), .A(n14107), .B(n19820), .ZN(
        n14113) );
  NAND3_X1 U17540 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n19771), .ZN(n15699) );
  NOR2_X1 U17541 ( .A1(n14109), .A2(n15699), .ZN(n14111) );
  AOI21_X1 U17542 ( .B1(n15623), .B2(n14109), .A(n15696), .ZN(n15691) );
  INV_X1 U17543 ( .A(n15691), .ZN(n14110) );
  MUX2_X1 U17544 ( .A(n14111), .B(n14110), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14112) );
  AOI211_X1 U17545 ( .C1(n14644), .C2(n19766), .A(n14113), .B(n14112), .ZN(
        n14114) );
  OAI21_X1 U17546 ( .B1(n14647), .B2(n15655), .A(n14114), .ZN(P1_U2827) );
  AOI22_X1 U17547 ( .A1(n15815), .A2(n19846), .B1(n14446), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14115) );
  OAI21_X1 U17548 ( .B1(n14647), .B2(n14463), .A(n14115), .ZN(P1_U2859) );
  INV_X1 U17549 ( .A(n14116), .ZN(n14117) );
  AOI21_X1 U17550 ( .B1(n14118), .B2(n14070), .A(n14117), .ZN(n15726) );
  INV_X1 U17551 ( .A(n15726), .ZN(n14132) );
  AOI21_X1 U17552 ( .B1(n14121), .B2(n14120), .A(n14119), .ZN(n14122) );
  NOR2_X1 U17553 ( .A1(n14122), .A2(n14154), .ZN(n15795) );
  AOI22_X1 U17554 ( .A1(n15795), .A2(n19846), .B1(n14446), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14123) );
  OAI21_X1 U17555 ( .B1(n14132), .B2(n14463), .A(n14123), .ZN(P1_U2857) );
  OR2_X1 U17556 ( .A1(n14125), .A2(n14124), .ZN(n14126) );
  NAND2_X1 U17557 ( .A1(n14127), .A2(n14126), .ZN(n15685) );
  INV_X1 U17558 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14129) );
  OAI222_X1 U17559 ( .A1(n15685), .A2(n14465), .B1(n14129), .B2(n19851), .C1(
        n14128), .C2(n14463), .ZN(P1_U2860) );
  OAI222_X1 U17560 ( .A1(n14132), .A2(n14493), .B1(n14137), .B2(n14131), .C1(
        n14482), .C2(n14130), .ZN(P1_U2889) );
  INV_X1 U17561 ( .A(DATAI_13_), .ZN(n14134) );
  NAND2_X1 U17562 ( .A1(n19957), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14133) );
  OAI21_X1 U17563 ( .B1(n19957), .B2(n14134), .A(n14133), .ZN(n19887) );
  INV_X1 U17564 ( .A(n19887), .ZN(n14136) );
  OAI222_X1 U17565 ( .A1(n14647), .A2(n14493), .B1(n14137), .B2(n14136), .C1(
        n14135), .C2(n14482), .ZN(P1_U2891) );
  INV_X1 U17566 ( .A(n14138), .ZN(n15256) );
  NAND2_X1 U17567 ( .A1(n15283), .A2(n14139), .ZN(n14140) );
  NAND2_X1 U17568 ( .A1(n15256), .A2(n14140), .ZN(n18689) );
  INV_X1 U17569 ( .A(n18689), .ZN(n14145) );
  INV_X1 U17570 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n18970) );
  OAI22_X1 U17571 ( .A1(n14928), .A2(n19030), .B1(n18922), .B2(n18970), .ZN(
        n14144) );
  INV_X1 U17572 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14142) );
  INV_X1 U17573 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14141) );
  OAI22_X1 U17574 ( .A1(n14932), .A2(n14142), .B1(n14930), .B2(n14141), .ZN(
        n14143) );
  AOI211_X1 U17575 ( .C1(n18932), .C2(n14145), .A(n14144), .B(n14143), .ZN(
        n14146) );
  OAI21_X1 U17576 ( .B1(n14147), .B2(n18936), .A(n14146), .ZN(P2_U2900) );
  AOI21_X1 U17577 ( .B1(n14149), .B2(n14116), .A(n14148), .ZN(n14150) );
  INV_X1 U17578 ( .A(n14150), .ZN(n14622) );
  INV_X1 U17579 ( .A(n14151), .ZN(n14152) );
  OAI21_X1 U17580 ( .B1(n14154), .B2(n14153), .A(n14152), .ZN(n14164) );
  INV_X1 U17581 ( .A(n14164), .ZN(n15789) );
  AOI22_X1 U17582 ( .A1(n15789), .A2(n19846), .B1(n14446), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14155) );
  OAI21_X1 U17583 ( .B1(n14622), .B2(n14463), .A(n14155), .ZN(P1_U2856) );
  AOI22_X1 U17584 ( .A1(n14507), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14506), .ZN(n14159) );
  AND2_X1 U17585 ( .A1(n14482), .A2(n14156), .ZN(n14509) );
  AOI22_X1 U17586 ( .A1(n14510), .A2(DATAI_16_), .B1(n14509), .B2(n14157), 
        .ZN(n14158) );
  OAI211_X1 U17587 ( .C1(n14622), .C2(n14493), .A(n14159), .B(n14158), .ZN(
        P1_U2888) );
  INV_X1 U17588 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15670) );
  NAND2_X1 U17589 ( .A1(n15623), .A2(n14167), .ZN(n15639) );
  NOR2_X1 U17590 ( .A1(n15670), .A2(n15639), .ZN(n15658) );
  INV_X1 U17591 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14166) );
  AOI21_X1 U17592 ( .B1(n19823), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19775), .ZN(n14160) );
  OAI21_X1 U17593 ( .B1(n19825), .B2(n14161), .A(n14160), .ZN(n14162) );
  AOI21_X1 U17594 ( .B1(n14619), .B2(n19766), .A(n14162), .ZN(n14163) );
  OAI21_X1 U17595 ( .B1(n14164), .B2(n19793), .A(n14163), .ZN(n14165) );
  AOI21_X1 U17596 ( .B1(n15658), .B2(n14166), .A(n14165), .ZN(n14169) );
  NOR2_X1 U17597 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15639), .ZN(n15665) );
  OAI21_X1 U17598 ( .B1(n15677), .B2(n14167), .A(n14405), .ZN(n15679) );
  OAI21_X1 U17599 ( .B1(n15665), .B2(n15679), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14168) );
  OAI211_X1 U17600 ( .C1(n14622), .C2(n15655), .A(n14169), .B(n14168), .ZN(
        P1_U2824) );
  INV_X1 U17601 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16386) );
  INV_X1 U17602 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16409) );
  INV_X1 U17603 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16730) );
  NOR3_X1 U17604 ( .A1(n16386), .A2(n16409), .A3(n16730), .ZN(n14170) );
  NAND3_X1 U17605 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n14170), .ZN(n15410) );
  NAND2_X1 U17606 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n15411) );
  INV_X1 U17607 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16911) );
  INV_X1 U17608 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16931) );
  NOR2_X1 U17609 ( .A1(n15510), .A2(n17077), .ZN(n14172) );
  NAND3_X1 U17610 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16974) );
  NOR3_X1 U17611 ( .A1(n20743), .A2(n16968), .A3(n16974), .ZN(n16954) );
  NAND2_X1 U17612 ( .A1(n16990), .A2(n16954), .ZN(n16964) );
  NAND3_X1 U17613 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(n16959), .ZN(n16956) );
  NOR3_X2 U17614 ( .A1(n16534), .A2(n16911), .A3(n16929), .ZN(n16884) );
  NAND4_X1 U17615 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .A4(n16884), .ZN(n16835) );
  NAND4_X1 U17616 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .A4(n16811), .ZN(n16794) );
  NAND4_X1 U17617 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(P3_EBX_REG_20__SCAN_IN), .A4(n16783), .ZN(n14174) );
  NOR3_X1 U17618 ( .A1(n15410), .A2(n15411), .A3(n14174), .ZN(n16695) );
  NAND2_X1 U17619 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16695), .ZN(n14175) );
  NOR2_X1 U17620 ( .A1(n17077), .A2(n14175), .ZN(n14177) );
  NAND2_X1 U17621 ( .A1(n16972), .A2(n14175), .ZN(n16696) );
  INV_X1 U17622 ( .A(n16696), .ZN(n14176) );
  MUX2_X1 U17623 ( .A(n14177), .B(n14176), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  AOI21_X1 U17624 ( .B1(n18401), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15498) );
  NAND2_X1 U17625 ( .A1(n15498), .A2(n15453), .ZN(n17938) );
  NOR2_X1 U17626 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17938), .ZN(n14178) );
  NAND3_X1 U17627 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n18553)
         );
  OAI21_X1 U17628 ( .B1(n14178), .B2(n18553), .A(n18147), .ZN(n17948) );
  INV_X1 U17629 ( .A(n17948), .ZN(n14179) );
  NOR2_X1 U17630 ( .A1(n18602), .A2(n17512), .ZN(n17942) );
  AOI21_X1 U17631 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n17942), .ZN(n17943) );
  NOR2_X1 U17632 ( .A1(n14179), .A2(n17943), .ZN(n14181) );
  NOR2_X1 U17633 ( .A1(n18555), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17993) );
  OR2_X1 U17634 ( .A1(n17993), .A2(n14179), .ZN(n17941) );
  OR2_X1 U17635 ( .A1(n18191), .A2(n17941), .ZN(n14180) );
  MUX2_X1 U17636 ( .A(n14181), .B(n14180), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AOI21_X1 U17637 ( .B1(n13690), .B2(n20333), .A(n14182), .ZN(n14184) );
  AOI22_X1 U17638 ( .A1(n14185), .A2(n14184), .B1(n14183), .B2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n14186) );
  OAI21_X1 U17639 ( .B1(n13417), .B2(n14187), .A(n14186), .ZN(P1_U3476) );
  OAI21_X1 U17640 ( .B1(n14190), .B2(n14189), .A(n14188), .ZN(n14206) );
  NAND2_X1 U17641 ( .A1(n15127), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14205) );
  OAI21_X1 U17642 ( .B1(n15996), .B2(n14206), .A(n14205), .ZN(n14199) );
  INV_X1 U17643 ( .A(n14191), .ZN(n14192) );
  AOI21_X1 U17644 ( .B1(n14194), .B2(n14193), .A(n14192), .ZN(n14203) );
  INV_X1 U17645 ( .A(n14203), .ZN(n14197) );
  INV_X1 U17646 ( .A(n14195), .ZN(n14196) );
  OAI22_X1 U17647 ( .A1(n14197), .A2(n15995), .B1(n15144), .B2(n14196), .ZN(
        n14198) );
  AOI211_X1 U17648 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n15105), .A(
        n14199), .B(n14198), .ZN(n14200) );
  OAI21_X1 U17649 ( .B1(n14217), .B2(n19057), .A(n14200), .ZN(P2_U3012) );
  AOI22_X1 U17650 ( .A1(n16044), .A2(n14203), .B1(n14202), .B2(n14201), .ZN(
        n14216) );
  INV_X1 U17651 ( .A(n14204), .ZN(n14214) );
  OAI21_X1 U17652 ( .B1(n16040), .B2(n14206), .A(n14205), .ZN(n14213) );
  OAI21_X1 U17653 ( .B1(n14209), .B2(n14208), .A(n14207), .ZN(n14210) );
  OAI21_X1 U17654 ( .B1(n14211), .B2(n16036), .A(n14210), .ZN(n14212) );
  AOI211_X1 U17655 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n14214), .A(
        n14213), .B(n14212), .ZN(n14215) );
  OAI211_X1 U17656 ( .C1(n14217), .C2(n16008), .A(n14216), .B(n14215), .ZN(
        P2_U3044) );
  INV_X1 U17657 ( .A(n15140), .ZN(n14220) );
  NOR2_X1 U17658 ( .A1(n14220), .A2(n14219), .ZN(n14221) );
  XNOR2_X1 U17659 ( .A(n14218), .B(n14221), .ZN(n14241) );
  OR2_X1 U17660 ( .A1(n14222), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14236) );
  NAND2_X1 U17661 ( .A1(n14222), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15987) );
  NAND3_X1 U17662 ( .A1(n14236), .A2(n15987), .A3(n10731), .ZN(n14235) );
  OAI21_X1 U17663 ( .B1(n14225), .B2(n14224), .A(n13509), .ZN(n18815) );
  NOR2_X1 U17664 ( .A1(n10750), .A2(n14056), .ZN(n14231) );
  OR2_X1 U17665 ( .A1(n14227), .A2(n14226), .ZN(n14229) );
  NAND2_X1 U17666 ( .A1(n14229), .A2(n14228), .ZN(n18911) );
  NOR2_X1 U17667 ( .A1(n16036), .A2(n18911), .ZN(n14230) );
  AOI211_X1 U17668 ( .C1(n16024), .C2(n16021), .A(n14231), .B(n14230), .ZN(
        n14232) );
  OAI21_X1 U17669 ( .B1(n18815), .B2(n16008), .A(n14232), .ZN(n14233) );
  AOI21_X1 U17670 ( .B1(n16025), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n14233), .ZN(n14234) );
  OAI211_X1 U17671 ( .C1(n14241), .C2(n16034), .A(n14235), .B(n14234), .ZN(
        P2_U3039) );
  NAND3_X1 U17672 ( .A1(n14236), .A2(n15987), .A3(n19052), .ZN(n14240) );
  OAI22_X1 U17673 ( .A1(n19061), .A2(n9802), .B1(n15144), .B2(n18812), .ZN(
        n14238) );
  NOR2_X1 U17674 ( .A1(n18815), .A2(n19057), .ZN(n14237) );
  AOI211_X1 U17675 ( .C1(n15392), .C2(P2_REIP_REG_7__SCAN_IN), .A(n14238), .B(
        n14237), .ZN(n14239) );
  OAI211_X1 U17676 ( .C1(n14241), .C2(n15995), .A(n14240), .B(n14239), .ZN(
        P2_U3007) );
  AOI22_X1 U17677 ( .A1(n14507), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14506), .ZN(n14243) );
  AOI22_X1 U17678 ( .A1(n14510), .A2(DATAI_30_), .B1(n14509), .B2(n19889), 
        .ZN(n14242) );
  OAI211_X1 U17679 ( .C1(n14250), .C2(n14493), .A(n14243), .B(n14242), .ZN(
        P1_U2874) );
  INV_X1 U17680 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14526) );
  INV_X1 U17681 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14244) );
  OAI21_X1 U17682 ( .B1(n14315), .B2(n14526), .A(n14244), .ZN(n14248) );
  AOI22_X1 U17683 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19823), .B1(
        n19766), .B2(n14517), .ZN(n14245) );
  OAI21_X1 U17684 ( .B1(n19825), .B2(n14246), .A(n14245), .ZN(n14247) );
  NAND2_X1 U17685 ( .A1(n15735), .A2(n14698), .ZN(n14252) );
  NAND2_X1 U17686 ( .A1(n14251), .A2(n14252), .ZN(n14256) );
  NAND2_X1 U17687 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14253) );
  NOR2_X1 U17688 ( .A1(n14256), .A2(n14253), .ZN(n14258) );
  NOR4_X1 U17689 ( .A1(n14254), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14255) );
  AND2_X1 U17690 ( .A1(n14256), .A2(n14255), .ZN(n14257) );
  MUX2_X1 U17691 ( .A(n14258), .B(n14257), .S(n15702), .Z(n14259) );
  XNOR2_X1 U17692 ( .A(n14259), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14686) );
  NAND2_X1 U17693 ( .A1(n12105), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14680) );
  OAI21_X1 U17694 ( .B1(n14653), .B2(n14260), .A(n14680), .ZN(n14264) );
  OR2_X1 U17695 ( .A1(n14336), .A2(n14261), .ZN(n14262) );
  NAND2_X2 U17696 ( .A1(n14309), .A2(n14262), .ZN(n14471) );
  NOR2_X1 U17697 ( .A1(n14471), .A2(n19960), .ZN(n14263) );
  OAI21_X1 U17698 ( .B1(n19746), .B2(n14686), .A(n14265), .ZN(P1_U2971) );
  NAND2_X1 U17699 ( .A1(n14873), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14266) );
  OAI21_X1 U17700 ( .B1(n14271), .B2(n14873), .A(n14266), .ZN(P2_U2856) );
  NAND2_X1 U17701 ( .A1(n15105), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14267) );
  OAI211_X1 U17702 ( .C1(n15144), .C2(n14269), .A(n14268), .B(n14267), .ZN(
        n14270) );
  NAND2_X1 U17703 ( .A1(n14273), .A2(n19052), .ZN(n14274) );
  XNOR2_X1 U17704 ( .A(n13649), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14276) );
  MUX2_X1 U17705 ( .A(n10479), .B(n18815), .S(n14840), .Z(n14275) );
  OAI21_X1 U17706 ( .B1(n14276), .B2(n14880), .A(n14275), .ZN(P2_U2880) );
  NOR2_X1 U17707 ( .A1(n14277), .A2(n14873), .ZN(n14278) );
  AOI21_X1 U17708 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14873), .A(n14278), .ZN(
        n14279) );
  OAI21_X1 U17709 ( .B1(n14280), .B2(n14880), .A(n14279), .ZN(P2_U2857) );
  NAND2_X1 U17710 ( .A1(n14281), .A2(n18890), .ZN(n14291) );
  OR2_X1 U17711 ( .A1(n14881), .A2(n14282), .ZN(n14283) );
  NAND2_X1 U17712 ( .A1(n14284), .A2(n14283), .ZN(n15910) );
  INV_X1 U17713 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14285) );
  OR2_X1 U17714 ( .A1(n18891), .A2(n14285), .ZN(n14287) );
  NAND2_X1 U17715 ( .A1(n18891), .A2(BUF2_REG_13__SCAN_IN), .ZN(n14286) );
  AND2_X1 U17716 ( .A1(n14287), .A2(n14286), .ZN(n19042) );
  INV_X1 U17717 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n18950) );
  OAI22_X1 U17718 ( .A1(n14928), .A2(n19042), .B1(n18922), .B2(n18950), .ZN(
        n14288) );
  AOI21_X1 U17719 ( .B1(n15155), .B2(n18932), .A(n14288), .ZN(n14290) );
  AOI22_X1 U17720 ( .A1(n18884), .A2(BUF2_REG_29__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14289) );
  OAI211_X1 U17721 ( .C1(n12928), .C2(n14291), .A(n14290), .B(n14289), .ZN(
        P2_U2890) );
  NAND2_X1 U17722 ( .A1(n14292), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14294)
         );
  NAND3_X1 U17723 ( .A1(n14294), .A2(n14293), .A3(n19743), .ZN(P1_U2801) );
  MUX2_X1 U17724 ( .A(n14296), .B(n14295), .S(n14301), .Z(n14299) );
  NAND2_X1 U17725 ( .A1(n12492), .A2(n14297), .ZN(n14298) );
  OAI211_X1 U17726 ( .C1(n14301), .C2(n14300), .A(n14299), .B(n14298), .ZN(
        n15567) );
  OAI22_X1 U17727 ( .A1(n14303), .A2(n12494), .B1(n14302), .B2(n14301), .ZN(
        n19741) );
  NAND3_X1 U17728 ( .A1(n14305), .A2(n14304), .A3(n12520), .ZN(n14306) );
  AND2_X1 U17729 ( .A1(n14306), .A2(n20647), .ZN(n20638) );
  OR2_X1 U17730 ( .A1(n19741), .A2(n20638), .ZN(n15565) );
  AND2_X1 U17731 ( .A1(n15565), .A2(n14307), .ZN(n19748) );
  MUX2_X1 U17732 ( .A(P1_MORE_REG_SCAN_IN), .B(n15567), .S(n19748), .Z(
        P1_U3484) );
  AOI21_X1 U17733 ( .B1(n14310), .B2(n14309), .A(n14308), .ZN(n14530) );
  INV_X1 U17734 ( .A(n14530), .ZN(n14468) );
  INV_X1 U17735 ( .A(n14311), .ZN(n14324) );
  OAI22_X1 U17736 ( .A1(n14312), .A2(n19769), .B1(n19821), .B2(n14528), .ZN(
        n14313) );
  AOI21_X1 U17737 ( .B1(n19797), .B2(P1_EBX_REG_29__SCAN_IN), .A(n14313), .ZN(
        n14314) );
  OAI21_X1 U17738 ( .B1(n14315), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14314), 
        .ZN(n14320) );
  AND2_X1 U17739 ( .A1(n14322), .A2(n14316), .ZN(n14317) );
  NOR2_X1 U17740 ( .A1(n14674), .A2(n19793), .ZN(n14319) );
  AOI211_X1 U17741 ( .C1(n14324), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14320), 
        .B(n14319), .ZN(n14321) );
  OAI21_X1 U17742 ( .B1(n14468), .B2(n15655), .A(n14321), .ZN(P1_U2811) );
  OAI21_X1 U17743 ( .B1(n14334), .B2(n14323), .A(n14322), .ZN(n14421) );
  INV_X1 U17744 ( .A(n14421), .ZN(n14684) );
  INV_X1 U17745 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14422) );
  INV_X1 U17746 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20604) );
  NOR3_X1 U17747 ( .A1(n15677), .A2(n20604), .A3(n14340), .ZN(n14325) );
  OAI21_X1 U17748 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14325), .A(n14324), 
        .ZN(n14328) );
  AOI22_X1 U17749 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19823), .B1(
        n19766), .B2(n14326), .ZN(n14327) );
  OAI211_X1 U17750 ( .C1(n14422), .C2(n19825), .A(n14328), .B(n14327), .ZN(
        n14329) );
  AOI21_X1 U17751 ( .B1(n14684), .B2(n19828), .A(n14329), .ZN(n14330) );
  OAI21_X1 U17752 ( .B1(n14471), .B2(n15655), .A(n14330), .ZN(P1_U2812) );
  NOR2_X1 U17753 ( .A1(n14331), .A2(n14332), .ZN(n14333) );
  AOI21_X1 U17754 ( .B1(n14337), .B2(n14335), .A(n14336), .ZN(n14540) );
  NAND2_X1 U17755 ( .A1(n14540), .A2(n19809), .ZN(n14347) );
  INV_X1 U17756 ( .A(n14340), .ZN(n14338) );
  OR2_X1 U17757 ( .A1(n15677), .A2(n14338), .ZN(n14339) );
  NAND2_X1 U17758 ( .A1(n14339), .A2(n14405), .ZN(n14352) );
  INV_X1 U17759 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14423) );
  OR3_X1 U17760 ( .A1(n15677), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14340), .ZN(
        n14344) );
  OAI22_X1 U17761 ( .A1(n14341), .A2(n19769), .B1(n19821), .B2(n14538), .ZN(
        n14342) );
  INV_X1 U17762 ( .A(n14342), .ZN(n14343) );
  OAI211_X1 U17763 ( .C1(n14423), .C2(n19825), .A(n14344), .B(n14343), .ZN(
        n14345) );
  AOI21_X1 U17764 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14352), .A(n14345), 
        .ZN(n14346) );
  OAI211_X1 U17765 ( .C1(n19793), .C2(n14692), .A(n14347), .B(n14346), .ZN(
        P1_U2813) );
  OAI21_X1 U17766 ( .B1(n14349), .B2(n14350), .A(n14335), .ZN(n14546) );
  AOI21_X1 U17767 ( .B1(n14351), .B2(n14364), .A(n14331), .ZN(n14702) );
  INV_X1 U17768 ( .A(n14352), .ZN(n14357) );
  AOI21_X1 U17769 ( .B1(n15623), .B2(n14353), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14356) );
  AOI22_X1 U17770 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19823), .B1(
        n19766), .B2(n14549), .ZN(n14355) );
  NAND2_X1 U17771 ( .A1(n19797), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14354) );
  OAI211_X1 U17772 ( .C1(n14357), .C2(n14356), .A(n14355), .B(n14354), .ZN(
        n14358) );
  AOI21_X1 U17773 ( .B1(n14702), .B2(n19828), .A(n14358), .ZN(n14359) );
  OAI21_X1 U17774 ( .B1(n14546), .B2(n15655), .A(n14359), .ZN(P1_U2814) );
  AOI21_X1 U17775 ( .B1(n14361), .B2(n14360), .A(n14349), .ZN(n14559) );
  INV_X1 U17776 ( .A(n14559), .ZN(n14479) );
  NAND2_X1 U17777 ( .A1(n14374), .A2(n14362), .ZN(n14363) );
  AND2_X1 U17778 ( .A1(n14364), .A2(n14363), .ZN(n14712) );
  AOI21_X1 U17779 ( .B1(n15623), .B2(n14382), .A(n14365), .ZN(n14380) );
  INV_X1 U17780 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14555) );
  OAI22_X1 U17781 ( .A1(n14366), .A2(n19769), .B1(n19821), .B2(n14557), .ZN(
        n14367) );
  AOI21_X1 U17782 ( .B1(n19797), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14367), .ZN(
        n14370) );
  OAI21_X1 U17783 ( .B1(n14382), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14368) );
  OAI211_X1 U17784 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(P1_REIP_REG_24__SCAN_IN), .A(n15623), .B(n14368), .ZN(n14369) );
  OAI211_X1 U17785 ( .C1(n14380), .C2(n14555), .A(n14370), .B(n14369), .ZN(
        n14371) );
  AOI21_X1 U17786 ( .B1(n14712), .B2(n19828), .A(n14371), .ZN(n14372) );
  OAI21_X1 U17787 ( .B1(n14479), .B2(n15655), .A(n14372), .ZN(P1_U2815) );
  OAI21_X1 U17788 ( .B1(n14373), .B2(n14375), .A(n14374), .ZN(n14717) );
  OAI21_X1 U17789 ( .B1(n14377), .B2(n14378), .A(n14360), .ZN(n14566) );
  INV_X1 U17790 ( .A(n14566), .ZN(n14379) );
  NAND2_X1 U17791 ( .A1(n14379), .A2(n19809), .ZN(n14386) );
  INV_X1 U17792 ( .A(n14380), .ZN(n14396) );
  INV_X1 U17793 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U17794 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19823), .B1(
        n19766), .B2(n14569), .ZN(n14381) );
  OAI21_X1 U17795 ( .B1(n19825), .B2(n14426), .A(n14381), .ZN(n14384) );
  NOR3_X1 U17796 ( .A1(n15677), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14382), 
        .ZN(n14383) );
  AOI211_X1 U17797 ( .C1(n14396), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14384), 
        .B(n14383), .ZN(n14385) );
  OAI211_X1 U17798 ( .C1(n19793), .C2(n14717), .A(n14386), .B(n14385), .ZN(
        P1_U2816) );
  AND2_X1 U17799 ( .A1(n14404), .A2(n14387), .ZN(n14388) );
  OR2_X1 U17800 ( .A1(n14388), .A2(n14373), .ZN(n14730) );
  AOI21_X1 U17801 ( .B1(n14390), .B2(n14389), .A(n14377), .ZN(n14576) );
  NAND2_X1 U17802 ( .A1(n14576), .A2(n19809), .ZN(n14398) );
  OAI21_X1 U17803 ( .B1(n15677), .B2(n14391), .A(n14572), .ZN(n14395) );
  INV_X1 U17804 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14427) );
  NOR2_X1 U17805 ( .A1(n19825), .A2(n14427), .ZN(n14394) );
  OAI22_X1 U17806 ( .A1(n14392), .A2(n19769), .B1(n19821), .B2(n14574), .ZN(
        n14393) );
  AOI211_X1 U17807 ( .C1(n14396), .C2(n14395), .A(n14394), .B(n14393), .ZN(
        n14397) );
  OAI211_X1 U17808 ( .C1(n19793), .C2(n14730), .A(n14398), .B(n14397), .ZN(
        P1_U2817) );
  OAI21_X1 U17809 ( .B1(n14399), .B2(n14400), .A(n14389), .ZN(n14586) );
  INV_X1 U17810 ( .A(n14401), .ZN(n14433) );
  NAND2_X1 U17811 ( .A1(n14433), .A2(n14402), .ZN(n14403) );
  AND2_X1 U17812 ( .A1(n14404), .A2(n14403), .ZN(n15761) );
  AND2_X1 U17813 ( .A1(n15622), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15610) );
  NAND2_X1 U17814 ( .A1(n14405), .A2(n15610), .ZN(n14406) );
  NAND2_X1 U17815 ( .A1(n19789), .A2(n14406), .ZN(n15634) );
  INV_X1 U17816 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20691) );
  INV_X1 U17817 ( .A(n14580), .ZN(n14407) );
  OAI22_X1 U17818 ( .A1(n14578), .A2(n19769), .B1(n19821), .B2(n14407), .ZN(
        n14408) );
  AOI21_X1 U17819 ( .B1(n19797), .B2(P1_EBX_REG_22__SCAN_IN), .A(n14408), .ZN(
        n14415) );
  NAND2_X1 U17820 ( .A1(n15622), .A2(n14409), .ZN(n14410) );
  NAND2_X1 U17821 ( .A1(n14410), .A2(n20691), .ZN(n14412) );
  NAND2_X1 U17822 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14411) );
  NAND2_X1 U17823 ( .A1(n14412), .A2(n14411), .ZN(n14413) );
  OR2_X1 U17824 ( .A1(n15677), .A2(n14413), .ZN(n14414) );
  OAI211_X1 U17825 ( .C1(n15634), .C2(n20691), .A(n14415), .B(n14414), .ZN(
        n14416) );
  AOI21_X1 U17826 ( .B1(n15761), .B2(n19828), .A(n14416), .ZN(n14417) );
  OAI21_X1 U17827 ( .B1(n14586), .B2(n15655), .A(n14417), .ZN(P1_U2818) );
  OAI22_X1 U17828 ( .A1(n14419), .A2(n14465), .B1(n14418), .B2(n19851), .ZN(
        P1_U2841) );
  OAI222_X1 U17829 ( .A1(n14420), .A2(n19851), .B1(n14465), .B2(n14674), .C1(
        n14468), .C2(n14463), .ZN(P1_U2843) );
  OAI222_X1 U17830 ( .A1(n14422), .A2(n19851), .B1(n14465), .B2(n14421), .C1(
        n14471), .C2(n14463), .ZN(P1_U2844) );
  INV_X1 U17831 ( .A(n14540), .ZN(n14474) );
  OAI222_X1 U17832 ( .A1(n14423), .A2(n19851), .B1(n14465), .B2(n14692), .C1(
        n14474), .C2(n14463), .ZN(P1_U2845) );
  AOI22_X1 U17833 ( .A1(n14702), .A2(n19846), .B1(n14446), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n14424) );
  OAI21_X1 U17834 ( .B1(n14546), .B2(n14463), .A(n14424), .ZN(P1_U2846) );
  AOI22_X1 U17835 ( .A1(n14712), .A2(n19846), .B1(n14446), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14425) );
  OAI21_X1 U17836 ( .B1(n14479), .B2(n14463), .A(n14425), .ZN(P1_U2847) );
  OAI222_X1 U17837 ( .A1(n14426), .A2(n19851), .B1(n14465), .B2(n14717), .C1(
        n14566), .C2(n14463), .ZN(P1_U2848) );
  INV_X1 U17838 ( .A(n14576), .ZN(n14489) );
  OAI222_X1 U17839 ( .A1(n14427), .A2(n19851), .B1(n14465), .B2(n14730), .C1(
        n14489), .C2(n14463), .ZN(P1_U2849) );
  NOR2_X1 U17840 ( .A1(n19851), .A2(n14428), .ZN(n14429) );
  AOI21_X1 U17841 ( .B1(n15761), .B2(n19846), .A(n14429), .ZN(n14430) );
  OAI21_X1 U17842 ( .B1(n14586), .B2(n14463), .A(n14430), .ZN(P1_U2850) );
  INV_X1 U17843 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15614) );
  NAND2_X1 U17844 ( .A1(n14440), .A2(n14431), .ZN(n14432) );
  NAND2_X1 U17845 ( .A1(n14433), .A2(n14432), .ZN(n15617) );
  OR2_X1 U17846 ( .A1(n14434), .A2(n14439), .ZN(n14437) );
  AND2_X1 U17847 ( .A1(n14437), .A2(n14435), .ZN(n14436) );
  OR2_X1 U17848 ( .A1(n14436), .A2(n14399), .ZN(n15618) );
  OAI222_X1 U17849 ( .A1(n15614), .A2(n19851), .B1(n14465), .B2(n15617), .C1(
        n15618), .C2(n14463), .ZN(P1_U2851) );
  INV_X1 U17850 ( .A(n14437), .ZN(n14438) );
  AOI21_X1 U17851 ( .B1(n14439), .B2(n14434), .A(n14438), .ZN(n14599) );
  INV_X1 U17852 ( .A(n14599), .ZN(n15627) );
  INV_X1 U17853 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15625) );
  OAI21_X1 U17854 ( .B1(n14444), .B2(n14441), .A(n14440), .ZN(n15626) );
  OAI222_X1 U17855 ( .A1(n14463), .A2(n15627), .B1(n19851), .B2(n15625), .C1(
        n15626), .C2(n14465), .ZN(P1_U2852) );
  OAI21_X1 U17856 ( .B1(n14442), .B2(n14443), .A(n14434), .ZN(n15638) );
  AOI21_X1 U17857 ( .B1(n14445), .B2(n14454), .A(n14444), .ZN(n15771) );
  AOI22_X1 U17858 ( .A1(n15771), .A2(n19846), .B1(n14446), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n14447) );
  OAI21_X1 U17859 ( .B1(n15638), .B2(n14463), .A(n14447), .ZN(P1_U2853) );
  INV_X1 U17860 ( .A(n14448), .ZN(n14449) );
  INV_X1 U17861 ( .A(n14442), .ZN(n14450) );
  OAI21_X1 U17862 ( .B1(n14451), .B2(n14449), .A(n14450), .ZN(n15651) );
  NAND2_X1 U17863 ( .A1(n14460), .A2(n14452), .ZN(n14453) );
  NAND2_X1 U17864 ( .A1(n14454), .A2(n14453), .ZN(n15654) );
  OAI22_X1 U17865 ( .A1(n15654), .A2(n14465), .B1(n14455), .B2(n19851), .ZN(
        n14456) );
  INV_X1 U17866 ( .A(n14456), .ZN(n14457) );
  OAI21_X1 U17867 ( .B1(n15651), .B2(n14463), .A(n14457), .ZN(P1_U2854) );
  OR2_X1 U17868 ( .A1(n14151), .A2(n14458), .ZN(n14459) );
  NAND2_X1 U17869 ( .A1(n14460), .A2(n14459), .ZN(n15779) );
  INV_X1 U17870 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14464) );
  NOR2_X1 U17871 ( .A1(n14148), .A2(n14461), .ZN(n14462) );
  OR2_X1 U17872 ( .A1(n14449), .A2(n14462), .ZN(n15717) );
  OAI222_X1 U17873 ( .A1(n15779), .A2(n14465), .B1(n14464), .B2(n19851), .C1(
        n15717), .C2(n14463), .ZN(P1_U2855) );
  AOI22_X1 U17874 ( .A1(n14507), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14506), .ZN(n14467) );
  AOI22_X1 U17875 ( .A1(n14510), .A2(DATAI_29_), .B1(n14509), .B2(n19887), 
        .ZN(n14466) );
  OAI211_X1 U17876 ( .C1(n14468), .C2(n14493), .A(n14467), .B(n14466), .ZN(
        P1_U2875) );
  AOI22_X1 U17877 ( .A1(n14507), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14506), .ZN(n14470) );
  AOI22_X1 U17878 ( .A1(n14510), .A2(DATAI_28_), .B1(n14509), .B2(n19885), 
        .ZN(n14469) );
  OAI211_X1 U17879 ( .C1(n14471), .C2(n14493), .A(n14470), .B(n14469), .ZN(
        P1_U2876) );
  AOI22_X1 U17880 ( .A1(n14507), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14506), .ZN(n14473) );
  AOI22_X1 U17881 ( .A1(n14510), .A2(DATAI_27_), .B1(n14509), .B2(n19883), 
        .ZN(n14472) );
  OAI211_X1 U17882 ( .C1(n14474), .C2(n14493), .A(n14473), .B(n14472), .ZN(
        P1_U2877) );
  AOI22_X1 U17883 ( .A1(n14507), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14506), .ZN(n14476) );
  AOI22_X1 U17884 ( .A1(n14510), .A2(DATAI_26_), .B1(n14509), .B2(n19881), 
        .ZN(n14475) );
  OAI211_X1 U17885 ( .C1(n14546), .C2(n14493), .A(n14476), .B(n14475), .ZN(
        P1_U2878) );
  AOI22_X1 U17886 ( .A1(n14507), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14506), .ZN(n14478) );
  AOI22_X1 U17887 ( .A1(n14510), .A2(DATAI_25_), .B1(n14509), .B2(n19879), 
        .ZN(n14477) );
  OAI211_X1 U17888 ( .C1(n14479), .C2(n14493), .A(n14478), .B(n14477), .ZN(
        P1_U2879) );
  AOI22_X1 U17889 ( .A1(n14507), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14506), .ZN(n14481) );
  AOI22_X1 U17890 ( .A1(n14510), .A2(DATAI_24_), .B1(n14509), .B2(n19877), 
        .ZN(n14480) );
  OAI211_X1 U17891 ( .C1(n14566), .C2(n14493), .A(n14481), .B(n14480), .ZN(
        P1_U2880) );
  INV_X1 U17892 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16189) );
  OAI22_X1 U17893 ( .A1(n14484), .A2(n16189), .B1(n14483), .B2(n14482), .ZN(
        n14485) );
  INV_X1 U17894 ( .A(n14485), .ZN(n14488) );
  AOI22_X1 U17895 ( .A1(n14510), .A2(DATAI_23_), .B1(n14509), .B2(n14486), 
        .ZN(n14487) );
  OAI211_X1 U17896 ( .C1(n14489), .C2(n14493), .A(n14488), .B(n14487), .ZN(
        P1_U2881) );
  AOI22_X1 U17897 ( .A1(n14507), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14506), .ZN(n14492) );
  AOI22_X1 U17898 ( .A1(n14510), .A2(DATAI_22_), .B1(n14509), .B2(n14490), 
        .ZN(n14491) );
  OAI211_X1 U17899 ( .C1(n14586), .C2(n14493), .A(n14492), .B(n14491), .ZN(
        P1_U2882) );
  AOI22_X1 U17900 ( .A1(n14507), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14506), .ZN(n14496) );
  AOI22_X1 U17901 ( .A1(n14510), .A2(DATAI_21_), .B1(n14509), .B2(n14494), 
        .ZN(n14495) );
  OAI211_X1 U17902 ( .C1(n15618), .C2(n14493), .A(n14496), .B(n14495), .ZN(
        P1_U2883) );
  AOI22_X1 U17903 ( .A1(n14507), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14506), .ZN(n14499) );
  AOI22_X1 U17904 ( .A1(n14510), .A2(DATAI_20_), .B1(n14509), .B2(n14497), 
        .ZN(n14498) );
  OAI211_X1 U17905 ( .C1(n15627), .C2(n14493), .A(n14499), .B(n14498), .ZN(
        P1_U2884) );
  AOI22_X1 U17906 ( .A1(n14507), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14506), .ZN(n14502) );
  AOI22_X1 U17907 ( .A1(n14510), .A2(DATAI_19_), .B1(n14509), .B2(n14500), 
        .ZN(n14501) );
  OAI211_X1 U17908 ( .C1(n15638), .C2(n14493), .A(n14502), .B(n14501), .ZN(
        P1_U2885) );
  AOI22_X1 U17909 ( .A1(n14507), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14506), .ZN(n14505) );
  AOI22_X1 U17910 ( .A1(n14510), .A2(DATAI_18_), .B1(n14509), .B2(n14503), 
        .ZN(n14504) );
  OAI211_X1 U17911 ( .C1(n15651), .C2(n14493), .A(n14505), .B(n14504), .ZN(
        P1_U2886) );
  AOI22_X1 U17912 ( .A1(n14507), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14506), .ZN(n14512) );
  AOI22_X1 U17913 ( .A1(n14510), .A2(DATAI_17_), .B1(n14509), .B2(n14508), 
        .ZN(n14511) );
  OAI211_X1 U17914 ( .C1(n15717), .C2(n14493), .A(n14512), .B(n14511), .ZN(
        P1_U2887) );
  INV_X1 U17915 ( .A(n14513), .ZN(n14515) );
  NAND2_X1 U17916 ( .A1(n14515), .A2(n14514), .ZN(n14516) );
  XNOR2_X1 U17917 ( .A(n14516), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14668) );
  NAND2_X1 U17918 ( .A1(n15731), .A2(n14517), .ZN(n14518) );
  NAND2_X1 U17919 ( .A1(n12105), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14660) );
  OAI211_X1 U17920 ( .C1(n14653), .C2(n14519), .A(n14518), .B(n14660), .ZN(
        n14520) );
  AOI21_X1 U17921 ( .B1(n14521), .B2(n19911), .A(n14520), .ZN(n14522) );
  OAI21_X1 U17922 ( .B1(n14668), .B2(n19746), .A(n14522), .ZN(P1_U2969) );
  INV_X1 U17923 ( .A(n14523), .ZN(n14524) );
  NOR2_X1 U17924 ( .A1(n19942), .A2(n14526), .ZN(n14669) );
  AOI21_X1 U17925 ( .B1(n19908), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14669), .ZN(n14527) );
  OAI21_X1 U17926 ( .B1(n19916), .B2(n14528), .A(n14527), .ZN(n14529) );
  AOI21_X1 U17927 ( .B1(n14530), .B2(n19911), .A(n14529), .ZN(n14531) );
  OAI21_X1 U17928 ( .B1(n14677), .B2(n19746), .A(n14531), .ZN(P1_U2970) );
  INV_X1 U17929 ( .A(n11536), .ZN(n14532) );
  NAND2_X1 U17930 ( .A1(n14533), .A2(n14532), .ZN(n14534) );
  MUX2_X1 U17931 ( .A(n14535), .B(n14534), .S(n15735), .Z(n14536) );
  XNOR2_X1 U17932 ( .A(n14536), .B(n14690), .ZN(n14696) );
  NOR2_X1 U17933 ( .A1(n19942), .A2(n20604), .ZN(n14688) );
  AOI21_X1 U17934 ( .B1(n19908), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14688), .ZN(n14537) );
  OAI21_X1 U17935 ( .B1(n19916), .B2(n14538), .A(n14537), .ZN(n14539) );
  AOI21_X1 U17936 ( .B1(n14540), .B2(n19911), .A(n14539), .ZN(n14541) );
  OAI21_X1 U17937 ( .B1(n19746), .B2(n14696), .A(n14541), .ZN(P1_U2972) );
  INV_X1 U17938 ( .A(n14251), .ZN(n14561) );
  OAI21_X1 U17939 ( .B1(n14561), .B2(n14698), .A(n15735), .ZN(n14542) );
  NAND2_X1 U17940 ( .A1(n14543), .A2(n14542), .ZN(n14544) );
  XOR2_X1 U17941 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14544), .Z(
        n14708) );
  NAND2_X1 U17942 ( .A1(n12105), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14697) );
  OAI21_X1 U17943 ( .B1(n14653), .B2(n14545), .A(n14697), .ZN(n14548) );
  NOR2_X1 U17944 ( .A1(n14546), .A2(n19960), .ZN(n14547) );
  OAI21_X1 U17945 ( .B1(n19746), .B2(n14708), .A(n14550), .ZN(P1_U2973) );
  NAND2_X1 U17946 ( .A1(n14551), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14563) );
  MUX2_X1 U17947 ( .A(n14723), .B(n14552), .S(n15702), .Z(n14553) );
  AOI21_X1 U17948 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14563), .A(
        n14553), .ZN(n14554) );
  XNOR2_X1 U17949 ( .A(n14554), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14709) );
  NOR2_X1 U17950 ( .A1(n19942), .A2(n14555), .ZN(n14710) );
  AOI21_X1 U17951 ( .B1(n19908), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14710), .ZN(n14556) );
  OAI21_X1 U17952 ( .B1(n19916), .B2(n14557), .A(n14556), .ZN(n14558) );
  AOI21_X1 U17953 ( .B1(n14559), .B2(n19911), .A(n14558), .ZN(n14560) );
  OAI21_X1 U17954 ( .B1(n19746), .B2(n14709), .A(n14560), .ZN(P1_U2974) );
  NAND2_X1 U17955 ( .A1(n14561), .A2(n14563), .ZN(n14562) );
  MUX2_X1 U17956 ( .A(n14563), .B(n14562), .S(n15702), .Z(n14564) );
  XNOR2_X1 U17957 ( .A(n14564), .B(n14723), .ZN(n14726) );
  NAND2_X1 U17958 ( .A1(n12105), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14719) );
  OAI21_X1 U17959 ( .B1(n14653), .B2(n14565), .A(n14719), .ZN(n14568) );
  NOR2_X1 U17960 ( .A1(n14566), .A2(n19960), .ZN(n14567) );
  AOI211_X1 U17961 ( .C1(n15731), .C2(n14569), .A(n14568), .B(n14567), .ZN(
        n14570) );
  OAI21_X1 U17962 ( .B1(n19746), .B2(n14726), .A(n14570), .ZN(P1_U2975) );
  XNOR2_X1 U17963 ( .A(n15735), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14571) );
  XNOR2_X1 U17964 ( .A(n14251), .B(n14571), .ZN(n14731) );
  NOR2_X1 U17965 ( .A1(n19942), .A2(n14572), .ZN(n14727) );
  AOI21_X1 U17966 ( .B1(n19908), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14727), .ZN(n14573) );
  OAI21_X1 U17967 ( .B1(n19916), .B2(n14574), .A(n14573), .ZN(n14575) );
  AOI21_X1 U17968 ( .B1(n14576), .B2(n19911), .A(n14575), .ZN(n14577) );
  OAI21_X1 U17969 ( .B1(n14731), .B2(n19746), .A(n14577), .ZN(P1_U2976) );
  OAI22_X1 U17970 ( .A1(n14653), .A2(n14578), .B1(n19942), .B2(n20691), .ZN(
        n14579) );
  AOI21_X1 U17971 ( .B1(n14580), .B2(n15731), .A(n14579), .ZN(n14585) );
  NAND2_X1 U17972 ( .A1(n14582), .A2(n14581), .ZN(n14583) );
  XNOR2_X1 U17973 ( .A(n14583), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15766) );
  NAND2_X1 U17974 ( .A1(n15766), .A2(n19912), .ZN(n14584) );
  OAI211_X1 U17975 ( .C1(n14586), .C2(n19960), .A(n14585), .B(n14584), .ZN(
        P1_U2977) );
  NOR2_X1 U17976 ( .A1(n14587), .A2(n15702), .ZN(n14595) );
  NOR2_X1 U17977 ( .A1(n14588), .A2(n15735), .ZN(n14594) );
  AOI22_X1 U17978 ( .A1(n14595), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n14594), .B2(n14751), .ZN(n14589) );
  XNOR2_X1 U17979 ( .A(n14589), .B(n14743), .ZN(n14747) );
  NAND2_X1 U17980 ( .A1(n12105), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14741) );
  OAI21_X1 U17981 ( .B1(n14653), .B2(n14590), .A(n14741), .ZN(n14592) );
  NOR2_X1 U17982 ( .A1(n15618), .A2(n19960), .ZN(n14591) );
  AOI211_X1 U17983 ( .C1(n15731), .C2(n15611), .A(n14592), .B(n14591), .ZN(
        n14593) );
  OAI21_X1 U17984 ( .B1(n14747), .B2(n19746), .A(n14593), .ZN(P1_U2978) );
  NOR2_X1 U17985 ( .A1(n14595), .A2(n14594), .ZN(n14596) );
  XNOR2_X1 U17986 ( .A(n14596), .B(n14751), .ZN(n14758) );
  NAND2_X1 U17987 ( .A1(n15731), .A2(n15630), .ZN(n14597) );
  NAND2_X1 U17988 ( .A1(n12105), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14753) );
  OAI211_X1 U17989 ( .C1(n14653), .C2(n15624), .A(n14597), .B(n14753), .ZN(
        n14598) );
  AOI21_X1 U17990 ( .B1(n14599), .B2(n19911), .A(n14598), .ZN(n14600) );
  OAI21_X1 U17991 ( .B1(n14758), .B2(n19746), .A(n14600), .ZN(P1_U2979) );
  NAND2_X1 U17992 ( .A1(n12105), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14768) );
  OAI21_X1 U17993 ( .B1(n14653), .B2(n14601), .A(n14768), .ZN(n14602) );
  AOI21_X1 U17994 ( .B1(n15649), .B2(n15731), .A(n14602), .ZN(n14607) );
  OR2_X1 U17995 ( .A1(n9625), .A2(n14603), .ZN(n14759) );
  NAND3_X1 U17996 ( .A1(n14759), .A2(n14605), .A3(n19912), .ZN(n14606) );
  OAI211_X1 U17997 ( .C1(n15651), .C2(n19960), .A(n14607), .B(n14606), .ZN(
        P1_U2981) );
  INV_X1 U17998 ( .A(n14608), .ZN(n14637) );
  INV_X1 U17999 ( .A(n14609), .ZN(n14611) );
  AOI21_X1 U18000 ( .B1(n14637), .B2(n14611), .A(n14610), .ZN(n15723) );
  INV_X1 U18001 ( .A(n14614), .ZN(n14612) );
  NOR2_X1 U18002 ( .A1(n14613), .A2(n14612), .ZN(n15722) );
  NAND2_X1 U18003 ( .A1(n15723), .A2(n15722), .ZN(n15721) );
  NAND2_X1 U18004 ( .A1(n15721), .A2(n14614), .ZN(n14616) );
  XNOR2_X1 U18005 ( .A(n14616), .B(n14615), .ZN(n15791) );
  NAND2_X1 U18006 ( .A1(n15791), .A2(n19912), .ZN(n14621) );
  NAND2_X1 U18007 ( .A1(n12105), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15787) );
  OAI21_X1 U18008 ( .B1(n14653), .B2(n14617), .A(n15787), .ZN(n14618) );
  AOI21_X1 U18009 ( .B1(n14619), .B2(n15731), .A(n14618), .ZN(n14620) );
  OAI211_X1 U18010 ( .C1(n19960), .C2(n14622), .A(n14621), .B(n14620), .ZN(
        P1_U2983) );
  NOR2_X1 U18011 ( .A1(n14637), .A2(n14623), .ZN(n15711) );
  NAND2_X1 U18012 ( .A1(n14624), .A2(n14639), .ZN(n14626) );
  OAI21_X1 U18013 ( .B1(n15711), .B2(n14626), .A(n14625), .ZN(n14628) );
  XNOR2_X1 U18014 ( .A(n14633), .B(n15809), .ZN(n14627) );
  XNOR2_X1 U18015 ( .A(n14628), .B(n14627), .ZN(n15806) );
  NAND2_X1 U18016 ( .A1(n15806), .A2(n19912), .ZN(n14631) );
  NOR2_X1 U18017 ( .A1(n19942), .A2(n15675), .ZN(n15803) );
  NOR2_X1 U18018 ( .A1(n19916), .A2(n15672), .ZN(n14629) );
  AOI211_X1 U18019 ( .C1(n19908), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15803), .B(n14629), .ZN(n14630) );
  OAI211_X1 U18020 ( .C1(n19960), .C2(n15674), .A(n14631), .B(n14630), .ZN(
        P1_U2985) );
  INV_X1 U18021 ( .A(n14632), .ZN(n14636) );
  AOI21_X1 U18022 ( .B1(n14634), .B2(n15738), .A(n15735), .ZN(n14635) );
  AOI21_X1 U18023 ( .B1(n14637), .B2(n14636), .A(n14635), .ZN(n14776) );
  INV_X1 U18024 ( .A(n14639), .ZN(n14638) );
  AOI21_X1 U18025 ( .B1(n15702), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14638), .ZN(n14775) );
  NAND2_X1 U18026 ( .A1(n14776), .A2(n14775), .ZN(n14774) );
  NAND2_X1 U18027 ( .A1(n14774), .A2(n14639), .ZN(n14640) );
  XOR2_X1 U18028 ( .A(n14641), .B(n14640), .Z(n15817) );
  NAND2_X1 U18029 ( .A1(n15817), .A2(n19912), .ZN(n14646) );
  INV_X1 U18030 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14642) );
  OAI22_X1 U18031 ( .A1(n14653), .A2(n14108), .B1(n19942), .B2(n14642), .ZN(
        n14643) );
  AOI21_X1 U18032 ( .B1(n15731), .B2(n14644), .A(n14643), .ZN(n14645) );
  OAI211_X1 U18033 ( .C1(n19960), .C2(n14647), .A(n14646), .B(n14645), .ZN(
        P1_U2986) );
  MUX2_X1 U18034 ( .A(n14649), .B(n14608), .S(n14633), .Z(n14650) );
  XOR2_X1 U18035 ( .A(n14634), .B(n14650), .Z(n15834) );
  NAND2_X1 U18036 ( .A1(n15834), .A2(n19912), .ZN(n14657) );
  INV_X1 U18037 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14651) );
  OAI22_X1 U18038 ( .A1(n14653), .A2(n14652), .B1(n19942), .B2(n14651), .ZN(
        n14654) );
  AOI21_X1 U18039 ( .B1(n14655), .B2(n15731), .A(n14654), .ZN(n14656) );
  OAI211_X1 U18040 ( .C1(n19960), .C2(n14658), .A(n14657), .B(n14656), .ZN(
        P1_U2989) );
  INV_X1 U18041 ( .A(n14659), .ZN(n14666) );
  INV_X1 U18042 ( .A(n14660), .ZN(n14665) );
  AOI21_X1 U18043 ( .B1(n14663), .B2(n14662), .A(n14661), .ZN(n14664) );
  AOI211_X1 U18044 ( .C1(n14666), .C2(n19925), .A(n14665), .B(n14664), .ZN(
        n14667) );
  OAI21_X1 U18045 ( .B1(n14668), .B2(n19946), .A(n14667), .ZN(P1_U3001) );
  AOI21_X1 U18046 ( .B1(n14670), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14669), .ZN(n14673) );
  NAND2_X1 U18047 ( .A1(n14671), .A2(n9649), .ZN(n14672) );
  OAI211_X1 U18048 ( .C1(n14674), .C2(n19945), .A(n14673), .B(n14672), .ZN(
        n14675) );
  INV_X1 U18049 ( .A(n14675), .ZN(n14676) );
  OAI21_X1 U18050 ( .B1(n14677), .B2(n19946), .A(n14676), .ZN(P1_U3002) );
  NAND3_X1 U18051 ( .A1(n14691), .A2(n14679), .A3(n14678), .ZN(n14681) );
  OAI211_X1 U18052 ( .C1(n14687), .C2(n14682), .A(n14681), .B(n14680), .ZN(
        n14683) );
  AOI21_X1 U18053 ( .B1(n14684), .B2(n19925), .A(n14683), .ZN(n14685) );
  OAI21_X1 U18054 ( .B1(n14686), .B2(n19946), .A(n14685), .ZN(P1_U3003) );
  NOR2_X1 U18055 ( .A1(n14687), .A2(n14690), .ZN(n14689) );
  AOI211_X1 U18056 ( .C1(n14691), .C2(n14690), .A(n14689), .B(n14688), .ZN(
        n14695) );
  INV_X1 U18057 ( .A(n14692), .ZN(n14693) );
  NAND2_X1 U18058 ( .A1(n14693), .A2(n19925), .ZN(n14694) );
  OAI211_X1 U18059 ( .C1(n14696), .C2(n19946), .A(n14695), .B(n14694), .ZN(
        P1_U3004) );
  INV_X1 U18060 ( .A(n14697), .ZN(n14701) );
  INV_X1 U18061 ( .A(n14734), .ZN(n14699) );
  NOR3_X1 U18062 ( .A1(n14699), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14698), .ZN(n14700) );
  AOI211_X1 U18063 ( .C1(n14702), .C2(n19925), .A(n14701), .B(n14700), .ZN(
        n14707) );
  AND3_X1 U18064 ( .A1(n14703), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14704) );
  NAND2_X1 U18065 ( .A1(n14734), .A2(n14704), .ZN(n14714) );
  INV_X1 U18066 ( .A(n14714), .ZN(n14705) );
  OAI21_X1 U18067 ( .B1(n14705), .B2(n14711), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14706) );
  OAI211_X1 U18068 ( .C1(n14708), .C2(n19946), .A(n14707), .B(n14706), .ZN(
        P1_U3005) );
  OR2_X1 U18069 ( .A1(n14709), .A2(n19946), .ZN(n14716) );
  AOI21_X1 U18070 ( .B1(n14711), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14710), .ZN(n14715) );
  NAND2_X1 U18071 ( .A1(n14712), .A2(n19925), .ZN(n14713) );
  NAND4_X1 U18072 ( .A1(n14716), .A2(n14715), .A3(n14714), .A4(n14713), .ZN(
        P1_U3006) );
  INV_X1 U18073 ( .A(n14717), .ZN(n14722) );
  AOI21_X1 U18074 ( .B1(n19935), .B2(n11535), .A(n14718), .ZN(n14720) );
  OAI21_X1 U18075 ( .B1(n14720), .B2(n14723), .A(n14719), .ZN(n14721) );
  AOI21_X1 U18076 ( .B1(n14722), .B2(n19925), .A(n14721), .ZN(n14725) );
  NAND3_X1 U18077 ( .A1(n14734), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14723), .ZN(n14724) );
  OAI211_X1 U18078 ( .C1(n14726), .C2(n19946), .A(n14725), .B(n14724), .ZN(
        P1_U3007) );
  AOI21_X1 U18079 ( .B1(n14728), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14727), .ZN(n14729) );
  OAI21_X1 U18080 ( .B1(n14730), .B2(n19945), .A(n14729), .ZN(n14733) );
  NOR2_X1 U18081 ( .A1(n14731), .A2(n19946), .ZN(n14732) );
  AOI211_X1 U18082 ( .C1(n14734), .C2(n11535), .A(n14733), .B(n14732), .ZN(
        n14735) );
  INV_X1 U18083 ( .A(n14735), .ZN(P1_U3008) );
  INV_X1 U18084 ( .A(n15617), .ZN(n14745) );
  NAND2_X1 U18085 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15812), .ZN(
        n14762) );
  INV_X1 U18086 ( .A(n14766), .ZN(n14736) );
  OAI22_X1 U18087 ( .A1(n14737), .A2(n14762), .B1(n14736), .B2(n19936), .ZN(
        n15813) );
  NAND2_X1 U18088 ( .A1(n15813), .A2(n14738), .ZN(n14748) );
  OAI21_X1 U18089 ( .B1(n14739), .B2(n14761), .A(n14748), .ZN(n15774) );
  AND2_X1 U18090 ( .A1(n15774), .A2(n14740), .ZN(n15768) );
  NAND2_X1 U18091 ( .A1(n15768), .A2(n14743), .ZN(n14742) );
  OAI211_X1 U18092 ( .C1(n15762), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        n14744) );
  AOI21_X1 U18093 ( .B1(n14745), .B2(n19925), .A(n14744), .ZN(n14746) );
  OAI21_X1 U18094 ( .B1(n14747), .B2(n19946), .A(n14746), .ZN(P1_U3010) );
  INV_X1 U18095 ( .A(n15626), .ZN(n14756) );
  AOI21_X1 U18096 ( .B1(n14748), .B2(n14761), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14750) );
  INV_X1 U18097 ( .A(n14749), .ZN(n15775) );
  OAI21_X1 U18098 ( .B1(n14750), .B2(n15775), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14754) );
  NAND3_X1 U18099 ( .A1(n15774), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14751), .ZN(n14752) );
  NAND3_X1 U18100 ( .A1(n14754), .A2(n14753), .A3(n14752), .ZN(n14755) );
  AOI21_X1 U18101 ( .B1(n14756), .B2(n19925), .A(n14755), .ZN(n14757) );
  OAI21_X1 U18102 ( .B1(n14758), .B2(n19946), .A(n14757), .ZN(P1_U3011) );
  NAND3_X1 U18103 ( .A1(n14759), .A2(n14605), .A3(n19929), .ZN(n14773) );
  NAND2_X1 U18104 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15786) );
  NOR3_X1 U18105 ( .A1(n15872), .A2(n14760), .A3(n15814), .ZN(n15805) );
  NAND2_X1 U18106 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15805), .ZN(
        n15796) );
  NOR2_X1 U18107 ( .A1(n15786), .A2(n15796), .ZN(n15782) );
  NOR2_X1 U18108 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11521), .ZN(
        n14771) );
  AOI21_X1 U18109 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15812), .A(
        n14761), .ZN(n15811) );
  AOI21_X1 U18110 ( .B1(n14763), .B2(n14762), .A(n15811), .ZN(n14765) );
  OAI211_X1 U18111 ( .C1(n14766), .C2(n19936), .A(n14765), .B(n14764), .ZN(
        n15816) );
  AOI21_X1 U18112 ( .B1(n15814), .B2(n15813), .A(n15816), .ZN(n15810) );
  OAI21_X1 U18113 ( .B1(n15790), .B2(n14767), .A(n15810), .ZN(n15781) );
  NAND2_X1 U18114 ( .A1(n15781), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14769) );
  OAI211_X1 U18115 ( .C1(n19945), .C2(n15654), .A(n14769), .B(n14768), .ZN(
        n14770) );
  AOI21_X1 U18116 ( .B1(n15782), .B2(n14771), .A(n14770), .ZN(n14772) );
  NAND2_X1 U18117 ( .A1(n14773), .A2(n14772), .ZN(P1_U3013) );
  NOR2_X1 U18118 ( .A1(n15872), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14786) );
  OAI21_X1 U18119 ( .B1(n14776), .B2(n14775), .A(n14774), .ZN(n14777) );
  INV_X1 U18120 ( .A(n14777), .ZN(n15734) );
  NOR2_X1 U18121 ( .A1(n14778), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15821) );
  INV_X1 U18122 ( .A(n19936), .ZN(n19951) );
  AOI21_X1 U18123 ( .B1(n19951), .B2(n15847), .A(n19938), .ZN(n14781) );
  OAI21_X1 U18124 ( .B1(n14779), .B2(n14778), .A(n19940), .ZN(n14780) );
  OAI211_X1 U18125 ( .C1(n14785), .C2(n19936), .A(n14781), .B(n14780), .ZN(
        n15825) );
  AOI21_X1 U18126 ( .B1(n19935), .B2(n15821), .A(n15825), .ZN(n14783) );
  OAI22_X1 U18127 ( .A1(n15734), .A2(n19946), .B1(n14783), .B2(n14782), .ZN(
        n14784) );
  AOI21_X1 U18128 ( .B1(n14786), .B2(n14785), .A(n14784), .ZN(n14788) );
  NAND2_X1 U18129 ( .A1(n12105), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14787) );
  OAI211_X1 U18130 ( .C1(n19945), .C2(n15685), .A(n14788), .B(n14787), .ZN(
        P1_U3019) );
  NAND3_X1 U18131 ( .A1(n14790), .A2(n15572), .A3(n14789), .ZN(n15587) );
  AOI22_X1 U18132 ( .A1(n19962), .A2(n20418), .B1(n11614), .B2(n14791), .ZN(
        n14792) );
  NAND2_X1 U18133 ( .A1(n15587), .A2(n14792), .ZN(n14793) );
  MUX2_X1 U18134 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n14793), .S(
        n19956), .Z(P1_U3478) );
  OR2_X1 U18135 ( .A1(n13694), .A2(n14794), .ZN(n14799) );
  NAND2_X1 U18136 ( .A1(n14803), .A2(n14802), .ZN(n14795) );
  NOR2_X1 U18137 ( .A1(n14796), .A2(n14795), .ZN(n14797) );
  AOI21_X1 U18138 ( .B1(n15550), .B2(n11314), .A(n14797), .ZN(n14798) );
  NAND2_X1 U18139 ( .A1(n14799), .A2(n14798), .ZN(n15549) );
  NAND2_X1 U18140 ( .A1(n15549), .A2(n14800), .ZN(n14805) );
  NAND3_X1 U18141 ( .A1(n14803), .A2(n14802), .A3(n14801), .ZN(n14804) );
  OAI211_X1 U18142 ( .C1(n14807), .C2(n14806), .A(n14805), .B(n14804), .ZN(
        n14809) );
  MUX2_X1 U18143 ( .A(n14809), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n14808), .Z(P1_U3473) );
  NAND2_X1 U18144 ( .A1(n12869), .A2(n14810), .ZN(n14812) );
  XNOR2_X1 U18145 ( .A(n14812), .B(n14811), .ZN(n14887) );
  INV_X1 U18146 ( .A(n14813), .ZN(n14814) );
  OAI21_X1 U18147 ( .B1(n13210), .B2(n14815), .A(n14814), .ZN(n15921) );
  NOR2_X1 U18148 ( .A1(n15921), .A2(n14873), .ZN(n14816) );
  AOI21_X1 U18149 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14873), .A(n14816), .ZN(
        n14817) );
  OAI21_X1 U18150 ( .B1(n14887), .B2(n14880), .A(n14817), .ZN(P2_U2859) );
  AOI21_X1 U18151 ( .B1(n14820), .B2(n14819), .A(n14818), .ZN(n14888) );
  NAND2_X1 U18152 ( .A1(n14888), .A2(n14870), .ZN(n14822) );
  NAND2_X1 U18153 ( .A1(n14873), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14821) );
  OAI211_X1 U18154 ( .C1(n14873), .C2(n15172), .A(n14822), .B(n14821), .ZN(
        P2_U2860) );
  OAI21_X1 U18155 ( .B1(n14825), .B2(n14824), .A(n14823), .ZN(n14904) );
  AND2_X1 U18156 ( .A1(n14835), .A2(n14826), .ZN(n14828) );
  OR2_X1 U18157 ( .A1(n14828), .A2(n14827), .ZN(n15928) );
  NOR2_X1 U18158 ( .A1(n15928), .A2(n14873), .ZN(n14829) );
  AOI21_X1 U18159 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14873), .A(n14829), .ZN(
        n14830) );
  OAI21_X1 U18160 ( .B1(n14904), .B2(n14880), .A(n14830), .ZN(P2_U2861) );
  OAI21_X1 U18161 ( .B1(n14833), .B2(n14832), .A(n14831), .ZN(n14910) );
  INV_X1 U18162 ( .A(n14834), .ZN(n14848) );
  INV_X1 U18163 ( .A(n14835), .ZN(n14836) );
  AOI21_X1 U18164 ( .B1(n14837), .B2(n14848), .A(n14836), .ZN(n15936) );
  NOR2_X1 U18165 ( .A1(n14840), .A2(n14838), .ZN(n14839) );
  AOI21_X1 U18166 ( .B1(n15936), .B2(n14840), .A(n14839), .ZN(n14841) );
  OAI21_X1 U18167 ( .B1(n14910), .B2(n14880), .A(n14841), .ZN(P2_U2862) );
  AOI21_X1 U18168 ( .B1(n14842), .B2(n14844), .A(n14843), .ZN(n14845) );
  XOR2_X1 U18169 ( .A(n14846), .B(n14845), .Z(n14917) );
  INV_X1 U18170 ( .A(n13194), .ZN(n14850) );
  INV_X1 U18171 ( .A(n14847), .ZN(n14849) );
  OAI21_X1 U18172 ( .B1(n14850), .B2(n14849), .A(n14848), .ZN(n15952) );
  MUX2_X1 U18173 ( .A(n9914), .B(n15952), .S(n14840), .Z(n14851) );
  OAI21_X1 U18174 ( .B1(n14917), .B2(n14880), .A(n14851), .ZN(P2_U2863) );
  AOI21_X1 U18175 ( .B1(n14852), .B2(n14854), .A(n14853), .ZN(n14855) );
  INV_X1 U18176 ( .A(n14855), .ZN(n14923) );
  NOR2_X1 U18177 ( .A1(n15218), .A2(n14873), .ZN(n14856) );
  AOI21_X1 U18178 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n14873), .A(n14856), .ZN(
        n14857) );
  OAI21_X1 U18179 ( .B1(n14923), .B2(n14880), .A(n14857), .ZN(P2_U2864) );
  NOR2_X1 U18180 ( .A1(n14864), .A2(n14858), .ZN(n14859) );
  OR2_X1 U18181 ( .A1(n13195), .A2(n14859), .ZN(n15537) );
  AOI21_X1 U18182 ( .B1(n14860), .B2(n14867), .A(n9674), .ZN(n15959) );
  NAND2_X1 U18183 ( .A1(n15959), .A2(n14870), .ZN(n14862) );
  NAND2_X1 U18184 ( .A1(n14873), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14861) );
  OAI211_X1 U18185 ( .C1(n15537), .C2(n14873), .A(n14862), .B(n14861), .ZN(
        P2_U2865) );
  AND2_X1 U18186 ( .A1(n14876), .A2(n14863), .ZN(n14865) );
  OR2_X1 U18187 ( .A1(n14865), .A2(n14864), .ZN(n18661) );
  INV_X1 U18188 ( .A(n14867), .ZN(n14868) );
  AOI21_X1 U18189 ( .B1(n14869), .B2(n14866), .A(n14868), .ZN(n14924) );
  NAND2_X1 U18190 ( .A1(n14924), .A2(n14870), .ZN(n14872) );
  NAND2_X1 U18191 ( .A1(n14873), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14871) );
  OAI211_X1 U18192 ( .C1(n18661), .C2(n14873), .A(n14872), .B(n14871), .ZN(
        P2_U2866) );
  OAI21_X1 U18193 ( .B1(n14084), .B2(n14874), .A(n14866), .ZN(n15964) );
  INV_X1 U18194 ( .A(n14087), .ZN(n14877) );
  OAI21_X1 U18195 ( .B1(n14877), .B2(n9738), .A(n14876), .ZN(n18678) );
  NOR2_X1 U18196 ( .A1(n18678), .A2(n14873), .ZN(n14878) );
  AOI21_X1 U18197 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n14873), .A(n14878), .ZN(
        n14879) );
  OAI21_X1 U18198 ( .B1(n14880), .B2(n15964), .A(n14879), .ZN(P2_U2867) );
  AOI21_X1 U18199 ( .B1(n14882), .B2(n13213), .A(n14881), .ZN(n15918) );
  INV_X1 U18200 ( .A(n18898), .ZN(n14883) );
  OAI22_X1 U18201 ( .A1(n14928), .A2(n14883), .B1(n18922), .B2(n18952), .ZN(
        n14884) );
  AOI21_X1 U18202 ( .B1(n15918), .B2(n18932), .A(n14884), .ZN(n14886) );
  AOI22_X1 U18203 ( .A1(n18884), .A2(BUF2_REG_28__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14885) );
  OAI211_X1 U18204 ( .C1(n14887), .C2(n18936), .A(n14886), .B(n14885), .ZN(
        P2_U2891) );
  INV_X1 U18205 ( .A(n14888), .ZN(n14896) );
  INV_X1 U18206 ( .A(n15177), .ZN(n14893) );
  INV_X1 U18207 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14889) );
  OR2_X1 U18208 ( .A1(n18891), .A2(n14889), .ZN(n14891) );
  NAND2_X1 U18209 ( .A1(n18891), .A2(BUF2_REG_11__SCAN_IN), .ZN(n14890) );
  AND2_X1 U18210 ( .A1(n14891), .A2(n14890), .ZN(n19040) );
  INV_X1 U18211 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n18954) );
  OAI22_X1 U18212 ( .A1(n14928), .A2(n19040), .B1(n18922), .B2(n18954), .ZN(
        n14892) );
  AOI21_X1 U18213 ( .B1(n14893), .B2(n18932), .A(n14892), .ZN(n14895) );
  AOI22_X1 U18214 ( .A1(n18884), .A2(BUF2_REG_27__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14894) );
  OAI211_X1 U18215 ( .C1(n14896), .C2(n18936), .A(n14895), .B(n14894), .ZN(
        P2_U2892) );
  NOR2_X1 U18216 ( .A1(n14898), .A2(n14897), .ZN(n14899) );
  OR2_X1 U18217 ( .A1(n13214), .A2(n14899), .ZN(n15185) );
  INV_X1 U18218 ( .A(n18932), .ZN(n18923) );
  INV_X1 U18219 ( .A(n14928), .ZN(n18882) );
  AOI22_X1 U18220 ( .A1(n18882), .A2(n18902), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n18931), .ZN(n14901) );
  AOI22_X1 U18221 ( .A1(n18884), .A2(BUF2_REG_26__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14900) );
  OAI211_X1 U18222 ( .C1(n15185), .C2(n18923), .A(n14901), .B(n14900), .ZN(
        n14902) );
  INV_X1 U18223 ( .A(n14902), .ZN(n14903) );
  OAI21_X1 U18224 ( .B1(n14904), .B2(n18936), .A(n14903), .ZN(P2_U2893) );
  XOR2_X1 U18225 ( .A(n14905), .B(n14911), .Z(n15935) );
  INV_X1 U18226 ( .A(n18905), .ZN(n14906) );
  OAI22_X1 U18227 ( .A1(n14928), .A2(n14906), .B1(n18922), .B2(n18958), .ZN(
        n14907) );
  AOI21_X1 U18228 ( .B1(n15935), .B2(n18932), .A(n14907), .ZN(n14909) );
  AOI22_X1 U18229 ( .A1(n18884), .A2(BUF2_REG_25__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14908) );
  OAI211_X1 U18230 ( .C1(n14910), .C2(n18936), .A(n14909), .B(n14908), .ZN(
        P2_U2894) );
  AOI21_X1 U18231 ( .B1(n14912), .B2(n13198), .A(n9897), .ZN(n15955) );
  INV_X1 U18232 ( .A(n18908), .ZN(n14913) );
  OAI22_X1 U18233 ( .A1(n14928), .A2(n14913), .B1(n18922), .B2(n18960), .ZN(
        n14914) );
  AOI21_X1 U18234 ( .B1(n15955), .B2(n18932), .A(n14914), .ZN(n14916) );
  AOI22_X1 U18235 ( .A1(n18884), .A2(BUF2_REG_24__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14915) );
  OAI211_X1 U18236 ( .C1(n14917), .C2(n18936), .A(n14916), .B(n14915), .ZN(
        P2_U2895) );
  INV_X1 U18237 ( .A(n15224), .ZN(n14921) );
  OAI22_X1 U18238 ( .A1(n14928), .A2(n19038), .B1(n18922), .B2(n18962), .ZN(
        n14920) );
  INV_X1 U18239 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n14918) );
  OAI22_X1 U18240 ( .A1(n14932), .A2(n14918), .B1(n14930), .B2(n16189), .ZN(
        n14919) );
  AOI211_X1 U18241 ( .C1(n18932), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14922) );
  OAI21_X1 U18242 ( .B1(n14923), .B2(n18936), .A(n14922), .ZN(P2_U2896) );
  INV_X1 U18243 ( .A(n14924), .ZN(n14936) );
  NAND2_X1 U18244 ( .A1(n14925), .A2(n14926), .ZN(n14927) );
  AND2_X1 U18245 ( .A1(n9671), .A2(n14927), .ZN(n18662) );
  INV_X1 U18246 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n18966) );
  OAI22_X1 U18247 ( .A1(n14928), .A2(n19034), .B1(n18922), .B2(n18966), .ZN(
        n14934) );
  INV_X1 U18248 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14931) );
  INV_X1 U18249 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14929) );
  OAI22_X1 U18250 ( .A1(n14932), .A2(n14931), .B1(n14930), .B2(n14929), .ZN(
        n14933) );
  AOI211_X1 U18251 ( .C1(n18932), .C2(n18662), .A(n14934), .B(n14933), .ZN(
        n14935) );
  OAI21_X1 U18252 ( .B1(n14936), .B2(n18936), .A(n14935), .ZN(P2_U2898) );
  NAND2_X1 U18253 ( .A1(n14938), .A2(n14937), .ZN(n14940) );
  XOR2_X1 U18254 ( .A(n14940), .B(n14939), .Z(n15159) );
  NAND2_X1 U18255 ( .A1(n15392), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15151) );
  OAI21_X1 U18256 ( .B1(n19061), .B2(n14942), .A(n15151), .ZN(n14943) );
  AOI21_X1 U18257 ( .B1(n19049), .B2(n15901), .A(n14943), .ZN(n14944) );
  OAI21_X1 U18258 ( .B1(n15906), .B2(n19057), .A(n14944), .ZN(n14945) );
  AOI21_X1 U18259 ( .B1(n9694), .B2(n19052), .A(n14945), .ZN(n14946) );
  OAI21_X1 U18260 ( .B1(n15159), .B2(n15995), .A(n14946), .ZN(P2_U2985) );
  INV_X1 U18261 ( .A(n14950), .ZN(n14952) );
  OAI22_X1 U18262 ( .A1(n14963), .A2(n15173), .B1(n14952), .B2(n14951), .ZN(
        n14955) );
  XNOR2_X1 U18263 ( .A(n14953), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14954) );
  XNOR2_X1 U18264 ( .A(n14955), .B(n14954), .ZN(n15171) );
  INV_X1 U18265 ( .A(n15921), .ZN(n14962) );
  NOR2_X1 U18266 ( .A1(n14056), .A2(n14956), .ZN(n15160) );
  AOI21_X1 U18267 ( .B1(n15105), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15160), .ZN(n14957) );
  OAI21_X1 U18268 ( .B1(n15144), .B2(n14958), .A(n14957), .ZN(n14961) );
  OR2_X2 U18269 ( .A1(n14964), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14960) );
  XNOR2_X1 U18270 ( .A(n14963), .B(n15173), .ZN(n15184) );
  AOI21_X1 U18271 ( .B1(n15173), .B2(n14972), .A(n14964), .ZN(n15181) );
  NAND2_X1 U18272 ( .A1(n15392), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15175) );
  OAI21_X1 U18273 ( .B1(n19061), .B2(n14965), .A(n15175), .ZN(n14966) );
  AOI21_X1 U18274 ( .B1(n19049), .B2(n14967), .A(n14966), .ZN(n14968) );
  OAI21_X1 U18275 ( .B1(n15172), .B2(n19057), .A(n14968), .ZN(n14969) );
  AOI21_X1 U18276 ( .B1(n15181), .B2(n19052), .A(n14969), .ZN(n14970) );
  OAI21_X1 U18277 ( .B1(n15184), .B2(n15995), .A(n14970), .ZN(P2_U2987) );
  NOR2_X1 U18278 ( .A1(n14991), .A2(n15199), .ZN(n14988) );
  OAI21_X1 U18279 ( .B1(n14988), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14972), .ZN(n15194) );
  OAI21_X1 U18280 ( .B1(n14973), .B2(n14983), .A(n14981), .ZN(n14975) );
  XNOR2_X1 U18281 ( .A(n14975), .B(n14974), .ZN(n15192) );
  NOR2_X1 U18282 ( .A1(n14056), .A2(n19649), .ZN(n15187) );
  NOR2_X1 U18283 ( .A1(n15144), .A2(n14976), .ZN(n14977) );
  AOI211_X1 U18284 ( .C1(n15105), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15187), .B(n14977), .ZN(n14978) );
  OAI21_X1 U18285 ( .B1(n15928), .B2(n19057), .A(n14978), .ZN(n14979) );
  AOI21_X1 U18286 ( .B1(n15192), .B2(n19050), .A(n14979), .ZN(n14980) );
  OAI21_X1 U18287 ( .B1(n15996), .B2(n15194), .A(n14980), .ZN(P2_U2988) );
  INV_X1 U18288 ( .A(n14981), .ZN(n14982) );
  NOR2_X1 U18289 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  XNOR2_X1 U18290 ( .A(n14973), .B(n14984), .ZN(n15206) );
  NAND2_X1 U18291 ( .A1(n19049), .A2(n15938), .ZN(n14985) );
  NAND2_X1 U18292 ( .A1(n15392), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15195) );
  OAI211_X1 U18293 ( .C1(n19061), .C2(n14986), .A(n14985), .B(n15195), .ZN(
        n14987) );
  AOI21_X1 U18294 ( .B1(n15936), .B2(n16001), .A(n14987), .ZN(n14990) );
  INV_X1 U18295 ( .A(n14988), .ZN(n15203) );
  NAND2_X1 U18296 ( .A1(n14991), .A2(n15199), .ZN(n15202) );
  NAND3_X1 U18297 ( .A1(n15203), .A2(n19052), .A3(n15202), .ZN(n14989) );
  OAI211_X1 U18298 ( .C1(n15206), .C2(n15995), .A(n14990), .B(n14989), .ZN(
        P2_U2989) );
  OAI21_X1 U18299 ( .B1(n15000), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14991), .ZN(n15216) );
  XNOR2_X1 U18300 ( .A(n14992), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14993) );
  XNOR2_X1 U18301 ( .A(n14994), .B(n14993), .ZN(n15214) );
  NOR2_X1 U18302 ( .A1(n15952), .A2(n19057), .ZN(n14998) );
  NAND2_X1 U18303 ( .A1(n15127), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15209) );
  NAND2_X1 U18304 ( .A1(n15105), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14995) );
  OAI211_X1 U18305 ( .C1(n15144), .C2(n14996), .A(n15209), .B(n14995), .ZN(
        n14997) );
  AOI211_X1 U18306 ( .C1(n15214), .C2(n19050), .A(n14998), .B(n14997), .ZN(
        n14999) );
  OAI21_X1 U18307 ( .B1(n15996), .B2(n15216), .A(n14999), .ZN(P2_U2990) );
  INV_X1 U18308 ( .A(n15000), .ZN(n15001) );
  OAI21_X1 U18309 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15012), .A(
        n15001), .ZN(n15230) );
  XOR2_X1 U18310 ( .A(n15003), .B(n15002), .Z(n15217) );
  NAND2_X1 U18311 ( .A1(n15392), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15223) );
  OAI21_X1 U18312 ( .B1(n19061), .B2(n15004), .A(n15223), .ZN(n15005) );
  AOI21_X1 U18313 ( .B1(n19049), .B2(n15006), .A(n15005), .ZN(n15007) );
  OAI21_X1 U18314 ( .B1(n15218), .B2(n19057), .A(n15007), .ZN(n15008) );
  AOI21_X1 U18315 ( .B1(n15217), .B2(n19050), .A(n15008), .ZN(n15009) );
  OAI21_X1 U18316 ( .B1(n15996), .B2(n15230), .A(n15009), .ZN(P2_U2991) );
  NOR2_X1 U18317 ( .A1(n15010), .A2(n15011), .ZN(n15032) );
  OAI21_X1 U18318 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15032), .A(
        n9877), .ZN(n15242) );
  NAND2_X1 U18319 ( .A1(n9699), .A2(n15014), .ZN(n15015) );
  XNOR2_X1 U18320 ( .A(n15013), .B(n15015), .ZN(n15240) );
  NOR2_X1 U18321 ( .A1(n15537), .A2(n19057), .ZN(n15019) );
  NAND2_X1 U18322 ( .A1(n15127), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n15232) );
  NAND2_X1 U18323 ( .A1(n15105), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15016) );
  OAI211_X1 U18324 ( .C1(n15144), .C2(n15017), .A(n15232), .B(n15016), .ZN(
        n15018) );
  AOI211_X1 U18325 ( .C1(n15240), .C2(n19050), .A(n15019), .B(n15018), .ZN(
        n15020) );
  OAI21_X1 U18326 ( .B1(n15242), .B2(n15996), .A(n15020), .ZN(P2_U2992) );
  NAND2_X1 U18327 ( .A1(n15022), .A2(n15021), .ZN(n15031) );
  OAI21_X2 U18328 ( .B1(n15025), .B2(n15024), .A(n15023), .ZN(n15063) );
  INV_X1 U18329 ( .A(n15063), .ZN(n15028) );
  INV_X1 U18330 ( .A(n15026), .ZN(n15049) );
  INV_X1 U18331 ( .A(n15037), .ZN(n15029) );
  OAI21_X1 U18332 ( .B1(n15040), .B2(n15029), .A(n15038), .ZN(n15030) );
  XOR2_X1 U18333 ( .A(n15031), .B(n15030), .Z(n15253) );
  OR2_X1 U18334 ( .A1(n15010), .A2(n15261), .ZN(n15041) );
  AOI21_X1 U18335 ( .B1(n15245), .B2(n15041), .A(n15032), .ZN(n15251) );
  NAND2_X1 U18336 ( .A1(n15127), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15243) );
  OAI21_X1 U18337 ( .B1(n19061), .B2(n18659), .A(n15243), .ZN(n15033) );
  AOI21_X1 U18338 ( .B1(n19049), .B2(n18656), .A(n15033), .ZN(n15034) );
  OAI21_X1 U18339 ( .B1(n18661), .B2(n19057), .A(n15034), .ZN(n15035) );
  AOI21_X1 U18340 ( .B1(n15251), .B2(n19052), .A(n15035), .ZN(n15036) );
  OAI21_X1 U18341 ( .B1(n15253), .B2(n15995), .A(n15036), .ZN(P2_U2993) );
  NAND2_X1 U18342 ( .A1(n15038), .A2(n15037), .ZN(n15039) );
  XNOR2_X1 U18343 ( .A(n15040), .B(n15039), .ZN(n15268) );
  INV_X1 U18344 ( .A(n15041), .ZN(n15042) );
  AOI21_X1 U18345 ( .B1(n15261), .B2(n15010), .A(n15042), .ZN(n15266) );
  NOR2_X1 U18346 ( .A1(n18678), .A2(n19057), .ZN(n15046) );
  NAND2_X1 U18347 ( .A1(n15127), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15258) );
  NAND2_X1 U18348 ( .A1(n15105), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15043) );
  OAI211_X1 U18349 ( .C1(n15144), .C2(n15044), .A(n15258), .B(n15043), .ZN(
        n15045) );
  AOI211_X1 U18350 ( .C1(n15266), .C2(n19052), .A(n15046), .B(n15045), .ZN(
        n15047) );
  OAI21_X1 U18351 ( .B1(n15268), .B2(n15995), .A(n15047), .ZN(P2_U2994) );
  NAND2_X1 U18352 ( .A1(n15049), .A2(n15048), .ZN(n15052) );
  INV_X1 U18353 ( .A(n15061), .ZN(n15050) );
  OAI21_X1 U18354 ( .B1(n15063), .B2(n15050), .A(n15060), .ZN(n15051) );
  XOR2_X1 U18355 ( .A(n15052), .B(n15051), .Z(n15279) );
  INV_X1 U18356 ( .A(n15053), .ZN(n18687) );
  NOR2_X1 U18357 ( .A1(n14056), .A2(n19637), .ZN(n15270) );
  AOI21_X1 U18358 ( .B1(n15105), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15270), .ZN(n15054) );
  OAI21_X1 U18359 ( .B1(n15055), .B2(n15144), .A(n15054), .ZN(n15058) );
  AND2_X1 U18360 ( .A1(n12470), .A2(n15056), .ZN(n15064) );
  OAI21_X1 U18361 ( .B1(n15064), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15010), .ZN(n15275) );
  NOR2_X1 U18362 ( .A1(n15275), .A2(n15996), .ZN(n15057) );
  AOI211_X1 U18363 ( .C1(n16001), .C2(n18687), .A(n15058), .B(n15057), .ZN(
        n15059) );
  OAI21_X1 U18364 ( .B1(n15279), .B2(n15995), .A(n15059), .ZN(P2_U2995) );
  NAND2_X1 U18365 ( .A1(n15061), .A2(n15060), .ZN(n15062) );
  XNOR2_X1 U18366 ( .A(n15063), .B(n15062), .ZN(n15295) );
  INV_X1 U18367 ( .A(n15284), .ZN(n15288) );
  NAND2_X1 U18368 ( .A1(n9678), .A2(n15288), .ZN(n15075) );
  AOI21_X1 U18369 ( .B1(n15075), .B2(n15065), .A(n15064), .ZN(n15293) );
  NOR2_X1 U18370 ( .A1(n14056), .A2(n15066), .ZN(n15286) );
  NOR2_X1 U18371 ( .A1(n15144), .A2(n15067), .ZN(n15068) );
  AOI211_X1 U18372 ( .C1(n15105), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15286), .B(n15068), .ZN(n15069) );
  OAI21_X1 U18373 ( .B1(n18698), .B2(n19057), .A(n15069), .ZN(n15070) );
  AOI21_X1 U18374 ( .B1(n15293), .B2(n19052), .A(n15070), .ZN(n15071) );
  OAI21_X1 U18375 ( .B1(n15295), .B2(n15995), .A(n15071), .ZN(P2_U2996) );
  NAND2_X1 U18376 ( .A1(n15105), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15072) );
  OAI211_X1 U18377 ( .C1(n15144), .C2(n18705), .A(n15073), .B(n15072), .ZN(
        n15074) );
  AOI21_X1 U18378 ( .B1(n18703), .B2(n16001), .A(n15074), .ZN(n15077) );
  OAI211_X1 U18379 ( .C1(n15084), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19052), .B(n15075), .ZN(n15076) );
  OAI211_X1 U18380 ( .C1(n15078), .C2(n15995), .A(n15077), .B(n15076), .ZN(
        P2_U2997) );
  XOR2_X1 U18381 ( .A(n15080), .B(n15079), .Z(n15309) );
  INV_X1 U18382 ( .A(n15309), .ZN(n15089) );
  INV_X1 U18383 ( .A(n18712), .ZN(n15082) );
  INV_X1 U18384 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19632) );
  NOR2_X1 U18385 ( .A1(n14056), .A2(n19632), .ZN(n15304) );
  AOI21_X1 U18386 ( .B1(n15105), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15304), .ZN(n15081) );
  OAI21_X1 U18387 ( .B1(n15144), .B2(n15082), .A(n15081), .ZN(n15087) );
  INV_X1 U18388 ( .A(n15298), .ZN(n15083) );
  AOI21_X1 U18389 ( .B1(n15083), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15085) );
  NOR3_X1 U18390 ( .A1(n15085), .A2(n15084), .A3(n15996), .ZN(n15086) );
  AOI211_X1 U18391 ( .C1(n18716), .C2(n16001), .A(n15087), .B(n15086), .ZN(
        n15088) );
  OAI21_X1 U18392 ( .B1(n15089), .B2(n15995), .A(n15088), .ZN(P2_U2998) );
  XNOR2_X1 U18393 ( .A(n15298), .B(n15090), .ZN(n15326) );
  NAND2_X1 U18394 ( .A1(n15092), .A2(n15091), .ZN(n15093) );
  XNOR2_X1 U18395 ( .A(n15094), .B(n15093), .ZN(n15324) );
  NOR2_X1 U18396 ( .A1(n18725), .A2(n19057), .ZN(n15097) );
  NAND2_X1 U18397 ( .A1(n15127), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15317) );
  NAND2_X1 U18398 ( .A1(n15105), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15095) );
  OAI211_X1 U18399 ( .C1(n15144), .C2(n18722), .A(n15317), .B(n15095), .ZN(
        n15096) );
  AOI211_X1 U18400 ( .C1(n15324), .C2(n19050), .A(n15097), .B(n15096), .ZN(
        n15098) );
  OAI21_X1 U18401 ( .B1(n15996), .B2(n15326), .A(n15098), .ZN(P2_U2999) );
  NAND2_X1 U18402 ( .A1(n9678), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15357) );
  OAI21_X1 U18403 ( .B1(n15357), .B2(n15346), .A(n15335), .ZN(n15099) );
  NAND2_X1 U18404 ( .A1(n15099), .A2(n15298), .ZN(n15340) );
  NAND2_X1 U18405 ( .A1(n15101), .A2(n15100), .ZN(n15103) );
  XOR2_X1 U18406 ( .A(n15103), .B(n15102), .Z(n15338) );
  NOR2_X1 U18407 ( .A1(n14056), .A2(n19628), .ZN(n15333) );
  NOR2_X1 U18408 ( .A1(n15144), .A2(n18735), .ZN(n15104) );
  AOI211_X1 U18409 ( .C1(n15105), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15333), .B(n15104), .ZN(n15106) );
  OAI21_X1 U18410 ( .B1(n18740), .B2(n19057), .A(n15106), .ZN(n15107) );
  AOI21_X1 U18411 ( .B1(n15338), .B2(n19050), .A(n15107), .ZN(n15108) );
  OAI21_X1 U18412 ( .B1(n15996), .B2(n15340), .A(n15108), .ZN(P2_U3000) );
  NOR2_X1 U18413 ( .A1(n15109), .A2(n15122), .ZN(n15113) );
  NOR2_X1 U18414 ( .A1(n15111), .A2(n15110), .ZN(n15112) );
  XNOR2_X1 U18415 ( .A(n15113), .B(n15112), .ZN(n15345) );
  XNOR2_X1 U18416 ( .A(n15357), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15341) );
  NAND2_X1 U18417 ( .A1(n15341), .A2(n19052), .ZN(n15117) );
  NAND2_X1 U18418 ( .A1(n15127), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15351) );
  OAI21_X1 U18419 ( .B1(n19061), .B2(n18742), .A(n15351), .ZN(n15115) );
  NOR2_X1 U18420 ( .A1(n18747), .A2(n19057), .ZN(n15114) );
  AOI211_X1 U18421 ( .C1(n19049), .C2(n18746), .A(n15115), .B(n15114), .ZN(
        n15116) );
  OAI211_X1 U18422 ( .C1(n15995), .C2(n15345), .A(n15117), .B(n15116), .ZN(
        P2_U3001) );
  NAND2_X1 U18423 ( .A1(n15118), .A2(n15119), .ZN(n15121) );
  NAND2_X1 U18424 ( .A1(n15121), .A2(n15120), .ZN(n15125) );
  NAND2_X1 U18425 ( .A1(n10512), .A2(n15123), .ZN(n15124) );
  XNOR2_X1 U18426 ( .A(n15125), .B(n15124), .ZN(n15370) );
  INV_X1 U18427 ( .A(n9678), .ZN(n15132) );
  NAND2_X1 U18428 ( .A1(n15132), .A2(n15126), .ZN(n15358) );
  NAND3_X1 U18429 ( .A1(n15358), .A2(n19052), .A3(n15357), .ZN(n15131) );
  NAND2_X1 U18430 ( .A1(n15127), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n15364) );
  OAI21_X1 U18431 ( .B1(n19061), .B2(n18753), .A(n15364), .ZN(n15129) );
  NOR2_X1 U18432 ( .A1(n18762), .A2(n19057), .ZN(n15128) );
  AOI211_X1 U18433 ( .C1(n19049), .C2(n18757), .A(n15129), .B(n15128), .ZN(
        n15130) );
  OAI211_X1 U18434 ( .C1(n15995), .C2(n15370), .A(n15131), .B(n15130), .ZN(
        P2_U3002) );
  NOR2_X1 U18435 ( .A1(n9669), .A2(n16012), .ZN(n15982) );
  OAI21_X1 U18436 ( .B1(n15982), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15132), .ZN(n15384) );
  AND2_X1 U18437 ( .A1(n15392), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n15375) );
  OAI22_X1 U18438 ( .A1(n19061), .A2(n10766), .B1(n15144), .B2(n18775), .ZN(
        n15133) );
  AOI211_X1 U18439 ( .C1(n18769), .C2(n16001), .A(n15375), .B(n15133), .ZN(
        n15139) );
  NAND2_X1 U18440 ( .A1(n15118), .A2(n15134), .ZN(n15137) );
  XNOR2_X1 U18441 ( .A(n15135), .B(n15371), .ZN(n15136) );
  XNOR2_X1 U18442 ( .A(n15137), .B(n15136), .ZN(n15381) );
  NAND2_X1 U18443 ( .A1(n15381), .A2(n19050), .ZN(n15138) );
  OAI211_X1 U18444 ( .C1(n15384), .C2(n15996), .A(n15139), .B(n15138), .ZN(
        P2_U3003) );
  OAI21_X1 U18445 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n12470), .A(
        n9669), .ZN(n15397) );
  NAND2_X1 U18446 ( .A1(n15141), .A2(n15140), .ZN(n15993) );
  INV_X1 U18447 ( .A(n15142), .ZN(n15992) );
  AOI21_X1 U18448 ( .B1(n15993), .B2(n9947), .A(n15992), .ZN(n15977) );
  NAND2_X1 U18449 ( .A1(n15974), .A2(n15976), .ZN(n15143) );
  XNOR2_X1 U18450 ( .A(n15977), .B(n15143), .ZN(n15395) );
  INV_X1 U18451 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15145) );
  OAI22_X1 U18452 ( .A1(n19061), .A2(n15145), .B1(n15144), .B2(n18790), .ZN(
        n15146) );
  AOI21_X1 U18453 ( .B1(n15392), .B2(P2_REIP_REG_9__SCAN_IN), .A(n15146), .ZN(
        n15147) );
  OAI21_X1 U18454 ( .B1(n18793), .B2(n19057), .A(n15147), .ZN(n15148) );
  AOI21_X1 U18455 ( .B1(n15395), .B2(n19050), .A(n15148), .ZN(n15149) );
  OAI21_X1 U18456 ( .B1(n15397), .B2(n15996), .A(n15149), .ZN(P2_U3005) );
  NOR2_X1 U18457 ( .A1(n15906), .A2(n16008), .ZN(n15157) );
  OR2_X1 U18458 ( .A1(n15153), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15176) );
  AND2_X1 U18459 ( .A1(n15174), .A2(n15176), .ZN(n15165) );
  OAI21_X1 U18460 ( .B1(n15173), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15150) );
  OAI21_X1 U18461 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n15150), .ZN(n15152) );
  OAI21_X1 U18462 ( .B1(n15153), .B2(n15152), .A(n15151), .ZN(n15154) );
  OAI21_X1 U18463 ( .B1(n15159), .B2(n16034), .A(n15158), .ZN(P2_U3017) );
  AOI21_X1 U18464 ( .B1(n15161), .B2(n15164), .A(n15160), .ZN(n15163) );
  NAND2_X1 U18465 ( .A1(n15918), .A2(n15354), .ZN(n15162) );
  OAI211_X1 U18466 ( .C1(n15165), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15166) );
  INV_X1 U18467 ( .A(n15166), .ZN(n15168) );
  INV_X1 U18468 ( .A(n15169), .ZN(n15170) );
  OAI21_X1 U18469 ( .B1(n15171), .B2(n16034), .A(n15170), .ZN(P2_U3018) );
  INV_X1 U18470 ( .A(n15172), .ZN(n15180) );
  NOR2_X1 U18471 ( .A1(n15174), .A2(n15173), .ZN(n15179) );
  OAI211_X1 U18472 ( .C1(n15177), .C2(n16036), .A(n15176), .B(n15175), .ZN(
        n15178) );
  AOI211_X1 U18473 ( .C1(n15180), .C2(n16038), .A(n15179), .B(n15178), .ZN(
        n15183) );
  NAND2_X1 U18474 ( .A1(n15181), .A2(n10731), .ZN(n15182) );
  OAI211_X1 U18475 ( .C1(n15184), .C2(n16034), .A(n15183), .B(n15182), .ZN(
        P2_U3019) );
  NOR2_X1 U18476 ( .A1(n15928), .A2(n16008), .ZN(n15191) );
  INV_X1 U18477 ( .A(n15185), .ZN(n15931) );
  AOI211_X1 U18478 ( .C1(n15189), .C2(n15199), .A(n15196), .B(n10728), .ZN(
        n15186) );
  AOI211_X1 U18479 ( .C1(n15931), .C2(n15354), .A(n15187), .B(n15186), .ZN(
        n15188) );
  OAI21_X1 U18480 ( .B1(n15200), .B2(n15189), .A(n15188), .ZN(n15190) );
  AOI211_X1 U18481 ( .C1(n15192), .C2(n16044), .A(n15191), .B(n15190), .ZN(
        n15193) );
  OAI21_X1 U18482 ( .B1(n16040), .B2(n15194), .A(n15193), .ZN(P2_U3020) );
  OAI21_X1 U18483 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15196), .A(
        n15195), .ZN(n15197) );
  AOI21_X1 U18484 ( .B1(n15935), .B2(n15354), .A(n15197), .ZN(n15198) );
  OAI21_X1 U18485 ( .B1(n15200), .B2(n15199), .A(n15198), .ZN(n15201) );
  AOI21_X1 U18486 ( .B1(n15936), .B2(n16038), .A(n15201), .ZN(n15205) );
  NAND3_X1 U18487 ( .A1(n15203), .A2(n10731), .A3(n15202), .ZN(n15204) );
  OAI211_X1 U18488 ( .C1(n15206), .C2(n16034), .A(n15205), .B(n15204), .ZN(
        P2_U3021) );
  NOR2_X1 U18489 ( .A1(n15952), .A2(n16008), .ZN(n15213) );
  INV_X1 U18490 ( .A(n15955), .ZN(n15211) );
  OAI21_X1 U18491 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15208), .A(
        n15207), .ZN(n15210) );
  OAI211_X1 U18492 ( .C1(n16036), .C2(n15211), .A(n15210), .B(n15209), .ZN(
        n15212) );
  AOI211_X1 U18493 ( .C1(n15214), .C2(n16044), .A(n15213), .B(n15212), .ZN(
        n15215) );
  OAI21_X1 U18494 ( .B1(n16040), .B2(n15216), .A(n15215), .ZN(P2_U3022) );
  NAND2_X1 U18495 ( .A1(n15217), .A2(n16044), .ZN(n15229) );
  INV_X1 U18496 ( .A(n15218), .ZN(n15227) );
  NOR2_X1 U18497 ( .A1(n15235), .A2(n15219), .ZN(n15226) );
  INV_X1 U18498 ( .A(n15233), .ZN(n15221) );
  OAI211_X1 U18499 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15221), .B(n15220), .ZN(
        n15222) );
  OAI211_X1 U18500 ( .C1(n16036), .C2(n15224), .A(n15223), .B(n15222), .ZN(
        n15225) );
  AOI211_X1 U18501 ( .C1(n15227), .C2(n16038), .A(n15226), .B(n15225), .ZN(
        n15228) );
  OAI211_X1 U18502 ( .C1(n15230), .C2(n16040), .A(n15229), .B(n15228), .ZN(
        P2_U3023) );
  AOI21_X1 U18503 ( .B1(n15231), .B2(n9671), .A(n13199), .ZN(n15958) );
  OAI21_X1 U18504 ( .B1(n15233), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15232), .ZN(n15237) );
  NOR2_X1 U18505 ( .A1(n15235), .A2(n15234), .ZN(n15236) );
  AOI211_X1 U18506 ( .C1(n15354), .C2(n15958), .A(n15237), .B(n15236), .ZN(
        n15238) );
  OAI21_X1 U18507 ( .B1(n16008), .B2(n15537), .A(n15238), .ZN(n15239) );
  AOI21_X1 U18508 ( .B1(n15240), .B2(n16044), .A(n15239), .ZN(n15241) );
  OAI21_X1 U18509 ( .B1(n15242), .B2(n16040), .A(n15241), .ZN(P2_U3024) );
  OAI21_X1 U18510 ( .B1(n15244), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15243), .ZN(n15248) );
  NOR2_X1 U18511 ( .A1(n15246), .A2(n15245), .ZN(n15247) );
  AOI211_X1 U18512 ( .C1(n15354), .C2(n18662), .A(n15248), .B(n15247), .ZN(
        n15249) );
  OAI21_X1 U18513 ( .B1(n16008), .B2(n18661), .A(n15249), .ZN(n15250) );
  AOI21_X1 U18514 ( .B1(n15251), .B2(n10731), .A(n15250), .ZN(n15252) );
  OAI21_X1 U18515 ( .B1(n15253), .B2(n16034), .A(n15252), .ZN(P2_U3025) );
  INV_X1 U18516 ( .A(n15254), .ZN(n15257) );
  INV_X1 U18517 ( .A(n14925), .ZN(n15255) );
  AOI21_X1 U18518 ( .B1(n15257), .B2(n15256), .A(n15255), .ZN(n18676) );
  INV_X1 U18519 ( .A(n15271), .ZN(n15260) );
  XNOR2_X1 U18520 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15259) );
  OAI21_X1 U18521 ( .B1(n15260), .B2(n15259), .A(n15258), .ZN(n15263) );
  NOR2_X1 U18522 ( .A1(n15274), .A2(n15261), .ZN(n15262) );
  AOI211_X1 U18523 ( .C1(n15354), .C2(n18676), .A(n15263), .B(n15262), .ZN(
        n15264) );
  OAI21_X1 U18524 ( .B1(n18678), .B2(n16008), .A(n15264), .ZN(n15265) );
  AOI21_X1 U18525 ( .B1(n15266), .B2(n10731), .A(n15265), .ZN(n15267) );
  OAI21_X1 U18526 ( .B1(n15268), .B2(n16034), .A(n15267), .ZN(P2_U3026) );
  NOR2_X1 U18527 ( .A1(n16036), .A2(n18689), .ZN(n15269) );
  AOI211_X1 U18528 ( .C1(n15271), .C2(n15273), .A(n15270), .B(n15269), .ZN(
        n15272) );
  OAI21_X1 U18529 ( .B1(n15274), .B2(n15273), .A(n15272), .ZN(n15277) );
  NOR2_X1 U18530 ( .A1(n15275), .A2(n16040), .ZN(n15276) );
  AOI211_X1 U18531 ( .C1(n18687), .C2(n16038), .A(n15277), .B(n15276), .ZN(
        n15278) );
  OAI21_X1 U18532 ( .B1(n15279), .B2(n16034), .A(n15278), .ZN(P2_U3027) );
  NAND2_X1 U18533 ( .A1(n15281), .A2(n15280), .ZN(n15282) );
  NOR3_X1 U18534 ( .A1(n15284), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15344), .ZN(n15285) );
  AOI211_X1 U18535 ( .C1(n15354), .C2(n9995), .A(n15286), .B(n15285), .ZN(
        n15291) );
  NOR2_X1 U18536 ( .A1(n16014), .A2(n15287), .ZN(n15367) );
  NOR2_X1 U18537 ( .A1(n16014), .A2(n15288), .ZN(n15289) );
  OAI21_X1 U18538 ( .B1(n15367), .B2(n15289), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15290) );
  OAI211_X1 U18539 ( .C1(n18698), .C2(n16008), .A(n15291), .B(n15290), .ZN(
        n15292) );
  AOI21_X1 U18540 ( .B1(n15293), .B2(n10731), .A(n15292), .ZN(n15294) );
  OAI21_X1 U18541 ( .B1(n15295), .B2(n16034), .A(n15294), .ZN(P2_U3028) );
  NAND2_X1 U18542 ( .A1(n15297), .A2(n15296), .ZN(n15318) );
  OAI21_X1 U18543 ( .B1(n15298), .B2(n16040), .A(n15318), .ZN(n15299) );
  NAND3_X1 U18544 ( .A1(n15299), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n15311), .ZN(n15306) );
  OR2_X1 U18545 ( .A1(n15301), .A2(n15300), .ZN(n15302) );
  AND2_X1 U18546 ( .A1(n15303), .A2(n15302), .ZN(n18885) );
  AOI21_X1 U18547 ( .B1(n15354), .B2(n18885), .A(n15304), .ZN(n15305) );
  OAI211_X1 U18548 ( .C1(n16008), .C2(n15307), .A(n15306), .B(n15305), .ZN(
        n15308) );
  AOI21_X1 U18549 ( .B1(n15309), .B2(n16044), .A(n15308), .ZN(n15310) );
  OAI21_X1 U18550 ( .B1(n15312), .B2(n15311), .A(n15310), .ZN(P2_U3030) );
  OR2_X1 U18551 ( .A1(n15313), .A2(n15314), .ZN(n15316) );
  NAND2_X1 U18552 ( .A1(n15316), .A2(n15315), .ZN(n18893) );
  NOR2_X1 U18553 ( .A1(n16036), .A2(n18893), .ZN(n15320) );
  OAI21_X1 U18554 ( .B1(n15318), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15317), .ZN(n15319) );
  AOI211_X1 U18555 ( .C1(n15321), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15320), .B(n15319), .ZN(n15322) );
  OAI21_X1 U18556 ( .B1(n18725), .B2(n16008), .A(n15322), .ZN(n15323) );
  AOI21_X1 U18557 ( .B1(n15324), .B2(n16044), .A(n15323), .ZN(n15325) );
  OAI21_X1 U18558 ( .B1(n16040), .B2(n15326), .A(n15325), .ZN(P2_U3031) );
  NOR2_X1 U18559 ( .A1(n18740), .A2(n16008), .ZN(n15337) );
  NOR2_X1 U18560 ( .A1(n15344), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15362) );
  NOR2_X1 U18561 ( .A1(n15367), .A2(n15362), .ZN(n15347) );
  NOR2_X1 U18562 ( .A1(n15327), .A2(n15328), .ZN(n15329) );
  OR2_X1 U18563 ( .A1(n15313), .A2(n15329), .ZN(n18896) );
  INV_X1 U18564 ( .A(n18896), .ZN(n18737) );
  NAND2_X1 U18565 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15331) );
  NOR2_X1 U18566 ( .A1(n15346), .A2(n15335), .ZN(n15330) );
  AOI211_X1 U18567 ( .C1(n15331), .C2(n15335), .A(n15330), .B(n15344), .ZN(
        n15332) );
  AOI211_X1 U18568 ( .C1(n15354), .C2(n18737), .A(n15333), .B(n15332), .ZN(
        n15334) );
  OAI21_X1 U18569 ( .B1(n15347), .B2(n15335), .A(n15334), .ZN(n15336) );
  AOI211_X1 U18570 ( .C1(n15338), .C2(n16044), .A(n15337), .B(n15336), .ZN(
        n15339) );
  OAI21_X1 U18571 ( .B1(n16040), .B2(n15340), .A(n15339), .ZN(P2_U3032) );
  NAND2_X1 U18572 ( .A1(n15341), .A2(n10731), .ZN(n15356) );
  AND2_X1 U18573 ( .A1(n9665), .A2(n15342), .ZN(n15343) );
  OR2_X1 U18574 ( .A1(n15343), .A2(n15327), .ZN(n18897) );
  INV_X1 U18575 ( .A(n18897), .ZN(n15353) );
  NOR2_X1 U18576 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15344), .ZN(
        n15349) );
  OAI22_X1 U18577 ( .A1(n15347), .A2(n15346), .B1(n16034), .B2(n15345), .ZN(
        n15348) );
  AOI21_X1 U18578 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15349), .A(
        n15348), .ZN(n15350) );
  NAND2_X1 U18579 ( .A1(n15351), .A2(n15350), .ZN(n15352) );
  AOI21_X1 U18580 ( .B1(n15354), .B2(n15353), .A(n15352), .ZN(n15355) );
  OAI211_X1 U18581 ( .C1(n18747), .C2(n16008), .A(n15356), .B(n15355), .ZN(
        P2_U3033) );
  NAND3_X1 U18582 ( .A1(n15358), .A2(n10731), .A3(n15357), .ZN(n15369) );
  NAND2_X1 U18583 ( .A1(n15360), .A2(n15359), .ZN(n15361) );
  AND2_X1 U18584 ( .A1(n9665), .A2(n15361), .ZN(n18759) );
  INV_X1 U18585 ( .A(n18759), .ZN(n18900) );
  INV_X1 U18586 ( .A(n15362), .ZN(n15363) );
  OAI211_X1 U18587 ( .C1(n16036), .C2(n18900), .A(n15364), .B(n15363), .ZN(
        n15366) );
  NOR2_X1 U18588 ( .A1(n18762), .A2(n16008), .ZN(n15365) );
  AOI211_X1 U18589 ( .C1(n15367), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15366), .B(n15365), .ZN(n15368) );
  OAI211_X1 U18590 ( .C1(n15370), .C2(n16034), .A(n15369), .B(n15368), .ZN(
        P2_U3034) );
  NOR3_X1 U18591 ( .A1(n16014), .A2(n16013), .A3(n15371), .ZN(n15380) );
  OR2_X1 U18592 ( .A1(n15373), .A2(n15372), .ZN(n15374) );
  NAND2_X1 U18593 ( .A1(n15359), .A2(n15374), .ZN(n18901) );
  INV_X1 U18594 ( .A(n15375), .ZN(n15378) );
  OAI211_X1 U18595 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n9793), .B(n16011), .ZN(n15377) );
  OAI211_X1 U18596 ( .C1(n16036), .C2(n18901), .A(n15378), .B(n15377), .ZN(
        n15379) );
  AOI211_X1 U18597 ( .C1(n18769), .C2(n16038), .A(n15380), .B(n15379), .ZN(
        n15383) );
  NAND2_X1 U18598 ( .A1(n15381), .A2(n16044), .ZN(n15382) );
  OAI211_X1 U18599 ( .C1(n15384), .C2(n16040), .A(n15383), .B(n15382), .ZN(
        P2_U3035) );
  AOI21_X1 U18600 ( .B1(n9792), .B2(n15385), .A(n16013), .ZN(n15391) );
  OR2_X1 U18601 ( .A1(n15387), .A2(n15386), .ZN(n15389) );
  NAND2_X1 U18602 ( .A1(n15389), .A2(n15388), .ZN(n18907) );
  NOR2_X1 U18603 ( .A1(n16036), .A2(n18907), .ZN(n15390) );
  AOI211_X1 U18604 ( .C1(n15392), .C2(P2_REIP_REG_9__SCAN_IN), .A(n15391), .B(
        n15390), .ZN(n15393) );
  OAI21_X1 U18605 ( .B1(n18793), .B2(n16008), .A(n15393), .ZN(n15394) );
  AOI21_X1 U18606 ( .B1(n15395), .B2(n16044), .A(n15394), .ZN(n15396) );
  OAI21_X1 U18607 ( .B1(n15397), .B2(n16040), .A(n15396), .ZN(P2_U3037) );
  OR2_X1 U18608 ( .A1(n15399), .A2(n15398), .ZN(n15403) );
  MUX2_X1 U18609 ( .A(n15400), .B(n13450), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15401) );
  INV_X1 U18610 ( .A(n15401), .ZN(n15402) );
  NAND2_X1 U18611 ( .A1(n15403), .A2(n15402), .ZN(n16075) );
  AOI21_X1 U18612 ( .B1(n16075), .B2(n19697), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n15406) );
  INV_X1 U18613 ( .A(n16049), .ZN(n15404) );
  OAI22_X1 U18614 ( .A1(n15407), .A2(n15406), .B1(n15405), .B2(n15404), .ZN(
        n15408) );
  MUX2_X1 U18615 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15408), .S(
        n15504), .Z(P2_U3601) );
  NAND2_X1 U18616 ( .A1(n17989), .A2(n16783), .ZN(n16766) );
  NAND2_X1 U18617 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16715), .ZN(n16702) );
  INV_X1 U18618 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n20777) );
  NAND2_X1 U18619 ( .A1(n17989), .A2(n9588), .ZN(n16973) );
  INV_X1 U18620 ( .A(n16973), .ZN(n16986) );
  NOR2_X1 U18621 ( .A1(n16715), .A2(n16987), .ZN(n16713) );
  AOI21_X1 U18622 ( .B1(n16986), .B2(n15411), .A(n16713), .ZN(n16701) );
  AOI22_X1 U18623 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15415) );
  AOI22_X1 U18624 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U18625 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12172), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U18626 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15412) );
  NAND4_X1 U18627 ( .A1(n15415), .A2(n15414), .A3(n15413), .A4(n15412), .ZN(
        n15421) );
  AOI22_X1 U18628 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U18629 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U18630 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U18631 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15416) );
  NAND4_X1 U18632 ( .A1(n15419), .A2(n15418), .A3(n15417), .A4(n15416), .ZN(
        n15420) );
  NOR2_X1 U18633 ( .A1(n15421), .A2(n15420), .ZN(n15485) );
  AOI22_X1 U18634 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12172), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15425) );
  AOI22_X1 U18635 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15424) );
  AOI22_X1 U18636 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15423) );
  AOI22_X1 U18637 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15422) );
  NAND4_X1 U18638 ( .A1(n15425), .A2(n15424), .A3(n15423), .A4(n15422), .ZN(
        n15431) );
  AOI22_X1 U18639 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15429) );
  AOI22_X1 U18640 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12207), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U18641 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9601), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15427) );
  AOI22_X1 U18642 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15426) );
  NAND4_X1 U18643 ( .A1(n15429), .A2(n15428), .A3(n15427), .A4(n15426), .ZN(
        n15430) );
  NOR2_X1 U18644 ( .A1(n15431), .A2(n15430), .ZN(n16712) );
  AOI22_X1 U18645 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n16922), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n15435) );
  AOI22_X1 U18646 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12172), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15434) );
  AOI22_X1 U18647 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9602), .ZN(n15433) );
  AOI22_X1 U18648 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16933), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16936), .ZN(n15432) );
  NAND4_X1 U18649 ( .A1(n15435), .A2(n15434), .A3(n15433), .A4(n15432), .ZN(
        n15441) );
  AOI22_X1 U18650 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n9586), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n16915), .ZN(n15439) );
  AOI22_X1 U18651 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15438) );
  AOI22_X1 U18652 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15437) );
  AOI22_X1 U18653 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16917), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15436) );
  NAND4_X1 U18654 ( .A1(n15439), .A2(n15438), .A3(n15437), .A4(n15436), .ZN(
        n15440) );
  NOR2_X1 U18655 ( .A1(n15441), .A2(n15440), .ZN(n16721) );
  AOI22_X1 U18656 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U18657 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15450) );
  AOI22_X1 U18658 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15442) );
  OAI21_X1 U18659 ( .B1(n16840), .B2(n16813), .A(n15442), .ZN(n15448) );
  AOI22_X1 U18660 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15446) );
  AOI22_X1 U18661 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15445) );
  AOI22_X1 U18662 ( .A1(n16877), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15444) );
  AOI22_X1 U18663 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15443) );
  NAND4_X1 U18664 ( .A1(n15446), .A2(n15445), .A3(n15444), .A4(n15443), .ZN(
        n15447) );
  AOI211_X1 U18665 ( .C1(n16917), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n15448), .B(n15447), .ZN(n15449) );
  NAND3_X1 U18666 ( .A1(n15451), .A2(n15450), .A3(n15449), .ZN(n16725) );
  AOI22_X1 U18667 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9601), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15462) );
  AOI22_X1 U18668 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15461) );
  INV_X1 U18669 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U18670 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15452) );
  OAI21_X1 U18671 ( .B1(n15453), .B2(n16958), .A(n15452), .ZN(n15459) );
  AOI22_X1 U18672 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U18673 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U18674 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U18675 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15454) );
  NAND4_X1 U18676 ( .A1(n15457), .A2(n15456), .A3(n15455), .A4(n15454), .ZN(
        n15458) );
  AOI211_X1 U18677 ( .C1(n16945), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n15459), .B(n15458), .ZN(n15460) );
  NAND3_X1 U18678 ( .A1(n15462), .A2(n15461), .A3(n15460), .ZN(n16726) );
  NAND2_X1 U18679 ( .A1(n16725), .A2(n16726), .ZN(n16724) );
  NOR2_X1 U18680 ( .A1(n16721), .A2(n16724), .ZN(n16718) );
  AOI22_X1 U18681 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U18682 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U18683 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12172), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15463) );
  OAI21_X1 U18684 ( .B1(n16840), .B2(n16982), .A(n15463), .ZN(n15469) );
  AOI22_X1 U18685 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15467) );
  AOI22_X1 U18686 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U18687 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15465) );
  AOI22_X1 U18688 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15464) );
  NAND4_X1 U18689 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        n15468) );
  AOI211_X1 U18690 ( .C1(n16917), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n15469), .B(n15468), .ZN(n15470) );
  NAND3_X1 U18691 ( .A1(n15472), .A2(n15471), .A3(n15470), .ZN(n16717) );
  NAND2_X1 U18692 ( .A1(n16718), .A2(n16717), .ZN(n16716) );
  NOR2_X1 U18693 ( .A1(n16712), .A2(n16716), .ZN(n16711) );
  AOI22_X1 U18694 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12207), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15484) );
  AOI22_X1 U18695 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U18696 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15474) );
  OAI21_X1 U18697 ( .B1(n12127), .B2(n20786), .A(n15474), .ZN(n15481) );
  AOI22_X1 U18698 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15479) );
  AOI22_X1 U18699 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U18700 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16917), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U18701 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15475), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15476) );
  NAND4_X1 U18702 ( .A1(n15479), .A2(n15478), .A3(n15477), .A4(n15476), .ZN(
        n15480) );
  AOI211_X1 U18703 ( .C1(n12206), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n15481), .B(n15480), .ZN(n15482) );
  NAND3_X1 U18704 ( .A1(n15484), .A2(n15483), .A3(n15482), .ZN(n16708) );
  NAND2_X1 U18705 ( .A1(n16711), .A2(n16708), .ZN(n16707) );
  NOR2_X1 U18706 ( .A1(n15485), .A2(n16707), .ZN(n16700) );
  AOI21_X1 U18707 ( .B1(n15485), .B2(n16707), .A(n16700), .ZN(n17007) );
  NAND2_X1 U18708 ( .A1(n16987), .A2(n17007), .ZN(n15486) );
  OAI221_X1 U18709 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16702), .C1(n20777), 
        .C2(n16701), .A(n15486), .ZN(P3_U2675) );
  NAND2_X1 U18710 ( .A1(n17960), .A2(n17208), .ZN(n18446) );
  INV_X1 U18711 ( .A(n18446), .ZN(n15487) );
  INV_X1 U18712 ( .A(n15508), .ZN(n18389) );
  NAND2_X1 U18713 ( .A1(n18389), .A2(n18599), .ZN(n15496) );
  AOI211_X1 U18714 ( .C1(n15492), .C2(n15491), .A(n15490), .B(n15489), .ZN(
        n15516) );
  NOR2_X1 U18715 ( .A1(n15606), .A2(n15494), .ZN(n15495) );
  OAI211_X1 U18716 ( .C1(n17142), .C2(n15496), .A(n15516), .B(n15495), .ZN(
        n18421) );
  INV_X1 U18717 ( .A(n18421), .ZN(n18431) );
  NAND2_X1 U18718 ( .A1(n18608), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17953) );
  INV_X1 U18719 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17939) );
  OR2_X1 U18720 ( .A1(n17939), .A2(n18553), .ZN(n15497) );
  INV_X1 U18721 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18395) );
  NOR2_X1 U18722 ( .A1(n15498), .A2(n18408), .ZN(n18443) );
  NAND3_X1 U18723 ( .A1(n18584), .A2(n18618), .A3(n18443), .ZN(n15499) );
  OAI21_X1 U18724 ( .B1(n18584), .B2(n18395), .A(n15499), .ZN(P3_U3284) );
  NAND4_X1 U18725 ( .A1(n15500), .A2(n16067), .A3(n19669), .A4(n16066), .ZN(
        n15501) );
  OR2_X1 U18726 ( .A1(n15502), .A2(n15501), .ZN(n15503) );
  OAI21_X1 U18727 ( .B1(n15504), .B2(n16073), .A(n15503), .ZN(P2_U3595) );
  INV_X1 U18728 ( .A(n18385), .ZN(n18416) );
  INV_X1 U18729 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17875) );
  INV_X1 U18730 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17898) );
  INV_X1 U18731 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17889) );
  NOR3_X1 U18732 ( .A1(n17875), .A2(n17898), .A3(n17889), .ZN(n17857) );
  NAND3_X1 U18733 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n17857), .ZN(n17731) );
  NOR2_X1 U18734 ( .A1(n17846), .A2(n17731), .ZN(n15505) );
  INV_X1 U18735 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18568) );
  OAI21_X1 U18736 ( .B1(n18583), .B2(n18568), .A(n17914), .ZN(n17899) );
  NAND2_X1 U18737 ( .A1(n15505), .A2(n17899), .ZN(n17743) );
  NOR2_X1 U18738 ( .A1(n17733), .A2(n17384), .ZN(n16149) );
  INV_X1 U18739 ( .A(n16149), .ZN(n16150) );
  NOR2_X1 U18740 ( .A1(n17743), .A2(n16150), .ZN(n17725) );
  NAND2_X1 U18741 ( .A1(n15506), .A2(n17725), .ZN(n15525) );
  NAND3_X1 U18742 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n15505), .ZN(n17769) );
  NOR2_X1 U18743 ( .A1(n17733), .A2(n17769), .ZN(n17678) );
  NAND2_X1 U18744 ( .A1(n15506), .A2(n17678), .ZN(n15523) );
  NAND2_X1 U18745 ( .A1(n18424), .A2(n18583), .ZN(n17916) );
  INV_X1 U18746 ( .A(n18424), .ZN(n18396) );
  NOR2_X1 U18747 ( .A1(n18409), .A2(n18396), .ZN(n17841) );
  NAND2_X1 U18748 ( .A1(n17916), .A2(n17903), .ZN(n17900) );
  OAI22_X1 U18749 ( .A1(n18416), .A2(n15525), .B1(n15523), .B2(n17900), .ZN(
        n16136) );
  NAND2_X1 U18750 ( .A1(n17108), .A2(n16156), .ZN(n17807) );
  OAI22_X1 U18751 ( .A1(n17806), .A2(n17616), .B1(n17807), .B2(n17615), .ZN(
        n15521) );
  OAI21_X1 U18752 ( .B1(n18604), .B2(n15507), .A(n18599), .ZN(n16276) );
  AOI211_X1 U18753 ( .C1(n17965), .C2(n15509), .A(n15508), .B(n16276), .ZN(
        n15520) );
  AOI21_X1 U18754 ( .B1(n17965), .B2(n15511), .A(n15510), .ZN(n15518) );
  NOR2_X1 U18755 ( .A1(n17960), .A2(n15512), .ZN(n15514) );
  NAND3_X1 U18756 ( .A1(n15514), .A2(n18390), .A3(n15513), .ZN(n15515) );
  OAI211_X1 U18757 ( .C1(n15518), .C2(n15517), .A(n15516), .B(n15515), .ZN(
        n15519) );
  OAI211_X1 U18758 ( .C1(n16136), .C2(n15521), .A(n17928), .B(n16116), .ZN(
        n15598) );
  NAND2_X1 U18759 ( .A1(n17882), .A2(n17928), .ZN(n17844) );
  INV_X1 U18760 ( .A(n17844), .ZN(n17917) );
  NOR2_X1 U18761 ( .A1(n17616), .A2(n16134), .ZN(n16117) );
  NOR2_X1 U18762 ( .A1(n17806), .A2(n17922), .ZN(n17921) );
  NAND2_X1 U18763 ( .A1(n17839), .A2(n17928), .ZN(n15522) );
  OAI22_X1 U18764 ( .A1(n16117), .A2(n17936), .B1(n16129), .B2(n15522), .ZN(
        n15595) );
  NOR2_X1 U18765 ( .A1(n18396), .A2(n18385), .ZN(n17788) );
  INV_X1 U18766 ( .A(n17788), .ZN(n17821) );
  INV_X1 U18767 ( .A(n15523), .ZN(n15527) );
  NOR2_X1 U18768 ( .A1(n18583), .A2(n17769), .ZN(n17830) );
  NAND2_X1 U18769 ( .A1(n17401), .A2(n17830), .ZN(n17698) );
  INV_X1 U18770 ( .A(n17698), .ZN(n17745) );
  NAND2_X1 U18771 ( .A1(n17618), .A2(n17745), .ZN(n17683) );
  NAND2_X1 U18772 ( .A1(n15524), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16151) );
  OAI21_X1 U18773 ( .B1(n17683), .B2(n16151), .A(n18409), .ZN(n15526) );
  NAND2_X1 U18774 ( .A1(n18385), .A2(n15525), .ZN(n17620) );
  OAI211_X1 U18775 ( .C1(n18424), .C2(n15527), .A(n15526), .B(n17620), .ZN(
        n15593) );
  AOI21_X1 U18776 ( .B1(n20690), .B2(n17821), .A(n15593), .ZN(n16159) );
  INV_X1 U18777 ( .A(n17930), .ZN(n17627) );
  OAI21_X1 U18778 ( .B1(n16159), .B2(n17922), .A(n17915), .ZN(n15528) );
  AOI211_X1 U18779 ( .C1(n17917), .C2(n16153), .A(n15595), .B(n15528), .ZN(
        n15535) );
  NOR2_X1 U18780 ( .A1(n15529), .A2(n16157), .ZN(n15531) );
  NOR2_X1 U18781 ( .A1(n15531), .A2(n15530), .ZN(n15532) );
  XNOR2_X1 U18782 ( .A(n15532), .B(n15536), .ZN(n16133) );
  INV_X1 U18783 ( .A(n16133), .ZN(n15533) );
  AOI22_X1 U18784 ( .A1(n17932), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17850), 
        .B2(n15533), .ZN(n15534) );
  OAI221_X1 U18785 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15598), 
        .C1(n15536), .C2(n15535), .A(n15534), .ZN(P3_U2833) );
  INV_X1 U18786 ( .A(n15537), .ZN(n15538) );
  AOI22_X1 U18787 ( .A1(n15538), .A2(n18868), .B1(n15958), .B2(n18859), .ZN(
        n15547) );
  AOI211_X1 U18788 ( .C1(n15541), .C2(n15540), .A(n15539), .B(n19582), .ZN(
        n15545) );
  AOI22_X1 U18789 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n18861), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18862), .ZN(n15542) );
  OAI21_X1 U18790 ( .B1(n15543), .B2(n18865), .A(n15542), .ZN(n15544) );
  AOI211_X1 U18791 ( .C1(n18842), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15545), .B(n15544), .ZN(n15546) );
  NAND2_X1 U18792 ( .A1(n15547), .A2(n15546), .ZN(P2_U2833) );
  NAND2_X1 U18793 ( .A1(n15549), .A2(n15548), .ZN(n15556) );
  AOI21_X1 U18794 ( .B1(n15550), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20416), .ZN(n15551) );
  AND2_X1 U18795 ( .A1(n15552), .A2(n15551), .ZN(n15554) );
  INV_X1 U18796 ( .A(n15554), .ZN(n15553) );
  NAND2_X1 U18797 ( .A1(n15553), .A2(n11542), .ZN(n15555) );
  AOI22_X1 U18798 ( .A1(n15556), .A2(n15555), .B1(n15554), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15559) );
  OAI21_X1 U18799 ( .B1(n15559), .B2(n15558), .A(n15557), .ZN(n15561) );
  NAND2_X1 U18800 ( .A1(n15559), .A2(n15558), .ZN(n15560) );
  NAND2_X1 U18801 ( .A1(n15561), .A2(n15560), .ZN(n15563) );
  AOI222_X1 U18802 ( .A1(n15563), .A2(n20363), .B1(n15563), .B2(n15562), .C1(
        n20363), .C2(n15562), .ZN(n15573) );
  INV_X1 U18803 ( .A(n15564), .ZN(n15569) );
  INV_X1 U18804 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15566) );
  AOI21_X1 U18805 ( .B1(n19747), .B2(n15566), .A(n15565), .ZN(n15568) );
  NOR4_X1 U18806 ( .A1(n15570), .A2(n15569), .A3(n15568), .A4(n15567), .ZN(
        n15571) );
  OAI211_X1 U18807 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15573), .A(
        n15572), .B(n15571), .ZN(n15582) );
  NAND2_X1 U18808 ( .A1(n15575), .A2(n15574), .ZN(n15579) );
  OAI21_X1 U18809 ( .B1(n20647), .B2(n15577), .A(n15576), .ZN(n15578) );
  OAI21_X1 U18810 ( .B1(n15580), .B2(n15579), .A(n15578), .ZN(n15886) );
  AOI221_X1 U18811 ( .B1(n20790), .B2(n20553), .C1(n15582), .C2(n20553), .A(
        n15886), .ZN(n15584) );
  NOR2_X1 U18812 ( .A1(n15584), .A2(n20790), .ZN(n15889) );
  OAI211_X1 U18813 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20647), .A(n15889), 
        .B(n15581), .ZN(n15887) );
  AOI21_X1 U18814 ( .B1(n15583), .B2(n15582), .A(n15887), .ZN(n15588) );
  INV_X1 U18815 ( .A(n15584), .ZN(n15585) );
  OAI21_X1 U18816 ( .B1(n20643), .B2(n20623), .A(n15585), .ZN(n15586) );
  AOI22_X1 U18817 ( .A1(n15588), .A2(n15587), .B1(n20790), .B2(n15586), .ZN(
        P1_U3161) );
  OR2_X1 U18818 ( .A1(n16134), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16114) );
  INV_X2 U18819 ( .A(n17930), .ZN(n17932) );
  INV_X1 U18820 ( .A(n15589), .ZN(n15591) );
  NAND2_X1 U18821 ( .A1(n15591), .A2(n15590), .ZN(n15592) );
  XOR2_X1 U18822 ( .A(n15592), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16110) );
  AOI22_X1 U18823 ( .A1(n17932), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n17850), 
        .B2(n16110), .ZN(n15597) );
  AOI22_X1 U18824 ( .A1(n17928), .A2(n15593), .B1(n17917), .B2(n16134), .ZN(
        n15594) );
  NAND2_X1 U18825 ( .A1(n15594), .A2(n17915), .ZN(n16143) );
  OAI21_X1 U18826 ( .B1(n16143), .B2(n15595), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15596) );
  OAI211_X1 U18827 ( .C1(n16114), .C2(n15598), .A(n15597), .B(n15596), .ZN(
        P3_U2832) );
  NAND2_X1 U18828 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20558) );
  INV_X1 U18829 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20562) );
  NOR2_X1 U18830 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20562), .ZN(n20566) );
  NOR2_X1 U18831 ( .A1(n20562), .A2(n20647), .ZN(n20564) );
  AOI211_X1 U18832 ( .C1(HOLD), .C2(n20566), .A(n15599), .B(n20564), .ZN(
        n15600) );
  OAI221_X1 U18833 ( .B1(n20558), .B2(HOLD), .C1(n20558), .C2(
        P1_STATE_REG_2__SCAN_IN), .A(n15600), .ZN(P1_U3195) );
  AND2_X1 U18834 ( .A1(n19872), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U18835 ( .A1(n19722), .A2(n19729), .ZN(n19578) );
  NAND2_X1 U18836 ( .A1(n19578), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15602) );
  AOI21_X1 U18837 ( .B1(n19688), .B2(n19729), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15601) );
  AOI21_X1 U18838 ( .B1(n15602), .B2(n15601), .A(n16103), .ZN(P2_U3178) );
  INV_X1 U18839 ( .A(n19712), .ZN(n16098) );
  AOI221_X1 U18840 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16103), .C1(n16098), .C2(
        n16103), .A(n19515), .ZN(n19704) );
  INV_X1 U18841 ( .A(n19704), .ZN(n19701) );
  NOR2_X1 U18842 ( .A1(n15603), .A2(n19701), .ZN(P2_U3047) );
  NOR3_X1 U18843 ( .A1(n15604), .A2(n17955), .A3(n18605), .ZN(n15605) );
  NOR2_X1 U18844 ( .A1(n17077), .A2(n17135), .ZN(n17138) );
  INV_X1 U18845 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17206) );
  AOI22_X1 U18846 ( .A1(n17136), .A2(BUF2_REG_0__SCAN_IN), .B1(n17079), .B2(
        n15607), .ZN(n15608) );
  OAI221_X1 U18847 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17126), .C1(n17206), 
        .C2(n16992), .A(n15608), .ZN(P3_U2735) );
  INV_X1 U18848 ( .A(n15634), .ZN(n15616) );
  NAND3_X1 U18849 ( .A1(n15623), .A2(n15610), .A3(n15609), .ZN(n15613) );
  AOI22_X1 U18850 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n19823), .B1(
        n19766), .B2(n15611), .ZN(n15612) );
  OAI211_X1 U18851 ( .C1(n15614), .C2(n19825), .A(n15613), .B(n15612), .ZN(
        n15615) );
  AOI21_X1 U18852 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15616), .A(n15615), 
        .ZN(n15621) );
  OAI22_X1 U18853 ( .A1(n15618), .A2(n15655), .B1(n15617), .B2(n19793), .ZN(
        n15619) );
  INV_X1 U18854 ( .A(n15619), .ZN(n15620) );
  NAND2_X1 U18855 ( .A1(n15621), .A2(n15620), .ZN(P1_U2819) );
  NAND2_X1 U18856 ( .A1(n15623), .A2(n15622), .ZN(n15632) );
  OAI22_X1 U18857 ( .A1(n19825), .A2(n15625), .B1(n15624), .B2(n19769), .ZN(
        n15629) );
  OAI22_X1 U18858 ( .A1(n15627), .A2(n15655), .B1(n19793), .B2(n15626), .ZN(
        n15628) );
  AOI211_X1 U18859 ( .C1(n15630), .C2(n19766), .A(n15629), .B(n15628), .ZN(
        n15631) );
  OAI221_X1 U18860 ( .B1(n15634), .B2(n15633), .C1(n15634), .C2(n15632), .A(
        n15631), .ZN(P1_U2820) );
  INV_X1 U18861 ( .A(n15707), .ZN(n15635) );
  AOI22_X1 U18862 ( .A1(n19797), .A2(P1_EBX_REG_19__SCAN_IN), .B1(n15635), 
        .B2(n19766), .ZN(n15645) );
  NOR3_X1 U18863 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n15677), .A3(n15636), 
        .ZN(n15637) );
  AOI211_X1 U18864 ( .C1(n19823), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15637), .B(n19775), .ZN(n15644) );
  INV_X1 U18865 ( .A(n15638), .ZN(n15704) );
  AOI22_X1 U18866 ( .A1(n15704), .A2(n19809), .B1(n15771), .B2(n19828), .ZN(
        n15643) );
  NOR3_X1 U18867 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15640), .A3(n15639), 
        .ZN(n15647) );
  INV_X1 U18868 ( .A(n15679), .ZN(n15671) );
  OAI21_X1 U18869 ( .B1(n15641), .B2(n15677), .A(n15671), .ZN(n15657) );
  OAI21_X1 U18870 ( .B1(n15647), .B2(n15657), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15642) );
  NAND4_X1 U18871 ( .A1(n15645), .A2(n15644), .A3(n15643), .A4(n15642), .ZN(
        P1_U2821) );
  NAND2_X1 U18872 ( .A1(n19823), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15646) );
  OAI211_X1 U18873 ( .C1(n19825), .C2(n14455), .A(n15646), .B(n19820), .ZN(
        n15648) );
  AOI211_X1 U18874 ( .C1(n19766), .C2(n15649), .A(n15648), .B(n15647), .ZN(
        n15650) );
  OAI21_X1 U18875 ( .B1(n15651), .B2(n15655), .A(n15650), .ZN(n15652) );
  AOI21_X1 U18876 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15657), .A(n15652), 
        .ZN(n15653) );
  OAI21_X1 U18877 ( .B1(n19793), .B2(n15654), .A(n15653), .ZN(P1_U2822) );
  AOI22_X1 U18878 ( .A1(n19797), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19823), .ZN(n15662) );
  AOI21_X1 U18879 ( .B1(n19766), .B2(n15715), .A(n19775), .ZN(n15661) );
  OAI22_X1 U18880 ( .A1(n15717), .A2(n15655), .B1(n19793), .B2(n15779), .ZN(
        n15656) );
  INV_X1 U18881 ( .A(n15656), .ZN(n15660) );
  OAI221_X1 U18882 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), .C1(P1_REIP_REG_17__SCAN_IN), .C2(n15658), .A(n15657), .ZN(n15659) );
  NAND4_X1 U18883 ( .A1(n15662), .A2(n15661), .A3(n15660), .A4(n15659), .ZN(
        P1_U2823) );
  AOI22_X1 U18884 ( .A1(n15725), .A2(n19766), .B1(n19828), .B2(n15795), .ZN(
        n15663) );
  OAI211_X1 U18885 ( .C1(n19769), .C2(n15664), .A(n15663), .B(n19820), .ZN(
        n15666) );
  AOI211_X1 U18886 ( .C1(n19797), .C2(P1_EBX_REG_15__SCAN_IN), .A(n15666), .B(
        n15665), .ZN(n15667) );
  INV_X1 U18887 ( .A(n15667), .ZN(n15668) );
  AOI21_X1 U18888 ( .B1(n15726), .B2(n19809), .A(n15668), .ZN(n15669) );
  OAI21_X1 U18889 ( .B1(n15671), .B2(n15670), .A(n15669), .ZN(P1_U2825) );
  INV_X1 U18890 ( .A(n15672), .ZN(n15673) );
  AOI22_X1 U18891 ( .A1(n19797), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n15673), 
        .B2(n19766), .ZN(n15683) );
  AOI22_X1 U18892 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19823), .B1(
        n19828), .B2(n15804), .ZN(n15682) );
  INV_X1 U18893 ( .A(n15674), .ZN(n15680) );
  OAI21_X1 U18894 ( .B1(n15677), .B2(n15676), .A(n15675), .ZN(n15678) );
  AOI22_X1 U18895 ( .A1(n15680), .A2(n19809), .B1(n15679), .B2(n15678), .ZN(
        n15681) );
  NAND4_X1 U18896 ( .A1(n15683), .A2(n15682), .A3(n15681), .A4(n19820), .ZN(
        P1_U2826) );
  INV_X1 U18897 ( .A(n15699), .ZN(n15684) );
  AOI21_X1 U18898 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15684), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15690) );
  AOI22_X1 U18899 ( .A1(n19797), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n15730), 
        .B2(n19766), .ZN(n15689) );
  OAI22_X1 U18900 ( .A1(n15686), .A2(n19769), .B1(n19793), .B2(n15685), .ZN(
        n15687) );
  AOI211_X1 U18901 ( .C1(n15729), .C2(n19809), .A(n19775), .B(n15687), .ZN(
        n15688) );
  OAI211_X1 U18902 ( .C1(n15691), .C2(n15690), .A(n15689), .B(n15688), .ZN(
        P1_U2828) );
  OAI22_X1 U18903 ( .A1(n15822), .A2(n19793), .B1(n19825), .B2(n15692), .ZN(
        n15693) );
  INV_X1 U18904 ( .A(n15693), .ZN(n15694) );
  OAI21_X1 U18905 ( .B1(n15743), .B2(n19821), .A(n15694), .ZN(n15695) );
  AOI211_X1 U18906 ( .C1(n19823), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19775), .B(n15695), .ZN(n15698) );
  AOI22_X1 U18907 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15696), .B1(n19809), 
        .B2(n15740), .ZN(n15697) );
  OAI211_X1 U18908 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15699), .A(n15698), 
        .B(n15697), .ZN(P1_U2829) );
  AOI22_X1 U18909 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15706) );
  NAND2_X1 U18910 ( .A1(n15702), .A2(n15700), .ZN(n15701) );
  MUX2_X1 U18911 ( .A(n15702), .B(n15701), .S(n14605), .Z(n15703) );
  XNOR2_X1 U18912 ( .A(n15703), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15772) );
  AOI22_X1 U18913 ( .A1(n19912), .A2(n15772), .B1(n15704), .B2(n19911), .ZN(
        n15705) );
  OAI211_X1 U18914 ( .C1(n19916), .C2(n15707), .A(n15706), .B(n15705), .ZN(
        P1_U2980) );
  INV_X1 U18915 ( .A(n15708), .ZN(n15709) );
  AOI21_X1 U18916 ( .B1(n15711), .B2(n15710), .A(n15709), .ZN(n15713) );
  NOR2_X1 U18917 ( .A1(n15713), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15712) );
  MUX2_X1 U18918 ( .A(n15713), .B(n15712), .S(n15702), .Z(n15714) );
  XNOR2_X1 U18919 ( .A(n15714), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15785) );
  AOI22_X1 U18920 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15720) );
  INV_X1 U18921 ( .A(n15715), .ZN(n15716) );
  OAI22_X1 U18922 ( .A1(n15717), .A2(n19960), .B1(n15716), .B2(n19916), .ZN(
        n15718) );
  INV_X1 U18923 ( .A(n15718), .ZN(n15719) );
  OAI211_X1 U18924 ( .C1(n19746), .C2(n15785), .A(n15720), .B(n15719), .ZN(
        P1_U2982) );
  OAI21_X1 U18925 ( .B1(n15723), .B2(n15722), .A(n15721), .ZN(n15724) );
  INV_X1 U18926 ( .A(n15724), .ZN(n15802) );
  AOI22_X1 U18927 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15728) );
  AOI22_X1 U18928 ( .A1(n15726), .A2(n19911), .B1(n15725), .B2(n15731), .ZN(
        n15727) );
  OAI211_X1 U18929 ( .C1(n15802), .C2(n19746), .A(n15728), .B(n15727), .ZN(
        P1_U2984) );
  AOI22_X1 U18930 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15733) );
  AOI22_X1 U18931 ( .A1(n15731), .A2(n15730), .B1(n19911), .B2(n15729), .ZN(
        n15732) );
  OAI211_X1 U18932 ( .C1(n15734), .C2(n19746), .A(n15733), .B(n15732), .ZN(
        P1_U2987) );
  AOI22_X1 U18933 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15742) );
  NOR2_X1 U18934 ( .A1(n14649), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15737) );
  NOR2_X1 U18935 ( .A1(n14608), .A2(n14634), .ZN(n15736) );
  MUX2_X1 U18936 ( .A(n15737), .B(n15736), .S(n14633), .Z(n15739) );
  XNOR2_X1 U18937 ( .A(n15739), .B(n15738), .ZN(n15824) );
  AOI22_X1 U18938 ( .A1(n19912), .A2(n15824), .B1(n19911), .B2(n15740), .ZN(
        n15741) );
  OAI211_X1 U18939 ( .C1(n19916), .C2(n15743), .A(n15742), .B(n15741), .ZN(
        P1_U2988) );
  AOI22_X1 U18940 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15749) );
  NAND2_X1 U18941 ( .A1(n15746), .A2(n15745), .ZN(n15747) );
  XNOR2_X1 U18942 ( .A(n15744), .B(n15747), .ZN(n15863) );
  AOI22_X1 U18943 ( .A1(n15863), .A2(n19912), .B1(n19911), .B2(n19801), .ZN(
        n15748) );
  OAI211_X1 U18944 ( .C1(n19916), .C2(n19791), .A(n15749), .B(n15748), .ZN(
        P1_U2992) );
  AOI22_X1 U18945 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15754) );
  XNOR2_X1 U18946 ( .A(n15751), .B(n15855), .ZN(n15752) );
  XNOR2_X1 U18947 ( .A(n15750), .B(n15752), .ZN(n15869) );
  AOI22_X1 U18948 ( .A1(n15869), .A2(n19912), .B1(n19911), .B2(n19842), .ZN(
        n15753) );
  OAI211_X1 U18949 ( .C1(n19916), .C2(n19805), .A(n15754), .B(n15753), .ZN(
        P1_U2993) );
  AOI22_X1 U18950 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15760) );
  OAI21_X1 U18951 ( .B1(n15757), .B2(n15756), .A(n15755), .ZN(n15758) );
  INV_X1 U18952 ( .A(n15758), .ZN(n15878) );
  AOI22_X1 U18953 ( .A1(n15878), .A2(n19912), .B1(n19911), .B2(n19848), .ZN(
        n15759) );
  OAI211_X1 U18954 ( .C1(n19916), .C2(n19812), .A(n15760), .B(n15759), .ZN(
        P1_U2994) );
  INV_X1 U18955 ( .A(n15761), .ZN(n15764) );
  OAI22_X1 U18956 ( .A1(n15764), .A2(n19945), .B1(n15763), .B2(n15762), .ZN(
        n15765) );
  AOI21_X1 U18957 ( .B1(n19929), .B2(n15766), .A(n15765), .ZN(n15770) );
  OAI211_X1 U18958 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15768), .B(n15767), .ZN(
        n15769) );
  OAI211_X1 U18959 ( .C1(n20691), .C2(n19942), .A(n15770), .B(n15769), .ZN(
        P1_U3009) );
  AOI22_X1 U18960 ( .A1(n15772), .A2(n19929), .B1(n19925), .B2(n15771), .ZN(
        n15777) );
  NOR2_X1 U18961 ( .A1(n19942), .A2(n20722), .ZN(n15773) );
  AOI221_X1 U18962 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15775), 
        .C1(n20747), .C2(n15774), .A(n15773), .ZN(n15776) );
  NAND2_X1 U18963 ( .A1(n15777), .A2(n15776), .ZN(P1_U3012) );
  INV_X1 U18964 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15778) );
  OAI22_X1 U18965 ( .A1(n15779), .A2(n19945), .B1(n19942), .B2(n15778), .ZN(
        n15780) );
  INV_X1 U18966 ( .A(n15780), .ZN(n15784) );
  OAI21_X1 U18967 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15782), .A(
        n15781), .ZN(n15783) );
  OAI211_X1 U18968 ( .C1(n15785), .C2(n19946), .A(n15784), .B(n15783), .ZN(
        P1_U3014) );
  OAI21_X1 U18969 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15786), .ZN(n15794) );
  INV_X1 U18970 ( .A(n15787), .ZN(n15788) );
  AOI21_X1 U18971 ( .B1(n15789), .B2(n19925), .A(n15788), .ZN(n15793) );
  OAI21_X1 U18972 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15790), .A(
        n15810), .ZN(n15799) );
  AOI22_X1 U18973 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15799), .B1(
        n19929), .B2(n15791), .ZN(n15792) );
  OAI211_X1 U18974 ( .C1(n15796), .C2(n15794), .A(n15793), .B(n15792), .ZN(
        P1_U3015) );
  AOI22_X1 U18975 ( .A1(n15795), .A2(n19925), .B1(n12105), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n15801) );
  INV_X1 U18976 ( .A(n15796), .ZN(n15798) );
  AOI22_X1 U18977 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15799), .B1(
        n15798), .B2(n15797), .ZN(n15800) );
  OAI211_X1 U18978 ( .C1(n15802), .C2(n19946), .A(n15801), .B(n15800), .ZN(
        P1_U3016) );
  AOI21_X1 U18979 ( .B1(n15804), .B2(n19925), .A(n15803), .ZN(n15808) );
  AOI22_X1 U18980 ( .A1(n19929), .A2(n15806), .B1(n15805), .B2(n15809), .ZN(
        n15807) );
  OAI211_X1 U18981 ( .C1(n15810), .C2(n15809), .A(n15808), .B(n15807), .ZN(
        P1_U3017) );
  AOI22_X1 U18982 ( .A1(n12105), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n15812), 
        .B2(n15811), .ZN(n15820) );
  AOI22_X1 U18983 ( .A1(n15815), .A2(n19925), .B1(n15814), .B2(n15813), .ZN(
        n15819) );
  AOI22_X1 U18984 ( .A1(n15817), .A2(n19929), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15816), .ZN(n15818) );
  NAND3_X1 U18985 ( .A1(n15820), .A2(n15819), .A3(n15818), .ZN(P1_U3018) );
  INV_X1 U18986 ( .A(n15821), .ZN(n15828) );
  OAI22_X1 U18987 ( .A1(n15822), .A2(n19945), .B1(n19942), .B2(n20588), .ZN(
        n15823) );
  INV_X1 U18988 ( .A(n15823), .ZN(n15827) );
  AOI22_X1 U18989 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15825), .B1(
        n19929), .B2(n15824), .ZN(n15826) );
  OAI211_X1 U18990 ( .C1(n15872), .C2(n15828), .A(n15827), .B(n15826), .ZN(
        P1_U3020) );
  OAI21_X1 U18991 ( .B1(n15850), .B2(n15849), .A(n15830), .ZN(n15829) );
  AOI221_X1 U18992 ( .B1(n15847), .B2(n15854), .C1(n15829), .C2(n15854), .A(
        n19938), .ZN(n15846) );
  INV_X1 U18993 ( .A(n15872), .ZN(n15857) );
  NAND2_X1 U18994 ( .A1(n15830), .A2(n15857), .ZN(n15842) );
  AOI221_X1 U18995 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14634), .C2(n14025), .A(
        n15842), .ZN(n15833) );
  OAI22_X1 U18996 ( .A1(n15831), .A2(n19945), .B1(n14651), .B2(n19942), .ZN(
        n15832) );
  AOI211_X1 U18997 ( .C1(n15834), .C2(n19929), .A(n15833), .B(n15832), .ZN(
        n15835) );
  OAI21_X1 U18998 ( .B1(n14634), .B2(n15846), .A(n15835), .ZN(P1_U3021) );
  INV_X1 U18999 ( .A(n15836), .ZN(n15844) );
  NAND2_X1 U19000 ( .A1(n15838), .A2(n15837), .ZN(n15839) );
  AND2_X1 U19001 ( .A1(n15840), .A2(n15839), .ZN(n19837) );
  AOI22_X1 U19002 ( .A1(n19837), .A2(n19925), .B1(n12105), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n15841) );
  OAI21_X1 U19003 ( .B1(n15842), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15841), .ZN(n15843) );
  AOI21_X1 U19004 ( .B1(n15844), .B2(n19929), .A(n15843), .ZN(n15845) );
  OAI21_X1 U19005 ( .B1(n14025), .B2(n15846), .A(n15845), .ZN(P1_U3022) );
  NOR2_X1 U19006 ( .A1(n19919), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15877) );
  INV_X1 U19007 ( .A(n15877), .ZN(n15852) );
  AND2_X1 U19008 ( .A1(n15847), .A2(n19951), .ZN(n15851) );
  OAI21_X1 U19009 ( .B1(n15850), .B2(n15849), .A(n15848), .ZN(n19917) );
  AOI211_X1 U19010 ( .C1(n19940), .C2(n19919), .A(n15851), .B(n19917), .ZN(
        n15881) );
  OAI21_X1 U19011 ( .B1(n15853), .B2(n15852), .A(n15881), .ZN(n15868) );
  AOI21_X1 U19012 ( .B1(n15855), .B2(n15854), .A(n15868), .ZN(n15865) );
  INV_X1 U19013 ( .A(n15856), .ZN(n15860) );
  NAND2_X1 U19014 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15857), .ZN(
        n15867) );
  AOI221_X1 U19015 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15862), .C2(n15866), .A(
        n15867), .ZN(n15859) );
  OAI22_X1 U19016 ( .A1(n19780), .A2(n19945), .B1(n19786), .B2(n19942), .ZN(
        n15858) );
  AOI211_X1 U19017 ( .C1(n15860), .C2(n19929), .A(n15859), .B(n15858), .ZN(
        n15861) );
  OAI21_X1 U19018 ( .B1(n15865), .B2(n15862), .A(n15861), .ZN(P1_U3023) );
  AOI222_X1 U19019 ( .A1(n15863), .A2(n19929), .B1(n19925), .B2(n19792), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(n12105), .ZN(n15864) );
  OAI221_X1 U19020 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15867), .C1(
        n15866), .C2(n15865), .A(n15864), .ZN(P1_U3024) );
  XNOR2_X1 U19021 ( .A(n15876), .B(n10005), .ZN(n19841) );
  AOI22_X1 U19022 ( .A1(n19841), .A2(n19925), .B1(n12105), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15871) );
  AOI22_X1 U19023 ( .A1(n15869), .A2(n19929), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15868), .ZN(n15870) );
  OAI211_X1 U19024 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15872), .A(
        n15871), .B(n15870), .ZN(P1_U3025) );
  OR2_X1 U19025 ( .A1(n15874), .A2(n15873), .ZN(n15875) );
  AND2_X1 U19026 ( .A1(n15876), .A2(n15875), .ZN(n19845) );
  AOI22_X1 U19027 ( .A1(n19845), .A2(n19925), .B1(n12105), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n15880) );
  AOI22_X1 U19028 ( .A1(n15878), .A2(n19929), .B1(n15877), .B2(n19928), .ZN(
        n15879) );
  OAI211_X1 U19029 ( .C1(n15881), .C2(n20699), .A(n15880), .B(n15879), .ZN(
        P1_U3026) );
  NAND4_X1 U19030 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20640), .A4(n20647), .ZN(n15882) );
  AND2_X1 U19031 ( .A1(n15883), .A2(n15882), .ZN(n20554) );
  NAND2_X1 U19032 ( .A1(n20554), .A2(n15884), .ZN(n15885) );
  AOI22_X1 U19033 ( .A1(n20553), .A2(n15887), .B1(n15886), .B2(n15885), .ZN(
        P1_U3162) );
  OAI21_X1 U19034 ( .B1(n15889), .B2(n20371), .A(n15888), .ZN(P1_U3466) );
  INV_X1 U19035 ( .A(n15891), .ZN(n15892) );
  INV_X1 U19036 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19659) );
  OAI22_X1 U19037 ( .A1(n15892), .A2(n18865), .B1(n19659), .B2(n18845), .ZN(
        n15896) );
  OAI22_X1 U19038 ( .A1(n13102), .A2(n18871), .B1(n15894), .B2(n15893), .ZN(
        n15895) );
  AOI211_X1 U19039 ( .C1(n18859), .C2(n15890), .A(n15896), .B(n15895), .ZN(
        n15899) );
  NAND4_X1 U19040 ( .A1(n18838), .A2(n15900), .A3(n15897), .A4(n13108), .ZN(
        n15898) );
  OAI211_X1 U19041 ( .C1(n14271), .C2(n18858), .A(n15899), .B(n15898), .ZN(
        P2_U2824) );
  AOI21_X1 U19042 ( .B1(n15902), .B2(n15901), .A(n15900), .ZN(n15908) );
  AOI22_X1 U19043 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n18862), .B1(n15903), 
        .B2(n18847), .ZN(n15905) );
  AOI22_X1 U19044 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18842), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n18861), .ZN(n15904) );
  OAI211_X1 U19045 ( .C1(n15906), .C2(n18858), .A(n15905), .B(n15904), .ZN(
        n15907) );
  AOI21_X1 U19046 ( .B1(n18838), .B2(n15908), .A(n15907), .ZN(n15909) );
  OAI21_X1 U19047 ( .B1(n15910), .B2(n18841), .A(n15909), .ZN(P2_U2826) );
  AOI22_X1 U19048 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18861), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18862), .ZN(n15911) );
  OAI21_X1 U19049 ( .B1(n15912), .B2(n18865), .A(n15911), .ZN(n15913) );
  AOI21_X1 U19050 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18842), .A(
        n15913), .ZN(n15920) );
  AOI21_X1 U19051 ( .B1(n15916), .B2(n15915), .A(n15914), .ZN(n15917) );
  AOI22_X1 U19052 ( .A1(n15918), .A2(n18859), .B1(n18838), .B2(n15917), .ZN(
        n15919) );
  OAI211_X1 U19053 ( .C1(n15921), .C2(n18858), .A(n15920), .B(n15919), .ZN(
        P2_U2827) );
  AOI211_X1 U19054 ( .C1(n15924), .C2(n15923), .A(n15922), .B(n19582), .ZN(
        n15930) );
  AOI22_X1 U19055 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n18862), .B1(n15925), 
        .B2(n18847), .ZN(n15927) );
  AOI22_X1 U19056 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18842), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n18861), .ZN(n15926) );
  OAI211_X1 U19057 ( .C1(n15928), .C2(n18858), .A(n15927), .B(n15926), .ZN(
        n15929) );
  AOI211_X1 U19058 ( .C1(n18859), .C2(n15931), .A(n15930), .B(n15929), .ZN(
        n15932) );
  INV_X1 U19059 ( .A(n15932), .ZN(P2_U2829) );
  OAI22_X1 U19060 ( .A1(n15933), .A2(n18865), .B1(n19647), .B2(n18845), .ZN(
        n15934) );
  INV_X1 U19061 ( .A(n15934), .ZN(n15943) );
  AOI22_X1 U19062 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n18861), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18842), .ZN(n15942) );
  AOI22_X1 U19063 ( .A1(n15936), .A2(n18868), .B1(n15935), .B2(n18859), .ZN(
        n15941) );
  AOI21_X1 U19064 ( .B1(n15938), .B2(n9666), .A(n15937), .ZN(n15939) );
  NAND2_X1 U19065 ( .A1(n18838), .A2(n15939), .ZN(n15940) );
  NAND4_X1 U19066 ( .A1(n15943), .A2(n15942), .A3(n15941), .A4(n15940), .ZN(
        P2_U2830) );
  AOI211_X1 U19067 ( .C1(n15946), .C2(n15945), .A(n15944), .B(n19582), .ZN(
        n15954) );
  INV_X1 U19068 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n15947) );
  OAI22_X1 U19069 ( .A1(n15948), .A2(n18865), .B1(n15947), .B2(n18845), .ZN(
        n15949) );
  INV_X1 U19070 ( .A(n15949), .ZN(n15951) );
  AOI22_X1 U19071 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18861), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18842), .ZN(n15950) );
  OAI211_X1 U19072 ( .C1(n15952), .C2(n18858), .A(n15951), .B(n15950), .ZN(
        n15953) );
  AOI211_X1 U19073 ( .C1(n18859), .C2(n15955), .A(n15954), .B(n15953), .ZN(
        n15956) );
  INV_X1 U19074 ( .A(n15956), .ZN(P2_U2831) );
  AOI22_X1 U19075 ( .A1(n18882), .A2(n15957), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n18931), .ZN(n15962) );
  AOI22_X1 U19076 ( .A1(n18884), .A2(BUF2_REG_22__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U19077 ( .A1(n15959), .A2(n18890), .B1(n18932), .B2(n15958), .ZN(
        n15960) );
  NAND3_X1 U19078 ( .A1(n15962), .A2(n15961), .A3(n15960), .ZN(P2_U2897) );
  AOI22_X1 U19079 ( .A1(n18882), .A2(n15963), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n18931), .ZN(n15968) );
  AOI22_X1 U19080 ( .A1(n18884), .A2(BUF2_REG_20__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15967) );
  INV_X1 U19081 ( .A(n15964), .ZN(n15965) );
  AOI22_X1 U19082 ( .A1(n15965), .A2(n18890), .B1(n18932), .B2(n18676), .ZN(
        n15966) );
  NAND3_X1 U19083 ( .A1(n15968), .A2(n15967), .A3(n15966), .ZN(P2_U2899) );
  AOI22_X1 U19084 ( .A1(n18882), .A2(n15969), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n18931), .ZN(n15973) );
  AOI22_X1 U19085 ( .A1(n18884), .A2(BUF2_REG_18__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15972) );
  AOI22_X1 U19086 ( .A1(n15970), .A2(n18890), .B1(n18932), .B2(n9995), .ZN(
        n15971) );
  NAND3_X1 U19087 ( .A1(n15973), .A2(n15972), .A3(n15971), .ZN(P2_U2901) );
  AOI22_X1 U19088 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n15127), .B1(n19049), 
        .B2(n18781), .ZN(n15985) );
  INV_X1 U19089 ( .A(n15974), .ZN(n15975) );
  AOI21_X1 U19090 ( .B1(n15977), .B2(n15976), .A(n15975), .ZN(n15981) );
  NAND2_X1 U19091 ( .A1(n15979), .A2(n15978), .ZN(n15980) );
  XNOR2_X1 U19092 ( .A(n15981), .B(n15980), .ZN(n16019) );
  INV_X1 U19093 ( .A(n16019), .ZN(n15983) );
  AOI21_X1 U19094 ( .B1(n16012), .B2(n9669), .A(n15982), .ZN(n16016) );
  AOI222_X1 U19095 ( .A1(n15983), .A2(n19050), .B1(n16001), .B2(n16006), .C1(
        n19052), .C2(n16016), .ZN(n15984) );
  OAI211_X1 U19096 ( .C1(n19061), .C2(n18787), .A(n15985), .B(n15984), .ZN(
        P2_U3004) );
  AOI22_X1 U19097 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n15127), .B1(n19049), 
        .B2(n18804), .ZN(n15999) );
  NAND2_X1 U19098 ( .A1(n15987), .A2(n15986), .ZN(n15990) );
  OAI21_X1 U19099 ( .B1(n15990), .B2(n15989), .A(n15988), .ZN(n16028) );
  NOR2_X1 U19100 ( .A1(n15992), .A2(n15991), .ZN(n15994) );
  XOR2_X1 U19101 ( .A(n15994), .B(n15993), .Z(n16033) );
  OAI222_X1 U19102 ( .A1(n16026), .A2(n19057), .B1(n16028), .B2(n15996), .C1(
        n15995), .C2(n16033), .ZN(n15997) );
  INV_X1 U19103 ( .A(n15997), .ZN(n15998) );
  OAI211_X1 U19104 ( .C1(n19061), .C2(n18799), .A(n15999), .B(n15998), .ZN(
        P2_U3006) );
  AOI22_X1 U19105 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n15127), .B1(n19049), 
        .B2(n18826), .ZN(n16005) );
  INV_X1 U19106 ( .A(n16000), .ZN(n16003) );
  AOI222_X1 U19107 ( .A1(n19052), .A2(n16003), .B1(n16002), .B2(n19050), .C1(
        n16001), .C2(n9716), .ZN(n16004) );
  OAI211_X1 U19108 ( .C1(n19061), .C2(n18821), .A(n16005), .B(n16004), .ZN(
        P2_U3008) );
  INV_X1 U19109 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19622) );
  NOR2_X1 U19110 ( .A1(n19622), .A2(n14056), .ZN(n16010) );
  INV_X1 U19111 ( .A(n16006), .ZN(n18782) );
  XNOR2_X1 U19112 ( .A(n15388), .B(n16007), .ZN(n18904) );
  OAI22_X1 U19113 ( .A1(n18782), .A2(n16008), .B1(n16036), .B2(n18904), .ZN(
        n16009) );
  AOI211_X1 U19114 ( .C1(n16011), .C2(n16012), .A(n16010), .B(n16009), .ZN(
        n16018) );
  NOR3_X1 U19115 ( .A1(n16014), .A2(n16013), .A3(n16012), .ZN(n16015) );
  AOI21_X1 U19116 ( .B1(n16016), .B2(n10731), .A(n16015), .ZN(n16017) );
  OAI211_X1 U19117 ( .C1(n16019), .C2(n16034), .A(n16018), .B(n16017), .ZN(
        P2_U3036) );
  AOI21_X1 U19118 ( .B1(n16022), .B2(n16021), .A(n16020), .ZN(n16023) );
  AOI22_X1 U19119 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16025), .B1(
        n16024), .B2(n16023), .ZN(n16032) );
  INV_X1 U19120 ( .A(n16026), .ZN(n18805) );
  XNOR2_X1 U19121 ( .A(n14228), .B(n16027), .ZN(n18910) );
  INV_X1 U19122 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19619) );
  OAI22_X1 U19123 ( .A1(n16036), .A2(n18910), .B1(n19619), .B2(n14056), .ZN(
        n16030) );
  NOR2_X1 U19124 ( .A1(n16028), .A2(n16040), .ZN(n16029) );
  AOI211_X1 U19125 ( .C1(n18805), .C2(n16038), .A(n16030), .B(n16029), .ZN(
        n16031) );
  OAI211_X1 U19126 ( .C1(n16034), .C2(n16033), .A(n16032), .B(n16031), .ZN(
        P2_U3038) );
  OAI21_X1 U19127 ( .B1(n19676), .B2(n16036), .A(n16035), .ZN(n16037) );
  AOI21_X1 U19128 ( .B1(n13444), .B2(n16038), .A(n16037), .ZN(n16039) );
  OAI21_X1 U19129 ( .B1(n16041), .B2(n16040), .A(n16039), .ZN(n16042) );
  AOI21_X1 U19130 ( .B1(n16044), .B2(n16043), .A(n16042), .ZN(n16045) );
  OAI221_X1 U19131 ( .B1(n16048), .B2(n16047), .C1(n16048), .C2(n16046), .A(
        n16045), .ZN(P2_U3043) );
  NAND2_X1 U19132 ( .A1(n16049), .A2(n19729), .ZN(n16094) );
  INV_X1 U19133 ( .A(n16050), .ZN(n16092) );
  MUX2_X1 U19134 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16051), .S(
        n16077), .Z(n16091) );
  INV_X1 U19135 ( .A(n16052), .ZN(n16053) );
  MUX2_X1 U19136 ( .A(n16054), .B(n16053), .S(n16077), .Z(n16074) );
  INV_X1 U19137 ( .A(n16074), .ZN(n16090) );
  INV_X1 U19138 ( .A(n16055), .ZN(n16061) );
  AOI22_X1 U19139 ( .A1(n16061), .A2(n16058), .B1(n16057), .B2(n16056), .ZN(
        n16059) );
  OAI21_X1 U19140 ( .B1(n16061), .B2(n16060), .A(n16059), .ZN(n19714) );
  INV_X1 U19141 ( .A(n16062), .ZN(n16064) );
  NOR3_X1 U19142 ( .A1(n16065), .A2(n16064), .A3(n16063), .ZN(n18632) );
  OAI21_X1 U19143 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n18632), .ZN(n16069) );
  NAND3_X1 U19144 ( .A1(n15500), .A2(n16067), .A3(n16066), .ZN(n16068) );
  OAI211_X1 U19145 ( .C1(n10121), .C2(n16070), .A(n16069), .B(n16068), .ZN(
        n16071) );
  NOR2_X1 U19146 ( .A1(n19714), .A2(n16071), .ZN(n16072) );
  OAI21_X1 U19147 ( .B1(n16077), .B2(n16073), .A(n16072), .ZN(n16089) );
  NAND2_X1 U19148 ( .A1(n16074), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n16084) );
  INV_X1 U19149 ( .A(n16075), .ZN(n16076) );
  NAND2_X1 U19150 ( .A1(n16076), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16079) );
  INV_X1 U19151 ( .A(n16079), .ZN(n16082) );
  INV_X1 U19152 ( .A(n16077), .ZN(n16081) );
  AOI21_X1 U19153 ( .B1(n19696), .B2(n16079), .A(n16078), .ZN(n16080) );
  AOI211_X1 U19154 ( .C1(n16082), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16081), .B(n16080), .ZN(n16083) );
  OAI211_X1 U19155 ( .C1(n16091), .C2(n19680), .A(n16084), .B(n16083), .ZN(
        n16087) );
  INV_X1 U19156 ( .A(n19131), .ZN(n16085) );
  AOI22_X1 U19157 ( .A1(n16090), .A2(n16085), .B1(n16091), .B2(n19680), .ZN(
        n16086) );
  AOI21_X1 U19158 ( .B1(n16087), .B2(n16086), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16088) );
  AOI211_X1 U19159 ( .C1(n16091), .C2(n16090), .A(n16089), .B(n16088), .ZN(
        n16096) );
  OAI211_X1 U19160 ( .C1(n10138), .C2(n16092), .A(n16096), .B(n19720), .ZN(
        n19579) );
  NAND2_X1 U19161 ( .A1(n19579), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16104) );
  AOI21_X1 U19162 ( .B1(n16094), .B2(n16104), .A(n16093), .ZN(n16102) );
  INV_X1 U19163 ( .A(n19008), .ZN(n19721) );
  INV_X2 U19164 ( .A(n19721), .ZN(n18988) );
  NOR2_X1 U19165 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19729), .ZN(n19580) );
  OAI22_X1 U19166 ( .A1(n16098), .A2(n16097), .B1(n16096), .B2(n18631), .ZN(
        n16099) );
  AOI211_X1 U19167 ( .C1(n19722), .C2(n19580), .A(n16100), .B(n16099), .ZN(
        n16101) );
  OAI221_X1 U19168 ( .B1(n16102), .B2(n19722), .C1(n16102), .C2(n18988), .A(
        n16101), .ZN(P2_U3176) );
  AOI21_X1 U19169 ( .B1(n16104), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16103), 
        .ZN(n16105) );
  INV_X1 U19170 ( .A(n16105), .ZN(P2_U3593) );
  INV_X1 U19171 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16325) );
  XNOR2_X1 U19172 ( .A(n16325), .B(n16119), .ZN(n16324) );
  NAND2_X1 U19173 ( .A1(n17932), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16106) );
  OAI221_X1 U19174 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16108), .C1(
        n16325), .C2(n16107), .A(n16106), .ZN(n16109) );
  AOI21_X1 U19175 ( .B1(n17465), .B2(n16324), .A(n16109), .ZN(n16113) );
  INV_X1 U19176 ( .A(n17520), .ZN(n17454) );
  OAI22_X1 U19177 ( .A1(n16129), .A2(n17454), .B1(n16117), .B2(n17613), .ZN(
        n16111) );
  AOI22_X1 U19178 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16111), .B1(
        n17519), .B2(n16110), .ZN(n16112) );
  OAI211_X1 U19179 ( .C1(n16115), .C2(n16114), .A(n16113), .B(n16112), .ZN(
        P3_U2800) );
  INV_X1 U19180 ( .A(n16116), .ZN(n16128) );
  NOR2_X1 U19181 ( .A1(n17616), .A2(n16128), .ZN(n16162) );
  NOR2_X1 U19182 ( .A1(n16117), .A2(n17613), .ZN(n16127) );
  AOI22_X1 U19183 ( .A1(n17932), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16118), .ZN(n16123) );
  AOI21_X1 U19184 ( .B1(n16337), .B2(n16120), .A(n16119), .ZN(n16336) );
  OAI21_X1 U19185 ( .B1(n16121), .B2(n17465), .A(n16336), .ZN(n16122) );
  OAI211_X1 U19186 ( .C1(n16125), .C2(n16124), .A(n16123), .B(n16122), .ZN(
        n16126) );
  AOI221_X1 U19187 ( .B1(n16162), .B2(n16127), .C1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16127), .A(n16126), .ZN(
        n16132) );
  NOR2_X1 U19188 ( .A1(n16128), .A2(n17615), .ZN(n16161) );
  NOR2_X1 U19189 ( .A1(n16129), .A2(n17454), .ZN(n16130) );
  OAI21_X1 U19190 ( .B1(n16161), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16130), .ZN(n16131) );
  OAI211_X1 U19191 ( .C1(n16133), .C2(n17498), .A(n16132), .B(n16131), .ZN(
        P3_U2801) );
  NOR3_X1 U19192 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16135), .A3(
        n16134), .ZN(n16137) );
  AOI22_X1 U19193 ( .A1(n17839), .A2(n16138), .B1(n16137), .B2(n16136), .ZN(
        n16139) );
  OAI21_X1 U19194 ( .B1(n16140), .B2(n17806), .A(n16139), .ZN(n16141) );
  AOI21_X1 U19195 ( .B1(n16142), .B2(n17882), .A(n16141), .ZN(n16147) );
  AOI22_X1 U19196 ( .A1(n17850), .A2(n16144), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16143), .ZN(n16146) );
  OAI211_X1 U19197 ( .C1(n16147), .C2(n17922), .A(n16146), .B(n16145), .ZN(
        P3_U2831) );
  INV_X1 U19198 ( .A(n17640), .ZN(n17304) );
  AOI22_X1 U19199 ( .A1(n18384), .A2(n17805), .B1(n17839), .B2(n17808), .ZN(
        n17732) );
  NOR2_X1 U19200 ( .A1(n17769), .A2(n17900), .ZN(n16148) );
  AOI22_X1 U19201 ( .A1(n18385), .A2(n17725), .B1(n16149), .B2(n16148), .ZN(
        n17647) );
  OAI21_X1 U19202 ( .B1(n17732), .B2(n16150), .A(n17647), .ZN(n17674) );
  NAND2_X1 U19203 ( .A1(n17304), .A2(n17674), .ZN(n17669) );
  AOI22_X1 U19204 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n17932), .B1(n16153), 
        .B2(n16152), .ZN(n16169) );
  INV_X1 U19205 ( .A(n16154), .ZN(n16155) );
  OAI211_X1 U19206 ( .C1(n16158), .C2(n16157), .A(n16156), .B(n16155), .ZN(
        n16160) );
  OAI211_X1 U19207 ( .C1(n17108), .C2(n16160), .A(n17928), .B(n16159), .ZN(
        n16164) );
  OAI22_X1 U19208 ( .A1(n16162), .A2(n17806), .B1(n16161), .B2(n17807), .ZN(
        n16163) );
  OAI211_X1 U19209 ( .C1(n16164), .C2(n16163), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17930), .ZN(n16168) );
  NAND3_X1 U19210 ( .A1(n16166), .A2(n17850), .A3(n16165), .ZN(n16167) );
  NAND3_X1 U19211 ( .A1(n16169), .A2(n16168), .A3(n16167), .ZN(P3_U2834) );
  NOR3_X1 U19212 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16171) );
  NOR4_X1 U19213 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16170) );
  NAND4_X1 U19214 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16171), .A3(n16170), .A4(
        U215), .ZN(U213) );
  INV_X1 U19215 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16264) );
  NOR2_X1 U19216 ( .A1(n16224), .A2(n16172), .ZN(n16225) );
  INV_X1 U19217 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16265) );
  OAI222_X1 U19218 ( .A1(U212), .A2(n16264), .B1(n16229), .B2(n16173), .C1(
        U214), .C2(n16265), .ZN(U216) );
  INV_X1 U19219 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16175) );
  INV_X1 U19220 ( .A(U212), .ZN(n16227) );
  AOI22_X1 U19221 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16227), .ZN(n16174) );
  OAI21_X1 U19222 ( .B1(n16175), .B2(n16229), .A(n16174), .ZN(U217) );
  INV_X1 U19223 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16177) );
  AOI22_X1 U19224 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16227), .ZN(n16176) );
  OAI21_X1 U19225 ( .B1(n16177), .B2(n16229), .A(n16176), .ZN(U218) );
  INV_X1 U19226 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16179) );
  AOI22_X1 U19227 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16227), .ZN(n16178) );
  OAI21_X1 U19228 ( .B1(n16179), .B2(n16229), .A(n16178), .ZN(U219) );
  INV_X1 U19229 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16181) );
  AOI22_X1 U19230 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16227), .ZN(n16180) );
  OAI21_X1 U19231 ( .B1(n16181), .B2(n16229), .A(n16180), .ZN(U220) );
  AOI22_X1 U19232 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16227), .ZN(n16182) );
  OAI21_X1 U19233 ( .B1(n16183), .B2(n16229), .A(n16182), .ZN(U221) );
  AOI22_X1 U19234 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16227), .ZN(n16184) );
  OAI21_X1 U19235 ( .B1(n16185), .B2(n16229), .A(n16184), .ZN(U222) );
  INV_X1 U19236 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16187) );
  AOI22_X1 U19237 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16227), .ZN(n16186) );
  OAI21_X1 U19238 ( .B1(n16187), .B2(n16229), .A(n16186), .ZN(U223) );
  AOI22_X1 U19239 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16227), .ZN(n16188) );
  OAI21_X1 U19240 ( .B1(n16189), .B2(n16229), .A(n16188), .ZN(U224) );
  AOI22_X1 U19241 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16227), .ZN(n16190) );
  OAI21_X1 U19242 ( .B1(n16191), .B2(n16229), .A(n16190), .ZN(U225) );
  AOI22_X1 U19243 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16227), .ZN(n16192) );
  OAI21_X1 U19244 ( .B1(n14929), .B2(n16229), .A(n16192), .ZN(U226) );
  INV_X1 U19245 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16194) );
  AOI22_X1 U19246 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16227), .ZN(n16193) );
  OAI21_X1 U19247 ( .B1(n16194), .B2(n16229), .A(n16193), .ZN(U227) );
  INV_X1 U19248 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n20696) );
  AOI22_X1 U19249 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n16225), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16224), .ZN(n16195) );
  OAI21_X1 U19250 ( .B1(n20696), .B2(U212), .A(n16195), .ZN(U228) );
  INV_X1 U19251 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16197) );
  AOI22_X1 U19252 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16227), .ZN(n16196) );
  OAI21_X1 U19253 ( .B1(n16197), .B2(n16229), .A(n16196), .ZN(U229) );
  AOI22_X1 U19254 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16227), .ZN(n16198) );
  OAI21_X1 U19255 ( .B1(n14032), .B2(n16229), .A(n16198), .ZN(U230) );
  AOI22_X1 U19256 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16227), .ZN(n16199) );
  OAI21_X1 U19257 ( .B1(n16200), .B2(n16229), .A(n16199), .ZN(U231) );
  INV_X1 U19258 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16202) );
  AOI22_X1 U19259 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16225), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16224), .ZN(n16201) );
  OAI21_X1 U19260 ( .B1(n16202), .B2(U212), .A(n16201), .ZN(U232) );
  INV_X1 U19261 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16204) );
  AOI22_X1 U19262 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16225), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16224), .ZN(n16203) );
  OAI21_X1 U19263 ( .B1(n16204), .B2(U212), .A(n16203), .ZN(U233) );
  INV_X1 U19264 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n20681) );
  AOI22_X1 U19265 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16225), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16227), .ZN(n16205) );
  OAI21_X1 U19266 ( .B1(n20681), .B2(U214), .A(n16205), .ZN(U234) );
  AOI22_X1 U19267 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16227), .ZN(n16206) );
  OAI21_X1 U19268 ( .B1(n16207), .B2(n16229), .A(n16206), .ZN(U235) );
  INV_X1 U19269 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16242) );
  AOI22_X1 U19270 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16225), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16224), .ZN(n16208) );
  OAI21_X1 U19271 ( .B1(n16242), .B2(U212), .A(n16208), .ZN(U236) );
  AOI22_X1 U19272 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16227), .ZN(n16209) );
  OAI21_X1 U19273 ( .B1(n16210), .B2(n16229), .A(n16209), .ZN(U237) );
  AOI22_X1 U19274 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16227), .ZN(n16211) );
  OAI21_X1 U19275 ( .B1(n16212), .B2(n16229), .A(n16211), .ZN(U238) );
  AOI22_X1 U19276 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16227), .ZN(n16213) );
  OAI21_X1 U19277 ( .B1(n16214), .B2(n16229), .A(n16213), .ZN(U239) );
  INV_X1 U19278 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16238) );
  AOI22_X1 U19279 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16225), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16224), .ZN(n16215) );
  OAI21_X1 U19280 ( .B1(n16238), .B2(U212), .A(n16215), .ZN(U240) );
  INV_X1 U19281 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16217) );
  AOI22_X1 U19282 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16227), .ZN(n16216) );
  OAI21_X1 U19283 ( .B1(n16217), .B2(n16229), .A(n16216), .ZN(U241) );
  INV_X1 U19284 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16236) );
  AOI22_X1 U19285 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16225), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16224), .ZN(n16218) );
  OAI21_X1 U19286 ( .B1(n16236), .B2(U212), .A(n16218), .ZN(U242) );
  INV_X1 U19287 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16220) );
  AOI22_X1 U19288 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16227), .ZN(n16219) );
  OAI21_X1 U19289 ( .B1(n16220), .B2(n16229), .A(n16219), .ZN(U243) );
  INV_X1 U19290 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16234) );
  AOI22_X1 U19291 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16225), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16224), .ZN(n16221) );
  OAI21_X1 U19292 ( .B1(n16234), .B2(U212), .A(n16221), .ZN(U244) );
  INV_X1 U19293 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16223) );
  AOI22_X1 U19294 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16227), .ZN(n16222) );
  OAI21_X1 U19295 ( .B1(n16223), .B2(n16229), .A(n16222), .ZN(U245) );
  INV_X1 U19296 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16232) );
  AOI22_X1 U19297 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16225), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16224), .ZN(n16226) );
  OAI21_X1 U19298 ( .B1(n16232), .B2(U212), .A(n16226), .ZN(U246) );
  INV_X1 U19299 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16230) );
  AOI22_X1 U19300 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16224), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16227), .ZN(n16228) );
  OAI21_X1 U19301 ( .B1(n16230), .B2(n16229), .A(n16228), .ZN(U247) );
  OAI22_X1 U19302 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16262), .ZN(n16231) );
  INV_X1 U19303 ( .A(n16231), .ZN(U251) );
  INV_X1 U19304 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U19305 ( .A1(n16262), .A2(n16232), .B1(n17958), .B2(U215), .ZN(U252) );
  OAI22_X1 U19306 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16249), .ZN(n16233) );
  INV_X1 U19307 ( .A(n16233), .ZN(U253) );
  INV_X1 U19308 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n17968) );
  AOI22_X1 U19309 ( .A1(n16262), .A2(n16234), .B1(n17968), .B2(U215), .ZN(U254) );
  OAI22_X1 U19310 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16249), .ZN(n16235) );
  INV_X1 U19311 ( .A(n16235), .ZN(U255) );
  INV_X1 U19312 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n17976) );
  AOI22_X1 U19313 ( .A1(n16262), .A2(n16236), .B1(n17976), .B2(U215), .ZN(U256) );
  OAI22_X1 U19314 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16249), .ZN(n16237) );
  INV_X1 U19315 ( .A(n16237), .ZN(U257) );
  INV_X1 U19316 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U19317 ( .A1(n16262), .A2(n16238), .B1(n17986), .B2(U215), .ZN(U258) );
  OAI22_X1 U19318 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16249), .ZN(n16239) );
  INV_X1 U19319 ( .A(n16239), .ZN(U259) );
  OAI22_X1 U19320 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16249), .ZN(n16240) );
  INV_X1 U19321 ( .A(n16240), .ZN(U260) );
  OAI22_X1 U19322 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16249), .ZN(n16241) );
  INV_X1 U19323 ( .A(n16241), .ZN(U261) );
  INV_X1 U19324 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U19325 ( .A1(n16262), .A2(n16242), .B1(n17242), .B2(U215), .ZN(U262) );
  OAI22_X1 U19326 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16249), .ZN(n16243) );
  INV_X1 U19327 ( .A(n16243), .ZN(U263) );
  OAI22_X1 U19328 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16262), .ZN(n16244) );
  INV_X1 U19329 ( .A(n16244), .ZN(U264) );
  OAI22_X1 U19330 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16249), .ZN(n16245) );
  INV_X1 U19331 ( .A(n16245), .ZN(U265) );
  OAI22_X1 U19332 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16262), .ZN(n16246) );
  INV_X1 U19333 ( .A(n16246), .ZN(U266) );
  OAI22_X1 U19334 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16249), .ZN(n16247) );
  INV_X1 U19335 ( .A(n16247), .ZN(U267) );
  OAI22_X1 U19336 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16262), .ZN(n16248) );
  INV_X1 U19337 ( .A(n16248), .ZN(U268) );
  OAI22_X1 U19338 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16249), .ZN(n16250) );
  INV_X1 U19339 ( .A(n16250), .ZN(U269) );
  AOI22_X1 U19340 ( .A1(n16262), .A2(n20696), .B1(n14142), .B2(U215), .ZN(U270) );
  OAI22_X1 U19341 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16262), .ZN(n16251) );
  INV_X1 U19342 ( .A(n16251), .ZN(U271) );
  OAI22_X1 U19343 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16262), .ZN(n16252) );
  INV_X1 U19344 ( .A(n16252), .ZN(U272) );
  OAI22_X1 U19345 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16262), .ZN(n16253) );
  INV_X1 U19346 ( .A(n16253), .ZN(U273) );
  OAI22_X1 U19347 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16262), .ZN(n16254) );
  INV_X1 U19348 ( .A(n16254), .ZN(U274) );
  OAI22_X1 U19349 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16262), .ZN(n16255) );
  INV_X1 U19350 ( .A(n16255), .ZN(U275) );
  OAI22_X1 U19351 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16262), .ZN(n16256) );
  INV_X1 U19352 ( .A(n16256), .ZN(U276) );
  OAI22_X1 U19353 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16262), .ZN(n16257) );
  INV_X1 U19354 ( .A(n16257), .ZN(U277) );
  OAI22_X1 U19355 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16262), .ZN(n16258) );
  INV_X1 U19356 ( .A(n16258), .ZN(U278) );
  OAI22_X1 U19357 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16262), .ZN(n16259) );
  INV_X1 U19358 ( .A(n16259), .ZN(U279) );
  OAI22_X1 U19359 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16262), .ZN(n16260) );
  INV_X1 U19360 ( .A(n16260), .ZN(U280) );
  OAI22_X1 U19361 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16262), .ZN(n16261) );
  INV_X1 U19362 ( .A(n16261), .ZN(U281) );
  AOI22_X1 U19363 ( .A1(n16262), .A2(n16264), .B1(n16997), .B2(U215), .ZN(U282) );
  INV_X1 U19364 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16263) );
  AOI222_X1 U19365 ( .A1(n16265), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16264), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16263), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16266) );
  INV_X2 U19366 ( .A(n16268), .ZN(n16267) );
  INV_X1 U19367 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18501) );
  INV_X1 U19368 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19623) );
  AOI22_X1 U19369 ( .A1(n16267), .A2(n18501), .B1(n19623), .B2(n16268), .ZN(
        U347) );
  INV_X1 U19370 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18499) );
  INV_X1 U19371 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19621) );
  AOI22_X1 U19372 ( .A1(n16266), .A2(n18499), .B1(n19621), .B2(n16268), .ZN(
        U348) );
  INV_X1 U19373 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18496) );
  INV_X1 U19374 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20683) );
  AOI22_X1 U19375 ( .A1(n16267), .A2(n18496), .B1(n20683), .B2(n16268), .ZN(
        U349) );
  INV_X1 U19376 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18495) );
  INV_X1 U19377 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19618) );
  AOI22_X1 U19378 ( .A1(n16267), .A2(n18495), .B1(n19618), .B2(n16268), .ZN(
        U350) );
  INV_X1 U19379 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18493) );
  INV_X1 U19380 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19617) );
  AOI22_X1 U19381 ( .A1(n16267), .A2(n18493), .B1(n19617), .B2(n16268), .ZN(
        U351) );
  INV_X1 U19382 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18490) );
  INV_X1 U19383 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19615) );
  AOI22_X1 U19384 ( .A1(n16267), .A2(n18490), .B1(n19615), .B2(n16268), .ZN(
        U352) );
  INV_X1 U19385 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18489) );
  INV_X1 U19386 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19613) );
  AOI22_X1 U19387 ( .A1(n16267), .A2(n18489), .B1(n19613), .B2(n16268), .ZN(
        U353) );
  INV_X1 U19388 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18487) );
  AOI22_X1 U19389 ( .A1(n16267), .A2(n18487), .B1(n19611), .B2(n16268), .ZN(
        U354) );
  INV_X1 U19390 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18544) );
  INV_X1 U19391 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19658) );
  AOI22_X1 U19392 ( .A1(n16267), .A2(n18544), .B1(n19658), .B2(n16268), .ZN(
        U355) );
  INV_X1 U19393 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18539) );
  INV_X1 U19394 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19654) );
  AOI22_X1 U19395 ( .A1(n16267), .A2(n18539), .B1(n19654), .B2(n16268), .ZN(
        U356) );
  INV_X1 U19396 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18537) );
  INV_X1 U19397 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19652) );
  AOI22_X1 U19398 ( .A1(n16267), .A2(n18537), .B1(n19652), .B2(n16268), .ZN(
        U357) );
  INV_X1 U19399 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18534) );
  INV_X1 U19400 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20678) );
  AOI22_X1 U19401 ( .A1(n16267), .A2(n18534), .B1(n20678), .B2(n16268), .ZN(
        U358) );
  INV_X1 U19402 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18533) );
  INV_X1 U19403 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U19404 ( .A1(n16267), .A2(n18533), .B1(n19650), .B2(n16268), .ZN(
        U359) );
  INV_X1 U19405 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18531) );
  INV_X1 U19406 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19648) );
  AOI22_X1 U19407 ( .A1(n16267), .A2(n18531), .B1(n19648), .B2(n16268), .ZN(
        U360) );
  INV_X1 U19408 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18529) );
  INV_X1 U19409 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19646) );
  AOI22_X1 U19410 ( .A1(n16267), .A2(n18529), .B1(n19646), .B2(n16268), .ZN(
        U361) );
  INV_X1 U19411 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18527) );
  INV_X1 U19412 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19645) );
  AOI22_X1 U19413 ( .A1(n16267), .A2(n18527), .B1(n19645), .B2(n16268), .ZN(
        U362) );
  INV_X1 U19414 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18525) );
  INV_X1 U19415 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19643) );
  AOI22_X1 U19416 ( .A1(n16267), .A2(n18525), .B1(n19643), .B2(n16268), .ZN(
        U363) );
  INV_X1 U19417 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18523) );
  INV_X1 U19418 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19642) );
  AOI22_X1 U19419 ( .A1(n16267), .A2(n18523), .B1(n19642), .B2(n16268), .ZN(
        U364) );
  INV_X1 U19420 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18485) );
  INV_X1 U19421 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19610) );
  AOI22_X1 U19422 ( .A1(n16267), .A2(n18485), .B1(n19610), .B2(n16268), .ZN(
        U365) );
  INV_X1 U19423 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18520) );
  INV_X1 U19424 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U19425 ( .A1(n16267), .A2(n18520), .B1(n19640), .B2(n16268), .ZN(
        U366) );
  INV_X1 U19426 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18519) );
  INV_X1 U19427 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19638) );
  AOI22_X1 U19428 ( .A1(n16267), .A2(n18519), .B1(n19638), .B2(n16268), .ZN(
        U367) );
  INV_X1 U19429 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18517) );
  INV_X1 U19430 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19636) );
  AOI22_X1 U19431 ( .A1(n16267), .A2(n18517), .B1(n19636), .B2(n16268), .ZN(
        U368) );
  INV_X1 U19432 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18515) );
  INV_X1 U19433 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19635) );
  AOI22_X1 U19434 ( .A1(n16267), .A2(n18515), .B1(n19635), .B2(n16268), .ZN(
        U369) );
  INV_X1 U19435 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18513) );
  INV_X1 U19436 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19633) );
  AOI22_X1 U19437 ( .A1(n16267), .A2(n18513), .B1(n19633), .B2(n16268), .ZN(
        U370) );
  INV_X1 U19438 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18511) );
  INV_X1 U19439 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19631) );
  AOI22_X1 U19440 ( .A1(n16266), .A2(n18511), .B1(n19631), .B2(n16268), .ZN(
        U371) );
  INV_X1 U19441 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18508) );
  INV_X1 U19442 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19629) );
  AOI22_X1 U19443 ( .A1(n16267), .A2(n18508), .B1(n19629), .B2(n16268), .ZN(
        U372) );
  INV_X1 U19444 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18507) );
  INV_X1 U19445 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19627) );
  AOI22_X1 U19446 ( .A1(n16267), .A2(n18507), .B1(n19627), .B2(n16268), .ZN(
        U373) );
  INV_X1 U19447 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18505) );
  INV_X1 U19448 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19626) );
  AOI22_X1 U19449 ( .A1(n16267), .A2(n18505), .B1(n19626), .B2(n16268), .ZN(
        U374) );
  INV_X1 U19450 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18503) );
  INV_X1 U19451 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19624) );
  AOI22_X1 U19452 ( .A1(n16266), .A2(n18503), .B1(n19624), .B2(n16268), .ZN(
        U375) );
  INV_X1 U19453 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18483) );
  INV_X1 U19454 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19609) );
  AOI22_X1 U19455 ( .A1(n16266), .A2(n18483), .B1(n19609), .B2(n16268), .ZN(
        U376) );
  INV_X1 U19456 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18482) );
  NAND2_X1 U19457 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18482), .ZN(n18470) );
  AOI22_X1 U19458 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18470), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18480), .ZN(n18552) );
  AOI21_X1 U19459 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18552), .ZN(n16269) );
  INV_X1 U19460 ( .A(n16269), .ZN(P3_U2633) );
  NOR2_X1 U19461 ( .A1(n16277), .A2(n17208), .ZN(n16270) );
  OAI21_X1 U19462 ( .B1(n16270), .B2(n17143), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16271) );
  OAI21_X1 U19463 ( .B1(n16272), .B2(n18455), .A(n16271), .ZN(P3_U2634) );
  AOI21_X1 U19464 ( .B1(n18480), .B2(n18482), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16273) );
  AOI22_X1 U19465 ( .A1(n18543), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16273), 
        .B2(n18615), .ZN(P3_U2635) );
  OAI21_X1 U19466 ( .B1(n16274), .B2(BS16), .A(n18552), .ZN(n18550) );
  OAI21_X1 U19467 ( .B1(n18552), .B2(n16275), .A(n18550), .ZN(P3_U2636) );
  OAI211_X1 U19468 ( .C1(n16277), .C2(n17208), .A(n16276), .B(n18389), .ZN(
        n16278) );
  INV_X1 U19469 ( .A(n16278), .ZN(n18392) );
  NOR2_X1 U19470 ( .A1(n18392), .A2(n18452), .ZN(n18597) );
  OAI21_X1 U19471 ( .B1(n18597), .B2(n17939), .A(n16279), .ZN(P3_U2637) );
  NOR4_X1 U19472 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16283) );
  NOR4_X1 U19473 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16282) );
  NOR4_X1 U19474 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16281) );
  NOR4_X1 U19475 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16280) );
  NAND4_X1 U19476 ( .A1(n16283), .A2(n16282), .A3(n16281), .A4(n16280), .ZN(
        n16289) );
  NOR4_X1 U19477 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16287) );
  AOI211_X1 U19478 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_28__SCAN_IN), .B(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16286) );
  NOR4_X1 U19479 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16285) );
  NOR4_X1 U19480 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16284) );
  NAND4_X1 U19481 ( .A1(n16287), .A2(n16286), .A3(n16285), .A4(n16284), .ZN(
        n16288) );
  NOR2_X1 U19482 ( .A1(n16289), .A2(n16288), .ZN(n16295) );
  NOR2_X1 U19483 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18589) );
  INV_X1 U19484 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n16292) );
  AOI21_X1 U19485 ( .B1(n18589), .B2(n16292), .A(P3_REIP_REG_1__SCAN_IN), .ZN(
        n16291) );
  INV_X1 U19486 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16290) );
  INV_X1 U19487 ( .A(n16295), .ZN(n18595) );
  AOI22_X1 U19488 ( .A1(n16295), .A2(n16291), .B1(n16290), .B2(n18595), .ZN(
        P3_U2638) );
  INV_X1 U19489 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18588) );
  INV_X1 U19490 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18551) );
  AOI22_X1 U19491 ( .A1(n18589), .A2(n16292), .B1(n18588), .B2(n18551), .ZN(
        n16294) );
  INV_X1 U19492 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16293) );
  AOI22_X1 U19493 ( .A1(n16295), .A2(n16294), .B1(n16293), .B2(n18595), .ZN(
        P3_U2639) );
  INV_X1 U19494 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18542) );
  INV_X1 U19495 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18530) );
  INV_X1 U19496 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18526) );
  NAND3_X1 U19497 ( .A1(n16426), .A2(P3_REIP_REG_22__SCAN_IN), .A3(
        P3_REIP_REG_21__SCAN_IN), .ZN(n16405) );
  NOR2_X1 U19498 ( .A1(n18526), .A2(n16405), .ZN(n16403) );
  NAND2_X1 U19499 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16403), .ZN(n16380) );
  NOR2_X1 U19500 ( .A1(n18530), .A2(n16380), .ZN(n16367) );
  NAND2_X1 U19501 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16367), .ZN(n16312) );
  NOR2_X1 U19502 ( .A1(n16659), .A2(n16312), .ZN(n16363) );
  NAND4_X1 U19503 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16363), .ZN(n16314) );
  NOR3_X1 U19504 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18542), .A3(n16314), 
        .ZN(n16296) );
  AOI21_X1 U19505 ( .B1(n16646), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16296), .ZN(
        n16320) );
  INV_X1 U19506 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20744) );
  NAND2_X1 U19507 ( .A1(n16431), .A2(n20744), .ZN(n16430) );
  NAND2_X1 U19508 ( .A1(n16413), .A2(n16409), .ZN(n16408) );
  NAND2_X1 U19509 ( .A1(n16391), .A2(n16386), .ZN(n16385) );
  INV_X1 U19510 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16709) );
  NAND2_X1 U19511 ( .A1(n16368), .A2(n16709), .ZN(n16364) );
  NOR2_X1 U19512 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16364), .ZN(n16346) );
  INV_X1 U19513 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16705) );
  NAND2_X1 U19514 ( .A1(n16346), .A2(n16705), .ZN(n16322) );
  NOR2_X1 U19515 ( .A1(n16665), .A2(n16322), .ZN(n16329) );
  INV_X1 U19516 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16318) );
  OAI21_X1 U19517 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16307), .A(
        n16297), .ZN(n17259) );
  INV_X1 U19518 ( .A(n17259), .ZN(n16359) );
  INV_X1 U19519 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16381) );
  NAND2_X1 U19520 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17280), .ZN(
        n16299) );
  AOI21_X1 U19521 ( .B1(n16381), .B2(n16299), .A(n16298), .ZN(n17281) );
  INV_X1 U19522 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17297) );
  OAI22_X1 U19523 ( .A1(n17297), .A2(n16300), .B1(n17280), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17295) );
  INV_X1 U19524 ( .A(n17295), .ZN(n16394) );
  INV_X1 U19525 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17326) );
  NAND3_X1 U19526 ( .A1(n17325), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16301) );
  NOR2_X1 U19527 ( .A1(n17312), .A2(n17602), .ZN(n16304) );
  AOI21_X1 U19528 ( .B1(n17326), .B2(n16301), .A(n16304), .ZN(n17329) );
  NOR2_X1 U19529 ( .A1(n16302), .A2(n16599), .ZN(n16425) );
  INV_X1 U19530 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17341) );
  NAND2_X1 U19531 ( .A1(n17325), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16303) );
  XOR2_X1 U19532 ( .A(n17341), .B(n16303), .Z(n17344) );
  NOR2_X1 U19533 ( .A1(n16414), .A2(n16599), .ZN(n16402) );
  INV_X1 U19534 ( .A(n16402), .ZN(n16306) );
  NOR2_X1 U19535 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16304), .ZN(
        n17308) );
  NOR2_X1 U19536 ( .A1(n17280), .A2(n17308), .ZN(n17315) );
  NAND2_X1 U19537 ( .A1(n16306), .A2(n16305), .ZN(n16400) );
  NOR2_X1 U19538 ( .A1(n16392), .A2(n16599), .ZN(n16379) );
  NOR2_X1 U19539 ( .A1(n17281), .A2(n16379), .ZN(n16378) );
  NOR2_X1 U19540 ( .A1(n16378), .A2(n16599), .ZN(n16371) );
  AOI21_X1 U19541 ( .B1(n16309), .B2(n16308), .A(n16307), .ZN(n17272) );
  INV_X1 U19542 ( .A(n17272), .ZN(n16310) );
  NOR2_X1 U19543 ( .A1(n16357), .A2(n16599), .ZN(n16348) );
  NOR2_X1 U19544 ( .A1(n16349), .A2(n16348), .ZN(n16347) );
  OR2_X1 U19545 ( .A1(n16347), .A2(n16599), .ZN(n16332) );
  INV_X1 U19546 ( .A(n16336), .ZN(n16311) );
  NAND2_X1 U19547 ( .A1(n16332), .A2(n16311), .ZN(n16333) );
  NOR4_X1 U19548 ( .A1(n16324), .A2(n16323), .A3(n16599), .A4(n18460), .ZN(
        n16317) );
  NOR2_X1 U19549 ( .A1(n16653), .A2(n16648), .ZN(n16439) );
  INV_X1 U19550 ( .A(n16439), .ZN(n16667) );
  NAND3_X1 U19551 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16313) );
  AOI21_X1 U19552 ( .B1(n16312), .B2(n16648), .A(n16653), .ZN(n16376) );
  INV_X1 U19553 ( .A(n16376), .ZN(n16352) );
  AOI21_X1 U19554 ( .B1(n16667), .B2(n16313), .A(n16352), .ZN(n16345) );
  NOR2_X1 U19555 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16314), .ZN(n16327) );
  INV_X1 U19556 ( .A(n16327), .ZN(n16315) );
  INV_X1 U19557 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18545) );
  AOI21_X1 U19558 ( .B1(n16345), .B2(n16315), .A(n18545), .ZN(n16316) );
  AOI211_X1 U19559 ( .C1(n16329), .C2(n16318), .A(n16317), .B(n16316), .ZN(
        n16319) );
  OAI211_X1 U19560 ( .C1(n16321), .C2(n16656), .A(n16320), .B(n16319), .ZN(
        P3_U2640) );
  NAND2_X1 U19561 ( .A1(n16654), .A2(n16322), .ZN(n16341) );
  XOR2_X1 U19562 ( .A(n16324), .B(n16323), .Z(n16328) );
  INV_X1 U19563 ( .A(n18460), .ZN(n16655) );
  OAI22_X1 U19564 ( .A1(n16345), .A2(n18542), .B1(n16325), .B2(n16656), .ZN(
        n16326) );
  OAI21_X1 U19565 ( .B1(n16646), .B2(n16329), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16330) );
  OAI211_X1 U19566 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16341), .A(n16331), .B(
        n16330), .ZN(P3_U2641) );
  INV_X1 U19567 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18538) );
  INV_X1 U19568 ( .A(n16332), .ZN(n16335) );
  INV_X1 U19569 ( .A(n16333), .ZN(n16334) );
  AOI211_X1 U19570 ( .C1(n16336), .C2(n16335), .A(n16334), .B(n18460), .ZN(
        n16340) );
  NAND3_X1 U19571 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16363), .ZN(n16338) );
  OAI22_X1 U19572 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16338), .B1(n16337), 
        .B2(n16656), .ZN(n16339) );
  AOI211_X1 U19573 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16646), .A(n16340), .B(
        n16339), .ZN(n16344) );
  INV_X1 U19574 ( .A(n16341), .ZN(n16342) );
  OAI21_X1 U19575 ( .B1(n16346), .B2(n16705), .A(n16342), .ZN(n16343) );
  OAI211_X1 U19576 ( .C1(n16345), .C2(n18538), .A(n16344), .B(n16343), .ZN(
        P3_U2642) );
  AOI22_X1 U19577 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16610), .B1(
        n16646), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16356) );
  AOI211_X1 U19578 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16364), .A(n16346), .B(
        n16665), .ZN(n16351) );
  AOI211_X1 U19579 ( .C1(n16349), .C2(n16348), .A(n16347), .B(n18460), .ZN(
        n16350) );
  AOI211_X1 U19580 ( .C1(n16352), .C2(P3_REIP_REG_28__SCAN_IN), .A(n16351), 
        .B(n16350), .ZN(n16355) );
  NAND2_X1 U19581 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16353) );
  OAI211_X1 U19582 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16363), .B(n16353), .ZN(n16354) );
  NAND3_X1 U19583 ( .A1(n16356), .A2(n16355), .A3(n16354), .ZN(P3_U2643) );
  INV_X1 U19584 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18535) );
  AOI211_X1 U19585 ( .C1(n16359), .C2(n16358), .A(n16357), .B(n18460), .ZN(
        n16362) );
  OAI22_X1 U19586 ( .A1(n16360), .A2(n16656), .B1(n16666), .B2(n16709), .ZN(
        n16361) );
  AOI211_X1 U19587 ( .C1(n16363), .C2(n18535), .A(n16362), .B(n16361), .ZN(
        n16366) );
  OAI211_X1 U19588 ( .C1(n16368), .C2(n16709), .A(n16654), .B(n16364), .ZN(
        n16365) );
  OAI211_X1 U19589 ( .C1(n16376), .C2(n18535), .A(n16366), .B(n16365), .ZN(
        P3_U2644) );
  AOI21_X1 U19590 ( .B1(n16648), .B2(n16367), .A(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n16377) );
  AOI22_X1 U19591 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16610), .B1(
        n16646), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16375) );
  AOI211_X1 U19592 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16385), .A(n16368), .B(
        n16665), .ZN(n16373) );
  INV_X1 U19593 ( .A(n16369), .ZN(n16370) );
  AOI211_X1 U19594 ( .C1(n17272), .C2(n16371), .A(n16370), .B(n18460), .ZN(
        n16372) );
  NOR2_X1 U19595 ( .A1(n16373), .A2(n16372), .ZN(n16374) );
  OAI211_X1 U19596 ( .C1(n16377), .C2(n16376), .A(n16375), .B(n16374), .ZN(
        P3_U2645) );
  INV_X1 U19597 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18528) );
  OAI21_X1 U19598 ( .B1(n16403), .B2(n16659), .A(n16669), .ZN(n16399) );
  AOI21_X1 U19599 ( .B1(n16648), .B2(n18528), .A(n16399), .ZN(n16389) );
  AOI211_X1 U19600 ( .C1(n17281), .C2(n16379), .A(n16378), .B(n18460), .ZN(
        n16384) );
  NOR3_X1 U19601 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16659), .A3(n16380), 
        .ZN(n16383) );
  OAI22_X1 U19602 ( .A1(n16381), .A2(n16656), .B1(n16666), .B2(n16386), .ZN(
        n16382) );
  NOR3_X1 U19603 ( .A1(n16384), .A2(n16383), .A3(n16382), .ZN(n16388) );
  OAI211_X1 U19604 ( .C1(n16391), .C2(n16386), .A(n16654), .B(n16385), .ZN(
        n16387) );
  OAI211_X1 U19605 ( .C1(n16389), .C2(n18530), .A(n16388), .B(n16387), .ZN(
        P3_U2646) );
  NOR2_X1 U19606 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16659), .ZN(n16390) );
  AOI22_X1 U19607 ( .A1(n16646), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16403), 
        .B2(n16390), .ZN(n16398) );
  AOI211_X1 U19608 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16408), .A(n16391), .B(
        n16665), .ZN(n16396) );
  AOI211_X1 U19609 ( .C1(n16394), .C2(n16393), .A(n16392), .B(n18460), .ZN(
        n16395) );
  AOI211_X1 U19610 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16399), .A(n16396), 
        .B(n16395), .ZN(n16397) );
  OAI211_X1 U19611 ( .C1(n17297), .C2(n16656), .A(n16398), .B(n16397), .ZN(
        P3_U2647) );
  INV_X1 U19612 ( .A(n16399), .ZN(n16412) );
  INV_X1 U19613 ( .A(n16400), .ZN(n16401) );
  AOI211_X1 U19614 ( .C1(n17315), .C2(n16402), .A(n16401), .B(n18460), .ZN(
        n16407) );
  OR2_X1 U19615 ( .A1(n16659), .A2(n16403), .ZN(n16404) );
  OAI22_X1 U19616 ( .A1(n16666), .A2(n16409), .B1(n16405), .B2(n16404), .ZN(
        n16406) );
  AOI211_X1 U19617 ( .C1(n16610), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16407), .B(n16406), .ZN(n16411) );
  OAI211_X1 U19618 ( .C1(n16413), .C2(n16409), .A(n16654), .B(n16408), .ZN(
        n16410) );
  OAI211_X1 U19619 ( .C1(n16412), .C2(n18526), .A(n16411), .B(n16410), .ZN(
        P3_U2648) );
  INV_X1 U19620 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18524) );
  INV_X1 U19621 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18522) );
  NOR2_X1 U19622 ( .A1(n18524), .A2(n18522), .ZN(n16421) );
  OAI211_X1 U19623 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16426), .B(n16648), .ZN(n16420) );
  AOI22_X1 U19624 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16610), .B1(
        n16646), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16419) );
  AOI211_X1 U19625 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16430), .A(n16413), .B(
        n16665), .ZN(n16417) );
  AOI211_X1 U19626 ( .C1(n17329), .C2(n16415), .A(n16414), .B(n18460), .ZN(
        n16416) );
  AOI211_X1 U19627 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16422), .A(n16417), 
        .B(n16416), .ZN(n16418) );
  OAI211_X1 U19628 ( .C1(n16421), .C2(n16420), .A(n16419), .B(n16418), .ZN(
        P3_U2649) );
  INV_X1 U19629 ( .A(n16422), .ZN(n16434) );
  INV_X1 U19630 ( .A(n16423), .ZN(n16424) );
  AOI211_X1 U19631 ( .C1(n17344), .C2(n16425), .A(n16424), .B(n18460), .ZN(
        n16429) );
  NAND2_X1 U19632 ( .A1(n16648), .A2(n16426), .ZN(n16427) );
  OAI22_X1 U19633 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16427), .B1(n16666), 
        .B2(n20744), .ZN(n16428) );
  AOI211_X1 U19634 ( .C1(n16610), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16429), .B(n16428), .ZN(n16433) );
  OAI211_X1 U19635 ( .C1(n16431), .C2(n20744), .A(n16654), .B(n16430), .ZN(
        n16432) );
  OAI211_X1 U19636 ( .C1(n16434), .C2(n18522), .A(n16433), .B(n16432), .ZN(
        P3_U2650) );
  OAI21_X1 U19637 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16447), .A(
        n17323), .ZN(n17366) );
  OAI21_X1 U19638 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17404), .A(
        n9589), .ZN(n16478) );
  OAI21_X1 U19639 ( .B1(n16447), .B2(n16599), .A(n16478), .ZN(n16435) );
  XOR2_X1 U19640 ( .A(n17366), .B(n16435), .Z(n16444) );
  INV_X1 U19641 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17367) );
  OAI211_X1 U19642 ( .C1(n16445), .C2(n16770), .A(n16654), .B(n16436), .ZN(
        n16437) );
  OAI211_X1 U19643 ( .C1(n17367), .C2(n16656), .A(n17930), .B(n16437), .ZN(
        n16438) );
  AOI21_X1 U19644 ( .B1(n16646), .B2(P3_EBX_REG_19__SCAN_IN), .A(n16438), .ZN(
        n16443) );
  AOI21_X1 U19645 ( .B1(n16648), .B2(n16490), .A(n16653), .ZN(n16499) );
  OAI21_X1 U19646 ( .B1(n16439), .B2(n16440), .A(n16499), .ZN(n16458) );
  INV_X1 U19647 ( .A(n16487), .ZN(n16474) );
  AND2_X1 U19648 ( .A1(n16440), .A2(n16474), .ZN(n16451) );
  INV_X1 U19649 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18518) );
  INV_X1 U19650 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18516) );
  XOR2_X1 U19651 ( .A(n18518), .B(n18516), .Z(n16441) );
  AOI22_X1 U19652 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16458), .B1(n16451), 
        .B2(n16441), .ZN(n16442) );
  OAI211_X1 U19653 ( .C1(n18460), .C2(n16444), .A(n16443), .B(n16442), .ZN(
        P3_U2652) );
  AOI211_X1 U19654 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16460), .A(n16445), .B(
        n16665), .ZN(n16446) );
  AOI211_X1 U19655 ( .C1(n16646), .C2(P3_EBX_REG_18__SCAN_IN), .A(n17932), .B(
        n16446), .ZN(n16453) );
  AOI21_X1 U19656 ( .B1(n17377), .B2(n17365), .A(n16447), .ZN(n17380) );
  OAI21_X1 U19657 ( .B1(n17365), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n9589), .ZN(n16456) );
  INV_X1 U19658 ( .A(n16456), .ZN(n16449) );
  OAI21_X1 U19659 ( .B1(n17380), .B2(n16449), .A(n16655), .ZN(n16448) );
  AOI21_X1 U19660 ( .B1(n17380), .B2(n16449), .A(n16448), .ZN(n16450) );
  AOI221_X1 U19661 ( .B1(n16451), .B2(n18516), .C1(n16458), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n16450), .ZN(n16452) );
  OAI211_X1 U19662 ( .C1(n17377), .C2(n16656), .A(n16453), .B(n16452), .ZN(
        P3_U2653) );
  AOI22_X1 U19663 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16610), .B1(
        n16646), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16463) );
  NOR2_X1 U19664 ( .A1(n16473), .A2(n16487), .ZN(n16459) );
  OAI21_X1 U19665 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16464), .A(
        n17365), .ZN(n17394) );
  NAND2_X1 U19666 ( .A1(n16655), .A2(n16599), .ZN(n16643) );
  NOR2_X1 U19667 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17404), .ZN(
        n16454) );
  OAI221_X1 U19668 ( .B1(n17394), .B2(n17408), .C1(n17394), .C2(n16454), .A(
        n16655), .ZN(n16455) );
  AOI22_X1 U19669 ( .A1(n16456), .A2(n17394), .B1(n16643), .B2(n16455), .ZN(
        n16457) );
  AOI221_X1 U19670 ( .B1(n16459), .B2(n18514), .C1(n16458), .C2(
        P3_REIP_REG_17__SCAN_IN), .A(n16457), .ZN(n16462) );
  OAI211_X1 U19671 ( .C1(n16469), .C2(n16797), .A(n16654), .B(n16460), .ZN(
        n16461) );
  NAND4_X1 U19672 ( .A1(n16463), .A2(n16462), .A3(n17930), .A4(n16461), .ZN(
        P3_U2654) );
  INV_X1 U19673 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18512) );
  INV_X1 U19674 ( .A(n16464), .ZN(n16465) );
  OAI21_X1 U19675 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16477), .A(
        n16465), .ZN(n17405) );
  OR2_X1 U19676 ( .A1(n16466), .A2(n16599), .ZN(n16468) );
  OAI21_X1 U19677 ( .B1(n17405), .B2(n16468), .A(n16655), .ZN(n16467) );
  AOI21_X1 U19678 ( .B1(n17405), .B2(n16468), .A(n16467), .ZN(n16472) );
  AOI211_X1 U19679 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16481), .A(n16469), .B(
        n16665), .ZN(n16471) );
  INV_X1 U19680 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17406) );
  INV_X1 U19681 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16796) );
  OAI22_X1 U19682 ( .A1(n17406), .A2(n16656), .B1(n16666), .B2(n16796), .ZN(
        n16470) );
  NOR4_X1 U19683 ( .A1(n17627), .A2(n16472), .A3(n16471), .A4(n16470), .ZN(
        n16476) );
  OAI211_X1 U19684 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16474), .B(n16473), .ZN(n16475) );
  OAI211_X1 U19685 ( .C1(n16499), .C2(n18512), .A(n16476), .B(n16475), .ZN(
        P3_U2655) );
  INV_X1 U19686 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18510) );
  AOI21_X1 U19687 ( .B1(n17415), .B2(n17404), .A(n16477), .ZN(n17418) );
  INV_X1 U19688 ( .A(n16478), .ZN(n16480) );
  INV_X1 U19689 ( .A(n17418), .ZN(n16479) );
  AOI221_X1 U19690 ( .B1(n17418), .B2(n16480), .C1(n16479), .C2(n16478), .A(
        n18460), .ZN(n16485) );
  OAI211_X1 U19691 ( .C1(n16489), .C2(n16483), .A(n16654), .B(n16481), .ZN(
        n16482) );
  OAI211_X1 U19692 ( .C1(n16666), .C2(n16483), .A(n17930), .B(n16482), .ZN(
        n16484) );
  AOI211_X1 U19693 ( .C1(n16610), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16485), .B(n16484), .ZN(n16486) );
  OAI221_X1 U19694 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16487), .C1(n18510), 
        .C2(n16499), .A(n16486), .ZN(P3_U2656) );
  INV_X1 U19695 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18509) );
  AOI22_X1 U19696 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16610), .B1(
        n16646), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16498) );
  NOR2_X1 U19697 ( .A1(n17429), .A2(n17602), .ZN(n16502) );
  AOI21_X1 U19698 ( .B1(n16502), .B2(n16658), .A(n16599), .ZN(n16488) );
  OAI21_X1 U19699 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16502), .A(
        n17404), .ZN(n17441) );
  XNOR2_X1 U19700 ( .A(n16488), .B(n17441), .ZN(n16496) );
  AOI211_X1 U19701 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16504), .A(n16489), .B(
        n16665), .ZN(n16495) );
  INV_X1 U19702 ( .A(n16490), .ZN(n16493) );
  NAND2_X1 U19703 ( .A1(n16648), .A2(n16491), .ZN(n16492) );
  OAI21_X1 U19704 ( .B1(n16493), .B2(n16492), .A(n17930), .ZN(n16494) );
  AOI211_X1 U19705 ( .C1(n16496), .C2(n16655), .A(n16495), .B(n16494), .ZN(
        n16497) );
  OAI211_X1 U19706 ( .C1(n18509), .C2(n16499), .A(n16498), .B(n16497), .ZN(
        P3_U2657) );
  OR2_X1 U19707 ( .A1(n16500), .A2(n16653), .ZN(n16545) );
  OAI21_X1 U19708 ( .B1(n16501), .B2(n16545), .A(n16667), .ZN(n16530) );
  INV_X1 U19709 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18504) );
  NAND2_X1 U19710 ( .A1(n16648), .A2(n18504), .ZN(n16517) );
  INV_X1 U19711 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17448) );
  NAND2_X1 U19712 ( .A1(n17479), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17443) );
  NOR2_X1 U19713 ( .A1(n17448), .A2(n17443), .ZN(n16513) );
  AOI21_X1 U19714 ( .B1(n16513), .B2(n16658), .A(n16599), .ZN(n16514) );
  INV_X1 U19715 ( .A(n16502), .ZN(n16503) );
  OAI21_X1 U19716 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16513), .A(
        n16503), .ZN(n17449) );
  XNOR2_X1 U19717 ( .A(n16514), .B(n17449), .ZN(n16511) );
  INV_X1 U19718 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17447) );
  OAI22_X1 U19719 ( .A1(n17447), .A2(n16656), .B1(n16666), .B2(n16505), .ZN(
        n16510) );
  NAND2_X1 U19720 ( .A1(n16648), .A2(n18506), .ZN(n16507) );
  OAI211_X1 U19721 ( .C1(n16515), .C2(n16505), .A(n16654), .B(n16504), .ZN(
        n16506) );
  OAI211_X1 U19722 ( .C1(n16508), .C2(n16507), .A(n17930), .B(n16506), .ZN(
        n16509) );
  AOI211_X1 U19723 ( .C1(n16655), .C2(n16511), .A(n16510), .B(n16509), .ZN(
        n16512) );
  OAI221_X1 U19724 ( .B1(n18506), .B2(n16530), .C1(n18506), .C2(n16517), .A(
        n16512), .ZN(P3_U2658) );
  AOI21_X1 U19725 ( .B1(n17448), .B2(n17443), .A(n16513), .ZN(n17464) );
  NAND2_X1 U19726 ( .A1(n16655), .A2(n16514), .ZN(n16525) );
  AOI211_X1 U19727 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16533), .A(n16515), .B(
        n16665), .ZN(n16521) );
  INV_X1 U19728 ( .A(n16516), .ZN(n16518) );
  OAI22_X1 U19729 ( .A1(n17448), .A2(n16656), .B1(n16518), .B2(n16517), .ZN(
        n16520) );
  INV_X1 U19730 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16885) );
  OAI22_X1 U19731 ( .A1(n16666), .A2(n16885), .B1(n18504), .B2(n16530), .ZN(
        n16519) );
  NOR4_X1 U19732 ( .A1(n17627), .A2(n16521), .A3(n16520), .A4(n16519), .ZN(
        n16524) );
  INV_X1 U19733 ( .A(n17443), .ZN(n16522) );
  AOI21_X1 U19734 ( .B1(n9589), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18460), .ZN(n16662) );
  OAI211_X1 U19735 ( .C1(n16522), .C2(n16599), .A(n17464), .B(n16662), .ZN(
        n16523) );
  OAI211_X1 U19736 ( .C1(n17464), .C2(n16525), .A(n16524), .B(n16523), .ZN(
        P3_U2659) );
  INV_X1 U19737 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18500) );
  INV_X1 U19738 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18498) );
  NOR2_X1 U19739 ( .A1(n18500), .A2(n18498), .ZN(n16547) );
  INV_X1 U19740 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18497) );
  NOR4_X1 U19741 ( .A1(n16659), .A2(n18491), .A3(n18488), .A4(n16624), .ZN(
        n16592) );
  NAND3_X1 U19742 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(n16592), .ZN(n16569) );
  NOR2_X1 U19743 ( .A1(n18497), .A2(n16569), .ZN(n16559) );
  AOI21_X1 U19744 ( .B1(n16547), .B2(n16559), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16531) );
  NOR2_X1 U19745 ( .A1(n17476), .A2(n17602), .ZN(n16600) );
  NAND2_X1 U19746 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16600), .ZN(
        n16587) );
  NOR2_X1 U19747 ( .A1(n16527), .A2(n16587), .ZN(n16542) );
  OAI21_X1 U19748 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16542), .A(
        n17443), .ZN(n17480) );
  NOR2_X1 U19749 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17602), .ZN(
        n16640) );
  NAND2_X1 U19750 ( .A1(n16526), .A2(n16640), .ZN(n16577) );
  OAI21_X1 U19751 ( .B1(n16527), .B2(n16577), .A(n9589), .ZN(n16528) );
  XNOR2_X1 U19752 ( .A(n17480), .B(n16528), .ZN(n16529) );
  OAI22_X1 U19753 ( .A1(n16531), .A2(n16530), .B1(n18460), .B2(n16529), .ZN(
        n16532) );
  AOI211_X1 U19754 ( .C1(n16646), .C2(P3_EBX_REG_11__SCAN_IN), .A(n17932), .B(
        n16532), .ZN(n16536) );
  OAI211_X1 U19755 ( .C1(n16538), .C2(n16534), .A(n16654), .B(n16533), .ZN(
        n16535) );
  OAI211_X1 U19756 ( .C1(n16656), .C2(n16537), .A(n16536), .B(n16535), .ZN(
        P3_U2660) );
  AOI211_X1 U19757 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16539), .A(n16538), .B(
        n16665), .ZN(n16540) );
  AOI211_X1 U19758 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n16610), .A(
        n17932), .B(n16540), .ZN(n16551) );
  NAND2_X1 U19759 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16541) );
  INV_X1 U19760 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17526) );
  NOR2_X1 U19761 ( .A1(n17526), .A2(n16587), .ZN(n16575) );
  INV_X1 U19762 ( .A(n16575), .ZN(n16564) );
  NOR2_X1 U19763 ( .A1(n16541), .A2(n16564), .ZN(n16555) );
  INV_X1 U19764 ( .A(n16542), .ZN(n16543) );
  OAI21_X1 U19765 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16555), .A(
        n16543), .ZN(n17489) );
  AOI21_X1 U19766 ( .B1(n16555), .B2(n16658), .A(n16599), .ZN(n16544) );
  XNOR2_X1 U19767 ( .A(n17489), .B(n16544), .ZN(n16549) );
  OAI21_X1 U19768 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16559), .ZN(n16546) );
  NAND2_X1 U19769 ( .A1(n16667), .A2(n16545), .ZN(n16568) );
  OAI22_X1 U19770 ( .A1(n16547), .A2(n16546), .B1(n18500), .B2(n16568), .ZN(
        n16548) );
  AOI21_X1 U19771 ( .B1(n16549), .B2(n16655), .A(n16548), .ZN(n16550) );
  OAI211_X1 U19772 ( .C1(n16666), .C2(n16911), .A(n16551), .B(n16550), .ZN(
        P3_U2661) );
  NOR2_X1 U19773 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16564), .ZN(
        n16563) );
  INV_X1 U19774 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17502) );
  NOR2_X1 U19775 ( .A1(n17502), .A2(n16564), .ZN(n16553) );
  INV_X1 U19776 ( .A(n16555), .ZN(n16552) );
  OAI21_X1 U19777 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16553), .A(
        n16552), .ZN(n17504) );
  AOI22_X1 U19778 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16563), .B1(
        n9589), .B2(n17504), .ZN(n16554) );
  AOI211_X1 U19779 ( .C1(n16555), .C2(n16658), .A(n16554), .B(n18460), .ZN(
        n16558) );
  NOR2_X1 U19780 ( .A1(n16560), .A2(n16665), .ZN(n16567) );
  AOI22_X1 U19781 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16610), .B1(
        n16567), .B2(n16851), .ZN(n16556) );
  OAI211_X1 U19782 ( .C1(n17504), .C2(n16643), .A(n16556), .B(n17930), .ZN(
        n16557) );
  AOI211_X1 U19783 ( .C1(n16559), .C2(n18498), .A(n16558), .B(n16557), .ZN(
        n16562) );
  OAI221_X1 U19784 ( .B1(n16646), .B2(n16654), .C1(n16646), .C2(n16560), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n16561) );
  OAI211_X1 U19785 ( .C1(n16568), .C2(n18498), .A(n16562), .B(n16561), .ZN(
        P3_U2662) );
  NOR2_X1 U19786 ( .A1(n16563), .A2(n16599), .ZN(n16565) );
  AOI22_X1 U19787 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16564), .B1(
        n16575), .B2(n17502), .ZN(n17514) );
  XOR2_X1 U19788 ( .A(n16565), .B(n17514), .Z(n16573) );
  NAND2_X1 U19789 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16579), .ZN(n16566) );
  AOI22_X1 U19790 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16610), .B1(
        n16567), .B2(n16566), .ZN(n16572) );
  AOI21_X1 U19791 ( .B1(n18497), .B2(n16569), .A(n16568), .ZN(n16570) );
  AOI211_X1 U19792 ( .C1(n16646), .C2(P3_EBX_REG_8__SCAN_IN), .A(n17932), .B(
        n16570), .ZN(n16571) );
  OAI211_X1 U19793 ( .C1(n18460), .C2(n16573), .A(n16572), .B(n16571), .ZN(
        P3_U2663) );
  OAI21_X1 U19794 ( .B1(n16659), .B2(n16574), .A(n16669), .ZN(n16601) );
  INV_X1 U19795 ( .A(n16601), .ZN(n16586) );
  INV_X1 U19796 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18494) );
  AOI21_X1 U19797 ( .B1(n17526), .B2(n16587), .A(n16575), .ZN(n16576) );
  INV_X1 U19798 ( .A(n16576), .ZN(n17537) );
  NAND2_X1 U19799 ( .A1(n9589), .A2(n16577), .ZN(n16593) );
  OAI21_X1 U19800 ( .B1(n17537), .B2(n16593), .A(n16655), .ZN(n16578) );
  AOI21_X1 U19801 ( .B1(n17537), .B2(n16593), .A(n16578), .ZN(n16583) );
  OAI211_X1 U19802 ( .C1(n16588), .C2(n16581), .A(n16654), .B(n16579), .ZN(
        n16580) );
  OAI211_X1 U19803 ( .C1(n16666), .C2(n16581), .A(n17930), .B(n16580), .ZN(
        n16582) );
  AOI211_X1 U19804 ( .C1(n16610), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16583), .B(n16582), .ZN(n16585) );
  INV_X1 U19805 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18492) );
  OAI221_X1 U19806 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(P3_REIP_REG_6__SCAN_IN), 
        .C1(n18494), .C2(n18492), .A(n16592), .ZN(n16584) );
  OAI211_X1 U19807 ( .C1(n16586), .C2(n18494), .A(n16585), .B(n16584), .ZN(
        P3_U2664) );
  OAI21_X1 U19808 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16600), .A(
        n16587), .ZN(n17545) );
  OAI21_X1 U19809 ( .B1(n16600), .B2(n16599), .A(n16662), .ZN(n16597) );
  AOI211_X1 U19810 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16603), .A(n16588), .B(
        n16665), .ZN(n16589) );
  AOI211_X1 U19811 ( .C1(n16646), .C2(P3_EBX_REG_6__SCAN_IN), .A(n17932), .B(
        n16589), .ZN(n16590) );
  OAI21_X1 U19812 ( .B1(n20724), .B2(n16656), .A(n16590), .ZN(n16591) );
  AOI221_X1 U19813 ( .B1(n16592), .B2(n18492), .C1(n16601), .C2(
        P3_REIP_REG_6__SCAN_IN), .A(n16591), .ZN(n16596) );
  INV_X1 U19814 ( .A(n16593), .ZN(n16594) );
  NAND3_X1 U19815 ( .A1(n16655), .A2(n16594), .A3(n17545), .ZN(n16595) );
  OAI211_X1 U19816 ( .C1(n17545), .C2(n16597), .A(n16596), .B(n16595), .ZN(
        P3_U2665) );
  AOI21_X1 U19817 ( .B1(n16598), .B2(n16640), .A(n16599), .ZN(n16616) );
  INV_X1 U19818 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17554) );
  NAND2_X1 U19819 ( .A1(n16598), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16615) );
  AOI21_X1 U19820 ( .B1(n17554), .B2(n16615), .A(n16600), .ZN(n17561) );
  XNOR2_X1 U19821 ( .A(n16616), .B(n17561), .ZN(n16608) );
  NOR3_X1 U19822 ( .A1(n16659), .A2(n18488), .A3(n16624), .ZN(n16602) );
  OAI21_X1 U19823 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n16602), .A(n16601), .ZN(
        n16605) );
  OAI211_X1 U19824 ( .C1(n16611), .C2(n16955), .A(n16654), .B(n16603), .ZN(
        n16604) );
  OAI211_X1 U19825 ( .C1(n16656), .C2(n17554), .A(n16605), .B(n16604), .ZN(
        n16606) );
  AOI211_X1 U19826 ( .C1(n16646), .C2(P3_EBX_REG_5__SCAN_IN), .A(n17932), .B(
        n16606), .ZN(n16607) );
  OAI21_X1 U19827 ( .B1(n18460), .B2(n16608), .A(n16607), .ZN(P3_U2666) );
  NOR2_X1 U19828 ( .A1(n16659), .A2(n16624), .ZN(n16609) );
  AOI22_X1 U19829 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16610), .B1(
        n16609), .B2(n18488), .ZN(n16622) );
  AOI211_X1 U19830 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16631), .A(n16611), .B(
        n16665), .ZN(n16620) );
  AOI21_X1 U19831 ( .B1(n16648), .B2(n16624), .A(n16653), .ZN(n16628) );
  NAND2_X1 U19832 ( .A1(n16612), .A2(n18620), .ZN(n16672) );
  INV_X1 U19833 ( .A(n16672), .ZN(n18622) );
  OAI21_X1 U19834 ( .B1(n12110), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18622), .ZN(n16613) );
  OAI211_X1 U19835 ( .C1(n16628), .C2(n18488), .A(n17930), .B(n16613), .ZN(
        n16619) );
  NOR2_X1 U19836 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16614), .ZN(
        n17565) );
  NOR2_X1 U19837 ( .A1(n16614), .A2(n17602), .ZN(n16626) );
  OAI21_X1 U19838 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16626), .A(
        n16615), .ZN(n17571) );
  AOI22_X1 U19839 ( .A1(n16640), .A2(n17565), .B1(n16616), .B2(n17571), .ZN(
        n16617) );
  OAI22_X1 U19840 ( .A1(n16617), .A2(n18460), .B1(n17571), .B2(n16643), .ZN(
        n16618) );
  NOR3_X1 U19841 ( .A1(n16620), .A2(n16619), .A3(n16618), .ZN(n16621) );
  OAI211_X1 U19842 ( .C1(n16666), .C2(n20743), .A(n16622), .B(n16621), .ZN(
        P3_U2667) );
  INV_X1 U19843 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20684) );
  NOR2_X1 U19844 ( .A1(n18586), .A2(n18419), .ZN(n16635) );
  INV_X1 U19845 ( .A(n16635), .ZN(n18405) );
  AOI21_X1 U19846 ( .B1(n18405), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n16922), .ZN(n16623) );
  INV_X1 U19847 ( .A(n16623), .ZN(n18558) );
  NAND2_X1 U19848 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16647) );
  NAND2_X1 U19849 ( .A1(n16648), .A2(n16624), .ZN(n16625) );
  OAI22_X1 U19850 ( .A1(n16666), .A2(n16968), .B1(n16647), .B2(n16625), .ZN(
        n16630) );
  INV_X1 U19851 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18486) );
  NAND2_X1 U19852 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16639) );
  AOI21_X1 U19853 ( .B1(n20684), .B2(n16639), .A(n16626), .ZN(n17578) );
  OAI21_X1 U19854 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16639), .A(
        n9589), .ZN(n16642) );
  XOR2_X1 U19855 ( .A(n17578), .B(n16642), .Z(n16627) );
  OAI22_X1 U19856 ( .A1(n16628), .A2(n18486), .B1(n18460), .B2(n16627), .ZN(
        n16629) );
  AOI211_X1 U19857 ( .C1(n18622), .C2(n18558), .A(n16630), .B(n16629), .ZN(
        n16633) );
  OAI211_X1 U19858 ( .C1(n16638), .C2(n16968), .A(n16654), .B(n16631), .ZN(
        n16632) );
  OAI211_X1 U19859 ( .C1(n16656), .C2(n20684), .A(n16633), .B(n16632), .ZN(
        P3_U2668) );
  INV_X1 U19860 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17595) );
  NOR2_X1 U19861 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16652) );
  INV_X1 U19862 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16634) );
  OAI21_X1 U19863 ( .B1(n16652), .B2(n16634), .A(n16654), .ZN(n16637) );
  AOI21_X1 U19864 ( .B1(n18573), .B2(n18412), .A(n16635), .ZN(n18569) );
  AOI22_X1 U19865 ( .A1(n16653), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18569), 
        .B2(n18622), .ZN(n16636) );
  OAI21_X1 U19866 ( .B1(n16638), .B2(n16637), .A(n16636), .ZN(n16645) );
  OAI21_X1 U19867 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16639), .ZN(n17592) );
  OAI21_X1 U19868 ( .B1(n16640), .B2(n17592), .A(n16655), .ZN(n16641) );
  OAI22_X1 U19869 ( .A1(n17592), .A2(n16643), .B1(n16642), .B2(n16641), .ZN(
        n16644) );
  AOI211_X1 U19870 ( .C1(n16646), .C2(P3_EBX_REG_2__SCAN_IN), .A(n16645), .B(
        n16644), .ZN(n16650) );
  OAI211_X1 U19871 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16648), .B(n16647), .ZN(n16649) );
  OAI211_X1 U19872 ( .C1(n16656), .C2(n17595), .A(n16650), .B(n16649), .ZN(
        P3_U2669) );
  NAND2_X1 U19873 ( .A1(n16651), .A2(n18412), .ZN(n18574) );
  AOI21_X1 U19874 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n16652), .ZN(n16983) );
  AOI22_X1 U19875 ( .A1(n16654), .A2(n16983), .B1(n16653), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n16664) );
  NAND2_X1 U19876 ( .A1(n9589), .A2(n16655), .ZN(n16657) );
  OAI21_X1 U19877 ( .B1(n16658), .B2(n16657), .A(n16656), .ZN(n16661) );
  INV_X1 U19878 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n16985) );
  OAI22_X1 U19879 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16659), .B1(n16666), 
        .B2(n16985), .ZN(n16660) );
  AOI221_X1 U19880 ( .B1(n16662), .B2(n17602), .C1(n16661), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16660), .ZN(n16663) );
  OAI211_X1 U19881 ( .C1(n18574), .C2(n16672), .A(n16664), .B(n16663), .ZN(
        P3_U2670) );
  NAND2_X1 U19882 ( .A1(n16666), .A2(n16665), .ZN(n16668) );
  AOI22_X1 U19883 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16668), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16667), .ZN(n16671) );
  INV_X1 U19884 ( .A(n18618), .ZN(n18560) );
  NAND3_X1 U19885 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18560), .A3(
        n16669), .ZN(n16670) );
  OAI211_X1 U19886 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16672), .A(
        n16671), .B(n16670), .ZN(P3_U2671) );
  AOI22_X1 U19887 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12172), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16676) );
  AOI22_X1 U19888 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16675) );
  AOI22_X1 U19889 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16674) );
  AOI22_X1 U19890 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16673) );
  NAND4_X1 U19891 ( .A1(n16676), .A2(n16675), .A3(n16674), .A4(n16673), .ZN(
        n16682) );
  AOI22_X1 U19892 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16680) );
  AOI22_X1 U19893 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16679) );
  AOI22_X1 U19894 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16678) );
  AOI22_X1 U19895 ( .A1(n12206), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16677) );
  NAND4_X1 U19896 ( .A1(n16680), .A2(n16679), .A3(n16678), .A4(n16677), .ZN(
        n16681) );
  NOR2_X1 U19897 ( .A1(n16682), .A2(n16681), .ZN(n16694) );
  AOI22_X1 U19898 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16693) );
  AOI22_X1 U19899 ( .A1(n16683), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16692) );
  AOI22_X1 U19900 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16684) );
  OAI21_X1 U19901 ( .B1(n12127), .B2(n20774), .A(n16684), .ZN(n16690) );
  AOI22_X1 U19902 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16688) );
  AOI22_X1 U19903 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16687) );
  AOI22_X1 U19904 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16686) );
  AOI22_X1 U19905 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16685) );
  NAND4_X1 U19906 ( .A1(n16688), .A2(n16687), .A3(n16686), .A4(n16685), .ZN(
        n16689) );
  AOI211_X1 U19907 ( .C1(n16945), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n16690), .B(n16689), .ZN(n16691) );
  NAND3_X1 U19908 ( .A1(n16693), .A2(n16692), .A3(n16691), .ZN(n16699) );
  NAND2_X1 U19909 ( .A1(n16700), .A2(n16699), .ZN(n16698) );
  XNOR2_X1 U19910 ( .A(n16694), .B(n16698), .ZN(n16998) );
  NOR2_X1 U19911 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16695), .ZN(n16697) );
  OAI22_X1 U19912 ( .A1(n16998), .A2(n16975), .B1(n16697), .B2(n16696), .ZN(
        P3_U2673) );
  OAI21_X1 U19913 ( .B1(n16700), .B2(n16699), .A(n16698), .ZN(n17006) );
  INV_X1 U19914 ( .A(n16701), .ZN(n16704) );
  OAI21_X1 U19915 ( .B1(n20777), .B2(n16702), .A(n16705), .ZN(n16703) );
  OAI21_X1 U19916 ( .B1(n16705), .B2(n16704), .A(n16703), .ZN(n16706) );
  OAI21_X1 U19917 ( .B1(n16975), .B2(n17006), .A(n16706), .ZN(P3_U2674) );
  OAI21_X1 U19918 ( .B1(n16711), .B2(n16708), .A(n16707), .ZN(n17015) );
  AOI22_X1 U19919 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16713), .B1(n16715), 
        .B2(n16709), .ZN(n16710) );
  OAI21_X1 U19920 ( .B1(n16975), .B2(n17015), .A(n16710), .ZN(P3_U2676) );
  NAND2_X1 U19921 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16723), .ZN(n16719) );
  AOI21_X1 U19922 ( .B1(n16712), .B2(n16716), .A(n16711), .ZN(n17016) );
  AOI22_X1 U19923 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16713), .B1(n17016), 
        .B2(n16987), .ZN(n16714) );
  OAI21_X1 U19924 ( .B1(n16715), .B2(n16719), .A(n16714), .ZN(P3_U2677) );
  OAI21_X1 U19925 ( .B1(n16718), .B2(n16717), .A(n16716), .ZN(n17024) );
  OAI211_X1 U19926 ( .C1(n16723), .C2(P3_EBX_REG_25__SCAN_IN), .A(n16972), .B(
        n16719), .ZN(n16720) );
  OAI21_X1 U19927 ( .B1(n17024), .B2(n16972), .A(n16720), .ZN(P3_U2678) );
  AOI21_X1 U19928 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16975), .A(n16728), .ZN(
        n16722) );
  XNOR2_X1 U19929 ( .A(n16721), .B(n16724), .ZN(n17029) );
  OAI22_X1 U19930 ( .A1(n16723), .A2(n16722), .B1(n17029), .B2(n16975), .ZN(
        P3_U2679) );
  AOI21_X1 U19931 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16975), .A(n16743), .ZN(
        n16727) );
  OAI21_X1 U19932 ( .B1(n16726), .B2(n16725), .A(n16724), .ZN(n17035) );
  OAI22_X1 U19933 ( .A1(n16728), .A2(n16727), .B1(n17035), .B2(n16975), .ZN(
        P3_U2680) );
  OAI21_X1 U19934 ( .B1(n16730), .B2(n16987), .A(n16729), .ZN(n16731) );
  INV_X1 U19935 ( .A(n16731), .ZN(n16742) );
  AOI22_X1 U19936 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16735) );
  AOI22_X1 U19937 ( .A1(n12206), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16734) );
  AOI22_X1 U19938 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16733) );
  AOI22_X1 U19939 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16732) );
  NAND4_X1 U19940 ( .A1(n16735), .A2(n16734), .A3(n16733), .A4(n16732), .ZN(
        n16741) );
  AOI22_X1 U19941 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9601), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16739) );
  AOI22_X1 U19942 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16738) );
  AOI22_X1 U19943 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16737) );
  AOI22_X1 U19944 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16736) );
  NAND4_X1 U19945 ( .A1(n16739), .A2(n16738), .A3(n16737), .A4(n16736), .ZN(
        n16740) );
  NOR2_X1 U19946 ( .A1(n16741), .A2(n16740), .ZN(n17039) );
  OAI22_X1 U19947 ( .A1(n16743), .A2(n16742), .B1(n17039), .B2(n16975), .ZN(
        P3_U2681) );
  AOI22_X1 U19948 ( .A1(n12163), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16747) );
  AOI22_X1 U19949 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16746) );
  AOI22_X1 U19950 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16745) );
  AOI22_X1 U19951 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16744) );
  NAND4_X1 U19952 ( .A1(n16747), .A2(n16746), .A3(n16745), .A4(n16744), .ZN(
        n16753) );
  AOI22_X1 U19953 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16751) );
  AOI22_X1 U19954 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16750) );
  AOI22_X1 U19955 ( .A1(n12206), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16749) );
  AOI22_X1 U19956 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16748) );
  NAND4_X1 U19957 ( .A1(n16751), .A2(n16750), .A3(n16749), .A4(n16748), .ZN(
        n16752) );
  NOR2_X1 U19958 ( .A1(n16753), .A2(n16752), .ZN(n17046) );
  AOI21_X1 U19959 ( .B1(n16783), .B2(P3_EBX_REG_20__SCAN_IN), .A(n16987), .ZN(
        n16767) );
  AOI22_X1 U19960 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16767), .B1(n16754), 
        .B2(n20744), .ZN(n16755) );
  OAI21_X1 U19961 ( .B1(n17046), .B2(n16972), .A(n16755), .ZN(P3_U2682) );
  AOI22_X1 U19962 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16759) );
  AOI22_X1 U19963 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16758) );
  AOI22_X1 U19964 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12172), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16757) );
  AOI22_X1 U19965 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16756) );
  NAND4_X1 U19966 ( .A1(n16759), .A2(n16758), .A3(n16757), .A4(n16756), .ZN(
        n16765) );
  AOI22_X1 U19967 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12163), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16763) );
  AOI22_X1 U19968 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16762) );
  AOI22_X1 U19969 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12177), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16761) );
  AOI22_X1 U19970 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16760) );
  NAND4_X1 U19971 ( .A1(n16763), .A2(n16762), .A3(n16761), .A4(n16760), .ZN(
        n16764) );
  NOR2_X1 U19972 ( .A1(n16765), .A2(n16764), .ZN(n17051) );
  INV_X1 U19973 ( .A(n16766), .ZN(n16768) );
  OAI21_X1 U19974 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16768), .A(n16767), .ZN(
        n16769) );
  OAI21_X1 U19975 ( .B1(n17051), .B2(n16972), .A(n16769), .ZN(P3_U2683) );
  AOI21_X1 U19976 ( .B1(n16770), .B2(n16794), .A(n16987), .ZN(n16771) );
  INV_X1 U19977 ( .A(n16771), .ZN(n16782) );
  AOI22_X1 U19978 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16775) );
  AOI22_X1 U19979 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U19980 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16773) );
  AOI22_X1 U19981 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16772) );
  NAND4_X1 U19982 ( .A1(n16775), .A2(n16774), .A3(n16773), .A4(n16772), .ZN(
        n16781) );
  AOI22_X1 U19983 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16779) );
  AOI22_X1 U19984 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16778) );
  AOI22_X1 U19985 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16777) );
  AOI22_X1 U19986 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16776) );
  NAND4_X1 U19987 ( .A1(n16779), .A2(n16778), .A3(n16777), .A4(n16776), .ZN(
        n16780) );
  NOR2_X1 U19988 ( .A1(n16781), .A2(n16780), .ZN(n17055) );
  OAI22_X1 U19989 ( .A1(n16783), .A2(n16782), .B1(n17055), .B2(n16975), .ZN(
        P3_U2684) );
  AOI22_X1 U19990 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16787) );
  AOI22_X1 U19991 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16786) );
  AOI22_X1 U19992 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16785) );
  AOI22_X1 U19993 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16784) );
  NAND4_X1 U19994 ( .A1(n16787), .A2(n16786), .A3(n16785), .A4(n16784), .ZN(
        n16793) );
  AOI22_X1 U19995 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9601), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16791) );
  AOI22_X1 U19996 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16790) );
  AOI22_X1 U19997 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16789) );
  AOI22_X1 U19998 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16788) );
  NAND4_X1 U19999 ( .A1(n16791), .A2(n16790), .A3(n16789), .A4(n16788), .ZN(
        n16792) );
  NOR2_X1 U20000 ( .A1(n16793), .A2(n16792), .ZN(n17060) );
  NAND2_X1 U20001 ( .A1(n17989), .A2(n16811), .ZN(n16824) );
  NOR3_X1 U20002 ( .A1(n16797), .A2(n16796), .A3(n16824), .ZN(n16810) );
  OAI21_X1 U20003 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16810), .A(n16794), .ZN(
        n16795) );
  AOI22_X1 U20004 ( .A1(n16987), .A2(n17060), .B1(n16795), .B2(n16975), .ZN(
        P3_U2685) );
  OAI22_X1 U20005 ( .A1(n16797), .A2(n16987), .B1(n16796), .B2(n16824), .ZN(
        n16798) );
  INV_X1 U20006 ( .A(n16798), .ZN(n16809) );
  AOI22_X1 U20007 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16915), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16802) );
  AOI22_X1 U20008 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n16916), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U20009 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9601), .ZN(n16800) );
  AOI22_X1 U20010 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n16936), .ZN(n16799) );
  NAND4_X1 U20011 ( .A1(n16802), .A2(n16801), .A3(n16800), .A4(n16799), .ZN(
        n16808) );
  AOI22_X1 U20012 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n16934), .ZN(n16806) );
  AOI22_X1 U20013 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n16922), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n16933), .ZN(n16805) );
  AOI22_X1 U20014 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16804) );
  AOI22_X1 U20015 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9585), .ZN(n16803) );
  NAND4_X1 U20016 ( .A1(n16806), .A2(n16805), .A3(n16804), .A4(n16803), .ZN(
        n16807) );
  NOR2_X1 U20017 ( .A1(n16808), .A2(n16807), .ZN(n17066) );
  OAI22_X1 U20018 ( .A1(n16810), .A2(n16809), .B1(n17066), .B2(n16975), .ZN(
        P3_U2686) );
  NOR2_X1 U20019 ( .A1(n16811), .A2(n16987), .ZN(n16836) );
  AOI22_X1 U20020 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16822) );
  AOI22_X1 U20021 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16821) );
  AOI22_X1 U20022 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16812) );
  OAI21_X1 U20023 ( .B1(n15453), .B2(n16813), .A(n16812), .ZN(n16819) );
  AOI22_X1 U20024 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16817) );
  AOI22_X1 U20025 ( .A1(n16933), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16816) );
  AOI22_X1 U20026 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16815) );
  AOI22_X1 U20027 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16814) );
  NAND4_X1 U20028 ( .A1(n16817), .A2(n16816), .A3(n16815), .A4(n16814), .ZN(
        n16818) );
  AOI211_X1 U20029 ( .C1(n16945), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n16819), .B(n16818), .ZN(n16820) );
  NAND3_X1 U20030 ( .A1(n16822), .A2(n16821), .A3(n16820), .ZN(n17067) );
  AOI22_X1 U20031 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16836), .B1(n16987), 
        .B2(n17067), .ZN(n16823) );
  OAI21_X1 U20032 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n16824), .A(n16823), .ZN(
        P3_U2687) );
  AOI22_X1 U20033 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U20034 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16827) );
  AOI22_X1 U20035 ( .A1(n12163), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16922), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16826) );
  AOI22_X1 U20036 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16825) );
  NAND4_X1 U20037 ( .A1(n16828), .A2(n16827), .A3(n16826), .A4(n16825), .ZN(
        n16834) );
  AOI22_X1 U20038 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16832) );
  AOI22_X1 U20039 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16831) );
  AOI22_X1 U20040 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16830) );
  AOI22_X1 U20041 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16829) );
  NAND4_X1 U20042 ( .A1(n16832), .A2(n16831), .A3(n16830), .A4(n16829), .ZN(
        n16833) );
  NOR2_X1 U20043 ( .A1(n16834), .A2(n16833), .ZN(n17076) );
  INV_X1 U20044 ( .A(n16835), .ZN(n16837) );
  OAI21_X1 U20045 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16837), .A(n16836), .ZN(
        n16838) );
  OAI21_X1 U20046 ( .B1(n17076), .B2(n16972), .A(n16838), .ZN(P3_U2688) );
  AOI22_X1 U20047 ( .A1(n12206), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16849) );
  AOI22_X1 U20048 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U20049 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16839) );
  OAI21_X1 U20050 ( .B1(n16840), .B2(n20774), .A(n16839), .ZN(n16846) );
  AOI22_X1 U20051 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16844) );
  AOI22_X1 U20052 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16843) );
  AOI22_X1 U20053 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16922), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16842) );
  AOI22_X1 U20054 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16841) );
  NAND4_X1 U20055 ( .A1(n16844), .A2(n16843), .A3(n16842), .A4(n16841), .ZN(
        n16845) );
  AOI211_X1 U20056 ( .C1(n16916), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16846), .B(n16845), .ZN(n16847) );
  NAND3_X1 U20057 ( .A1(n16849), .A2(n16848), .A3(n16847), .ZN(n17078) );
  INV_X1 U20058 ( .A(n17078), .ZN(n16857) );
  NOR2_X1 U20059 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16973), .ZN(n16869) );
  NAND2_X1 U20060 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .ZN(n16850) );
  NOR4_X1 U20061 ( .A1(n16851), .A2(n16931), .A3(n16955), .A4(n16850), .ZN(
        n16852) );
  NAND4_X1 U20062 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n16954), .A4(n16852), .ZN(n16853) );
  NOR2_X1 U20063 ( .A1(n16885), .A2(n16853), .ZN(n16868) );
  OAI21_X1 U20064 ( .B1(n16868), .B2(n17077), .A(n9588), .ZN(n16870) );
  OAI21_X1 U20065 ( .B1(n16869), .B2(n16870), .A(P3_EBX_REG_14__SCAN_IN), .ZN(
        n16856) );
  NOR2_X1 U20066 ( .A1(n16973), .A2(n16853), .ZN(n16886) );
  INV_X1 U20067 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16854) );
  NAND4_X1 U20068 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n16886), .A4(n16854), .ZN(n16855) );
  OAI211_X1 U20069 ( .C1(n16857), .C2(n16975), .A(n16856), .B(n16855), .ZN(
        P3_U2689) );
  AOI22_X1 U20070 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16922), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20071 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16860) );
  AOI22_X1 U20072 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20073 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16858) );
  NAND4_X1 U20074 ( .A1(n16861), .A2(n16860), .A3(n16859), .A4(n16858), .ZN(
        n16867) );
  AOI22_X1 U20075 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16865) );
  AOI22_X1 U20076 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16864) );
  AOI22_X1 U20077 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16863) );
  AOI22_X1 U20078 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16862) );
  NAND4_X1 U20079 ( .A1(n16865), .A2(n16864), .A3(n16863), .A4(n16862), .ZN(
        n16866) );
  NOR2_X1 U20080 ( .A1(n16867), .A2(n16866), .ZN(n17084) );
  AOI22_X1 U20081 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16870), .B1(n16869), 
        .B2(n16868), .ZN(n16871) );
  OAI21_X1 U20082 ( .B1(n17084), .B2(n16972), .A(n16871), .ZN(P3_U2690) );
  AOI22_X1 U20083 ( .A1(n9586), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16876) );
  AOI22_X1 U20084 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U20085 ( .A1(n12206), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U20086 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16873) );
  NAND4_X1 U20087 ( .A1(n16876), .A2(n16875), .A3(n16874), .A4(n16873), .ZN(
        n16883) );
  AOI22_X1 U20088 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16881) );
  AOI22_X1 U20089 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20090 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16922), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20091 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16877), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16878) );
  NAND4_X1 U20092 ( .A1(n16881), .A2(n16880), .A3(n16879), .A4(n16878), .ZN(
        n16882) );
  NOR2_X1 U20093 ( .A1(n16883), .A2(n16882), .ZN(n17088) );
  NOR2_X1 U20094 ( .A1(n16884), .A2(n16987), .ZN(n16898) );
  AOI22_X1 U20095 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16898), .B1(n16886), 
        .B2(n16885), .ZN(n16887) );
  OAI21_X1 U20096 ( .B1(n17088), .B2(n16972), .A(n16887), .ZN(P3_U2691) );
  AOI22_X1 U20097 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20098 ( .A1(n16917), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16890) );
  AOI22_X1 U20099 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16922), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20100 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16888) );
  NAND4_X1 U20101 ( .A1(n16891), .A2(n16890), .A3(n16889), .A4(n16888), .ZN(
        n16897) );
  AOI22_X1 U20102 ( .A1(n12206), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16895) );
  AOI22_X1 U20103 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12172), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16894) );
  AOI22_X1 U20104 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20105 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16892) );
  NAND4_X1 U20106 ( .A1(n16895), .A2(n16894), .A3(n16893), .A4(n16892), .ZN(
        n16896) );
  NOR2_X1 U20107 ( .A1(n16897), .A2(n16896), .ZN(n17091) );
  NOR2_X1 U20108 ( .A1(n16911), .A2(n16929), .ZN(n16914) );
  OAI21_X1 U20109 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16914), .A(n16898), .ZN(
        n16899) );
  OAI21_X1 U20110 ( .B1(n17091), .B2(n16972), .A(n16899), .ZN(P3_U2692) );
  AOI22_X1 U20111 ( .A1(n16900), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16922), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20112 ( .A1(n16941), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20113 ( .A1(n16916), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20114 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16936), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16901) );
  NAND4_X1 U20115 ( .A1(n16904), .A2(n16903), .A3(n16902), .A4(n16901), .ZN(
        n16910) );
  AOI22_X1 U20116 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16917), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16908) );
  AOI22_X1 U20117 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U20118 ( .A1(n9601), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16934), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16906) );
  AOI22_X1 U20119 ( .A1(n9595), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16905) );
  NAND4_X1 U20120 ( .A1(n16908), .A2(n16907), .A3(n16906), .A4(n16905), .ZN(
        n16909) );
  NOR2_X1 U20121 ( .A1(n16910), .A2(n16909), .ZN(n17098) );
  AOI21_X1 U20122 ( .B1(n16911), .B2(n16929), .A(n16987), .ZN(n16912) );
  INV_X1 U20123 ( .A(n16912), .ZN(n16913) );
  OAI22_X1 U20124 ( .A1(n17098), .A2(n16975), .B1(n16914), .B2(n16913), .ZN(
        P3_U2693) );
  AOI22_X1 U20125 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9602), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n16915), .ZN(n16921) );
  AOI22_X1 U20126 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9586), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20127 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U20128 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16936), .B1(
        n16917), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16918) );
  NAND4_X1 U20129 ( .A1(n16921), .A2(n16920), .A3(n16919), .A4(n16918), .ZN(
        n16928) );
  AOI22_X1 U20130 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12172), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16926) );
  AOI22_X1 U20131 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n16941), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n16922), .ZN(n16925) );
  AOI22_X1 U20132 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16934), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n16933), .ZN(n16924) );
  AOI22_X1 U20133 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9601), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16923) );
  NAND4_X1 U20134 ( .A1(n16926), .A2(n16925), .A3(n16924), .A4(n16923), .ZN(
        n16927) );
  NOR2_X1 U20135 ( .A1(n16928), .A2(n16927), .ZN(n17100) );
  OAI21_X1 U20136 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16953), .A(n16929), .ZN(
        n16930) );
  AOI22_X1 U20137 ( .A1(n16987), .A2(n17100), .B1(n16930), .B2(n16975), .ZN(
        P3_U2694) );
  AOI21_X1 U20138 ( .B1(n16931), .B2(n16956), .A(n16987), .ZN(n16932) );
  INV_X1 U20139 ( .A(n16932), .ZN(n16952) );
  AOI22_X1 U20140 ( .A1(n12172), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9601), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20141 ( .A1(n16934), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16933), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20142 ( .A1(n9602), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9585), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16938) );
  AOI22_X1 U20143 ( .A1(n16936), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16935), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16937) );
  NAND4_X1 U20144 ( .A1(n16940), .A2(n16939), .A3(n16938), .A4(n16937), .ZN(
        n16951) );
  AOI22_X1 U20145 ( .A1(n9594), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16941), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20146 ( .A1(n16942), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16915), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20147 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20148 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9595), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16946) );
  NAND4_X1 U20149 ( .A1(n16949), .A2(n16948), .A3(n16947), .A4(n16946), .ZN(
        n16950) );
  NOR2_X1 U20150 ( .A1(n16951), .A2(n16950), .ZN(n17106) );
  OAI22_X1 U20151 ( .A1(n16953), .A2(n16952), .B1(n17106), .B2(n16975), .ZN(
        P3_U2695) );
  NAND2_X1 U20152 ( .A1(n16954), .A2(n16986), .ZN(n16969) );
  NOR2_X1 U20153 ( .A1(n16955), .A2(n16969), .ZN(n16961) );
  OAI221_X1 U20154 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(P3_EBX_REG_6__SCAN_IN), 
        .C1(P3_EBX_REG_7__SCAN_IN), .C2(n16961), .A(n16956), .ZN(n16957) );
  AOI22_X1 U20155 ( .A1(n16987), .A2(n16958), .B1(n16957), .B2(n16975), .ZN(
        P3_U2696) );
  INV_X1 U20156 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16963) );
  NOR2_X1 U20157 ( .A1(n16959), .A2(n16987), .ZN(n16965) );
  INV_X1 U20158 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20159 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16965), .B1(n16961), .B2(
        n16960), .ZN(n16962) );
  OAI21_X1 U20160 ( .B1(n16963), .B2(n16972), .A(n16962), .ZN(P3_U2697) );
  INV_X1 U20161 ( .A(n16964), .ZN(n16966) );
  OAI21_X1 U20162 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n16966), .A(n16965), .ZN(
        n16967) );
  OAI21_X1 U20163 ( .B1(n16972), .B2(n20785), .A(n16967), .ZN(P3_U2698) );
  NOR3_X1 U20164 ( .A1(n16968), .A2(n16974), .A3(n16973), .ZN(n16978) );
  OAI211_X1 U20165 ( .C1(n16978), .C2(P3_EBX_REG_4__SCAN_IN), .A(n16972), .B(
        n16969), .ZN(n16970) );
  OAI21_X1 U20166 ( .B1(n16972), .B2(n16971), .A(n16970), .ZN(P3_U2699) );
  NOR2_X1 U20167 ( .A1(n16974), .A2(n16973), .ZN(n16980) );
  AOI21_X1 U20168 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n16975), .A(n16980), .ZN(
        n16977) );
  INV_X1 U20169 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16976) );
  OAI22_X1 U20170 ( .A1(n16978), .A2(n16977), .B1(n16976), .B2(n16975), .ZN(
        P3_U2700) );
  INV_X1 U20171 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n16989) );
  NOR2_X1 U20172 ( .A1(n16989), .A2(n16985), .ZN(n16979) );
  AOI221_X1 U20173 ( .B1(n16979), .B2(n9588), .C1(n17077), .C2(n9588), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n16981) );
  AOI211_X1 U20174 ( .C1(n16987), .C2(n16982), .A(n16981), .B(n16980), .ZN(
        P3_U2701) );
  AOI22_X1 U20175 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16987), .B1(
        n16986), .B2(n16983), .ZN(n16984) );
  OAI21_X1 U20176 ( .B1(n9588), .B2(n16985), .A(n16984), .ZN(P3_U2702) );
  AOI22_X1 U20177 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16987), .B1(
        n16986), .B2(n16989), .ZN(n16988) );
  OAI21_X1 U20178 ( .B1(n9588), .B2(n16989), .A(n16988), .ZN(P3_U2703) );
  NOR2_X2 U20179 ( .A1(n17128), .A2(n17983), .ZN(n17068) );
  INV_X1 U20180 ( .A(n17068), .ZN(n17037) );
  INV_X1 U20181 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17150) );
  INV_X1 U20182 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17154) );
  INV_X1 U20183 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17156) );
  INV_X1 U20184 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17158) );
  INV_X1 U20185 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17256) );
  INV_X1 U20186 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17198) );
  INV_X1 U20187 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17200) );
  NAND2_X1 U20188 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17137) );
  NAND2_X1 U20189 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n17107) );
  NOR4_X1 U20190 ( .A1(n17198), .A2(n17200), .A3(n17137), .A4(n17107), .ZN(
        n16991) );
  NAND4_X1 U20191 ( .A1(n16992), .A2(P3_EAX_REG_7__SCAN_IN), .A3(
        P3_EAX_REG_6__SCAN_IN), .A4(n16991), .ZN(n17103) );
  NAND4_X1 U20192 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n16993)
         );
  NOR2_X1 U20193 ( .A1(n17103), .A2(n16993), .ZN(n16994) );
  NAND4_X1 U20194 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n16994), .ZN(n17080) );
  NAND3_X1 U20195 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .ZN(n17036) );
  NAND2_X1 U20196 ( .A1(n17989), .A2(n17030), .ZN(n17025) );
  NAND2_X1 U20197 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17011), .ZN(n17008) );
  NOR2_X1 U20198 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17002), .ZN(n16995) );
  OAI21_X1 U20199 ( .B1(n16997), .B2(n17037), .A(n16996), .ZN(P3_U2704) );
  INV_X1 U20200 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17225) );
  NAND2_X1 U20201 ( .A1(n17977), .A2(n17095), .ZN(n17072) );
  INV_X1 U20202 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n17981) );
  OAI22_X1 U20203 ( .A1(n16998), .A2(n17131), .B1(n17981), .B2(n17037), .ZN(
        n16999) );
  AOI21_X1 U20204 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17061), .A(n16999), .ZN(
        n17000) );
  OAI221_X1 U20205 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17002), .C1(n17225), 
        .C2(n17001), .A(n17000), .ZN(P3_U2705) );
  AOI22_X1 U20206 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17068), .ZN(n17005) );
  OAI211_X1 U20207 ( .C1(n17003), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17128), .B(
        n17002), .ZN(n17004) );
  OAI211_X1 U20208 ( .C1(n17006), .C2(n17131), .A(n17005), .B(n17004), .ZN(
        P3_U2706) );
  INV_X1 U20209 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17244) );
  AOI22_X1 U20210 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17068), .B1(n17079), .B2(
        n17007), .ZN(n17010) );
  OAI211_X1 U20211 ( .C1(n17011), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17128), .B(
        n17008), .ZN(n17009) );
  OAI211_X1 U20212 ( .C1(n17072), .C2(n17244), .A(n17010), .B(n17009), .ZN(
        P3_U2707) );
  AOI22_X1 U20213 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17068), .ZN(n17014) );
  AOI211_X1 U20214 ( .C1(n17150), .C2(n17017), .A(n17011), .B(n17095), .ZN(
        n17012) );
  INV_X1 U20215 ( .A(n17012), .ZN(n17013) );
  OAI211_X1 U20216 ( .C1(n17015), .C2(n17131), .A(n17014), .B(n17013), .ZN(
        P3_U2708) );
  INV_X1 U20217 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U20218 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17068), .B1(n17079), .B2(
        n17016), .ZN(n17019) );
  OAI211_X1 U20219 ( .C1(n17020), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17128), .B(
        n17017), .ZN(n17018) );
  OAI211_X1 U20220 ( .C1(n17072), .C2(n17240), .A(n17019), .B(n17018), .ZN(
        P3_U2709) );
  AOI22_X1 U20221 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17068), .ZN(n17023) );
  AOI211_X1 U20222 ( .C1(n17154), .C2(n9673), .A(n17020), .B(n17095), .ZN(
        n17021) );
  INV_X1 U20223 ( .A(n17021), .ZN(n17022) );
  OAI211_X1 U20224 ( .C1(n17024), .C2(n17131), .A(n17023), .B(n17022), .ZN(
        P3_U2710) );
  AOI22_X1 U20225 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17068), .ZN(n17028) );
  OAI21_X1 U20226 ( .B1(n17156), .B2(n17095), .A(n17025), .ZN(n17026) );
  NAND2_X1 U20227 ( .A1(n17026), .A2(n9673), .ZN(n17027) );
  OAI211_X1 U20228 ( .C1(n17029), .C2(n17131), .A(n17028), .B(n17027), .ZN(
        P3_U2711) );
  AOI211_X1 U20229 ( .C1(n17158), .C2(n17031), .A(n17095), .B(n17030), .ZN(
        n17032) );
  AOI21_X1 U20230 ( .B1(n17068), .B2(BUF2_REG_23__SCAN_IN), .A(n17032), .ZN(
        n17034) );
  NAND2_X1 U20231 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17061), .ZN(n17033) );
  OAI211_X1 U20232 ( .C1(n17035), .C2(n17131), .A(n17034), .B(n17033), .ZN(
        P3_U2712) );
  NOR2_X1 U20233 ( .A1(n17077), .A2(n17069), .ZN(n17063) );
  NAND2_X1 U20234 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17063), .ZN(n17062) );
  NOR2_X1 U20235 ( .A1(n17036), .A2(n17062), .ZN(n17047) );
  NAND2_X1 U20236 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17047), .ZN(n17043) );
  NAND2_X1 U20237 ( .A1(n17043), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17042) );
  OAI22_X1 U20238 ( .A1(n17039), .A2(n17131), .B1(n17038), .B2(n17037), .ZN(
        n17040) );
  AOI21_X1 U20239 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17061), .A(n17040), .ZN(
        n17041) );
  OAI221_X1 U20240 ( .B1(n17043), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17042), 
        .C2(n17095), .A(n17041), .ZN(P3_U2713) );
  AOI22_X1 U20241 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17068), .ZN(n17045) );
  OAI211_X1 U20242 ( .C1(n17047), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17128), .B(
        n17043), .ZN(n17044) );
  OAI211_X1 U20243 ( .C1(n17046), .C2(n17131), .A(n17045), .B(n17044), .ZN(
        P3_U2714) );
  AOI22_X1 U20244 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17068), .ZN(n17050) );
  INV_X1 U20245 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17164) );
  INV_X1 U20246 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17168) );
  NOR2_X1 U20247 ( .A1(n17168), .A2(n17062), .ZN(n17056) );
  NAND2_X1 U20248 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17056), .ZN(n17052) );
  AOI211_X1 U20249 ( .C1(n17164), .C2(n17052), .A(n17047), .B(n17095), .ZN(
        n17048) );
  INV_X1 U20250 ( .A(n17048), .ZN(n17049) );
  OAI211_X1 U20251 ( .C1(n17051), .C2(n17131), .A(n17050), .B(n17049), .ZN(
        P3_U2715) );
  AOI22_X1 U20252 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17068), .ZN(n17054) );
  OAI211_X1 U20253 ( .C1(n17056), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17128), .B(
        n17052), .ZN(n17053) );
  OAI211_X1 U20254 ( .C1(n17055), .C2(n17131), .A(n17054), .B(n17053), .ZN(
        P3_U2716) );
  AOI22_X1 U20255 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17068), .ZN(n17059) );
  AOI211_X1 U20256 ( .C1(n17168), .C2(n17062), .A(n17056), .B(n17095), .ZN(
        n17057) );
  INV_X1 U20257 ( .A(n17057), .ZN(n17058) );
  OAI211_X1 U20258 ( .C1(n17060), .C2(n17131), .A(n17059), .B(n17058), .ZN(
        P3_U2717) );
  AOI22_X1 U20259 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17061), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17068), .ZN(n17065) );
  OAI211_X1 U20260 ( .C1(n17063), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17128), .B(
        n17062), .ZN(n17064) );
  OAI211_X1 U20261 ( .C1(n17066), .C2(n17131), .A(n17065), .B(n17064), .ZN(
        P3_U2718) );
  INV_X1 U20262 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n17950) );
  AOI22_X1 U20263 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17068), .B1(n17079), .B2(
        n17067), .ZN(n17071) );
  OAI211_X1 U20264 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17073), .A(n17128), .B(
        n17069), .ZN(n17070) );
  OAI211_X1 U20265 ( .C1(n17072), .C2(n17950), .A(n17071), .B(n17070), .ZN(
        P3_U2719) );
  AOI211_X1 U20266 ( .C1(n17256), .C2(n17080), .A(n17095), .B(n17073), .ZN(
        n17074) );
  AOI21_X1 U20267 ( .B1(n17136), .B2(BUF2_REG_15__SCAN_IN), .A(n17074), .ZN(
        n17075) );
  OAI21_X1 U20268 ( .B1(n17076), .B2(n17131), .A(n17075), .ZN(P3_U2720) );
  INV_X1 U20269 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17179) );
  INV_X1 U20270 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17183) );
  NOR2_X1 U20271 ( .A1(n17077), .A2(n17103), .ZN(n17110) );
  NAND3_X1 U20272 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17110), .ZN(n17099) );
  NAND2_X1 U20273 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17094), .ZN(n17087) );
  NOR2_X1 U20274 ( .A1(n17179), .A2(n17087), .ZN(n17090) );
  NAND2_X1 U20275 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17090), .ZN(n17083) );
  AOI22_X1 U20276 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17136), .B1(n17079), .B2(
        n17078), .ZN(n17082) );
  NAND3_X1 U20277 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17128), .A3(n17080), 
        .ZN(n17081) );
  OAI211_X1 U20278 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17083), .A(n17082), .B(
        n17081), .ZN(P3_U2721) );
  INV_X1 U20279 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17249) );
  INV_X1 U20280 ( .A(n17083), .ZN(n17086) );
  AOI21_X1 U20281 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17128), .A(n17090), .ZN(
        n17085) );
  OAI222_X1 U20282 ( .A1(n17134), .A2(n17249), .B1(n17086), .B2(n17085), .C1(
        n17131), .C2(n17084), .ZN(P3_U2722) );
  INV_X1 U20283 ( .A(n17087), .ZN(n17093) );
  AOI21_X1 U20284 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17128), .A(n17093), .ZN(
        n17089) );
  OAI222_X1 U20285 ( .A1(n17134), .A2(n17244), .B1(n17090), .B2(n17089), .C1(
        n17131), .C2(n17088), .ZN(P3_U2723) );
  AOI21_X1 U20286 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17128), .A(n17094), .ZN(
        n17092) );
  OAI222_X1 U20287 ( .A1(n17134), .A2(n17242), .B1(n17093), .B2(n17092), .C1(
        n17131), .C2(n17091), .ZN(P3_U2724) );
  AOI211_X1 U20288 ( .C1(n17183), .C2(n17099), .A(n17095), .B(n17094), .ZN(
        n17096) );
  AOI21_X1 U20289 ( .B1(n17136), .B2(BUF2_REG_10__SCAN_IN), .A(n17096), .ZN(
        n17097) );
  OAI21_X1 U20290 ( .B1(n17098), .B2(n17131), .A(n17097), .ZN(P3_U2725) );
  INV_X1 U20291 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17238) );
  INV_X1 U20292 ( .A(n17099), .ZN(n17102) );
  AOI22_X1 U20293 ( .A1(n17110), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17128), .ZN(n17101) );
  OAI222_X1 U20294 ( .A1(n17134), .A2(n17238), .B1(n17102), .B2(n17101), .C1(
        n17131), .C2(n17100), .ZN(P3_U2726) );
  INV_X1 U20295 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20296 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17136), .B1(n17110), .B2(
        n17187), .ZN(n17105) );
  NAND3_X1 U20297 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17128), .A3(n17103), .ZN(
        n17104) );
  OAI211_X1 U20298 ( .C1(n17106), .C2(n17131), .A(n17105), .B(n17104), .ZN(
        P3_U2727) );
  NAND2_X1 U20299 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17133), .ZN(n17118) );
  NOR2_X1 U20300 ( .A1(n17107), .A2(n17118), .ZN(n17117) );
  AOI22_X1 U20301 ( .A1(n17117), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17128), .ZN(n17109) );
  OAI222_X1 U20302 ( .A1(n17134), .A2(n17986), .B1(n17110), .B2(n17109), .C1(
        n17131), .C2(n17108), .ZN(P3_U2728) );
  INV_X1 U20303 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n17982) );
  AND2_X1 U20304 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17117), .ZN(n17114) );
  AOI21_X1 U20305 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17128), .A(n17117), .ZN(
        n17113) );
  INV_X1 U20306 ( .A(n17111), .ZN(n17112) );
  OAI222_X1 U20307 ( .A1(n17982), .A2(n17134), .B1(n17114), .B2(n17113), .C1(
        n17131), .C2(n17112), .ZN(P3_U2729) );
  INV_X1 U20308 ( .A(n17118), .ZN(n17125) );
  AOI22_X1 U20309 ( .A1(n17125), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17128), .ZN(n17116) );
  OAI222_X1 U20310 ( .A1(n17976), .A2(n17134), .B1(n17117), .B2(n17116), .C1(
        n17131), .C2(n17115), .ZN(P3_U2730) );
  INV_X1 U20311 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n17972) );
  INV_X1 U20312 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17196) );
  NOR2_X1 U20313 ( .A1(n17196), .A2(n17118), .ZN(n17122) );
  AOI21_X1 U20314 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17128), .A(n17125), .ZN(
        n17121) );
  INV_X1 U20315 ( .A(n17119), .ZN(n17120) );
  OAI222_X1 U20316 ( .A1(n17972), .A2(n17134), .B1(n17122), .B2(n17121), .C1(
        n17131), .C2(n17120), .ZN(P3_U2731) );
  AOI21_X1 U20317 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17128), .A(n17133), .ZN(
        n17124) );
  OAI222_X1 U20318 ( .A1(n17968), .A2(n17134), .B1(n17125), .B2(n17124), .C1(
        n17131), .C2(n17123), .ZN(P3_U2732) );
  INV_X1 U20319 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n17964) );
  NOR2_X1 U20320 ( .A1(n17137), .A2(n17126), .ZN(n17127) );
  AOI21_X1 U20321 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17128), .A(n17127), .ZN(
        n17132) );
  INV_X1 U20322 ( .A(n17129), .ZN(n17130) );
  OAI222_X1 U20323 ( .A1(n17964), .A2(n17134), .B1(n17133), .B2(n17132), .C1(
        n17131), .C2(n17130), .ZN(P3_U2733) );
  AOI22_X1 U20324 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17136), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n17135), .ZN(n17140) );
  OAI211_X1 U20325 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17138), .B(n17137), .ZN(n17139) );
  OAI211_X1 U20326 ( .C1(n17141), .C2(n17131), .A(n17140), .B(n17139), .ZN(
        P3_U2734) );
  AND2_X1 U20327 ( .A1(n17190), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20328 ( .A1(n17173), .A2(n17955), .ZN(n17171) );
  AOI22_X1 U20329 ( .A1(n18600), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17144) );
  OAI21_X1 U20330 ( .B1(n17225), .B2(n17171), .A(n17144), .ZN(P3_U2737) );
  INV_X1 U20331 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20332 ( .A1(n18600), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17145) );
  OAI21_X1 U20333 ( .B1(n17146), .B2(n17171), .A(n17145), .ZN(P3_U2738) );
  INV_X1 U20334 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20335 ( .A1(n18600), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17147) );
  OAI21_X1 U20336 ( .B1(n17148), .B2(n17171), .A(n17147), .ZN(P3_U2739) );
  AOI22_X1 U20337 ( .A1(n18600), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17149) );
  OAI21_X1 U20338 ( .B1(n17150), .B2(n17171), .A(n17149), .ZN(P3_U2740) );
  INV_X1 U20339 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17152) );
  AOI22_X1 U20340 ( .A1(n18600), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17151) );
  OAI21_X1 U20341 ( .B1(n17152), .B2(n17171), .A(n17151), .ZN(P3_U2741) );
  AOI22_X1 U20342 ( .A1(n18600), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17153) );
  OAI21_X1 U20343 ( .B1(n17154), .B2(n17171), .A(n17153), .ZN(P3_U2742) );
  AOI22_X1 U20344 ( .A1(n18600), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17155) );
  OAI21_X1 U20345 ( .B1(n17156), .B2(n17171), .A(n17155), .ZN(P3_U2743) );
  AOI22_X1 U20346 ( .A1(n17203), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17157) );
  OAI21_X1 U20347 ( .B1(n17158), .B2(n17171), .A(n17157), .ZN(P3_U2744) );
  INV_X1 U20348 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20349 ( .A1(n17203), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20350 ( .B1(n17160), .B2(n17171), .A(n17159), .ZN(P3_U2745) );
  INV_X1 U20351 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20352 ( .A1(n17203), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17161) );
  OAI21_X1 U20353 ( .B1(n17162), .B2(n17171), .A(n17161), .ZN(P3_U2746) );
  AOI22_X1 U20354 ( .A1(n17203), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17163) );
  OAI21_X1 U20355 ( .B1(n17164), .B2(n17171), .A(n17163), .ZN(P3_U2747) );
  INV_X1 U20356 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20357 ( .A1(n17203), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17165) );
  OAI21_X1 U20358 ( .B1(n17166), .B2(n17171), .A(n17165), .ZN(P3_U2748) );
  AOI22_X1 U20359 ( .A1(n17203), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17167) );
  OAI21_X1 U20360 ( .B1(n17168), .B2(n17171), .A(n17167), .ZN(P3_U2749) );
  INV_X1 U20361 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20362 ( .A1(n17203), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17169) );
  OAI21_X1 U20363 ( .B1(n17211), .B2(n17171), .A(n17169), .ZN(P3_U2750) );
  INV_X1 U20364 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17172) );
  AOI22_X1 U20365 ( .A1(n17203), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17170) );
  OAI21_X1 U20366 ( .B1(n17172), .B2(n17171), .A(n17170), .ZN(P3_U2751) );
  AOI22_X1 U20367 ( .A1(n17203), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17174) );
  OAI21_X1 U20368 ( .B1(n17256), .B2(n17205), .A(n17174), .ZN(P3_U2752) );
  INV_X1 U20369 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20370 ( .A1(n17203), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17175) );
  OAI21_X1 U20371 ( .B1(n17251), .B2(n17205), .A(n17175), .ZN(P3_U2753) );
  INV_X1 U20372 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20373 ( .A1(n17203), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17176) );
  OAI21_X1 U20374 ( .B1(n17177), .B2(n17205), .A(n17176), .ZN(P3_U2754) );
  AOI22_X1 U20375 ( .A1(n17203), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17178) );
  OAI21_X1 U20376 ( .B1(n17179), .B2(n17205), .A(n17178), .ZN(P3_U2755) );
  INV_X1 U20377 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17181) );
  AOI22_X1 U20378 ( .A1(n17203), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17180) );
  OAI21_X1 U20379 ( .B1(n17181), .B2(n17205), .A(n17180), .ZN(P3_U2756) );
  AOI22_X1 U20380 ( .A1(n17203), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17182) );
  OAI21_X1 U20381 ( .B1(n17183), .B2(n17205), .A(n17182), .ZN(P3_U2757) );
  INV_X1 U20382 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20383 ( .A1(n17203), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17184) );
  OAI21_X1 U20384 ( .B1(n17185), .B2(n17205), .A(n17184), .ZN(P3_U2758) );
  AOI22_X1 U20385 ( .A1(n17203), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17186) );
  OAI21_X1 U20386 ( .B1(n17187), .B2(n17205), .A(n17186), .ZN(P3_U2759) );
  INV_X1 U20387 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20388 ( .A1(n17203), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17188) );
  OAI21_X1 U20389 ( .B1(n17189), .B2(n17205), .A(n17188), .ZN(P3_U2760) );
  INV_X1 U20390 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U20391 ( .A1(n17203), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17190), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17191) );
  OAI21_X1 U20392 ( .B1(n17192), .B2(n17205), .A(n17191), .ZN(P3_U2761) );
  INV_X1 U20393 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20394 ( .A1(n17203), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17193) );
  OAI21_X1 U20395 ( .B1(n17194), .B2(n17205), .A(n17193), .ZN(P3_U2762) );
  AOI22_X1 U20396 ( .A1(n17203), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17195) );
  OAI21_X1 U20397 ( .B1(n17196), .B2(n17205), .A(n17195), .ZN(P3_U2763) );
  AOI22_X1 U20398 ( .A1(n17203), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17197) );
  OAI21_X1 U20399 ( .B1(n17198), .B2(n17205), .A(n17197), .ZN(P3_U2764) );
  AOI22_X1 U20400 ( .A1(n17203), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17199) );
  OAI21_X1 U20401 ( .B1(n17200), .B2(n17205), .A(n17199), .ZN(P3_U2765) );
  INV_X1 U20402 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20403 ( .A1(n17203), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17201) );
  OAI21_X1 U20404 ( .B1(n17228), .B2(n17205), .A(n17201), .ZN(P3_U2766) );
  AOI22_X1 U20405 ( .A1(n17203), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17202), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17204) );
  OAI21_X1 U20406 ( .B1(n17206), .B2(n17205), .A(n17204), .ZN(P3_U2767) );
  INV_X2 U20407 ( .A(n17253), .ZN(n17248) );
  NAND3_X1 U20408 ( .A1(n17960), .A2(n17208), .A3(n17207), .ZN(n17255) );
  INV_X2 U20409 ( .A(n17255), .ZN(n17246) );
  AOI22_X1 U20410 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17245), .ZN(n17209) );
  OAI21_X1 U20411 ( .B1(n17950), .B2(n17248), .A(n17209), .ZN(P3_U2768) );
  AOI22_X1 U20412 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17253), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17245), .ZN(n17210) );
  OAI21_X1 U20413 ( .B1(n17211), .B2(n17255), .A(n17210), .ZN(P3_U2769) );
  AOI22_X1 U20414 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17245), .ZN(n17212) );
  OAI21_X1 U20415 ( .B1(n17964), .B2(n17248), .A(n17212), .ZN(P3_U2770) );
  AOI22_X1 U20416 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17245), .ZN(n17213) );
  OAI21_X1 U20417 ( .B1(n17968), .B2(n17248), .A(n17213), .ZN(P3_U2771) );
  AOI22_X1 U20418 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17245), .ZN(n17214) );
  OAI21_X1 U20419 ( .B1(n17972), .B2(n17248), .A(n17214), .ZN(P3_U2772) );
  AOI22_X1 U20420 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17245), .ZN(n17215) );
  OAI21_X1 U20421 ( .B1(n17976), .B2(n17248), .A(n17215), .ZN(P3_U2773) );
  AOI22_X1 U20422 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17245), .ZN(n17216) );
  OAI21_X1 U20423 ( .B1(n17982), .B2(n17248), .A(n17216), .ZN(P3_U2774) );
  AOI22_X1 U20424 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17245), .ZN(n17217) );
  OAI21_X1 U20425 ( .B1(n17986), .B2(n17248), .A(n17217), .ZN(P3_U2775) );
  INV_X1 U20426 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20427 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17245), .ZN(n17218) );
  OAI21_X1 U20428 ( .B1(n17236), .B2(n17248), .A(n17218), .ZN(P3_U2776) );
  AOI22_X1 U20429 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17245), .ZN(n17219) );
  OAI21_X1 U20430 ( .B1(n17238), .B2(n17248), .A(n17219), .ZN(P3_U2777) );
  AOI22_X1 U20431 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17245), .ZN(n17220) );
  OAI21_X1 U20432 ( .B1(n17240), .B2(n17248), .A(n17220), .ZN(P3_U2778) );
  AOI22_X1 U20433 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17245), .ZN(n17221) );
  OAI21_X1 U20434 ( .B1(n17242), .B2(n17248), .A(n17221), .ZN(P3_U2779) );
  AOI22_X1 U20435 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17245), .ZN(n17222) );
  OAI21_X1 U20436 ( .B1(n17244), .B2(n17248), .A(n17222), .ZN(P3_U2780) );
  AOI22_X1 U20437 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17246), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17245), .ZN(n17223) );
  OAI21_X1 U20438 ( .B1(n17249), .B2(n17248), .A(n17223), .ZN(P3_U2781) );
  AOI22_X1 U20439 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17253), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17245), .ZN(n17224) );
  OAI21_X1 U20440 ( .B1(n17225), .B2(n17255), .A(n17224), .ZN(P3_U2782) );
  AOI22_X1 U20441 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17245), .ZN(n17226) );
  OAI21_X1 U20442 ( .B1(n17950), .B2(n17248), .A(n17226), .ZN(P3_U2783) );
  AOI22_X1 U20443 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17253), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17245), .ZN(n17227) );
  OAI21_X1 U20444 ( .B1(n17228), .B2(n17255), .A(n17227), .ZN(P3_U2784) );
  AOI22_X1 U20445 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17245), .ZN(n17229) );
  OAI21_X1 U20446 ( .B1(n17964), .B2(n17248), .A(n17229), .ZN(P3_U2785) );
  AOI22_X1 U20447 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17245), .ZN(n17230) );
  OAI21_X1 U20448 ( .B1(n17968), .B2(n17248), .A(n17230), .ZN(P3_U2786) );
  AOI22_X1 U20449 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17252), .ZN(n17231) );
  OAI21_X1 U20450 ( .B1(n17972), .B2(n17248), .A(n17231), .ZN(P3_U2787) );
  AOI22_X1 U20451 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17252), .ZN(n17232) );
  OAI21_X1 U20452 ( .B1(n17976), .B2(n17248), .A(n17232), .ZN(P3_U2788) );
  AOI22_X1 U20453 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17252), .ZN(n17233) );
  OAI21_X1 U20454 ( .B1(n17982), .B2(n17248), .A(n17233), .ZN(P3_U2789) );
  AOI22_X1 U20455 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17252), .ZN(n17234) );
  OAI21_X1 U20456 ( .B1(n17986), .B2(n17248), .A(n17234), .ZN(P3_U2790) );
  AOI22_X1 U20457 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17252), .ZN(n17235) );
  OAI21_X1 U20458 ( .B1(n17236), .B2(n17248), .A(n17235), .ZN(P3_U2791) );
  AOI22_X1 U20459 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17252), .ZN(n17237) );
  OAI21_X1 U20460 ( .B1(n17238), .B2(n17248), .A(n17237), .ZN(P3_U2792) );
  AOI22_X1 U20461 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17252), .ZN(n17239) );
  OAI21_X1 U20462 ( .B1(n17240), .B2(n17248), .A(n17239), .ZN(P3_U2793) );
  AOI22_X1 U20463 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17252), .ZN(n17241) );
  OAI21_X1 U20464 ( .B1(n17242), .B2(n17248), .A(n17241), .ZN(P3_U2794) );
  AOI22_X1 U20465 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17245), .ZN(n17243) );
  OAI21_X1 U20466 ( .B1(n17244), .B2(n17248), .A(n17243), .ZN(P3_U2795) );
  AOI22_X1 U20467 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17246), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17245), .ZN(n17247) );
  OAI21_X1 U20468 ( .B1(n17249), .B2(n17248), .A(n17247), .ZN(P3_U2796) );
  AOI22_X1 U20469 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17253), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17252), .ZN(n17250) );
  OAI21_X1 U20470 ( .B1(n17251), .B2(n17255), .A(n17250), .ZN(P3_U2797) );
  AOI22_X1 U20471 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17253), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17252), .ZN(n17254) );
  OAI21_X1 U20472 ( .B1(n17256), .B2(n17255), .A(n17254), .ZN(P3_U2798) );
  AOI21_X1 U20473 ( .B1(n9847), .B2(n17258), .A(n17257), .ZN(n17630) );
  OAI22_X1 U20474 ( .A1(n17930), .A2(n18535), .B1(n17450), .B2(n17259), .ZN(
        n17260) );
  AOI211_X1 U20475 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17262), .A(
        n17261), .B(n17260), .ZN(n17266) );
  OAI21_X1 U20476 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17264), .A(
        n17263), .ZN(n17265) );
  OAI211_X1 U20477 ( .C1(n17630), .C2(n17498), .A(n17266), .B(n17265), .ZN(
        P3_U2803) );
  INV_X1 U20478 ( .A(n17267), .ZN(n17268) );
  AOI21_X1 U20479 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17269), .A(
        n17268), .ZN(n17637) );
  INV_X1 U20480 ( .A(n17391), .ZN(n17413) );
  NOR4_X1 U20481 ( .A1(n17663), .A2(n17654), .A3(n17294), .A4(n17413), .ZN(
        n17278) );
  INV_X1 U20482 ( .A(n17270), .ZN(n17277) );
  AOI21_X1 U20483 ( .B1(n18329), .B2(n17271), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17274) );
  OAI21_X1 U20484 ( .B1(n17465), .B2(n17353), .A(n17272), .ZN(n17273) );
  NAND2_X1 U20485 ( .A1(n17627), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17635) );
  OAI211_X1 U20486 ( .C1(n17275), .C2(n17274), .A(n17273), .B(n17635), .ZN(
        n17276) );
  AOI221_X1 U20487 ( .B1(n17278), .B2(n12240), .C1(n17277), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17276), .ZN(n17279) );
  OAI21_X1 U20488 ( .B1(n17637), .B2(n17498), .A(n17279), .ZN(P3_U2804) );
  NAND2_X1 U20489 ( .A1(n18329), .A2(n17288), .ZN(n17311) );
  OAI211_X1 U20490 ( .C1(n17280), .C2(n18464), .A(n17609), .B(n17311), .ZN(
        n17307) );
  AOI22_X1 U20491 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17307), .B1(
        n17465), .B2(n17281), .ZN(n17293) );
  NOR2_X1 U20492 ( .A1(n17681), .A2(n17294), .ZN(n17659) );
  NAND2_X1 U20493 ( .A1(n17659), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17282) );
  XOR2_X1 U20494 ( .A(n17282), .B(n17654), .Z(n17643) );
  NOR2_X1 U20495 ( .A1(n17682), .A2(n17294), .ZN(n17316) );
  NAND2_X1 U20496 ( .A1(n17316), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17283) );
  XOR2_X1 U20497 ( .A(n17283), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17649) );
  OAI21_X1 U20498 ( .B1(n9847), .B2(n17285), .A(n17284), .ZN(n17286) );
  XOR2_X1 U20499 ( .A(n17286), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17648) );
  OAI22_X1 U20500 ( .A1(n17649), .A2(n17613), .B1(n17498), .B2(n17648), .ZN(
        n17287) );
  AOI21_X1 U20501 ( .B1(n17520), .B2(n17643), .A(n17287), .ZN(n17292) );
  NAND2_X1 U20502 ( .A1(n17627), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17652) );
  NOR2_X1 U20503 ( .A1(n17289), .A2(n17288), .ZN(n17298) );
  OAI211_X1 U20504 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17298), .B(n17290), .ZN(n17291) );
  NAND4_X1 U20505 ( .A1(n17293), .A2(n17292), .A3(n17652), .A4(n17291), .ZN(
        P3_U2805) );
  OR2_X1 U20506 ( .A1(n17294), .A2(n17413), .ZN(n17303) );
  OAI22_X1 U20507 ( .A1(n17930), .A2(n18528), .B1(n17450), .B2(n17295), .ZN(
        n17296) );
  AOI221_X1 U20508 ( .B1(n17298), .B2(n17297), .C1(n17307), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17296), .ZN(n17302) );
  OAI22_X1 U20509 ( .A1(n17659), .A2(n17454), .B1(n17316), .B2(n17613), .ZN(
        n17319) );
  OAI21_X1 U20510 ( .B1(n17300), .B2(n17663), .A(n17299), .ZN(n17655) );
  AOI22_X1 U20511 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17319), .B1(
        n17519), .B2(n17655), .ZN(n17301) );
  OAI211_X1 U20512 ( .C1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n17303), .A(
        n17302), .B(n17301), .ZN(P3_U2806) );
  AOI21_X1 U20513 ( .B1(n17304), .B2(n17383), .A(n17332), .ZN(n17305) );
  AOI211_X1 U20514 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n9847), .A(
        n17348), .B(n17305), .ZN(n17306) );
  XOR2_X1 U20515 ( .A(n17668), .B(n17306), .Z(n17673) );
  INV_X1 U20516 ( .A(n17307), .ZN(n17309) );
  AOI211_X1 U20517 ( .C1(n17354), .C2(n17310), .A(n17309), .B(n17308), .ZN(
        n17314) );
  OAI22_X1 U20518 ( .A1(n17930), .A2(n18526), .B1(n17312), .B2(n17311), .ZN(
        n17313) );
  AOI211_X1 U20519 ( .C1(n17315), .C2(n17465), .A(n17314), .B(n17313), .ZN(
        n17322) );
  INV_X1 U20520 ( .A(n17316), .ZN(n17657) );
  NAND2_X1 U20521 ( .A1(n17601), .A2(n17657), .ZN(n17318) );
  NAND3_X1 U20522 ( .A1(n17752), .A2(n17520), .A3(n17668), .ZN(n17317) );
  OAI21_X1 U20523 ( .B1(n17318), .B2(n17682), .A(n17317), .ZN(n17320) );
  AOI22_X1 U20524 ( .A1(n17618), .A2(n17320), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17319), .ZN(n17321) );
  OAI211_X1 U20525 ( .C1(n17498), .C2(n17673), .A(n17322), .B(n17321), .ZN(
        P3_U2807) );
  NAND2_X1 U20526 ( .A1(n17325), .A2(n17446), .ZN(n17342) );
  AOI221_X1 U20527 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17341), .C2(n17326), .A(
        n17342), .ZN(n17328) );
  INV_X1 U20528 ( .A(n18464), .ZN(n17444) );
  NAND2_X1 U20529 ( .A1(n17444), .A2(n17323), .ZN(n17324) );
  OAI211_X1 U20530 ( .C1(n17325), .C2(n17566), .A(n17609), .B(n17324), .ZN(
        n17358) );
  AOI21_X1 U20531 ( .B1(n17353), .B2(n17350), .A(n17358), .ZN(n17340) );
  NAND2_X1 U20532 ( .A1(n17932), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17689) );
  OAI21_X1 U20533 ( .B1(n17340), .B2(n17326), .A(n17689), .ZN(n17327) );
  AOI211_X1 U20534 ( .C1(n17329), .C2(n17465), .A(n17328), .B(n17327), .ZN(
        n17336) );
  OAI22_X1 U20535 ( .A1(n17454), .A2(n17752), .B1(n17613), .B2(n17760), .ZN(
        n17374) );
  INV_X1 U20536 ( .A(n17374), .ZN(n17412) );
  OAI21_X1 U20537 ( .B1(n17679), .B2(n17359), .A(n17412), .ZN(n17345) );
  INV_X1 U20538 ( .A(n17348), .ZN(n17330) );
  OAI221_X1 U20539 ( .B1(n17332), .B2(n17331), .C1(n17332), .C2(n17337), .A(
        n17330), .ZN(n17333) );
  XOR2_X1 U20540 ( .A(n17691), .B(n17333), .Z(n17688) );
  AOI22_X1 U20541 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17345), .B1(
        n17519), .B2(n17688), .ZN(n17335) );
  NAND3_X1 U20542 ( .A1(n17679), .A2(n17391), .A3(n17691), .ZN(n17334) );
  NAND3_X1 U20543 ( .A1(n17336), .A2(n17335), .A3(n17334), .ZN(P3_U2808) );
  NAND3_X1 U20544 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17518), .A3(
        n17337), .ZN(n17362) );
  OAI22_X1 U20545 ( .A1(n17695), .A2(n17362), .B1(n17338), .B2(n17383), .ZN(
        n17339) );
  XOR2_X1 U20546 ( .A(n17694), .B(n17339), .Z(n17706) );
  NAND2_X1 U20547 ( .A1(n17627), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17704) );
  OAI221_X1 U20548 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17342), .C1(
        n17341), .C2(n17340), .A(n17704), .ZN(n17343) );
  AOI21_X1 U20549 ( .B1(n17465), .B2(n17344), .A(n17343), .ZN(n17347) );
  NOR2_X1 U20550 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17695), .ZN(
        n17703) );
  NAND2_X1 U20551 ( .A1(n17729), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17697) );
  NOR2_X1 U20552 ( .A1(n17413), .A2(n17697), .ZN(n17370) );
  AOI22_X1 U20553 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17345), .B1(
        n17703), .B2(n17370), .ZN(n17346) );
  OAI211_X1 U20554 ( .C1(n17706), .C2(n17498), .A(n17347), .B(n17346), .ZN(
        P3_U2809) );
  INV_X1 U20555 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17723) );
  XOR2_X1 U20556 ( .A(n20755), .B(n17349), .Z(n17716) );
  OAI21_X1 U20557 ( .B1(n17351), .B2(n17980), .A(n17350), .ZN(n17357) );
  INV_X1 U20558 ( .A(n17352), .ZN(n17355) );
  INV_X1 U20559 ( .A(n17353), .ZN(n17354) );
  NAND2_X1 U20560 ( .A1(n17627), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17714) );
  OAI221_X1 U20561 ( .B1(n17355), .B2(n17450), .C1(n17355), .C2(n17354), .A(
        n17714), .ZN(n17356) );
  AOI21_X1 U20562 ( .B1(n17358), .B2(n17357), .A(n17356), .ZN(n17361) );
  NOR2_X1 U20563 ( .A1(n17723), .A2(n17697), .ZN(n17708) );
  OAI21_X1 U20564 ( .B1(n17359), .B2(n17708), .A(n17412), .ZN(n17371) );
  NOR2_X1 U20565 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17723), .ZN(
        n17712) );
  AOI22_X1 U20566 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17371), .B1(
        n17370), .B2(n17712), .ZN(n17360) );
  OAI211_X1 U20567 ( .C1(n17498), .C2(n17716), .A(n17361), .B(n17360), .ZN(
        P3_U2810) );
  OAI21_X1 U20568 ( .B1(n17383), .B2(n17381), .A(n17362), .ZN(n17363) );
  XOR2_X1 U20569 ( .A(n17363), .B(n17723), .Z(n17717) );
  NAND2_X1 U20570 ( .A1(n17364), .A2(n17446), .ZN(n17378) );
  AOI221_X1 U20571 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n17377), .C2(n17367), .A(
        n17378), .ZN(n17369) );
  OAI21_X1 U20572 ( .B1(n17364), .B2(n17566), .A(n17609), .ZN(n17398) );
  AOI21_X1 U20573 ( .B1(n17444), .B2(n17365), .A(n17398), .ZN(n17376) );
  OAI22_X1 U20574 ( .A1(n17376), .A2(n17367), .B1(n17450), .B2(n17366), .ZN(
        n17368) );
  AOI211_X1 U20575 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n17932), .A(n17369), 
        .B(n17368), .ZN(n17373) );
  AOI22_X1 U20576 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17371), .B1(
        n17370), .B2(n17723), .ZN(n17372) );
  OAI211_X1 U20577 ( .C1(n17717), .C2(n17498), .A(n17373), .B(n17372), .ZN(
        P3_U2811) );
  AOI21_X1 U20578 ( .B1(n17391), .B2(n17384), .A(n17374), .ZN(n17393) );
  NAND2_X1 U20579 ( .A1(n17627), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17375) );
  OAI221_X1 U20580 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17378), .C1(
        n17377), .C2(n17376), .A(n17375), .ZN(n17379) );
  AOI21_X1 U20581 ( .B1(n17465), .B2(n17380), .A(n17379), .ZN(n17386) );
  OAI21_X1 U20582 ( .B1(n17693), .B2(n9847), .A(n17381), .ZN(n17382) );
  XOR2_X1 U20583 ( .A(n17383), .B(n17382), .Z(n17735) );
  NOR2_X1 U20584 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17384), .ZN(
        n17734) );
  AOI22_X1 U20585 ( .A1(n17519), .A2(n17735), .B1(n17391), .B2(n17734), .ZN(
        n17385) );
  OAI211_X1 U20586 ( .C1(n17393), .C2(n17693), .A(n17386), .B(n17385), .ZN(
        P3_U2812) );
  AOI21_X1 U20587 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17388), .A(
        n17387), .ZN(n17742) );
  OAI21_X1 U20588 ( .B1(n17980), .B2(n17390), .A(n17389), .ZN(n17397) );
  NOR2_X1 U20589 ( .A1(n17930), .A2(n18514), .ZN(n17396) );
  AOI21_X1 U20590 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17391), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17392) );
  OAI22_X1 U20591 ( .A1(n17593), .A2(n17394), .B1(n17393), .B2(n17392), .ZN(
        n17395) );
  AOI211_X1 U20592 ( .C1(n17398), .C2(n17397), .A(n17396), .B(n17395), .ZN(
        n17399) );
  OAI21_X1 U20593 ( .B1(n17742), .B2(n17498), .A(n17399), .ZN(P3_U2813) );
  NAND2_X1 U20594 ( .A1(n17518), .A2(n17400), .ZN(n17499) );
  INV_X1 U20595 ( .A(n17499), .ZN(n17462) );
  AOI22_X1 U20596 ( .A1(n9847), .A2(n17402), .B1(n17401), .B2(n17462), .ZN(
        n17403) );
  XOR2_X1 U20597 ( .A(n17747), .B(n17403), .Z(n17749) );
  OAI21_X1 U20598 ( .B1(n13174), .B2(n17566), .A(n17609), .ZN(n17431) );
  AOI21_X1 U20599 ( .B1(n17444), .B2(n17404), .A(n17431), .ZN(n17414) );
  OAI22_X1 U20600 ( .A1(n17414), .A2(n17406), .B1(n17450), .B2(n17405), .ZN(
        n17410) );
  OAI211_X1 U20601 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n13174), .B(n17446), .ZN(n17407) );
  OAI22_X1 U20602 ( .A1(n17408), .A2(n17407), .B1(n17930), .B2(n18512), .ZN(
        n17409) );
  AOI211_X1 U20603 ( .C1(n17519), .C2(n17749), .A(n17410), .B(n17409), .ZN(
        n17411) );
  OAI221_X1 U20604 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17413), 
        .C1(n17747), .C2(n17412), .A(n17411), .ZN(P3_U2814) );
  INV_X1 U20605 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n20759) );
  INV_X1 U20606 ( .A(n17442), .ZN(n17793) );
  INV_X1 U20607 ( .A(n17805), .ZN(n17483) );
  NOR2_X1 U20608 ( .A1(n17793), .A2(n17483), .ZN(n17453) );
  INV_X1 U20609 ( .A(n17453), .ZN(n17786) );
  NOR3_X1 U20610 ( .A1(n17771), .A2(n20759), .A3(n17786), .ZN(n17432) );
  NOR2_X1 U20611 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17432), .ZN(
        n17759) );
  NAND2_X1 U20612 ( .A1(n17601), .A2(n17682), .ZN(n17427) );
  NAND2_X1 U20613 ( .A1(n13174), .A2(n17446), .ZN(n17416) );
  NAND2_X1 U20614 ( .A1(n17627), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17761) );
  OAI221_X1 U20615 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17416), .C1(
        n17415), .C2(n17414), .A(n17761), .ZN(n17417) );
  AOI21_X1 U20616 ( .B1(n17465), .B2(n17418), .A(n17417), .ZN(n17426) );
  NAND2_X1 U20617 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17518), .ZN(
        n17455) );
  NAND2_X1 U20618 ( .A1(n17419), .A2(n9847), .ZN(n17473) );
  OR3_X1 U20619 ( .A1(n17473), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17433) );
  NOR2_X1 U20620 ( .A1(n17783), .A2(n17420), .ZN(n17457) );
  NAND3_X1 U20621 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n17457), .ZN(n17421) );
  AOI22_X1 U20622 ( .A1(n17422), .A2(n17455), .B1(n17433), .B2(n17421), .ZN(
        n17423) );
  XOR2_X1 U20623 ( .A(n17423), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n17765) );
  NOR2_X1 U20624 ( .A1(n17752), .A2(n17454), .ZN(n17424) );
  INV_X1 U20625 ( .A(n17435), .ZN(n17770) );
  INV_X1 U20626 ( .A(n17808), .ZN(n17484) );
  INV_X1 U20627 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17762) );
  OAI21_X1 U20628 ( .B1(n17770), .B2(n17484), .A(n17762), .ZN(n17757) );
  AOI22_X1 U20629 ( .A1(n17519), .A2(n17765), .B1(n17424), .B2(n17757), .ZN(
        n17425) );
  OAI211_X1 U20630 ( .C1(n17759), .C2(n17427), .A(n17426), .B(n17425), .ZN(
        P3_U2815) );
  OAI21_X1 U20631 ( .B1(n17429), .B2(n17980), .A(n17428), .ZN(n17430) );
  AOI22_X1 U20632 ( .A1(n17932), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17431), 
        .B2(n17430), .ZN(n17440) );
  AOI221_X1 U20633 ( .B1(n20759), .B2(n17771), .C1(n17786), .C2(n17771), .A(
        n17432), .ZN(n17777) );
  OAI22_X1 U20634 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17433), .B1(
        n17499), .B2(n17754), .ZN(n17434) );
  XOR2_X1 U20635 ( .A(n17771), .B(n17434), .Z(n17781) );
  INV_X1 U20636 ( .A(n17754), .ZN(n17437) );
  NAND2_X1 U20637 ( .A1(n17435), .A2(n17808), .ZN(n17436) );
  OAI221_X1 U20638 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17437), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17808), .A(n17436), .ZN(
        n17774) );
  OAI22_X1 U20639 ( .A1(n17781), .A2(n17498), .B1(n17454), .B2(n17774), .ZN(
        n17438) );
  AOI21_X1 U20640 ( .B1(n17601), .B2(n17777), .A(n17438), .ZN(n17439) );
  OAI211_X1 U20641 ( .C1(n17593), .C2(n17441), .A(n17440), .B(n17439), .ZN(
        P3_U2816) );
  NAND2_X1 U20642 ( .A1(n17442), .A2(n20759), .ZN(n17792) );
  NAND2_X1 U20643 ( .A1(n17444), .A2(n17443), .ZN(n17445) );
  OAI211_X1 U20644 ( .C1(n17479), .C2(n17566), .A(n17609), .B(n17445), .ZN(
        n17466) );
  NAND2_X1 U20645 ( .A1(n17479), .A2(n17446), .ZN(n17468) );
  AOI221_X1 U20646 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C1(n17448), .C2(n17447), .A(
        n17468), .ZN(n17452) );
  OAI22_X1 U20647 ( .A1(n17930), .A2(n18506), .B1(n17450), .B2(n17449), .ZN(
        n17451) );
  AOI211_X1 U20648 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17466), .A(
        n17452), .B(n17451), .ZN(n17460) );
  NOR2_X1 U20649 ( .A1(n17793), .A2(n17484), .ZN(n17784) );
  OAI22_X1 U20650 ( .A1(n17784), .A2(n17454), .B1(n17453), .B2(n17613), .ZN(
        n17470) );
  NOR2_X1 U20651 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17473), .ZN(
        n17461) );
  INV_X1 U20652 ( .A(n17455), .ZN(n17456) );
  OAI22_X1 U20653 ( .A1(n17457), .A2(n17794), .B1(n17461), .B2(n17456), .ZN(
        n17458) );
  XOR2_X1 U20654 ( .A(n20759), .B(n17458), .Z(n17782) );
  AOI22_X1 U20655 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17470), .B1(
        n17519), .B2(n17782), .ZN(n17459) );
  OAI211_X1 U20656 ( .C1(n17511), .C2(n17792), .A(n17460), .B(n17459), .ZN(
        P3_U2817) );
  INV_X1 U20657 ( .A(n17783), .ZN(n17796) );
  AOI21_X1 U20658 ( .B1(n17462), .B2(n17796), .A(n17461), .ZN(n17463) );
  XOR2_X1 U20659 ( .A(n17463), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17803) );
  NOR2_X1 U20660 ( .A1(n17511), .A2(n17783), .ZN(n17471) );
  AOI22_X1 U20661 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17466), .B1(
        n17465), .B2(n17464), .ZN(n17467) );
  NAND2_X1 U20662 ( .A1(n17932), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17801) );
  OAI211_X1 U20663 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17468), .A(
        n17467), .B(n17801), .ZN(n17469) );
  AOI221_X1 U20664 ( .B1(n17471), .B2(n17794), .C1(n17470), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17469), .ZN(n17472) );
  OAI21_X1 U20665 ( .B1(n17803), .B2(n17498), .A(n17472), .ZN(P3_U2818) );
  INV_X1 U20666 ( .A(n17814), .ZN(n17474) );
  OR2_X1 U20667 ( .A1(n17474), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17819) );
  OAI21_X1 U20668 ( .B1(n17499), .B2(n17474), .A(n17473), .ZN(n17475) );
  XOR2_X1 U20669 ( .A(n17475), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n17804) );
  NAND3_X1 U20670 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17477) );
  INV_X1 U20671 ( .A(n17476), .ZN(n17538) );
  NAND4_X1 U20672 ( .A1(n18329), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n17538), .A4(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17513) );
  NOR2_X1 U20673 ( .A1(n17477), .A2(n17513), .ZN(n17491) );
  AOI21_X1 U20674 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17604), .A(
        n17491), .ZN(n17478) );
  AOI21_X1 U20675 ( .B1(n17479), .B2(n18329), .A(n17478), .ZN(n17482) );
  INV_X1 U20676 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18502) );
  OAI22_X1 U20677 ( .A1(n17593), .A2(n17480), .B1(n17930), .B2(n18502), .ZN(
        n17481) );
  AOI211_X1 U20678 ( .C1(n17519), .C2(n17804), .A(n17482), .B(n17481), .ZN(
        n17486) );
  NOR2_X1 U20679 ( .A1(n17814), .A2(n17511), .ZN(n17495) );
  AOI22_X1 U20680 ( .A1(n17484), .A2(n17520), .B1(n17483), .B2(n17601), .ZN(
        n17510) );
  INV_X1 U20681 ( .A(n17510), .ZN(n17494) );
  OAI21_X1 U20682 ( .B1(n17495), .B2(n17494), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17485) );
  OAI211_X1 U20683 ( .C1(n17511), .C2(n17819), .A(n17486), .B(n17485), .ZN(
        P3_U2819) );
  NAND2_X1 U20684 ( .A1(n17487), .A2(n17846), .ZN(n17500) );
  AOI22_X1 U20685 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17499), .B1(
        n17500), .B2(n17836), .ZN(n17488) );
  XOR2_X1 U20686 ( .A(n17822), .B(n17488), .Z(n17828) );
  NOR2_X1 U20687 ( .A1(n17930), .A2(n18500), .ZN(n17493) );
  INV_X1 U20688 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20793) );
  NOR3_X1 U20689 ( .A1(n20793), .A2(n17502), .A3(n17513), .ZN(n17506) );
  AOI21_X1 U20690 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17604), .A(
        n17506), .ZN(n17490) );
  OAI22_X1 U20691 ( .A1(n17491), .A2(n17490), .B1(n17593), .B2(n17489), .ZN(
        n17492) );
  AOI211_X1 U20692 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17494), .A(
        n17493), .B(n17492), .ZN(n17497) );
  OAI21_X1 U20693 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17495), .ZN(n17496) );
  OAI211_X1 U20694 ( .C1(n17828), .C2(n17498), .A(n17497), .B(n17496), .ZN(
        P3_U2820) );
  NAND2_X1 U20695 ( .A1(n17500), .A2(n17499), .ZN(n17501) );
  XOR2_X1 U20696 ( .A(n17501), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n17833) );
  NOR2_X1 U20697 ( .A1(n17930), .A2(n18498), .ZN(n17508) );
  NOR2_X1 U20698 ( .A1(n17502), .A2(n17513), .ZN(n17503) );
  AOI21_X1 U20699 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17604), .A(
        n17503), .ZN(n17505) );
  OAI22_X1 U20700 ( .A1(n17506), .A2(n17505), .B1(n17593), .B2(n17504), .ZN(
        n17507) );
  AOI211_X1 U20701 ( .C1(n17519), .C2(n17833), .A(n17508), .B(n17507), .ZN(
        n17509) );
  OAI221_X1 U20702 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17511), .C1(
        n17836), .C2(n17510), .A(n17509), .ZN(P3_U2821) );
  OAI21_X1 U20703 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17852), .A(
        n17851), .ZN(n17523) );
  AOI21_X1 U20704 ( .B1(n17512), .B2(n17525), .A(n17596), .ZN(n17527) );
  OAI21_X1 U20705 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17980), .A(
        n17527), .ZN(n17516) );
  NOR2_X1 U20706 ( .A1(n17930), .A2(n18497), .ZN(n17847) );
  OAI22_X1 U20707 ( .A1(n17593), .A2(n17514), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17513), .ZN(n17515) );
  AOI211_X1 U20708 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17516), .A(
        n17847), .B(n17515), .ZN(n17522) );
  OAI21_X1 U20709 ( .B1(n17518), .B2(n17840), .A(n17517), .ZN(n17849) );
  AOI22_X1 U20710 ( .A1(n17840), .A2(n17520), .B1(n17519), .B2(n17849), .ZN(
        n17521) );
  OAI211_X1 U20711 ( .C1(n17613), .C2(n17523), .A(n17522), .B(n17521), .ZN(
        P3_U2822) );
  NAND2_X1 U20712 ( .A1(n18329), .A2(n17526), .ZN(n17524) );
  OAI22_X1 U20713 ( .A1(n17527), .A2(n17526), .B1(n17525), .B2(n17524), .ZN(
        n17535) );
  OAI21_X1 U20714 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17529), .A(
        n17528), .ZN(n17858) );
  OAI21_X1 U20715 ( .B1(n17532), .B2(n17531), .A(n17530), .ZN(n17533) );
  XOR2_X1 U20716 ( .A(n17533), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n17864) );
  OAI22_X1 U20717 ( .A1(n17612), .A2(n17858), .B1(n17613), .B2(n17864), .ZN(
        n17534) );
  AOI211_X1 U20718 ( .C1(n17932), .C2(P3_REIP_REG_7__SCAN_IN), .A(n17535), .B(
        n17534), .ZN(n17536) );
  OAI21_X1 U20719 ( .B1(n17593), .B2(n17537), .A(n17536), .ZN(P3_U2823) );
  NAND2_X1 U20720 ( .A1(n18329), .A2(n17538), .ZN(n17542) );
  NAND2_X1 U20721 ( .A1(n17604), .A2(n17542), .ZN(n17552) );
  OAI21_X1 U20722 ( .B1(n17541), .B2(n17540), .A(n17539), .ZN(n17866) );
  OAI22_X1 U20723 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17542), .B1(
        n17612), .B2(n17866), .ZN(n17547) );
  OAI21_X1 U20724 ( .B1(n17544), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17543), .ZN(n17873) );
  OAI22_X1 U20725 ( .A1(n17593), .A2(n17545), .B1(n17613), .B2(n17873), .ZN(
        n17546) );
  AOI211_X1 U20726 ( .C1(n17932), .C2(P3_REIP_REG_6__SCAN_IN), .A(n17547), .B(
        n17546), .ZN(n17548) );
  OAI21_X1 U20727 ( .B1(n20724), .B2(n17552), .A(n17548), .ZN(P3_U2824) );
  OAI21_X1 U20728 ( .B1(n17551), .B2(n17550), .A(n17549), .ZN(n17874) );
  AOI221_X1 U20729 ( .B1(n17596), .B2(n17554), .C1(n17553), .C2(n17554), .A(
        n17552), .ZN(n17560) );
  INV_X1 U20730 ( .A(n17557), .ZN(n17556) );
  OAI222_X1 U20731 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17558), .B1(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17557), .C1(n17556), .C2(
        n17555), .ZN(n17880) );
  OAI22_X1 U20732 ( .A1(n17930), .A2(n18491), .B1(n17612), .B2(n17880), .ZN(
        n17559) );
  AOI211_X1 U20733 ( .C1(n17561), .C2(n17603), .A(n17560), .B(n17559), .ZN(
        n17562) );
  OAI21_X1 U20734 ( .B1(n17613), .B2(n17874), .A(n17562), .ZN(P3_U2825) );
  OAI21_X1 U20735 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17564), .A(
        n17563), .ZN(n17883) );
  AOI22_X1 U20736 ( .A1(n17932), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18329), 
        .B2(n17565), .ZN(n17574) );
  OAI21_X1 U20737 ( .B1(n17567), .B2(n17566), .A(n17609), .ZN(n17584) );
  OAI21_X1 U20738 ( .B1(n17570), .B2(n17569), .A(n17568), .ZN(n17884) );
  OAI22_X1 U20739 ( .A1(n17593), .A2(n17571), .B1(n17612), .B2(n17884), .ZN(
        n17572) );
  AOI21_X1 U20740 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17584), .A(
        n17572), .ZN(n17573) );
  OAI211_X1 U20741 ( .C1(n17613), .C2(n17883), .A(n17574), .B(n17573), .ZN(
        P3_U2826) );
  OAI21_X1 U20742 ( .B1(n17577), .B2(n17576), .A(n17575), .ZN(n17891) );
  NOR2_X1 U20743 ( .A1(n17596), .A2(n17595), .ZN(n17583) );
  INV_X1 U20744 ( .A(n17578), .ZN(n17581) );
  OAI21_X1 U20745 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17580), .A(
        n17579), .ZN(n17892) );
  OAI22_X1 U20746 ( .A1(n17593), .A2(n17581), .B1(n17612), .B2(n17892), .ZN(
        n17582) );
  AOI221_X1 U20747 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17584), .C1(
        n17583), .C2(n17584), .A(n17582), .ZN(n17585) );
  NAND2_X1 U20748 ( .A1(n17627), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n17896) );
  OAI211_X1 U20749 ( .C1(n17613), .C2(n17891), .A(n17585), .B(n17896), .ZN(
        P3_U2827) );
  OAI21_X1 U20750 ( .B1(n17588), .B2(n17587), .A(n17586), .ZN(n17907) );
  OAI21_X1 U20751 ( .B1(n17591), .B2(n17590), .A(n17589), .ZN(n17908) );
  OAI22_X1 U20752 ( .A1(n17593), .A2(n17592), .B1(n17612), .B2(n17908), .ZN(
        n17594) );
  AOI221_X1 U20753 ( .B1(n17596), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18329), .C2(n17595), .A(n17594), .ZN(n17597) );
  NAND2_X1 U20754 ( .A1(n17627), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n17912) );
  OAI211_X1 U20755 ( .C1(n17613), .C2(n17907), .A(n17597), .B(n17912), .ZN(
        P3_U2828) );
  OAI21_X1 U20756 ( .B1(n17599), .B2(n17607), .A(n17598), .ZN(n17927) );
  NAND2_X1 U20757 ( .A1(n18583), .A2(n17608), .ZN(n17600) );
  XNOR2_X1 U20758 ( .A(n17600), .B(n17599), .ZN(n17920) );
  AOI22_X1 U20759 ( .A1(n17932), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17601), 
        .B2(n17920), .ZN(n17606) );
  AOI22_X1 U20760 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17604), .B1(
        n17603), .B2(n17602), .ZN(n17605) );
  OAI211_X1 U20761 ( .C1(n17612), .C2(n17927), .A(n17606), .B(n17605), .ZN(
        P3_U2829) );
  AOI21_X1 U20762 ( .B1(n17608), .B2(n18583), .A(n17607), .ZN(n17937) );
  INV_X1 U20763 ( .A(n17937), .ZN(n17935) );
  NAND3_X1 U20764 ( .A1(n18566), .A2(n18464), .A3(n17609), .ZN(n17610) );
  AOI22_X1 U20765 ( .A1(n17932), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17610), .ZN(n17611) );
  OAI221_X1 U20766 ( .B1(n17937), .B2(n17613), .C1(n17935), .C2(n17612), .A(
        n17611), .ZN(P3_U2830) );
  NOR2_X1 U20767 ( .A1(n17668), .A2(n17669), .ZN(n17664) );
  NAND3_X1 U20768 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n17664), .ZN(n17632) );
  NOR2_X1 U20769 ( .A1(n12240), .A2(n17632), .ZN(n17625) );
  AOI22_X1 U20770 ( .A1(n18409), .A2(n17614), .B1(n18396), .B2(n17654), .ZN(
        n17622) );
  AOI22_X1 U20771 ( .A1(n18384), .A2(n17616), .B1(n17839), .B2(n17615), .ZN(
        n17621) );
  INV_X1 U20772 ( .A(n18409), .ZN(n18422) );
  NOR2_X1 U20773 ( .A1(n18422), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17901) );
  INV_X1 U20774 ( .A(n17678), .ZN(n17617) );
  NOR2_X1 U20775 ( .A1(n17901), .A2(n17617), .ZN(n17724) );
  NAND2_X1 U20776 ( .A1(n17618), .A2(n17724), .ZN(n17656) );
  OAI21_X1 U20777 ( .B1(n17619), .B2(n17656), .A(n17903), .ZN(n17641) );
  NAND4_X1 U20778 ( .A1(n17622), .A2(n17621), .A3(n17620), .A4(n17641), .ZN(
        n17631) );
  AOI21_X1 U20779 ( .B1(n18396), .B2(n12240), .A(n17631), .ZN(n17623) );
  INV_X1 U20780 ( .A(n17623), .ZN(n17624) );
  MUX2_X1 U20781 ( .A(n17625), .B(n17624), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17626) );
  AOI22_X1 U20782 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17924), .B1(
        n17928), .B2(n17626), .ZN(n17629) );
  NAND2_X1 U20783 ( .A1(n17627), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17628) );
  OAI211_X1 U20784 ( .C1(n17630), .C2(n17827), .A(n17629), .B(n17628), .ZN(
        P3_U2835) );
  INV_X1 U20785 ( .A(n17631), .ZN(n17633) );
  AOI221_X1 U20786 ( .B1(n17633), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n17632), .C2(n12240), .A(n17922), .ZN(n17634) );
  AOI21_X1 U20787 ( .B1(n17924), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17634), .ZN(n17636) );
  OAI211_X1 U20788 ( .C1(n17637), .C2(n17827), .A(n17636), .B(n17635), .ZN(
        P3_U2836) );
  NOR2_X1 U20789 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17663), .ZN(
        n17638) );
  NAND2_X1 U20790 ( .A1(n17639), .A2(n17638), .ZN(n17646) );
  INV_X1 U20791 ( .A(n17725), .ZN(n17676) );
  OAI21_X1 U20792 ( .B1(n17640), .B2(n17676), .A(n18385), .ZN(n17661) );
  OAI211_X1 U20793 ( .C1(n17642), .C2(n18416), .A(n17661), .B(n17641), .ZN(
        n17644) );
  AOI22_X1 U20794 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17644), .B1(
        n17839), .B2(n17643), .ZN(n17645) );
  OAI21_X1 U20795 ( .B1(n17647), .B2(n17646), .A(n17645), .ZN(n17651) );
  OAI22_X1 U20796 ( .A1(n17649), .A2(n17936), .B1(n17827), .B2(n17648), .ZN(
        n17650) );
  AOI21_X1 U20797 ( .B1(n17928), .B2(n17651), .A(n17650), .ZN(n17653) );
  OAI211_X1 U20798 ( .C1(n17915), .C2(n17654), .A(n17653), .B(n17652), .ZN(
        P3_U2837) );
  AOI22_X1 U20799 ( .A1(n17932), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17850), 
        .B2(n17655), .ZN(n17667) );
  AOI22_X1 U20800 ( .A1(n18384), .A2(n17657), .B1(n17903), .B2(n17656), .ZN(
        n17658) );
  OAI211_X1 U20801 ( .C1(n17659), .C2(n17807), .A(n17658), .B(n17915), .ZN(
        n17662) );
  NOR2_X1 U20802 ( .A1(n17668), .A2(n17662), .ZN(n17660) );
  AOI21_X1 U20803 ( .B1(n17661), .B2(n17660), .A(n17932), .ZN(n17671) );
  OAI211_X1 U20804 ( .C1(n17882), .C2(n17662), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17671), .ZN(n17666) );
  NAND3_X1 U20805 ( .A1(n17928), .A2(n17664), .A3(n17663), .ZN(n17665) );
  NAND3_X1 U20806 ( .A1(n17667), .A2(n17666), .A3(n17665), .ZN(P3_U2838) );
  OAI21_X1 U20807 ( .B1(n17924), .B2(n17669), .A(n17668), .ZN(n17670) );
  AOI22_X1 U20808 ( .A1(n17932), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17671), 
        .B2(n17670), .ZN(n17672) );
  OAI21_X1 U20809 ( .B1(n17827), .B2(n17673), .A(n17672), .ZN(P3_U2839) );
  NAND2_X1 U20810 ( .A1(n17928), .A2(n17674), .ZN(n17692) );
  OAI22_X1 U20811 ( .A1(n17675), .A2(n17692), .B1(n17691), .B2(n17922), .ZN(
        n17687) );
  OAI21_X1 U20812 ( .B1(n17693), .B2(n17676), .A(n18385), .ZN(n17677) );
  OAI221_X1 U20813 ( .B1(n18424), .B2(n17678), .C1(n18424), .C2(n17708), .A(
        n17677), .ZN(n17710) );
  NOR2_X1 U20814 ( .A1(n18384), .A2(n17839), .ZN(n17813) );
  OAI22_X1 U20815 ( .A1(n18424), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17679), .B2(n17813), .ZN(n17680) );
  NOR2_X1 U20816 ( .A1(n17710), .A2(n17680), .ZN(n17699) );
  AOI22_X1 U20817 ( .A1(n18384), .A2(n17682), .B1(n17839), .B2(n17681), .ZN(
        n17696) );
  AOI22_X1 U20818 ( .A1(n18385), .A2(n17695), .B1(n17694), .B2(n17821), .ZN(
        n17685) );
  OAI21_X1 U20819 ( .B1(n17691), .B2(n18409), .A(n17683), .ZN(n17684) );
  NAND4_X1 U20820 ( .A1(n17699), .A2(n17696), .A3(n17685), .A4(n17684), .ZN(
        n17686) );
  AOI22_X1 U20821 ( .A1(n17850), .A2(n17688), .B1(n17687), .B2(n17686), .ZN(
        n17690) );
  OAI211_X1 U20822 ( .C1(n17915), .C2(n17691), .A(n17690), .B(n17689), .ZN(
        P3_U2840) );
  NOR2_X1 U20823 ( .A1(n17693), .A2(n17692), .ZN(n17718) );
  NOR2_X1 U20824 ( .A1(n17932), .A2(n17694), .ZN(n17702) );
  INV_X1 U20825 ( .A(n17695), .ZN(n17700) );
  NAND2_X1 U20826 ( .A1(n17928), .A2(n17696), .ZN(n17746) );
  AOI221_X1 U20827 ( .B1(n17698), .B2(n18409), .C1(n17697), .C2(n18409), .A(
        n17746), .ZN(n17707) );
  OAI211_X1 U20828 ( .C1(n17923), .C2(n17700), .A(n17707), .B(n17699), .ZN(
        n17701) );
  AOI22_X1 U20829 ( .A1(n17703), .A2(n17718), .B1(n17702), .B2(n17701), .ZN(
        n17705) );
  OAI211_X1 U20830 ( .C1(n17706), .C2(n17827), .A(n17705), .B(n17704), .ZN(
        P3_U2841) );
  NAND2_X1 U20831 ( .A1(n17723), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17711) );
  OAI21_X1 U20832 ( .B1(n17708), .B2(n17813), .A(n17707), .ZN(n17709) );
  OAI21_X1 U20833 ( .B1(n17710), .B2(n17709), .A(n17930), .ZN(n17722) );
  OAI21_X1 U20834 ( .B1(n17923), .B2(n17711), .A(n17722), .ZN(n17713) );
  AOI22_X1 U20835 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17713), .B1(
        n17718), .B2(n17712), .ZN(n17715) );
  OAI211_X1 U20836 ( .C1(n17827), .C2(n17716), .A(n17715), .B(n17714), .ZN(
        P3_U2842) );
  INV_X1 U20837 ( .A(n17717), .ZN(n17719) );
  AOI22_X1 U20838 ( .A1(n17850), .A2(n17719), .B1(n17718), .B2(n17723), .ZN(
        n17721) );
  NAND2_X1 U20839 ( .A1(n17932), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17720) );
  OAI211_X1 U20840 ( .C1(n17723), .C2(n17722), .A(n17721), .B(n17720), .ZN(
        P3_U2843) );
  NAND2_X1 U20841 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17724), .ZN(
        n17727) );
  NOR2_X1 U20842 ( .A1(n17725), .A2(n18416), .ZN(n17726) );
  AOI211_X1 U20843 ( .C1(n17903), .C2(n17727), .A(n17726), .B(n17746), .ZN(
        n17728) );
  OAI21_X1 U20844 ( .B1(n17729), .B2(n17813), .A(n17728), .ZN(n17738) );
  INV_X1 U20845 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17739) );
  OAI221_X1 U20846 ( .B1(n17738), .B2(n17739), .C1(n17738), .C2(n17903), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17737) );
  NOR2_X1 U20847 ( .A1(n17914), .A2(n18568), .ZN(n17842) );
  INV_X1 U20848 ( .A(n17900), .ZN(n17730) );
  AOI22_X1 U20849 ( .A1(n18385), .A2(n17899), .B1(n17842), .B2(n17730), .ZN(
        n17856) );
  NOR2_X1 U20850 ( .A1(n17856), .A2(n17731), .ZN(n17838) );
  NAND2_X1 U20851 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17838), .ZN(
        n17753) );
  NAND2_X1 U20852 ( .A1(n17732), .A2(n17753), .ZN(n17795) );
  NAND2_X1 U20853 ( .A1(n17928), .A2(n17795), .ZN(n17837) );
  NOR2_X1 U20854 ( .A1(n17733), .A2(n17837), .ZN(n17748) );
  AOI22_X1 U20855 ( .A1(n17850), .A2(n17735), .B1(n17748), .B2(n17734), .ZN(
        n17736) );
  OAI221_X1 U20856 ( .B1(n17932), .B2(n17737), .C1(n17930), .C2(n18516), .A(
        n17736), .ZN(P3_U2844) );
  OAI221_X1 U20857 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n17930), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17932), .A(n17738), .ZN(
        n17741) );
  NAND3_X1 U20858 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17748), .A3(
        n17739), .ZN(n17740) );
  OAI211_X1 U20859 ( .C1(n17742), .C2(n17827), .A(n17741), .B(n17740), .ZN(
        P3_U2845) );
  AND2_X1 U20860 ( .A1(n18396), .A2(n17769), .ZN(n17832) );
  AND2_X1 U20861 ( .A1(n18385), .A2(n17743), .ZN(n17810) );
  AOI211_X1 U20862 ( .C1(n17770), .C2(n17821), .A(n17832), .B(n17810), .ZN(
        n17744) );
  OAI211_X1 U20863 ( .C1(n17745), .C2(n18422), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17744), .ZN(n17756) );
  OAI221_X1 U20864 ( .B1(n17746), .B2(n17882), .C1(n17746), .C2(n17756), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U20865 ( .A1(n17850), .A2(n17749), .B1(n17748), .B2(n17747), .ZN(
        n17750) );
  OAI221_X1 U20866 ( .B1(n17932), .B2(n17751), .C1(n17930), .C2(n18512), .A(
        n17750), .ZN(P3_U2846) );
  NOR2_X1 U20867 ( .A1(n17752), .A2(n17807), .ZN(n17758) );
  OR2_X1 U20868 ( .A1(n17754), .A2(n17753), .ZN(n17768) );
  OAI21_X1 U20869 ( .B1(n17771), .B2(n17768), .A(n17762), .ZN(n17755) );
  AOI22_X1 U20870 ( .A1(n17758), .A2(n17757), .B1(n17756), .B2(n17755), .ZN(
        n17767) );
  NOR3_X1 U20871 ( .A1(n17760), .A2(n17759), .A3(n17936), .ZN(n17764) );
  OAI21_X1 U20872 ( .B1(n17915), .B2(n17762), .A(n17761), .ZN(n17763) );
  AOI211_X1 U20873 ( .C1(n17765), .C2(n17850), .A(n17764), .B(n17763), .ZN(
        n17766) );
  OAI21_X1 U20874 ( .B1(n17767), .B2(n17922), .A(n17766), .ZN(P3_U2847) );
  AOI22_X1 U20875 ( .A1(n17932), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17924), .ZN(n17780) );
  AND2_X1 U20876 ( .A1(n17771), .A2(n17768), .ZN(n17776) );
  OAI22_X1 U20877 ( .A1(n18396), .A2(n17771), .B1(n17770), .B2(n17769), .ZN(
        n17772) );
  INV_X1 U20878 ( .A(n17830), .ZN(n17811) );
  OAI21_X1 U20879 ( .B1(n17793), .B2(n17811), .A(n18409), .ZN(n17787) );
  OAI211_X1 U20880 ( .C1(n17923), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n17772), .B(n17787), .ZN(n17773) );
  AOI211_X1 U20881 ( .C1(n18385), .C2(n17793), .A(n17810), .B(n17773), .ZN(
        n17775) );
  OAI22_X1 U20882 ( .A1(n17776), .A2(n17775), .B1(n17807), .B2(n17774), .ZN(
        n17778) );
  AOI22_X1 U20883 ( .A1(n17928), .A2(n17778), .B1(n17921), .B2(n17777), .ZN(
        n17779) );
  OAI211_X1 U20884 ( .C1(n17781), .C2(n17827), .A(n17780), .B(n17779), .ZN(
        P3_U2848) );
  AOI22_X1 U20885 ( .A1(n17932), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17850), 
        .B2(n17782), .ZN(n17791) );
  AOI21_X1 U20886 ( .B1(n17783), .B2(n17821), .A(n17832), .ZN(n17815) );
  OAI21_X1 U20887 ( .B1(n17784), .B2(n17807), .A(n17815), .ZN(n17785) );
  AOI211_X1 U20888 ( .C1(n18384), .C2(n17786), .A(n17810), .B(n17785), .ZN(
        n17799) );
  OAI211_X1 U20889 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17788), .A(
        n17799), .B(n17787), .ZN(n17789) );
  OAI211_X1 U20890 ( .C1(n17922), .C2(n17789), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17930), .ZN(n17790) );
  OAI211_X1 U20891 ( .C1(n17792), .C2(n17837), .A(n17791), .B(n17790), .ZN(
        P3_U2849) );
  OAI22_X1 U20892 ( .A1(n18409), .A2(n17794), .B1(n17793), .B2(n17811), .ZN(
        n17798) );
  AOI21_X1 U20893 ( .B1(n17796), .B2(n17795), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17797) );
  AOI211_X1 U20894 ( .C1(n17799), .C2(n17798), .A(n17797), .B(n17922), .ZN(
        n17800) );
  AOI21_X1 U20895 ( .B1(n17924), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17800), .ZN(n17802) );
  OAI211_X1 U20896 ( .C1(n17803), .C2(n17827), .A(n17802), .B(n17801), .ZN(
        P3_U2850) );
  AOI22_X1 U20897 ( .A1(n17932), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17850), 
        .B2(n17804), .ZN(n17818) );
  OAI22_X1 U20898 ( .A1(n17808), .A2(n17807), .B1(n17806), .B2(n17805), .ZN(
        n17809) );
  NOR3_X1 U20899 ( .A1(n17810), .A2(n17922), .A3(n17809), .ZN(n17829) );
  OAI21_X1 U20900 ( .B1(n17836), .B2(n17811), .A(n18409), .ZN(n17812) );
  OAI211_X1 U20901 ( .C1(n17814), .C2(n17813), .A(n17829), .B(n17812), .ZN(
        n17820) );
  OAI21_X1 U20902 ( .B1(n18422), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17815), .ZN(n17816) );
  OAI211_X1 U20903 ( .C1(n17820), .C2(n17816), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17930), .ZN(n17817) );
  OAI211_X1 U20904 ( .C1(n17819), .C2(n17837), .A(n17818), .B(n17817), .ZN(
        P3_U2851) );
  AOI211_X1 U20905 ( .C1(n17836), .C2(n17821), .A(n17832), .B(n17820), .ZN(
        n17823) );
  NOR2_X1 U20906 ( .A1(n17823), .A2(n17822), .ZN(n17825) );
  NOR3_X1 U20907 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17836), .A3(
        n17837), .ZN(n17824) );
  AOI221_X1 U20908 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17932), .C1(n17825), 
        .C2(n17930), .A(n17824), .ZN(n17826) );
  OAI21_X1 U20909 ( .B1(n17828), .B2(n17827), .A(n17826), .ZN(P3_U2852) );
  OAI21_X1 U20910 ( .B1(n18422), .B2(n17830), .A(n17829), .ZN(n17831) );
  OAI21_X1 U20911 ( .B1(n17832), .B2(n17831), .A(n17930), .ZN(n17835) );
  AOI22_X1 U20912 ( .A1(n17932), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17850), 
        .B2(n17833), .ZN(n17834) );
  OAI221_X1 U20913 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17837), .C1(
        n17836), .C2(n17835), .A(n17834), .ZN(P3_U2853) );
  AOI22_X1 U20914 ( .A1(n17840), .A2(n17839), .B1(n17838), .B2(n17846), .ZN(
        n17855) );
  NAND2_X1 U20915 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17845) );
  OAI22_X1 U20916 ( .A1(n17842), .A2(n17841), .B1(n18416), .B2(n17899), .ZN(
        n17843) );
  OAI21_X1 U20917 ( .B1(n17901), .B2(n17843), .A(n17928), .ZN(n17881) );
  OAI21_X1 U20918 ( .B1(n17857), .B2(n17844), .A(n17881), .ZN(n17865) );
  AOI21_X1 U20919 ( .B1(n17917), .B2(n17845), .A(n17865), .ZN(n17860) );
  AOI21_X1 U20920 ( .B1(n17860), .B2(n17915), .A(n17846), .ZN(n17848) );
  AOI211_X1 U20921 ( .C1(n17850), .C2(n17849), .A(n17848), .B(n17847), .ZN(
        n17854) );
  OAI211_X1 U20922 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n17852), .A(
        n17921), .B(n17851), .ZN(n17853) );
  OAI211_X1 U20923 ( .C1(n17855), .C2(n17922), .A(n17854), .B(n17853), .ZN(
        P3_U2854) );
  NOR2_X1 U20924 ( .A1(n17930), .A2(n18494), .ZN(n17862) );
  INV_X1 U20925 ( .A(n17856), .ZN(n17894) );
  AND2_X1 U20926 ( .A1(n17894), .A2(n17857), .ZN(n17871) );
  AOI21_X1 U20927 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17871), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17859) );
  OAI22_X1 U20928 ( .A1(n17860), .A2(n17859), .B1(n17934), .B2(n17858), .ZN(
        n17861) );
  AOI211_X1 U20929 ( .C1(n17924), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17862), .B(n17861), .ZN(n17863) );
  OAI21_X1 U20930 ( .B1(n17936), .B2(n17864), .A(n17863), .ZN(P3_U2855) );
  NOR2_X1 U20931 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17922), .ZN(
        n17870) );
  NOR2_X1 U20932 ( .A1(n17930), .A2(n18492), .ZN(n17869) );
  NOR2_X1 U20933 ( .A1(n17924), .A2(n17865), .ZN(n17876) );
  INV_X1 U20934 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17867) );
  OAI22_X1 U20935 ( .A1(n17876), .A2(n17867), .B1(n17934), .B2(n17866), .ZN(
        n17868) );
  AOI211_X1 U20936 ( .C1(n17871), .C2(n17870), .A(n17869), .B(n17868), .ZN(
        n17872) );
  OAI21_X1 U20937 ( .B1(n17936), .B2(n17873), .A(n17872), .ZN(P3_U2856) );
  NAND3_X1 U20938 ( .A1(n17928), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17894), .ZN(n17890) );
  NOR3_X1 U20939 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17889), .A3(
        n17890), .ZN(n17878) );
  OAI22_X1 U20940 ( .A1(n17876), .A2(n17875), .B1(n17936), .B2(n17874), .ZN(
        n17877) );
  AOI211_X1 U20941 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n17932), .A(n17878), .B(
        n17877), .ZN(n17879) );
  OAI21_X1 U20942 ( .B1(n17934), .B2(n17880), .A(n17879), .ZN(P3_U2857) );
  OAI21_X1 U20943 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17922), .A(
        n17881), .ZN(n17895) );
  AOI21_X1 U20944 ( .B1(n17882), .B2(n17895), .A(n17924), .ZN(n17888) );
  INV_X1 U20945 ( .A(n17883), .ZN(n17886) );
  OAI22_X1 U20946 ( .A1(n17930), .A2(n18488), .B1(n17934), .B2(n17884), .ZN(
        n17885) );
  AOI21_X1 U20947 ( .B1(n17921), .B2(n17886), .A(n17885), .ZN(n17887) );
  OAI221_X1 U20948 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17890), .C1(
        n17889), .C2(n17888), .A(n17887), .ZN(P3_U2858) );
  OAI22_X1 U20949 ( .A1(n17934), .A2(n17892), .B1(n17936), .B2(n17891), .ZN(
        n17893) );
  AOI221_X1 U20950 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17895), .C1(
        n17894), .C2(n17895), .A(n17893), .ZN(n17897) );
  OAI211_X1 U20951 ( .C1(n17915), .C2(n17898), .A(n17897), .B(n17896), .ZN(
        P3_U2859) );
  NOR2_X1 U20952 ( .A1(n18416), .A2(n17899), .ZN(n17911) );
  NOR2_X1 U20953 ( .A1(n18568), .A2(n17900), .ZN(n17906) );
  NOR3_X1 U20954 ( .A1(n18416), .A2(n18583), .A3(n18568), .ZN(n17902) );
  AOI211_X1 U20955 ( .C1(n18568), .C2(n17903), .A(n17902), .B(n17901), .ZN(
        n17904) );
  INV_X1 U20956 ( .A(n17904), .ZN(n17905) );
  MUX2_X1 U20957 ( .A(n17906), .B(n17905), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n17910) );
  OAI22_X1 U20958 ( .A1(n17934), .A2(n17908), .B1(n17936), .B2(n17907), .ZN(
        n17909) );
  AOI221_X1 U20959 ( .B1(n17911), .B2(n17928), .C1(n17910), .C2(n17928), .A(
        n17909), .ZN(n17913) );
  OAI211_X1 U20960 ( .C1(n17915), .C2(n17914), .A(n17913), .B(n17912), .ZN(
        P3_U2860) );
  NOR2_X1 U20961 ( .A1(n17930), .A2(n18588), .ZN(n17919) );
  AND3_X1 U20962 ( .A1(n17917), .A2(n18568), .A3(n17916), .ZN(n17918) );
  AOI211_X1 U20963 ( .C1(n17921), .C2(n17920), .A(n17919), .B(n17918), .ZN(
        n17926) );
  NOR3_X1 U20964 ( .A1(n17923), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n17922), .ZN(n17929) );
  OAI21_X1 U20965 ( .B1(n17924), .B2(n17929), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17925) );
  OAI211_X1 U20966 ( .C1(n17927), .C2(n17934), .A(n17926), .B(n17925), .ZN(
        P3_U2861) );
  AOI21_X1 U20967 ( .B1(n18424), .B2(n17928), .A(n18583), .ZN(n17931) );
  AOI221_X1 U20968 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n17932), .C1(n17931), 
        .C2(n17930), .A(n17929), .ZN(n17933) );
  OAI221_X1 U20969 ( .B1(n17937), .B2(n17936), .C1(n17935), .C2(n17934), .A(
        n17933), .ZN(P3_U2862) );
  INV_X1 U20970 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18234) );
  AOI211_X1 U20971 ( .C1(n17939), .C2(n17938), .A(n18566), .B(n18617), .ZN(
        n18447) );
  OAI21_X1 U20972 ( .B1(n18447), .B2(n17993), .A(n17948), .ZN(n17940) );
  OAI221_X1 U20973 ( .B1(n18234), .B2(n18602), .C1(n18234), .C2(n17948), .A(
        n17940), .ZN(P3_U2863) );
  NAND2_X1 U20974 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18165) );
  AOI221_X1 U20975 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18165), .C1(n17942), 
        .C2(n18165), .A(n17941), .ZN(n17947) );
  NOR2_X1 U20976 ( .A1(n17943), .A2(n18428), .ZN(n17944) );
  OAI21_X1 U20977 ( .B1(n17944), .B2(n18191), .A(n17948), .ZN(n17945) );
  AOI22_X1 U20978 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17947), .B1(
        n17945), .B2(n18433), .ZN(P3_U2865) );
  INV_X1 U20979 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18436) );
  NAND2_X1 U20980 ( .A1(n18436), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18123) );
  NAND2_X1 U20981 ( .A1(n18191), .A2(n18213), .ZN(n18235) );
  AND2_X1 U20982 ( .A1(n18123), .A2(n18235), .ZN(n17946) );
  OAI22_X1 U20983 ( .A1(n17947), .A2(n18436), .B1(n17946), .B2(n17945), .ZN(
        P3_U2866) );
  NOR2_X1 U20984 ( .A1(n18437), .A2(n17948), .ZN(P3_U2867) );
  NOR2_X1 U20985 ( .A1(n18433), .A2(n18436), .ZN(n18259) );
  INV_X1 U20986 ( .A(n18259), .ZN(n17951) );
  NOR2_X1 U20987 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17951), .ZN(
        n18328) );
  NAND2_X1 U20988 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18328), .ZN(
        n18382) );
  NAND2_X1 U20989 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18329), .ZN(n18264) );
  NOR2_X2 U20990 ( .A1(n17980), .A2(n17949), .ZN(n18330) );
  NOR2_X1 U20991 ( .A1(n18428), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18099) );
  NAND2_X1 U20992 ( .A1(n18099), .A2(n18259), .ZN(n18293) );
  NOR2_X2 U20993 ( .A1(n18147), .A2(n17950), .ZN(n18324) );
  INV_X1 U20994 ( .A(n18323), .ZN(n18456) );
  NAND2_X1 U20995 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18427) );
  NOR2_X2 U20996 ( .A1(n18427), .A2(n17951), .ZN(n18377) );
  NOR2_X1 U20997 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18144) );
  NOR2_X1 U20998 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18033) );
  NAND2_X1 U20999 ( .A1(n18144), .A2(n18033), .ZN(n18053) );
  NAND2_X1 U21000 ( .A1(n18334), .A2(n18053), .ZN(n17952) );
  INV_X1 U21001 ( .A(n17952), .ZN(n18012) );
  NOR2_X1 U21002 ( .A1(n18456), .A2(n18012), .ZN(n17987) );
  AOI22_X1 U21003 ( .A1(n18330), .A2(n18317), .B1(n18324), .B2(n17987), .ZN(
        n17957) );
  NOR2_X1 U21004 ( .A1(n18234), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18168) );
  NOR2_X1 U21005 ( .A1(n18168), .A2(n18099), .ZN(n18236) );
  NOR2_X1 U21006 ( .A1(n18236), .A2(n17951), .ZN(n18285) );
  AOI21_X1 U21007 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18147), .ZN(n18189) );
  AOI22_X1 U21008 ( .A1(n18329), .A2(n18285), .B1(n18189), .B2(n17952), .ZN(
        n17990) );
  NOR2_X1 U21009 ( .A1(n17954), .A2(n17953), .ZN(n17959) );
  NAND2_X1 U21010 ( .A1(n17955), .A2(n17959), .ZN(n18333) );
  INV_X1 U21011 ( .A(n18333), .ZN(n18261) );
  AOI22_X1 U21012 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17990), .B1(
        n18046), .B2(n18261), .ZN(n17956) );
  OAI211_X1 U21013 ( .C1(n18382), .C2(n18264), .A(n17957), .B(n17956), .ZN(
        P3_U2868) );
  NAND2_X1 U21014 ( .A1(n18329), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18297) );
  INV_X1 U21015 ( .A(n18382), .ZN(n18360) );
  NAND2_X1 U21016 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18329), .ZN(n18340) );
  INV_X1 U21017 ( .A(n18340), .ZN(n18294) );
  NOR2_X2 U21018 ( .A1(n18147), .A2(n17958), .ZN(n18335) );
  AOI22_X1 U21019 ( .A1(n18360), .A2(n18294), .B1(n17987), .B2(n18335), .ZN(
        n17962) );
  INV_X1 U21020 ( .A(n17959), .ZN(n17988) );
  NOR2_X2 U21021 ( .A1(n17960), .A2(n17988), .ZN(n18337) );
  AOI22_X1 U21022 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17990), .B1(
        n18046), .B2(n18337), .ZN(n17961) );
  OAI211_X1 U21023 ( .C1(n18293), .C2(n18297), .A(n17962), .B(n17961), .ZN(
        P3_U2869) );
  NOR2_X1 U21024 ( .A1(n17963), .A2(n17980), .ZN(n18267) );
  INV_X1 U21025 ( .A(n18267), .ZN(n18346) );
  NAND2_X1 U21026 ( .A1(n18329), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18270) );
  INV_X1 U21027 ( .A(n18270), .ZN(n18342) );
  NOR2_X2 U21028 ( .A1(n18147), .A2(n17964), .ZN(n18341) );
  AOI22_X1 U21029 ( .A1(n18317), .A2(n18342), .B1(n17987), .B2(n18341), .ZN(
        n17967) );
  NOR2_X2 U21030 ( .A1(n17965), .A2(n17988), .ZN(n18343) );
  AOI22_X1 U21031 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n17990), .B1(
        n18046), .B2(n18343), .ZN(n17966) );
  OAI211_X1 U21032 ( .C1(n18382), .C2(n18346), .A(n17967), .B(n17966), .ZN(
        P3_U2870) );
  NOR2_X1 U21033 ( .A1(n17980), .A2(n14142), .ZN(n18348) );
  INV_X1 U21034 ( .A(n18348), .ZN(n18303) );
  NAND2_X1 U21035 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18329), .ZN(n18352) );
  INV_X1 U21036 ( .A(n18352), .ZN(n18300) );
  NOR2_X2 U21037 ( .A1(n18147), .A2(n17968), .ZN(n18347) );
  AOI22_X1 U21038 ( .A1(n18360), .A2(n18300), .B1(n17987), .B2(n18347), .ZN(
        n17971) );
  NOR2_X2 U21039 ( .A1(n17969), .A2(n17988), .ZN(n18349) );
  AOI22_X1 U21040 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n17990), .B1(
        n18046), .B2(n18349), .ZN(n17970) );
  OAI211_X1 U21041 ( .C1(n18293), .C2(n18303), .A(n17971), .B(n17970), .ZN(
        P3_U2871) );
  NAND2_X1 U21042 ( .A1(n18329), .A2(BUF2_REG_20__SCAN_IN), .ZN(n20812) );
  NAND2_X1 U21043 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18329), .ZN(n18357) );
  INV_X1 U21044 ( .A(n18357), .ZN(n20809) );
  NOR2_X2 U21045 ( .A1(n18147), .A2(n17972), .ZN(n20806) );
  AOI22_X1 U21046 ( .A1(n20809), .A2(n18360), .B1(n20806), .B2(n17987), .ZN(
        n17975) );
  NOR2_X2 U21047 ( .A1(n17988), .A2(n17973), .ZN(n18354) );
  AOI22_X1 U21048 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n17990), .B1(
        n18354), .B2(n18046), .ZN(n17974) );
  OAI211_X1 U21049 ( .C1(n20812), .C2(n18293), .A(n17975), .B(n17974), .ZN(
        P3_U2872) );
  NAND2_X1 U21050 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18329), .ZN(n18365) );
  NAND2_X1 U21051 ( .A1(n18329), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18310) );
  INV_X1 U21052 ( .A(n18310), .ZN(n18359) );
  NOR2_X2 U21053 ( .A1(n18147), .A2(n17976), .ZN(n18358) );
  AOI22_X1 U21054 ( .A1(n18317), .A2(n18359), .B1(n17987), .B2(n18358), .ZN(
        n17979) );
  NOR2_X2 U21055 ( .A1(n17977), .A2(n17988), .ZN(n18361) );
  AOI22_X1 U21056 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n17990), .B1(
        n18046), .B2(n18361), .ZN(n17978) );
  OAI211_X1 U21057 ( .C1(n18382), .C2(n18365), .A(n17979), .B(n17978), .ZN(
        P3_U2873) );
  NOR2_X1 U21058 ( .A1(n17981), .A2(n17980), .ZN(n18367) );
  INV_X1 U21059 ( .A(n18367), .ZN(n18314) );
  NAND2_X1 U21060 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18329), .ZN(n18371) );
  INV_X1 U21061 ( .A(n18371), .ZN(n18311) );
  NOR2_X2 U21062 ( .A1(n17982), .A2(n18147), .ZN(n18366) );
  AOI22_X1 U21063 ( .A1(n18317), .A2(n18311), .B1(n17987), .B2(n18366), .ZN(
        n17985) );
  NOR2_X2 U21064 ( .A1(n17983), .A2(n17988), .ZN(n18368) );
  AOI22_X1 U21065 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17990), .B1(
        n18046), .B2(n18368), .ZN(n17984) );
  OAI211_X1 U21066 ( .C1(n18382), .C2(n18314), .A(n17985), .B(n17984), .ZN(
        P3_U2874) );
  NAND2_X1 U21067 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18329), .ZN(n18381) );
  NAND2_X1 U21068 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18329), .ZN(n18322) );
  INV_X1 U21069 ( .A(n18322), .ZN(n18375) );
  NOR2_X2 U21070 ( .A1(n17986), .A2(n18147), .ZN(n18373) );
  AOI22_X1 U21071 ( .A1(n18360), .A2(n18375), .B1(n17987), .B2(n18373), .ZN(
        n17992) );
  NOR2_X2 U21072 ( .A1(n17989), .A2(n17988), .ZN(n18376) );
  AOI22_X1 U21073 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17990), .B1(
        n18046), .B2(n18376), .ZN(n17991) );
  OAI211_X1 U21074 ( .C1(n18293), .C2(n18381), .A(n17992), .B(n17991), .ZN(
        P3_U2875) );
  INV_X1 U21075 ( .A(n18033), .ZN(n18077) );
  NAND2_X1 U21076 ( .A1(n18428), .A2(n18323), .ZN(n18164) );
  NOR2_X1 U21077 ( .A1(n18077), .A2(n18164), .ZN(n18008) );
  AOI22_X1 U21078 ( .A1(n18377), .A2(n18330), .B1(n18324), .B2(n18008), .ZN(
        n17995) );
  NOR2_X1 U21079 ( .A1(n18436), .A2(n18165), .ZN(n18326) );
  NOR2_X1 U21080 ( .A1(n18147), .A2(n17993), .ZN(n18327) );
  INV_X1 U21081 ( .A(n18327), .ZN(n18032) );
  NOR2_X1 U21082 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18032), .ZN(
        n18258) );
  AOI22_X1 U21083 ( .A1(n18329), .A2(n18326), .B1(n18033), .B2(n18258), .ZN(
        n18009) );
  NAND2_X1 U21084 ( .A1(n18168), .A2(n18033), .ZN(n18075) );
  AOI22_X1 U21085 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18009), .B1(
        n18261), .B2(n18068), .ZN(n17994) );
  OAI211_X1 U21086 ( .C1(n18264), .C2(n18293), .A(n17995), .B(n17994), .ZN(
        P3_U2876) );
  INV_X1 U21087 ( .A(n18297), .ZN(n18336) );
  AOI22_X1 U21088 ( .A1(n18377), .A2(n18336), .B1(n18335), .B2(n18008), .ZN(
        n17997) );
  AOI22_X1 U21089 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18009), .B1(
        n18337), .B2(n18068), .ZN(n17996) );
  OAI211_X1 U21090 ( .C1(n18293), .C2(n18340), .A(n17997), .B(n17996), .ZN(
        P3_U2877) );
  AOI22_X1 U21091 ( .A1(n18317), .A2(n18267), .B1(n18341), .B2(n18008), .ZN(
        n17999) );
  AOI22_X1 U21092 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18009), .B1(
        n18343), .B2(n18068), .ZN(n17998) );
  OAI211_X1 U21093 ( .C1(n18334), .C2(n18270), .A(n17999), .B(n17998), .ZN(
        P3_U2878) );
  AOI22_X1 U21094 ( .A1(n18377), .A2(n18348), .B1(n18347), .B2(n18008), .ZN(
        n18001) );
  AOI22_X1 U21095 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18009), .B1(
        n18349), .B2(n18068), .ZN(n18000) );
  OAI211_X1 U21096 ( .C1(n18293), .C2(n18352), .A(n18001), .B(n18000), .ZN(
        P3_U2879) );
  AOI22_X1 U21097 ( .A1(n18353), .A2(n18377), .B1(n20806), .B2(n18008), .ZN(
        n18003) );
  AOI22_X1 U21098 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18009), .B1(
        n18354), .B2(n18068), .ZN(n18002) );
  OAI211_X1 U21099 ( .C1(n18357), .C2(n18293), .A(n18003), .B(n18002), .ZN(
        P3_U2880) );
  AOI22_X1 U21100 ( .A1(n18377), .A2(n18359), .B1(n18358), .B2(n18008), .ZN(
        n18005) );
  AOI22_X1 U21101 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18009), .B1(
        n18361), .B2(n18068), .ZN(n18004) );
  OAI211_X1 U21102 ( .C1(n18293), .C2(n18365), .A(n18005), .B(n18004), .ZN(
        P3_U2881) );
  AOI22_X1 U21103 ( .A1(n18317), .A2(n18367), .B1(n18366), .B2(n18008), .ZN(
        n18007) );
  AOI22_X1 U21104 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18009), .B1(
        n18368), .B2(n18068), .ZN(n18006) );
  OAI211_X1 U21105 ( .C1(n18334), .C2(n18371), .A(n18007), .B(n18006), .ZN(
        P3_U2882) );
  AOI22_X1 U21106 ( .A1(n18317), .A2(n18375), .B1(n18373), .B2(n18008), .ZN(
        n18011) );
  AOI22_X1 U21107 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18009), .B1(
        n18376), .B2(n18068), .ZN(n18010) );
  OAI211_X1 U21108 ( .C1(n18334), .C2(n18381), .A(n18011), .B(n18010), .ZN(
        P3_U2883) );
  NAND2_X1 U21109 ( .A1(n18099), .A2(n18033), .ZN(n18098) );
  NOR2_X1 U21110 ( .A1(n18068), .A2(n18087), .ZN(n18054) );
  NOR2_X1 U21111 ( .A1(n18456), .A2(n18054), .ZN(n18028) );
  AOI22_X1 U21112 ( .A1(n18046), .A2(n18330), .B1(n18324), .B2(n18028), .ZN(
        n18015) );
  OAI21_X1 U21113 ( .B1(n18012), .B2(n18287), .A(n18054), .ZN(n18013) );
  OAI211_X1 U21114 ( .C1(n18087), .C2(n18555), .A(n18290), .B(n18013), .ZN(
        n18029) );
  AOI22_X1 U21115 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18029), .B1(
        n18261), .B2(n18087), .ZN(n18014) );
  OAI211_X1 U21116 ( .C1(n18264), .C2(n18334), .A(n18015), .B(n18014), .ZN(
        P3_U2884) );
  AOI22_X1 U21117 ( .A1(n18377), .A2(n18294), .B1(n18335), .B2(n18028), .ZN(
        n18017) );
  AOI22_X1 U21118 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18029), .B1(
        n18337), .B2(n18087), .ZN(n18016) );
  OAI211_X1 U21119 ( .C1(n18053), .C2(n18297), .A(n18017), .B(n18016), .ZN(
        P3_U2885) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18029), .B1(
        n18341), .B2(n18028), .ZN(n18019) );
  AOI22_X1 U21121 ( .A1(n18377), .A2(n18267), .B1(n18343), .B2(n18087), .ZN(
        n18018) );
  OAI211_X1 U21122 ( .C1(n18053), .C2(n18270), .A(n18019), .B(n18018), .ZN(
        P3_U2886) );
  AOI22_X1 U21123 ( .A1(n18377), .A2(n18300), .B1(n18347), .B2(n18028), .ZN(
        n18021) );
  AOI22_X1 U21124 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18029), .B1(
        n18349), .B2(n18087), .ZN(n18020) );
  OAI211_X1 U21125 ( .C1(n18053), .C2(n18303), .A(n18021), .B(n18020), .ZN(
        P3_U2887) );
  AOI22_X1 U21126 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18029), .B1(
        n20806), .B2(n18028), .ZN(n18023) );
  AOI22_X1 U21127 ( .A1(n18353), .A2(n18046), .B1(n18354), .B2(n18087), .ZN(
        n18022) );
  OAI211_X1 U21128 ( .C1(n18357), .C2(n18334), .A(n18023), .B(n18022), .ZN(
        P3_U2888) );
  AOI22_X1 U21129 ( .A1(n18046), .A2(n18359), .B1(n18358), .B2(n18028), .ZN(
        n18025) );
  AOI22_X1 U21130 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18029), .B1(
        n18361), .B2(n18087), .ZN(n18024) );
  OAI211_X1 U21131 ( .C1(n18334), .C2(n18365), .A(n18025), .B(n18024), .ZN(
        P3_U2889) );
  AOI22_X1 U21132 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18029), .B1(
        n18366), .B2(n18028), .ZN(n18027) );
  AOI22_X1 U21133 ( .A1(n18377), .A2(n18367), .B1(n18368), .B2(n18087), .ZN(
        n18026) );
  OAI211_X1 U21134 ( .C1(n18053), .C2(n18371), .A(n18027), .B(n18026), .ZN(
        P3_U2890) );
  AOI22_X1 U21135 ( .A1(n18377), .A2(n18375), .B1(n18373), .B2(n18028), .ZN(
        n18031) );
  AOI22_X1 U21136 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18029), .B1(
        n18376), .B2(n18087), .ZN(n18030) );
  OAI211_X1 U21137 ( .C1(n18053), .C2(n18381), .A(n18031), .B(n18030), .ZN(
        P3_U2891) );
  NOR2_X2 U21138 ( .A1(n18427), .A2(n18077), .ZN(n18111) );
  INV_X1 U21139 ( .A(n18264), .ZN(n18325) );
  AOI22_X1 U21140 ( .A1(n18325), .A2(n18046), .B1(n18324), .B2(n18049), .ZN(
        n18035) );
  AOI21_X1 U21141 ( .B1(n18428), .B2(n18287), .A(n18032), .ZN(n18121) );
  NAND2_X1 U21142 ( .A1(n18033), .A2(n18121), .ZN(n18050) );
  AOI22_X1 U21143 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18050), .B1(
        n18330), .B2(n18068), .ZN(n18034) );
  OAI211_X1 U21144 ( .C1(n18333), .C2(n18120), .A(n18035), .B(n18034), .ZN(
        P3_U2892) );
  AOI22_X1 U21145 ( .A1(n18336), .A2(n18068), .B1(n18335), .B2(n18049), .ZN(
        n18037) );
  AOI22_X1 U21146 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18050), .B1(
        n18337), .B2(n18111), .ZN(n18036) );
  OAI211_X1 U21147 ( .C1(n18053), .C2(n18340), .A(n18037), .B(n18036), .ZN(
        P3_U2893) );
  AOI22_X1 U21148 ( .A1(n18342), .A2(n18068), .B1(n18341), .B2(n18049), .ZN(
        n18039) );
  AOI22_X1 U21149 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18050), .B1(
        n18343), .B2(n18111), .ZN(n18038) );
  OAI211_X1 U21150 ( .C1(n18053), .C2(n18346), .A(n18039), .B(n18038), .ZN(
        P3_U2894) );
  AOI22_X1 U21151 ( .A1(n18348), .A2(n18068), .B1(n18347), .B2(n18049), .ZN(
        n18041) );
  AOI22_X1 U21152 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18050), .B1(
        n18349), .B2(n18111), .ZN(n18040) );
  OAI211_X1 U21153 ( .C1(n18053), .C2(n18352), .A(n18041), .B(n18040), .ZN(
        P3_U2895) );
  INV_X1 U21154 ( .A(n18354), .ZN(n20813) );
  AOI22_X1 U21155 ( .A1(n20809), .A2(n18046), .B1(n20806), .B2(n18049), .ZN(
        n18043) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18050), .B1(
        n18353), .B2(n18068), .ZN(n18042) );
  OAI211_X1 U21157 ( .C1(n20813), .C2(n18120), .A(n18043), .B(n18042), .ZN(
        P3_U2896) );
  AOI22_X1 U21158 ( .A1(n18359), .A2(n18068), .B1(n18358), .B2(n18049), .ZN(
        n18045) );
  AOI22_X1 U21159 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18050), .B1(
        n18361), .B2(n18111), .ZN(n18044) );
  OAI211_X1 U21160 ( .C1(n18053), .C2(n18365), .A(n18045), .B(n18044), .ZN(
        P3_U2897) );
  AOI22_X1 U21161 ( .A1(n18046), .A2(n18367), .B1(n18366), .B2(n18049), .ZN(
        n18048) );
  AOI22_X1 U21162 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18050), .B1(
        n18368), .B2(n18111), .ZN(n18047) );
  OAI211_X1 U21163 ( .C1(n18371), .C2(n18075), .A(n18048), .B(n18047), .ZN(
        P3_U2898) );
  INV_X1 U21164 ( .A(n18381), .ZN(n18316) );
  AOI22_X1 U21165 ( .A1(n18316), .A2(n18068), .B1(n18373), .B2(n18049), .ZN(
        n18052) );
  AOI22_X1 U21166 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18050), .B1(
        n18376), .B2(n18111), .ZN(n18051) );
  OAI211_X1 U21167 ( .C1(n18053), .C2(n18322), .A(n18052), .B(n18051), .ZN(
        P3_U2899) );
  INV_X1 U21168 ( .A(n18144), .ZN(n18429) );
  NOR2_X2 U21169 ( .A1(n18429), .A2(n18123), .ZN(n18140) );
  AOI21_X1 U21170 ( .B1(n18120), .B2(n18136), .A(n18456), .ZN(n18071) );
  AOI22_X1 U21171 ( .A1(n18325), .A2(n18068), .B1(n18324), .B2(n18071), .ZN(
        n18057) );
  AOI221_X1 U21172 ( .B1(n18054), .B2(n18120), .C1(n18287), .C2(n18120), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18055) );
  OAI21_X1 U21173 ( .B1(n18140), .B2(n18055), .A(n18290), .ZN(n18072) );
  AOI22_X1 U21174 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18072), .B1(
        n18330), .B2(n18087), .ZN(n18056) );
  OAI211_X1 U21175 ( .C1(n18333), .C2(n18136), .A(n18057), .B(n18056), .ZN(
        P3_U2900) );
  AOI22_X1 U21176 ( .A1(n18294), .A2(n18068), .B1(n18335), .B2(n18071), .ZN(
        n18059) );
  AOI22_X1 U21177 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18072), .B1(
        n18337), .B2(n18140), .ZN(n18058) );
  OAI211_X1 U21178 ( .C1(n18297), .C2(n18098), .A(n18059), .B(n18058), .ZN(
        P3_U2901) );
  AOI22_X1 U21179 ( .A1(n18342), .A2(n18087), .B1(n18341), .B2(n18071), .ZN(
        n18061) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18072), .B1(
        n18343), .B2(n18140), .ZN(n18060) );
  OAI211_X1 U21181 ( .C1(n18346), .C2(n18075), .A(n18061), .B(n18060), .ZN(
        P3_U2902) );
  AOI22_X1 U21182 ( .A1(n18348), .A2(n18087), .B1(n18347), .B2(n18071), .ZN(
        n18063) );
  AOI22_X1 U21183 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18072), .B1(
        n18349), .B2(n18140), .ZN(n18062) );
  OAI211_X1 U21184 ( .C1(n18352), .C2(n18075), .A(n18063), .B(n18062), .ZN(
        P3_U2903) );
  AOI22_X1 U21185 ( .A1(n18353), .A2(n18087), .B1(n20806), .B2(n18071), .ZN(
        n18065) );
  AOI22_X1 U21186 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18072), .B1(
        n18354), .B2(n18140), .ZN(n18064) );
  OAI211_X1 U21187 ( .C1(n18357), .C2(n18075), .A(n18065), .B(n18064), .ZN(
        P3_U2904) );
  AOI22_X1 U21188 ( .A1(n18359), .A2(n18087), .B1(n18358), .B2(n18071), .ZN(
        n18067) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18072), .B1(
        n18361), .B2(n18140), .ZN(n18066) );
  OAI211_X1 U21190 ( .C1(n18365), .C2(n18075), .A(n18067), .B(n18066), .ZN(
        P3_U2905) );
  AOI22_X1 U21191 ( .A1(n18367), .A2(n18068), .B1(n18366), .B2(n18071), .ZN(
        n18070) );
  AOI22_X1 U21192 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18072), .B1(
        n18368), .B2(n18140), .ZN(n18069) );
  OAI211_X1 U21193 ( .C1(n18371), .C2(n18098), .A(n18070), .B(n18069), .ZN(
        P3_U2906) );
  AOI22_X1 U21194 ( .A1(n18316), .A2(n18087), .B1(n18373), .B2(n18071), .ZN(
        n18074) );
  AOI22_X1 U21195 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18072), .B1(
        n18376), .B2(n18140), .ZN(n18073) );
  OAI211_X1 U21196 ( .C1(n18322), .C2(n18075), .A(n18074), .B(n18073), .ZN(
        P3_U2907) );
  INV_X1 U21197 ( .A(n18168), .ZN(n18076) );
  NOR2_X2 U21198 ( .A1(n18123), .A2(n18076), .ZN(n20808) );
  NOR2_X1 U21199 ( .A1(n18123), .A2(n18164), .ZN(n18094) );
  AOI22_X1 U21200 ( .A1(n18330), .A2(n18111), .B1(n18324), .B2(n18094), .ZN(
        n18080) );
  NOR2_X1 U21201 ( .A1(n18428), .A2(n18077), .ZN(n18078) );
  INV_X1 U21202 ( .A(n18123), .ZN(n18122) );
  AOI22_X1 U21203 ( .A1(n18329), .A2(n18078), .B1(n18122), .B2(n18258), .ZN(
        n18095) );
  AOI22_X1 U21204 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18095), .B1(
        n18325), .B2(n18087), .ZN(n18079) );
  OAI211_X1 U21205 ( .C1(n18163), .C2(n18333), .A(n18080), .B(n18079), .ZN(
        P3_U2908) );
  AOI22_X1 U21206 ( .A1(n18336), .A2(n18111), .B1(n18335), .B2(n18094), .ZN(
        n18082) );
  AOI22_X1 U21207 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18095), .B1(
        n20808), .B2(n18337), .ZN(n18081) );
  OAI211_X1 U21208 ( .C1(n18340), .C2(n18098), .A(n18082), .B(n18081), .ZN(
        P3_U2909) );
  AOI22_X1 U21209 ( .A1(n18267), .A2(n18087), .B1(n18341), .B2(n18094), .ZN(
        n18084) );
  AOI22_X1 U21210 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18095), .B1(
        n20808), .B2(n18343), .ZN(n18083) );
  OAI211_X1 U21211 ( .C1(n18270), .C2(n18120), .A(n18084), .B(n18083), .ZN(
        P3_U2910) );
  AOI22_X1 U21212 ( .A1(n18348), .A2(n18111), .B1(n18347), .B2(n18094), .ZN(
        n18086) );
  AOI22_X1 U21213 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18095), .B1(
        n20808), .B2(n18349), .ZN(n18085) );
  OAI211_X1 U21214 ( .C1(n18352), .C2(n18098), .A(n18086), .B(n18085), .ZN(
        P3_U2911) );
  AOI22_X1 U21215 ( .A1(n20809), .A2(n18087), .B1(n20806), .B2(n18094), .ZN(
        n18089) );
  AOI22_X1 U21216 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18095), .B1(
        n18354), .B2(n20808), .ZN(n18088) );
  OAI211_X1 U21217 ( .C1(n20812), .C2(n18120), .A(n18089), .B(n18088), .ZN(
        P3_U2912) );
  AOI22_X1 U21218 ( .A1(n18359), .A2(n18111), .B1(n18358), .B2(n18094), .ZN(
        n18091) );
  AOI22_X1 U21219 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18095), .B1(
        n20808), .B2(n18361), .ZN(n18090) );
  OAI211_X1 U21220 ( .C1(n18365), .C2(n18098), .A(n18091), .B(n18090), .ZN(
        P3_U2913) );
  AOI22_X1 U21221 ( .A1(n18366), .A2(n18094), .B1(n18311), .B2(n18111), .ZN(
        n18093) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18095), .B1(
        n20808), .B2(n18368), .ZN(n18092) );
  OAI211_X1 U21223 ( .C1(n18314), .C2(n18098), .A(n18093), .B(n18092), .ZN(
        P3_U2914) );
  AOI22_X1 U21224 ( .A1(n18316), .A2(n18111), .B1(n18373), .B2(n18094), .ZN(
        n18097) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18095), .B1(
        n20808), .B2(n18376), .ZN(n18096) );
  OAI211_X1 U21226 ( .C1(n18322), .C2(n18098), .A(n18097), .B(n18096), .ZN(
        P3_U2915) );
  INV_X1 U21227 ( .A(n18099), .ZN(n18188) );
  NOR2_X2 U21228 ( .A1(n18123), .A2(n18188), .ZN(n18179) );
  NOR2_X1 U21229 ( .A1(n18123), .A2(n18236), .ZN(n18145) );
  AND2_X1 U21230 ( .A1(n18323), .A2(n18145), .ZN(n18116) );
  AOI22_X1 U21231 ( .A1(n18330), .A2(n18140), .B1(n18324), .B2(n18116), .ZN(
        n18102) );
  NAND2_X1 U21232 ( .A1(n18120), .A2(n18136), .ZN(n18100) );
  OAI221_X1 U21233 ( .B1(n18145), .B2(n18191), .C1(n18145), .C2(n18100), .A(
        n18189), .ZN(n18117) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18117), .B1(
        n18325), .B2(n18111), .ZN(n18101) );
  OAI211_X1 U21235 ( .C1(n20811), .C2(n18333), .A(n18102), .B(n18101), .ZN(
        P3_U2916) );
  AOI22_X1 U21236 ( .A1(n18336), .A2(n18140), .B1(n18335), .B2(n18116), .ZN(
        n18104) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18117), .B1(
        n18179), .B2(n18337), .ZN(n18103) );
  OAI211_X1 U21238 ( .C1(n18340), .C2(n18120), .A(n18104), .B(n18103), .ZN(
        P3_U2917) );
  AOI22_X1 U21239 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18117), .B1(
        n18341), .B2(n18116), .ZN(n18106) );
  AOI22_X1 U21240 ( .A1(n18179), .A2(n18343), .B1(n18267), .B2(n18111), .ZN(
        n18105) );
  OAI211_X1 U21241 ( .C1(n18270), .C2(n18136), .A(n18106), .B(n18105), .ZN(
        P3_U2918) );
  AOI22_X1 U21242 ( .A1(n18348), .A2(n18140), .B1(n18347), .B2(n18116), .ZN(
        n18108) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18117), .B1(
        n18179), .B2(n18349), .ZN(n18107) );
  OAI211_X1 U21244 ( .C1(n18352), .C2(n18120), .A(n18108), .B(n18107), .ZN(
        P3_U2919) );
  AOI22_X1 U21245 ( .A1(n18353), .A2(n18140), .B1(n20806), .B2(n18116), .ZN(
        n18110) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18117), .B1(
        n18179), .B2(n18354), .ZN(n18109) );
  OAI211_X1 U21247 ( .C1(n18357), .C2(n18120), .A(n18110), .B(n18109), .ZN(
        P3_U2920) );
  INV_X1 U21248 ( .A(n18365), .ZN(n18307) );
  AOI22_X1 U21249 ( .A1(n18307), .A2(n18111), .B1(n18358), .B2(n18116), .ZN(
        n18113) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18117), .B1(
        n18179), .B2(n18361), .ZN(n18112) );
  OAI211_X1 U21251 ( .C1(n18310), .C2(n18136), .A(n18113), .B(n18112), .ZN(
        P3_U2921) );
  AOI22_X1 U21252 ( .A1(n18366), .A2(n18116), .B1(n18311), .B2(n18140), .ZN(
        n18115) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18117), .B1(
        n18179), .B2(n18368), .ZN(n18114) );
  OAI211_X1 U21254 ( .C1(n18314), .C2(n18120), .A(n18115), .B(n18114), .ZN(
        P3_U2922) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18117), .B1(
        n18373), .B2(n18116), .ZN(n18119) );
  AOI22_X1 U21256 ( .A1(n18179), .A2(n18376), .B1(n18316), .B2(n18140), .ZN(
        n18118) );
  OAI211_X1 U21257 ( .C1(n18322), .C2(n18120), .A(n18119), .B(n18118), .ZN(
        P3_U2923) );
  AOI22_X1 U21258 ( .A1(n20808), .A2(n18330), .B1(n18324), .B2(n18139), .ZN(
        n18125) );
  NAND2_X1 U21259 ( .A1(n18122), .A2(n18121), .ZN(n18141) );
  NOR2_X2 U21260 ( .A1(n18427), .A2(n18123), .ZN(n18205) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18141), .B1(
        n18205), .B2(n18261), .ZN(n18124) );
  OAI211_X1 U21262 ( .C1(n18264), .C2(n18136), .A(n18125), .B(n18124), .ZN(
        P3_U2924) );
  AOI22_X1 U21263 ( .A1(n18294), .A2(n18140), .B1(n18335), .B2(n18139), .ZN(
        n18127) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18141), .B1(
        n18205), .B2(n18337), .ZN(n18126) );
  OAI211_X1 U21265 ( .C1(n18163), .C2(n18297), .A(n18127), .B(n18126), .ZN(
        P3_U2925) );
  AOI22_X1 U21266 ( .A1(n20808), .A2(n18342), .B1(n18341), .B2(n18139), .ZN(
        n18129) );
  AOI22_X1 U21267 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18141), .B1(
        n18205), .B2(n18343), .ZN(n18128) );
  OAI211_X1 U21268 ( .C1(n18346), .C2(n18136), .A(n18129), .B(n18128), .ZN(
        P3_U2926) );
  AOI22_X1 U21269 ( .A1(n18300), .A2(n18140), .B1(n18347), .B2(n18139), .ZN(
        n18131) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18141), .B1(
        n18205), .B2(n18349), .ZN(n18130) );
  OAI211_X1 U21271 ( .C1(n18163), .C2(n18303), .A(n18131), .B(n18130), .ZN(
        P3_U2927) );
  AOI22_X1 U21272 ( .A1(n18353), .A2(n20808), .B1(n20806), .B2(n18139), .ZN(
        n18133) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18141), .B1(
        n18205), .B2(n18354), .ZN(n18132) );
  OAI211_X1 U21274 ( .C1(n18357), .C2(n18136), .A(n18133), .B(n18132), .ZN(
        P3_U2928) );
  AOI22_X1 U21275 ( .A1(n20808), .A2(n18359), .B1(n18358), .B2(n18139), .ZN(
        n18135) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18141), .B1(
        n18205), .B2(n18361), .ZN(n18134) );
  OAI211_X1 U21277 ( .C1(n18365), .C2(n18136), .A(n18135), .B(n18134), .ZN(
        P3_U2929) );
  AOI22_X1 U21278 ( .A1(n18367), .A2(n18140), .B1(n18366), .B2(n18139), .ZN(
        n18138) );
  AOI22_X1 U21279 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18141), .B1(
        n18205), .B2(n18368), .ZN(n18137) );
  OAI211_X1 U21280 ( .C1(n18163), .C2(n18371), .A(n18138), .B(n18137), .ZN(
        P3_U2930) );
  AOI22_X1 U21281 ( .A1(n18375), .A2(n18140), .B1(n18373), .B2(n18139), .ZN(
        n18143) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18141), .B1(
        n18205), .B2(n18376), .ZN(n18142) );
  OAI211_X1 U21283 ( .C1(n18163), .C2(n18381), .A(n18143), .B(n18142), .ZN(
        P3_U2931) );
  NAND2_X1 U21284 ( .A1(n18144), .A2(n18213), .ZN(n20814) );
  NAND2_X1 U21285 ( .A1(n20814), .A2(n18212), .ZN(n18190) );
  AND2_X1 U21286 ( .A1(n18323), .A2(n18190), .ZN(n20807) );
  AOI22_X1 U21287 ( .A1(n18179), .A2(n18330), .B1(n20807), .B2(n18324), .ZN(
        n18150) );
  AOI21_X1 U21288 ( .B1(n18191), .B2(n18145), .A(n18190), .ZN(n18146) );
  AOI211_X1 U21289 ( .C1(n20814), .C2(P3_STATE2_REG_3__SCAN_IN), .A(n18147), 
        .B(n18146), .ZN(n18148) );
  INV_X1 U21290 ( .A(n18148), .ZN(n20817) );
  INV_X1 U21291 ( .A(n20814), .ZN(n18219) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20817), .B1(
        n18219), .B2(n18261), .ZN(n18149) );
  OAI211_X1 U21293 ( .C1(n18163), .C2(n18264), .A(n18150), .B(n18149), .ZN(
        P3_U2932) );
  AOI22_X1 U21294 ( .A1(n18179), .A2(n18336), .B1(n20807), .B2(n18335), .ZN(
        n18152) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20817), .B1(
        n18219), .B2(n18337), .ZN(n18151) );
  OAI211_X1 U21296 ( .C1(n18163), .C2(n18340), .A(n18152), .B(n18151), .ZN(
        P3_U2933) );
  AOI22_X1 U21297 ( .A1(n20808), .A2(n18267), .B1(n20807), .B2(n18341), .ZN(
        n18154) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20817), .B1(
        n18219), .B2(n18343), .ZN(n18153) );
  OAI211_X1 U21299 ( .C1(n20811), .C2(n18270), .A(n18154), .B(n18153), .ZN(
        P3_U2934) );
  AOI22_X1 U21300 ( .A1(n18179), .A2(n18348), .B1(n20807), .B2(n18347), .ZN(
        n18156) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20817), .B1(
        n18219), .B2(n18349), .ZN(n18155) );
  OAI211_X1 U21302 ( .C1(n18163), .C2(n18352), .A(n18156), .B(n18155), .ZN(
        P3_U2935) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20817), .B1(
        n20807), .B2(n18358), .ZN(n18158) );
  AOI22_X1 U21304 ( .A1(n18219), .A2(n18361), .B1(n20808), .B2(n18307), .ZN(
        n18157) );
  OAI211_X1 U21305 ( .C1(n20811), .C2(n18310), .A(n18158), .B(n18157), .ZN(
        P3_U2937) );
  AOI22_X1 U21306 ( .A1(n18179), .A2(n18311), .B1(n20807), .B2(n18366), .ZN(
        n18160) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20817), .B1(
        n18219), .B2(n18368), .ZN(n18159) );
  OAI211_X1 U21308 ( .C1(n18163), .C2(n18314), .A(n18160), .B(n18159), .ZN(
        P3_U2938) );
  AOI22_X1 U21309 ( .A1(n18179), .A2(n18316), .B1(n20807), .B2(n18373), .ZN(
        n18162) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20817), .B1(
        n18219), .B2(n18376), .ZN(n18161) );
  OAI211_X1 U21311 ( .C1(n18163), .C2(n18322), .A(n18162), .B(n18161), .ZN(
        P3_U2939) );
  INV_X1 U21312 ( .A(n18213), .ZN(n18214) );
  NOR2_X1 U21313 ( .A1(n18214), .A2(n18164), .ZN(n18184) );
  AOI22_X1 U21314 ( .A1(n18205), .A2(n18330), .B1(n18324), .B2(n18184), .ZN(
        n18170) );
  NOR2_X1 U21315 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18165), .ZN(
        n18167) );
  NOR2_X1 U21316 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18214), .ZN(
        n18166) );
  AOI22_X1 U21317 ( .A1(n18329), .A2(n18167), .B1(n18327), .B2(n18166), .ZN(
        n18185) );
  NAND2_X1 U21318 ( .A1(n18168), .A2(n18213), .ZN(n18248) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18185), .B1(
        n18261), .B2(n18254), .ZN(n18169) );
  OAI211_X1 U21320 ( .C1(n20811), .C2(n18264), .A(n18170), .B(n18169), .ZN(
        P3_U2940) );
  AOI22_X1 U21321 ( .A1(n18205), .A2(n18336), .B1(n18335), .B2(n18184), .ZN(
        n18172) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18185), .B1(
        n18337), .B2(n18254), .ZN(n18171) );
  OAI211_X1 U21323 ( .C1(n20811), .C2(n18340), .A(n18172), .B(n18171), .ZN(
        P3_U2941) );
  AOI22_X1 U21324 ( .A1(n18179), .A2(n18267), .B1(n18341), .B2(n18184), .ZN(
        n18174) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18185), .B1(
        n18343), .B2(n18254), .ZN(n18173) );
  OAI211_X1 U21326 ( .C1(n18212), .C2(n18270), .A(n18174), .B(n18173), .ZN(
        P3_U2942) );
  AOI22_X1 U21327 ( .A1(n18205), .A2(n18348), .B1(n18347), .B2(n18184), .ZN(
        n18176) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18185), .B1(
        n18349), .B2(n18254), .ZN(n18175) );
  OAI211_X1 U21329 ( .C1(n20811), .C2(n18352), .A(n18176), .B(n18175), .ZN(
        P3_U2943) );
  AOI22_X1 U21330 ( .A1(n18179), .A2(n20809), .B1(n20806), .B2(n18184), .ZN(
        n18178) );
  AOI22_X1 U21331 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18185), .B1(
        n18354), .B2(n18254), .ZN(n18177) );
  OAI211_X1 U21332 ( .C1(n18212), .C2(n20812), .A(n18178), .B(n18177), .ZN(
        P3_U2944) );
  AOI22_X1 U21333 ( .A1(n18179), .A2(n18307), .B1(n18358), .B2(n18184), .ZN(
        n18181) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18185), .B1(
        n18361), .B2(n18254), .ZN(n18180) );
  OAI211_X1 U21335 ( .C1(n18212), .C2(n18310), .A(n18181), .B(n18180), .ZN(
        P3_U2945) );
  AOI22_X1 U21336 ( .A1(n18205), .A2(n18311), .B1(n18366), .B2(n18184), .ZN(
        n18183) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18185), .B1(
        n18368), .B2(n18254), .ZN(n18182) );
  OAI211_X1 U21338 ( .C1(n20811), .C2(n18314), .A(n18183), .B(n18182), .ZN(
        P3_U2946) );
  AOI22_X1 U21339 ( .A1(n18205), .A2(n18316), .B1(n18373), .B2(n18184), .ZN(
        n18187) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18185), .B1(
        n18376), .B2(n18254), .ZN(n18186) );
  OAI211_X1 U21341 ( .C1(n20811), .C2(n18322), .A(n18187), .B(n18186), .ZN(
        P3_U2947) );
  NOR2_X2 U21342 ( .A1(n18188), .A2(n18214), .ZN(n18281) );
  AOI21_X1 U21343 ( .B1(n18248), .B2(n18277), .A(n18456), .ZN(n18208) );
  AOI22_X1 U21344 ( .A1(n18205), .A2(n18325), .B1(n18324), .B2(n18208), .ZN(
        n18194) );
  NAND2_X1 U21345 ( .A1(n18248), .A2(n18277), .ZN(n18192) );
  OAI221_X1 U21346 ( .B1(n18192), .B2(n18191), .C1(n18192), .C2(n18190), .A(
        n18189), .ZN(n18209) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18209), .B1(
        n18219), .B2(n18330), .ZN(n18193) );
  OAI211_X1 U21348 ( .C1(n18333), .C2(n18277), .A(n18194), .B(n18193), .ZN(
        P3_U2948) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18209), .B1(
        n18335), .B2(n18208), .ZN(n18196) );
  AOI22_X1 U21350 ( .A1(n18205), .A2(n18294), .B1(n18337), .B2(n18281), .ZN(
        n18195) );
  OAI211_X1 U21351 ( .C1(n20814), .C2(n18297), .A(n18196), .B(n18195), .ZN(
        P3_U2949) );
  AOI22_X1 U21352 ( .A1(n18219), .A2(n18342), .B1(n18341), .B2(n18208), .ZN(
        n18198) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18209), .B1(
        n18343), .B2(n18281), .ZN(n18197) );
  OAI211_X1 U21354 ( .C1(n18212), .C2(n18346), .A(n18198), .B(n18197), .ZN(
        P3_U2950) );
  AOI22_X1 U21355 ( .A1(n18219), .A2(n18348), .B1(n18347), .B2(n18208), .ZN(
        n18200) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18209), .B1(
        n18349), .B2(n18281), .ZN(n18199) );
  OAI211_X1 U21357 ( .C1(n18212), .C2(n18352), .A(n18200), .B(n18199), .ZN(
        P3_U2951) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18209), .B1(
        n20806), .B2(n18208), .ZN(n18202) );
  AOI22_X1 U21359 ( .A1(n18205), .A2(n20809), .B1(n18354), .B2(n18281), .ZN(
        n18201) );
  OAI211_X1 U21360 ( .C1(n20814), .C2(n20812), .A(n18202), .B(n18201), .ZN(
        P3_U2952) );
  AOI22_X1 U21361 ( .A1(n18219), .A2(n18359), .B1(n18358), .B2(n18208), .ZN(
        n18204) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18209), .B1(
        n18361), .B2(n18281), .ZN(n18203) );
  OAI211_X1 U21363 ( .C1(n18212), .C2(n18365), .A(n18204), .B(n18203), .ZN(
        P3_U2953) );
  AOI22_X1 U21364 ( .A1(n18205), .A2(n18367), .B1(n18366), .B2(n18208), .ZN(
        n18207) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18209), .B1(
        n18368), .B2(n18281), .ZN(n18206) );
  OAI211_X1 U21366 ( .C1(n20814), .C2(n18371), .A(n18207), .B(n18206), .ZN(
        P3_U2954) );
  AOI22_X1 U21367 ( .A1(n18219), .A2(n18316), .B1(n18373), .B2(n18208), .ZN(
        n18211) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18209), .B1(
        n18376), .B2(n18281), .ZN(n18210) );
  OAI211_X1 U21369 ( .C1(n18212), .C2(n18322), .A(n18211), .B(n18210), .ZN(
        P3_U2955) );
  NOR2_X1 U21370 ( .A1(n18428), .A2(n18214), .ZN(n18260) );
  AND2_X1 U21371 ( .A1(n18323), .A2(n18260), .ZN(n18230) );
  AOI22_X1 U21372 ( .A1(n18330), .A2(n18254), .B1(n18324), .B2(n18230), .ZN(
        n18216) );
  OAI211_X1 U21373 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18329), .A(
        n18327), .B(n18213), .ZN(n18231) );
  NOR2_X2 U21374 ( .A1(n18427), .A2(n18214), .ZN(n18306) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18231), .B1(
        n18261), .B2(n18306), .ZN(n18215) );
  OAI211_X1 U21376 ( .C1(n20814), .C2(n18264), .A(n18216), .B(n18215), .ZN(
        P3_U2956) );
  AOI22_X1 U21377 ( .A1(n18336), .A2(n18254), .B1(n18335), .B2(n18230), .ZN(
        n18218) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18231), .B1(
        n18337), .B2(n18306), .ZN(n18217) );
  OAI211_X1 U21379 ( .C1(n20814), .C2(n18340), .A(n18218), .B(n18217), .ZN(
        P3_U2957) );
  AOI22_X1 U21380 ( .A1(n18219), .A2(n18267), .B1(n18341), .B2(n18230), .ZN(
        n18221) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18231), .B1(
        n18343), .B2(n18306), .ZN(n18220) );
  OAI211_X1 U21382 ( .C1(n18270), .C2(n18248), .A(n18221), .B(n18220), .ZN(
        P3_U2958) );
  AOI22_X1 U21383 ( .A1(n18348), .A2(n18254), .B1(n18347), .B2(n18230), .ZN(
        n18223) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18231), .B1(
        n18349), .B2(n18306), .ZN(n18222) );
  OAI211_X1 U21385 ( .C1(n20814), .C2(n18352), .A(n18223), .B(n18222), .ZN(
        P3_U2959) );
  AOI22_X1 U21386 ( .A1(n18353), .A2(n18254), .B1(n20806), .B2(n18230), .ZN(
        n18225) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18231), .B1(
        n18354), .B2(n18306), .ZN(n18224) );
  OAI211_X1 U21388 ( .C1(n20814), .C2(n18357), .A(n18225), .B(n18224), .ZN(
        P3_U2960) );
  AOI22_X1 U21389 ( .A1(n18359), .A2(n18254), .B1(n18358), .B2(n18230), .ZN(
        n18227) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18231), .B1(
        n18361), .B2(n18306), .ZN(n18226) );
  OAI211_X1 U21391 ( .C1(n20814), .C2(n18365), .A(n18227), .B(n18226), .ZN(
        P3_U2961) );
  AOI22_X1 U21392 ( .A1(n18366), .A2(n18230), .B1(n18311), .B2(n18254), .ZN(
        n18229) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18231), .B1(
        n18368), .B2(n18306), .ZN(n18228) );
  OAI211_X1 U21394 ( .C1(n20814), .C2(n18314), .A(n18229), .B(n18228), .ZN(
        P3_U2962) );
  AOI22_X1 U21395 ( .A1(n18316), .A2(n18254), .B1(n18373), .B2(n18230), .ZN(
        n18233) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18231), .B1(
        n18376), .B2(n18306), .ZN(n18232) );
  OAI211_X1 U21397 ( .C1(n20814), .C2(n18322), .A(n18233), .B(n18232), .ZN(
        P3_U2963) );
  NAND2_X1 U21398 ( .A1(n18328), .A2(n18234), .ZN(n18364) );
  INV_X1 U21399 ( .A(n18364), .ZN(n18374) );
  NOR2_X1 U21400 ( .A1(n18306), .A2(n18374), .ZN(n18288) );
  OAI21_X1 U21401 ( .B1(n18236), .B2(n18235), .A(n18288), .ZN(n18237) );
  OAI211_X1 U21402 ( .C1(n18374), .C2(n18555), .A(n18290), .B(n18237), .ZN(
        n18255) );
  NOR2_X1 U21403 ( .A1(n18456), .A2(n18288), .ZN(n18253) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18255), .B1(
        n18324), .B2(n18253), .ZN(n18239) );
  AOI22_X1 U21405 ( .A1(n18325), .A2(n18254), .B1(n18330), .B2(n18281), .ZN(
        n18238) );
  OAI211_X1 U21406 ( .C1(n18333), .C2(n18364), .A(n18239), .B(n18238), .ZN(
        P3_U2964) );
  AOI22_X1 U21407 ( .A1(n18336), .A2(n18281), .B1(n18335), .B2(n18253), .ZN(
        n18241) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18255), .B1(
        n18337), .B2(n18374), .ZN(n18240) );
  OAI211_X1 U21409 ( .C1(n18340), .C2(n18248), .A(n18241), .B(n18240), .ZN(
        P3_U2965) );
  AOI22_X1 U21410 ( .A1(n18267), .A2(n18254), .B1(n18341), .B2(n18253), .ZN(
        n18243) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18255), .B1(
        n18343), .B2(n18374), .ZN(n18242) );
  OAI211_X1 U21412 ( .C1(n18270), .C2(n18277), .A(n18243), .B(n18242), .ZN(
        P3_U2966) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18255), .B1(
        n18347), .B2(n18253), .ZN(n18245) );
  AOI22_X1 U21414 ( .A1(n18349), .A2(n18374), .B1(n18300), .B2(n18254), .ZN(
        n18244) );
  OAI211_X1 U21415 ( .C1(n18303), .C2(n18277), .A(n18245), .B(n18244), .ZN(
        P3_U2967) );
  AOI22_X1 U21416 ( .A1(n18353), .A2(n18281), .B1(n20806), .B2(n18253), .ZN(
        n18247) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18255), .B1(
        n18354), .B2(n18374), .ZN(n18246) );
  OAI211_X1 U21418 ( .C1(n18357), .C2(n18248), .A(n18247), .B(n18246), .ZN(
        P3_U2968) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18255), .B1(
        n18358), .B2(n18253), .ZN(n18250) );
  AOI22_X1 U21420 ( .A1(n18307), .A2(n18254), .B1(n18361), .B2(n18374), .ZN(
        n18249) );
  OAI211_X1 U21421 ( .C1(n18310), .C2(n18277), .A(n18250), .B(n18249), .ZN(
        P3_U2969) );
  AOI22_X1 U21422 ( .A1(n18367), .A2(n18254), .B1(n18366), .B2(n18253), .ZN(
        n18252) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18255), .B1(
        n18368), .B2(n18374), .ZN(n18251) );
  OAI211_X1 U21424 ( .C1(n18371), .C2(n18277), .A(n18252), .B(n18251), .ZN(
        P3_U2970) );
  AOI22_X1 U21425 ( .A1(n18375), .A2(n18254), .B1(n18373), .B2(n18253), .ZN(
        n18257) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18255), .B1(
        n18376), .B2(n18374), .ZN(n18256) );
  OAI211_X1 U21427 ( .C1(n18381), .C2(n18277), .A(n18257), .B(n18256), .ZN(
        P3_U2971) );
  AND2_X1 U21428 ( .A1(n18323), .A2(n18328), .ZN(n18280) );
  AOI22_X1 U21429 ( .A1(n18330), .A2(n18306), .B1(n18324), .B2(n18280), .ZN(
        n18263) );
  AOI22_X1 U21430 ( .A1(n18329), .A2(n18260), .B1(n18259), .B2(n18258), .ZN(
        n18282) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18282), .B1(
        n18360), .B2(n18261), .ZN(n18262) );
  OAI211_X1 U21432 ( .C1(n18264), .C2(n18277), .A(n18263), .B(n18262), .ZN(
        P3_U2972) );
  INV_X1 U21433 ( .A(n18306), .ZN(n18321) );
  AOI22_X1 U21434 ( .A1(n18294), .A2(n18281), .B1(n18335), .B2(n18280), .ZN(
        n18266) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18282), .B1(
        n18360), .B2(n18337), .ZN(n18265) );
  OAI211_X1 U21436 ( .C1(n18297), .C2(n18321), .A(n18266), .B(n18265), .ZN(
        P3_U2973) );
  AOI22_X1 U21437 ( .A1(n18267), .A2(n18281), .B1(n18341), .B2(n18280), .ZN(
        n18269) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18282), .B1(
        n18360), .B2(n18343), .ZN(n18268) );
  OAI211_X1 U21439 ( .C1(n18270), .C2(n18321), .A(n18269), .B(n18268), .ZN(
        P3_U2974) );
  AOI22_X1 U21440 ( .A1(n18300), .A2(n18281), .B1(n18347), .B2(n18280), .ZN(
        n18272) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18282), .B1(
        n18360), .B2(n18349), .ZN(n18271) );
  OAI211_X1 U21442 ( .C1(n18303), .C2(n18321), .A(n18272), .B(n18271), .ZN(
        P3_U2975) );
  AOI22_X1 U21443 ( .A1(n18353), .A2(n18306), .B1(n20806), .B2(n18280), .ZN(
        n18274) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18282), .B1(
        n18354), .B2(n18360), .ZN(n18273) );
  OAI211_X1 U21445 ( .C1(n18357), .C2(n18277), .A(n18274), .B(n18273), .ZN(
        P3_U2976) );
  AOI22_X1 U21446 ( .A1(n18359), .A2(n18306), .B1(n18358), .B2(n18280), .ZN(
        n18276) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18282), .B1(
        n18360), .B2(n18361), .ZN(n18275) );
  OAI211_X1 U21448 ( .C1(n18365), .C2(n18277), .A(n18276), .B(n18275), .ZN(
        P3_U2977) );
  AOI22_X1 U21449 ( .A1(n18367), .A2(n18281), .B1(n18366), .B2(n18280), .ZN(
        n18279) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18282), .B1(
        n18360), .B2(n18368), .ZN(n18278) );
  OAI211_X1 U21451 ( .C1(n18371), .C2(n18321), .A(n18279), .B(n18278), .ZN(
        P3_U2978) );
  AOI22_X1 U21452 ( .A1(n18375), .A2(n18281), .B1(n18373), .B2(n18280), .ZN(
        n18284) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18282), .B1(
        n18360), .B2(n18376), .ZN(n18283) );
  OAI211_X1 U21454 ( .C1(n18381), .C2(n18321), .A(n18284), .B(n18283), .ZN(
        P3_U2979) );
  INV_X1 U21455 ( .A(n18285), .ZN(n18286) );
  NOR2_X1 U21456 ( .A1(n18456), .A2(n18286), .ZN(n18315) );
  AOI22_X1 U21457 ( .A1(n18325), .A2(n18306), .B1(n18324), .B2(n18315), .ZN(
        n18292) );
  OAI21_X1 U21458 ( .B1(n18288), .B2(n18287), .A(n18286), .ZN(n18289) );
  OAI211_X1 U21459 ( .C1(n18317), .C2(n18555), .A(n18290), .B(n18289), .ZN(
        n18318) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18318), .B1(
        n18330), .B2(n18374), .ZN(n18291) );
  OAI211_X1 U21461 ( .C1(n18333), .C2(n18293), .A(n18292), .B(n18291), .ZN(
        P3_U2980) );
  AOI22_X1 U21462 ( .A1(n18294), .A2(n18306), .B1(n18335), .B2(n18315), .ZN(
        n18296) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18337), .ZN(n18295) );
  OAI211_X1 U21464 ( .C1(n18297), .C2(n18364), .A(n18296), .B(n18295), .ZN(
        P3_U2981) );
  AOI22_X1 U21465 ( .A1(n18342), .A2(n18374), .B1(n18341), .B2(n18315), .ZN(
        n18299) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18343), .ZN(n18298) );
  OAI211_X1 U21467 ( .C1(n18346), .C2(n18321), .A(n18299), .B(n18298), .ZN(
        P3_U2982) );
  AOI22_X1 U21468 ( .A1(n18300), .A2(n18306), .B1(n18347), .B2(n18315), .ZN(
        n18302) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18349), .ZN(n18301) );
  OAI211_X1 U21470 ( .C1(n18303), .C2(n18364), .A(n18302), .B(n18301), .ZN(
        P3_U2983) );
  AOI22_X1 U21471 ( .A1(n20809), .A2(n18306), .B1(n20806), .B2(n18315), .ZN(
        n18305) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18318), .B1(
        n18354), .B2(n18317), .ZN(n18304) );
  OAI211_X1 U21473 ( .C1(n20812), .C2(n18364), .A(n18305), .B(n18304), .ZN(
        P3_U2984) );
  AOI22_X1 U21474 ( .A1(n18307), .A2(n18306), .B1(n18358), .B2(n18315), .ZN(
        n18309) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18361), .ZN(n18308) );
  OAI211_X1 U21476 ( .C1(n18310), .C2(n18364), .A(n18309), .B(n18308), .ZN(
        P3_U2985) );
  AOI22_X1 U21477 ( .A1(n18366), .A2(n18315), .B1(n18311), .B2(n18374), .ZN(
        n18313) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18368), .ZN(n18312) );
  OAI211_X1 U21479 ( .C1(n18314), .C2(n18321), .A(n18313), .B(n18312), .ZN(
        P3_U2986) );
  AOI22_X1 U21480 ( .A1(n18316), .A2(n18374), .B1(n18373), .B2(n18315), .ZN(
        n18320) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18376), .ZN(n18319) );
  OAI211_X1 U21482 ( .C1(n18322), .C2(n18321), .A(n18320), .B(n18319), .ZN(
        P3_U2987) );
  AND2_X1 U21483 ( .A1(n18323), .A2(n18326), .ZN(n18372) );
  AOI22_X1 U21484 ( .A1(n18325), .A2(n18374), .B1(n18324), .B2(n18372), .ZN(
        n18332) );
  AOI22_X1 U21485 ( .A1(n18329), .A2(n18328), .B1(n18327), .B2(n18326), .ZN(
        n18378) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18378), .B1(
        n18360), .B2(n18330), .ZN(n18331) );
  OAI211_X1 U21487 ( .C1(n18334), .C2(n18333), .A(n18332), .B(n18331), .ZN(
        P3_U2988) );
  AOI22_X1 U21488 ( .A1(n18360), .A2(n18336), .B1(n18335), .B2(n18372), .ZN(
        n18339) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18378), .B1(
        n18377), .B2(n18337), .ZN(n18338) );
  OAI211_X1 U21490 ( .C1(n18340), .C2(n18364), .A(n18339), .B(n18338), .ZN(
        P3_U2989) );
  AOI22_X1 U21491 ( .A1(n18360), .A2(n18342), .B1(n18341), .B2(n18372), .ZN(
        n18345) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18378), .B1(
        n18377), .B2(n18343), .ZN(n18344) );
  OAI211_X1 U21493 ( .C1(n18346), .C2(n18364), .A(n18345), .B(n18344), .ZN(
        P3_U2990) );
  AOI22_X1 U21494 ( .A1(n18360), .A2(n18348), .B1(n18347), .B2(n18372), .ZN(
        n18351) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18378), .B1(
        n18377), .B2(n18349), .ZN(n18350) );
  OAI211_X1 U21496 ( .C1(n18352), .C2(n18364), .A(n18351), .B(n18350), .ZN(
        P3_U2991) );
  AOI22_X1 U21497 ( .A1(n18353), .A2(n18360), .B1(n20806), .B2(n18372), .ZN(
        n18356) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18378), .B1(
        n18354), .B2(n18377), .ZN(n18355) );
  OAI211_X1 U21499 ( .C1(n18357), .C2(n18364), .A(n18356), .B(n18355), .ZN(
        P3_U2992) );
  AOI22_X1 U21500 ( .A1(n18360), .A2(n18359), .B1(n18358), .B2(n18372), .ZN(
        n18363) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18378), .B1(
        n18377), .B2(n18361), .ZN(n18362) );
  OAI211_X1 U21502 ( .C1(n18365), .C2(n18364), .A(n18363), .B(n18362), .ZN(
        P3_U2993) );
  AOI22_X1 U21503 ( .A1(n18367), .A2(n18374), .B1(n18366), .B2(n18372), .ZN(
        n18370) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18378), .B1(
        n18377), .B2(n18368), .ZN(n18369) );
  OAI211_X1 U21505 ( .C1(n18382), .C2(n18371), .A(n18370), .B(n18369), .ZN(
        P3_U2994) );
  AOI22_X1 U21506 ( .A1(n18375), .A2(n18374), .B1(n18373), .B2(n18372), .ZN(
        n18380) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18378), .B1(
        n18377), .B2(n18376), .ZN(n18379) );
  OAI211_X1 U21508 ( .C1(n18382), .C2(n18381), .A(n18380), .B(n18379), .ZN(
        P3_U2995) );
  AND2_X1 U21509 ( .A1(n18408), .A2(n18383), .ZN(n18388) );
  NOR2_X1 U21510 ( .A1(n18385), .A2(n18384), .ZN(n18387) );
  OAI222_X1 U21511 ( .A1(n18391), .A2(n18390), .B1(n18389), .B2(n18388), .C1(
        n18387), .C2(n18386), .ZN(n18598) );
  OAI21_X1 U21512 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18392), .ZN(n18393) );
  OAI211_X1 U21513 ( .C1(n18395), .C2(n18421), .A(n18394), .B(n18393), .ZN(
        n18442) );
  NOR2_X1 U21514 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18396), .ZN(
        n18425) );
  AND2_X1 U21515 ( .A1(n18573), .A2(n18412), .ZN(n18404) );
  OAI22_X1 U21516 ( .A1(n18419), .A2(n18425), .B1(n18416), .B2(n18404), .ZN(
        n18397) );
  INV_X1 U21517 ( .A(n18397), .ZN(n18556) );
  NOR2_X1 U21518 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18556), .ZN(
        n18407) );
  OAI21_X1 U21519 ( .B1(n18400), .B2(n18399), .A(n18398), .ZN(n18414) );
  AOI21_X1 U21520 ( .B1(n18411), .B2(n18402), .A(n18401), .ZN(n18403) );
  AOI211_X1 U21521 ( .C1(n18414), .C2(n18405), .A(n18404), .B(n18403), .ZN(
        n18559) );
  NAND2_X1 U21522 ( .A1(n18421), .A2(n18559), .ZN(n18406) );
  AOI22_X1 U21523 ( .A1(n18421), .A2(n18407), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18406), .ZN(n18440) );
  AOI21_X1 U21524 ( .B1(n18573), .B2(n18580), .A(n18408), .ZN(n18420) );
  NAND2_X1 U21525 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18409), .ZN(
        n18410) );
  AOI211_X1 U21526 ( .C1(n18411), .C2(n18410), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18580), .ZN(n18418) );
  OAI221_X1 U21527 ( .B1(n18414), .B2(n18580), .C1(n18414), .C2(n18413), .A(
        n18412), .ZN(n18415) );
  OAI22_X1 U21528 ( .A1(n18569), .A2(n18416), .B1(n18573), .B2(n18415), .ZN(
        n18417) );
  AOI211_X1 U21529 ( .C1(n18420), .C2(n18419), .A(n18418), .B(n18417), .ZN(
        n18565) );
  AOI22_X1 U21530 ( .A1(n18431), .A2(n18573), .B1(n18565), .B2(n18421), .ZN(
        n18435) );
  AND2_X1 U21531 ( .A1(n18423), .A2(n18422), .ZN(n18426) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18424), .B1(
        n18426), .B2(n18586), .ZN(n18582) );
  OAI22_X1 U21533 ( .A1(n18426), .A2(n18574), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18425), .ZN(n18578) );
  AOI222_X1 U21534 ( .A1(n18582), .A2(n18578), .B1(n18582), .B2(n18428), .C1(
        n18578), .C2(n18427), .ZN(n18430) );
  OAI21_X1 U21535 ( .B1(n18431), .B2(n18430), .A(n18429), .ZN(n18434) );
  AND2_X1 U21536 ( .A1(n18435), .A2(n18434), .ZN(n18432) );
  OAI221_X1 U21537 ( .B1(n18435), .B2(n18434), .C1(n18433), .C2(n18432), .A(
        n18437), .ZN(n18439) );
  AOI21_X1 U21538 ( .B1(n18437), .B2(n18436), .A(n18435), .ZN(n18438) );
  AOI222_X1 U21539 ( .A1(n18440), .A2(n18439), .B1(n18440), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18439), .C2(n18438), .ZN(
        n18441) );
  NOR4_X1 U21540 ( .A1(n18443), .A2(n18598), .A3(n18442), .A4(n18441), .ZN(
        n18453) );
  NOR2_X1 U21541 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18611) );
  AOI22_X1 U21542 ( .A1(n18606), .A2(n18600), .B1(n18581), .B2(n18611), .ZN(
        n18444) );
  INV_X1 U21543 ( .A(n18444), .ZN(n18449) );
  OAI211_X1 U21544 ( .C1(n18446), .C2(n18445), .A(n18603), .B(n18453), .ZN(
        n18554) );
  OAI21_X1 U21545 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18599), .A(n18554), 
        .ZN(n18454) );
  NOR2_X1 U21546 ( .A1(n18447), .A2(n18454), .ZN(n18448) );
  MUX2_X1 U21547 ( .A(n18449), .B(n18448), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18451) );
  OAI211_X1 U21548 ( .C1(n18453), .C2(n18452), .A(n18451), .B(n18450), .ZN(
        P3_U2996) );
  NAND2_X1 U21549 ( .A1(n18606), .A2(n18600), .ZN(n18459) );
  NOR4_X1 U21550 ( .A1(n18608), .A2(n18566), .A3(n18599), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18462) );
  INV_X1 U21551 ( .A(n18462), .ZN(n18458) );
  OR3_X1 U21552 ( .A1(n18456), .A2(n18455), .A3(n18454), .ZN(n18457) );
  NAND4_X1 U21553 ( .A1(n18460), .A2(n18459), .A3(n18458), .A4(n18457), .ZN(
        P3_U2997) );
  OAI21_X1 U21554 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18461), .ZN(n18463) );
  AOI21_X1 U21555 ( .B1(n18464), .B2(n18463), .A(n18462), .ZN(P3_U2998) );
  AND2_X1 U21556 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18465), .ZN(
        P3_U2999) );
  AND2_X1 U21557 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18465), .ZN(
        P3_U3000) );
  AND2_X1 U21558 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18465), .ZN(
        P3_U3001) );
  AND2_X1 U21559 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18465), .ZN(
        P3_U3002) );
  AND2_X1 U21560 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18465), .ZN(
        P3_U3003) );
  AND2_X1 U21561 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18465), .ZN(
        P3_U3004) );
  AND2_X1 U21562 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18465), .ZN(
        P3_U3005) );
  AND2_X1 U21563 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18465), .ZN(
        P3_U3006) );
  AND2_X1 U21564 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18465), .ZN(
        P3_U3007) );
  AND2_X1 U21565 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18465), .ZN(
        P3_U3008) );
  AND2_X1 U21566 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18465), .ZN(
        P3_U3009) );
  AND2_X1 U21567 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18465), .ZN(
        P3_U3010) );
  AND2_X1 U21568 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18465), .ZN(
        P3_U3011) );
  AND2_X1 U21569 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18465), .ZN(
        P3_U3012) );
  AND2_X1 U21570 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18465), .ZN(
        P3_U3013) );
  AND2_X1 U21571 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18465), .ZN(
        P3_U3014) );
  AND2_X1 U21572 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18465), .ZN(
        P3_U3015) );
  AND2_X1 U21573 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18465), .ZN(
        P3_U3016) );
  AND2_X1 U21574 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18465), .ZN(
        P3_U3017) );
  AND2_X1 U21575 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18465), .ZN(
        P3_U3018) );
  AND2_X1 U21576 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18465), .ZN(
        P3_U3019) );
  AND2_X1 U21577 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18465), .ZN(
        P3_U3020) );
  AND2_X1 U21578 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18465), .ZN(P3_U3021) );
  AND2_X1 U21579 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18465), .ZN(P3_U3022) );
  AND2_X1 U21580 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18465), .ZN(P3_U3023) );
  AND2_X1 U21581 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18465), .ZN(P3_U3024) );
  AND2_X1 U21582 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18465), .ZN(P3_U3025) );
  AND2_X1 U21583 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18465), .ZN(P3_U3026) );
  AND2_X1 U21584 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18465), .ZN(P3_U3027) );
  AND2_X1 U21585 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18465), .ZN(P3_U3028) );
  INV_X1 U21586 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18613) );
  AOI21_X1 U21587 ( .B1(HOLD), .B2(n18466), .A(n18613), .ZN(n18469) );
  NAND2_X1 U21588 ( .A1(n18606), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18476) );
  INV_X1 U21589 ( .A(n18476), .ZN(n18474) );
  OAI21_X1 U21590 ( .B1(n18474), .B2(n18480), .A(n18482), .ZN(n18468) );
  NAND3_X1 U21591 ( .A1(NA), .A2(n18480), .A3(n18467), .ZN(n18475) );
  OAI211_X1 U21592 ( .C1(n18543), .C2(n18469), .A(n18468), .B(n18475), .ZN(
        P3_U3029) );
  INV_X1 U21593 ( .A(HOLD), .ZN(n19603) );
  NOR2_X1 U21594 ( .A1(n18482), .A2(n19603), .ZN(n18478) );
  OAI22_X1 U21595 ( .A1(n18478), .A2(n18613), .B1(n19603), .B2(n18470), .ZN(
        n18471) );
  NAND2_X1 U21596 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18471), .ZN(n18473) );
  NAND3_X1 U21597 ( .A1(n18473), .A2(n18476), .A3(n18472), .ZN(P3_U3030) );
  AOI21_X1 U21598 ( .B1(n18480), .B2(n18475), .A(n18474), .ZN(n18481) );
  OAI22_X1 U21599 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18476), .ZN(n18477) );
  OAI22_X1 U21600 ( .A1(n18478), .A2(n18477), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18479) );
  OAI22_X1 U21601 ( .A1(n18481), .A2(n18482), .B1(n18480), .B2(n18479), .ZN(
        P3_U3031) );
  INV_X1 U21602 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18484) );
  OAI222_X1 U21603 ( .A1(n18588), .A2(n18541), .B1(n18483), .B2(n18543), .C1(
        n18484), .C2(n18540), .ZN(P3_U3032) );
  OAI222_X1 U21604 ( .A1(n18540), .A2(n18486), .B1(n18485), .B2(n18543), .C1(
        n18484), .C2(n18541), .ZN(P3_U3033) );
  OAI222_X1 U21605 ( .A1(n18540), .A2(n18488), .B1(n18487), .B2(n18543), .C1(
        n18486), .C2(n18541), .ZN(P3_U3034) );
  OAI222_X1 U21606 ( .A1(n18540), .A2(n18491), .B1(n18489), .B2(n18543), .C1(
        n18488), .C2(n18541), .ZN(P3_U3035) );
  OAI222_X1 U21607 ( .A1(n18491), .A2(n18541), .B1(n18490), .B2(n18543), .C1(
        n18492), .C2(n18540), .ZN(P3_U3036) );
  OAI222_X1 U21608 ( .A1(n18540), .A2(n18494), .B1(n18493), .B2(n18543), .C1(
        n18492), .C2(n18541), .ZN(P3_U3037) );
  OAI222_X1 U21609 ( .A1(n18540), .A2(n18497), .B1(n18495), .B2(n18543), .C1(
        n18494), .C2(n18541), .ZN(P3_U3038) );
  OAI222_X1 U21610 ( .A1(n18497), .A2(n18541), .B1(n18496), .B2(n18543), .C1(
        n18498), .C2(n18540), .ZN(P3_U3039) );
  OAI222_X1 U21611 ( .A1(n18540), .A2(n18500), .B1(n18499), .B2(n18543), .C1(
        n18498), .C2(n18541), .ZN(P3_U3040) );
  OAI222_X1 U21612 ( .A1(n18540), .A2(n18502), .B1(n18501), .B2(n18543), .C1(
        n18500), .C2(n18541), .ZN(P3_U3041) );
  OAI222_X1 U21613 ( .A1(n18540), .A2(n18504), .B1(n18503), .B2(n18543), .C1(
        n18502), .C2(n18541), .ZN(P3_U3042) );
  OAI222_X1 U21614 ( .A1(n18540), .A2(n18506), .B1(n18505), .B2(n18543), .C1(
        n18504), .C2(n18541), .ZN(P3_U3043) );
  OAI222_X1 U21615 ( .A1(n18540), .A2(n18509), .B1(n18507), .B2(n18543), .C1(
        n18506), .C2(n18541), .ZN(P3_U3044) );
  OAI222_X1 U21616 ( .A1(n18509), .A2(n18541), .B1(n18508), .B2(n18543), .C1(
        n18510), .C2(n18540), .ZN(P3_U3045) );
  OAI222_X1 U21617 ( .A1(n18540), .A2(n18512), .B1(n18511), .B2(n18543), .C1(
        n18510), .C2(n18541), .ZN(P3_U3046) );
  OAI222_X1 U21618 ( .A1(n18540), .A2(n18514), .B1(n18513), .B2(n18543), .C1(
        n18512), .C2(n18541), .ZN(P3_U3047) );
  OAI222_X1 U21619 ( .A1(n18540), .A2(n18516), .B1(n18515), .B2(n18543), .C1(
        n18514), .C2(n18541), .ZN(P3_U3048) );
  OAI222_X1 U21620 ( .A1(n18540), .A2(n18518), .B1(n18517), .B2(n18543), .C1(
        n18516), .C2(n18541), .ZN(P3_U3049) );
  OAI222_X1 U21621 ( .A1(n18540), .A2(n18521), .B1(n18519), .B2(n18543), .C1(
        n18518), .C2(n18541), .ZN(P3_U3050) );
  OAI222_X1 U21622 ( .A1(n18521), .A2(n18541), .B1(n18520), .B2(n18543), .C1(
        n18522), .C2(n18540), .ZN(P3_U3051) );
  OAI222_X1 U21623 ( .A1(n18540), .A2(n18524), .B1(n18523), .B2(n18543), .C1(
        n18522), .C2(n18541), .ZN(P3_U3052) );
  OAI222_X1 U21624 ( .A1(n18540), .A2(n18526), .B1(n18525), .B2(n18543), .C1(
        n18524), .C2(n18541), .ZN(P3_U3053) );
  OAI222_X1 U21625 ( .A1(n18540), .A2(n18528), .B1(n18527), .B2(n18543), .C1(
        n18526), .C2(n18541), .ZN(P3_U3054) );
  OAI222_X1 U21626 ( .A1(n18540), .A2(n18530), .B1(n18529), .B2(n18543), .C1(
        n18528), .C2(n18541), .ZN(P3_U3055) );
  INV_X1 U21627 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18532) );
  OAI222_X1 U21628 ( .A1(n18540), .A2(n18532), .B1(n18531), .B2(n18543), .C1(
        n18530), .C2(n18541), .ZN(P3_U3056) );
  OAI222_X1 U21629 ( .A1(n18540), .A2(n18535), .B1(n18533), .B2(n18543), .C1(
        n18532), .C2(n18541), .ZN(P3_U3057) );
  INV_X1 U21630 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18536) );
  OAI222_X1 U21631 ( .A1(n18541), .A2(n18535), .B1(n18534), .B2(n18543), .C1(
        n18536), .C2(n18540), .ZN(P3_U3058) );
  OAI222_X1 U21632 ( .A1(n18540), .A2(n18538), .B1(n18537), .B2(n18543), .C1(
        n18536), .C2(n18541), .ZN(P3_U3059) );
  OAI222_X1 U21633 ( .A1(n18540), .A2(n18542), .B1(n18539), .B2(n18543), .C1(
        n18538), .C2(n18541), .ZN(P3_U3060) );
  OAI222_X1 U21634 ( .A1(n18540), .A2(n18545), .B1(n18544), .B2(n18543), .C1(
        n18542), .C2(n18541), .ZN(P3_U3061) );
  OAI22_X1 U21635 ( .A1(n18615), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18543), .ZN(n18546) );
  INV_X1 U21636 ( .A(n18546), .ZN(P3_U3274) );
  MUX2_X1 U21637 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n18615), .Z(P3_U3275) );
  OAI22_X1 U21638 ( .A1(n18615), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18543), .ZN(n18547) );
  INV_X1 U21639 ( .A(n18547), .ZN(P3_U3276) );
  OAI22_X1 U21640 ( .A1(n18615), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18543), .ZN(n18548) );
  INV_X1 U21641 ( .A(n18548), .ZN(P3_U3277) );
  OAI21_X1 U21642 ( .B1(n18552), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18550), 
        .ZN(n18549) );
  INV_X1 U21643 ( .A(n18549), .ZN(P3_U3280) );
  OAI21_X1 U21644 ( .B1(n18552), .B2(n18551), .A(n18550), .ZN(P3_U3281) );
  OAI221_X1 U21645 ( .B1(n18555), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18555), 
        .C2(n18554), .A(n18553), .ZN(P3_U3282) );
  INV_X1 U21646 ( .A(n18584), .ZN(n18587) );
  NOR3_X1 U21647 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18556), .A3(
        n18560), .ZN(n18557) );
  AOI21_X1 U21648 ( .B1(n18581), .B2(n18558), .A(n18557), .ZN(n18564) );
  OAI21_X1 U21649 ( .B1(n18560), .B2(n18559), .A(n18584), .ZN(n18561) );
  INV_X1 U21650 ( .A(n18561), .ZN(n18563) );
  OAI22_X1 U21651 ( .A1(n18587), .A2(n18564), .B1(n18563), .B2(n18562), .ZN(
        P3_U3285) );
  INV_X1 U21652 ( .A(n18565), .ZN(n18571) );
  NOR2_X1 U21653 ( .A1(n18566), .A2(n18583), .ZN(n18575) );
  OAI22_X1 U21654 ( .A1(n18568), .A2(n18567), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18576) );
  INV_X1 U21655 ( .A(n18576), .ZN(n18570) );
  AOI222_X1 U21656 ( .A1(n18571), .A2(n18618), .B1(n18575), .B2(n18570), .C1(
        n18581), .C2(n18569), .ZN(n18572) );
  AOI22_X1 U21657 ( .A1(n18587), .A2(n18573), .B1(n18572), .B2(n18584), .ZN(
        P3_U3288) );
  INV_X1 U21658 ( .A(n18574), .ZN(n18577) );
  AOI222_X1 U21659 ( .A1(n18578), .A2(n18618), .B1(n18581), .B2(n18577), .C1(
        n18576), .C2(n18575), .ZN(n18579) );
  AOI22_X1 U21660 ( .A1(n18587), .A2(n18580), .B1(n18579), .B2(n18584), .ZN(
        P3_U3289) );
  AOI222_X1 U21661 ( .A1(n18583), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18618), 
        .B2(n18582), .C1(n18586), .C2(n18581), .ZN(n18585) );
  AOI22_X1 U21662 ( .A1(n18587), .A2(n18586), .B1(n18585), .B2(n18584), .ZN(
        P3_U3290) );
  AOI22_X1 U21663 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18589), .B2(n18588), .ZN(n18592) );
  NOR3_X1 U21664 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .A3(n18595), .ZN(n18593) );
  NAND2_X1 U21665 ( .A1(P3_DATAWIDTH_REG_0__SCAN_IN), .A2(n18593), .ZN(n18591)
         );
  NAND2_X1 U21666 ( .A1(n18595), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18590) );
  OAI211_X1 U21667 ( .C1(n18595), .C2(n18592), .A(n18591), .B(n18590), .ZN(
        P3_U3292) );
  INV_X1 U21668 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18594) );
  AOI21_X1 U21669 ( .B1(n18595), .B2(n18594), .A(n18593), .ZN(P3_U3293) );
  INV_X1 U21670 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18621) );
  OAI22_X1 U21671 ( .A1(n18615), .A2(n18621), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18543), .ZN(n18596) );
  INV_X1 U21672 ( .A(n18596), .ZN(P3_U3294) );
  MUX2_X1 U21673 ( .A(P3_MORE_REG_SCAN_IN), .B(n18598), .S(n18597), .Z(
        P3_U3295) );
  AOI21_X1 U21674 ( .B1(n18600), .B2(n18599), .A(n18620), .ZN(n18601) );
  OAI21_X1 U21675 ( .B1(n18603), .B2(n18602), .A(n18601), .ZN(n18614) );
  OAI21_X1 U21676 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18605), .A(n18604), 
        .ZN(n18607) );
  AOI211_X1 U21677 ( .C1(n18619), .C2(n18607), .A(n18606), .B(n18617), .ZN(
        n18609) );
  NOR2_X1 U21678 ( .A1(n18609), .A2(n18608), .ZN(n18610) );
  OAI21_X1 U21679 ( .B1(n18611), .B2(n18610), .A(n18614), .ZN(n18612) );
  OAI21_X1 U21680 ( .B1(n18614), .B2(n18613), .A(n18612), .ZN(P3_U3296) );
  OAI22_X1 U21681 ( .A1(n18615), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18543), .ZN(n18616) );
  INV_X1 U21682 ( .A(n18616), .ZN(P3_U3297) );
  AOI21_X1 U21683 ( .B1(n18618), .B2(n18617), .A(n18620), .ZN(n18624) );
  AOI22_X1 U21684 ( .A1(n18624), .A2(n18621), .B1(n18620), .B2(n18619), .ZN(
        P3_U3298) );
  INV_X1 U21685 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18623) );
  AOI21_X1 U21686 ( .B1(n18624), .B2(n18623), .A(n18622), .ZN(P3_U3299) );
  INV_X1 U21687 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19602) );
  NAND2_X1 U21688 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19608), .ZN(n19595) );
  NAND2_X1 U21689 ( .A1(n19602), .A2(n19587), .ZN(n19591) );
  OAI21_X1 U21690 ( .B1(n19602), .B2(n19595), .A(n19591), .ZN(n19667) );
  AOI21_X1 U21691 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19667), .ZN(n18625) );
  INV_X1 U21692 ( .A(n18625), .ZN(P2_U2815) );
  INV_X1 U21693 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18629) );
  NAND2_X1 U21694 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19697), .ZN(n18628) );
  NAND2_X1 U21695 ( .A1(n18626), .A2(n19504), .ZN(n18627) );
  OAI22_X1 U21696 ( .A1(n19724), .A2(n18629), .B1(n18628), .B2(n18627), .ZN(
        P2_U2816) );
  INV_X2 U21697 ( .A(n19737), .ZN(n19736) );
  AOI21_X1 U21698 ( .B1(n19602), .B2(n19608), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18630) );
  AOI22_X1 U21699 ( .A1(n19736), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18630), 
        .B2(n19737), .ZN(P2_U2817) );
  OAI21_X1 U21700 ( .B1(n19600), .B2(BS16), .A(n19667), .ZN(n19665) );
  OAI21_X1 U21701 ( .B1(n19667), .B2(n19668), .A(n19665), .ZN(P2_U2818) );
  NOR2_X1 U21702 ( .A1(n18632), .A2(n18631), .ZN(n19706) );
  OAI21_X1 U21703 ( .B1(n19706), .B2(n18634), .A(n18633), .ZN(P2_U2819) );
  NOR4_X1 U21704 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18638) );
  NOR4_X1 U21705 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18637) );
  NOR4_X1 U21706 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18636) );
  NOR4_X1 U21707 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18635) );
  NAND4_X1 U21708 ( .A1(n18638), .A2(n18637), .A3(n18636), .A4(n18635), .ZN(
        n18644) );
  NOR4_X1 U21709 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18642) );
  AOI211_X1 U21710 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_3__SCAN_IN), .B(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18641) );
  NOR4_X1 U21711 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18640) );
  NOR4_X1 U21712 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18639) );
  NAND4_X1 U21713 ( .A1(n18642), .A2(n18641), .A3(n18640), .A4(n18639), .ZN(
        n18643) );
  NOR2_X1 U21714 ( .A1(n18644), .A2(n18643), .ZN(n18653) );
  INV_X1 U21715 ( .A(n18653), .ZN(n18652) );
  NOR2_X1 U21716 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18652), .ZN(n18647) );
  INV_X1 U21717 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18645) );
  AOI22_X1 U21718 ( .A1(n18647), .A2(n10156), .B1(n18652), .B2(n18645), .ZN(
        P2_U2820) );
  OR3_X1 U21719 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18651) );
  INV_X1 U21720 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18646) );
  AOI22_X1 U21721 ( .A1(n18647), .A2(n18651), .B1(n18652), .B2(n18646), .ZN(
        P2_U2821) );
  INV_X1 U21722 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19666) );
  NAND2_X1 U21723 ( .A1(n18647), .A2(n19666), .ZN(n18650) );
  OAI21_X1 U21724 ( .B1(n10168), .B2(n10156), .A(n18653), .ZN(n18648) );
  OAI21_X1 U21725 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18653), .A(n18648), 
        .ZN(n18649) );
  OAI221_X1 U21726 ( .B1(n18650), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18650), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18649), .ZN(P2_U2822) );
  INV_X1 U21727 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19661) );
  OAI221_X1 U21728 ( .B1(n18653), .B2(n19661), .C1(n18652), .C2(n18651), .A(
        n18650), .ZN(P2_U2823) );
  AOI211_X1 U21729 ( .C1(n18656), .C2(n18655), .A(n18654), .B(n19582), .ZN(
        n18657) );
  INV_X1 U21730 ( .A(n18657), .ZN(n18667) );
  AOI22_X1 U21731 ( .A1(n18861), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18862), .ZN(n18666) );
  OAI22_X1 U21732 ( .A1(n18659), .A2(n18871), .B1(n18658), .B2(n18865), .ZN(
        n18660) );
  INV_X1 U21733 ( .A(n18660), .ZN(n18665) );
  INV_X1 U21734 ( .A(n18661), .ZN(n18663) );
  AOI22_X1 U21735 ( .A1(n18663), .A2(n18868), .B1(n18662), .B2(n18859), .ZN(
        n18664) );
  NAND4_X1 U21736 ( .A1(n18667), .A2(n18666), .A3(n18665), .A4(n18664), .ZN(
        P2_U2834) );
  AOI211_X1 U21737 ( .C1(n18670), .C2(n18669), .A(n18668), .B(n19582), .ZN(
        n18675) );
  AOI22_X1 U21738 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n18861), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18862), .ZN(n18672) );
  NAND2_X1 U21739 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18842), .ZN(
        n18671) );
  OAI211_X1 U21740 ( .C1(n18673), .C2(n18865), .A(n18672), .B(n18671), .ZN(
        n18674) );
  AOI211_X1 U21741 ( .C1(n18859), .C2(n18676), .A(n18675), .B(n18674), .ZN(
        n18677) );
  OAI21_X1 U21742 ( .B1(n18678), .B2(n18858), .A(n18677), .ZN(P2_U2835) );
  AOI211_X1 U21743 ( .C1(n18681), .C2(n18680), .A(n18679), .B(n19582), .ZN(
        n18686) );
  AOI21_X1 U21744 ( .B1(P2_REIP_REG_19__SCAN_IN), .B2(n18862), .A(n15127), 
        .ZN(n18683) );
  AOI22_X1 U21745 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18842), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n18861), .ZN(n18682) );
  OAI211_X1 U21746 ( .C1(n18684), .C2(n18865), .A(n18683), .B(n18682), .ZN(
        n18685) );
  AOI211_X1 U21747 ( .C1(n18868), .C2(n18687), .A(n18686), .B(n18685), .ZN(
        n18688) );
  OAI21_X1 U21748 ( .B1(n18689), .B2(n18841), .A(n18688), .ZN(P2_U2836) );
  AOI211_X1 U21749 ( .C1(n18691), .C2(n18704), .A(n18690), .B(n19582), .ZN(
        n18696) );
  AOI21_X1 U21750 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n18862), .A(n15127), 
        .ZN(n18693) );
  AOI22_X1 U21751 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18842), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n18861), .ZN(n18692) );
  OAI211_X1 U21752 ( .C1(n18694), .C2(n18865), .A(n18693), .B(n18692), .ZN(
        n18695) );
  AOI211_X1 U21753 ( .C1(n18859), .C2(n9995), .A(n18696), .B(n18695), .ZN(
        n18697) );
  OAI21_X1 U21754 ( .B1(n18698), .B2(n18858), .A(n18697), .ZN(P2_U2837) );
  AOI22_X1 U21755 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n18861), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18842), .ZN(n18699) );
  OAI211_X1 U21756 ( .C1(n19634), .C2(n18845), .A(n18699), .B(n14056), .ZN(
        n18702) );
  OAI22_X1 U21757 ( .A1(n18700), .A2(n18865), .B1(n18705), .B2(n18870), .ZN(
        n18701) );
  AOI211_X1 U21758 ( .C1(n18703), .C2(n18868), .A(n18702), .B(n18701), .ZN(
        n18708) );
  OAI211_X1 U21759 ( .C1(n18706), .C2(n18705), .A(n18838), .B(n18704), .ZN(
        n18707) );
  OAI211_X1 U21760 ( .C1(n18841), .C2(n18709), .A(n18708), .B(n18707), .ZN(
        P2_U2838) );
  NAND2_X1 U21761 ( .A1(n13108), .A2(n18710), .ZN(n18711) );
  XOR2_X1 U21762 ( .A(n18712), .B(n18711), .Z(n18719) );
  AOI22_X1 U21763 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18842), .B1(
        n18713), .B2(n18847), .ZN(n18714) );
  OAI211_X1 U21764 ( .C1(n19632), .C2(n18845), .A(n18714), .B(n14056), .ZN(
        n18715) );
  AOI21_X1 U21765 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n18861), .A(n18715), .ZN(
        n18718) );
  AOI22_X1 U21766 ( .A1(n18716), .A2(n18868), .B1(n18885), .B2(n18859), .ZN(
        n18717) );
  OAI211_X1 U21767 ( .C1(n19582), .C2(n18719), .A(n18718), .B(n18717), .ZN(
        P2_U2839) );
  NOR2_X1 U21768 ( .A1(n18810), .A2(n18720), .ZN(n18721) );
  XOR2_X1 U21769 ( .A(n18722), .B(n18721), .Z(n18729) );
  AOI22_X1 U21770 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n18861), .B1(n18723), 
        .B2(n18847), .ZN(n18724) );
  OAI211_X1 U21771 ( .C1(n19630), .C2(n18845), .A(n18724), .B(n14056), .ZN(
        n18727) );
  OAI22_X1 U21772 ( .A1(n18725), .A2(n18858), .B1(n18893), .B2(n18841), .ZN(
        n18726) );
  AOI211_X1 U21773 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18842), .A(
        n18727), .B(n18726), .ZN(n18728) );
  OAI21_X1 U21774 ( .B1(n19582), .B2(n18729), .A(n18728), .ZN(P2_U2840) );
  AOI22_X1 U21775 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18842), .B1(
        n18730), .B2(n18847), .ZN(n18731) );
  OAI211_X1 U21776 ( .C1(n19628), .C2(n18845), .A(n18731), .B(n14056), .ZN(
        n18732) );
  AOI21_X1 U21777 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n18861), .A(n18732), .ZN(
        n18739) );
  NAND2_X1 U21778 ( .A1(n13108), .A2(n18733), .ZN(n18734) );
  XOR2_X1 U21779 ( .A(n18735), .B(n18734), .Z(n18736) );
  AOI22_X1 U21780 ( .A1(n18737), .A2(n18859), .B1(n18838), .B2(n18736), .ZN(
        n18738) );
  OAI211_X1 U21781 ( .C1(n18740), .C2(n18858), .A(n18739), .B(n18738), .ZN(
        P2_U2841) );
  OAI22_X1 U21782 ( .A1(n18742), .A2(n18871), .B1(n18741), .B2(n18865), .ZN(
        n18743) );
  AOI211_X1 U21783 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18862), .A(n15127), 
        .B(n18743), .ZN(n18751) );
  NOR2_X1 U21784 ( .A1(n18810), .A2(n18744), .ZN(n18745) );
  XOR2_X1 U21785 ( .A(n18746), .B(n18745), .Z(n18749) );
  OAI22_X1 U21786 ( .A1(n18747), .A2(n18858), .B1(n18897), .B2(n18841), .ZN(
        n18748) );
  AOI21_X1 U21787 ( .B1(n18749), .B2(n18838), .A(n18748), .ZN(n18750) );
  OAI211_X1 U21788 ( .C1(n18777), .C2(n10507), .A(n18751), .B(n18750), .ZN(
        P2_U2842) );
  INV_X1 U21789 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19625) );
  OAI21_X1 U21790 ( .B1(n19625), .B2(n18845), .A(n14056), .ZN(n18755) );
  OAI22_X1 U21791 ( .A1(n18753), .A2(n18871), .B1(n18752), .B2(n18865), .ZN(
        n18754) );
  AOI211_X1 U21792 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n18861), .A(n18755), .B(
        n18754), .ZN(n18761) );
  NAND2_X1 U21793 ( .A1(n13108), .A2(n18770), .ZN(n18756) );
  XNOR2_X1 U21794 ( .A(n18757), .B(n18756), .ZN(n18758) );
  AOI22_X1 U21795 ( .A1(n18859), .A2(n18759), .B1(n18838), .B2(n18758), .ZN(
        n18760) );
  OAI211_X1 U21796 ( .C1(n18858), .C2(n18762), .A(n18761), .B(n18760), .ZN(
        P2_U2843) );
  OAI22_X1 U21797 ( .A1(n18777), .A2(n18763), .B1(n10766), .B2(n18871), .ZN(
        n18768) );
  INV_X1 U21798 ( .A(n18901), .ZN(n18764) );
  AOI22_X1 U21799 ( .A1(n18765), .A2(n18847), .B1(n18859), .B2(n18764), .ZN(
        n18766) );
  OAI211_X1 U21800 ( .C1(n10767), .C2(n18845), .A(n18766), .B(n14056), .ZN(
        n18767) );
  AOI211_X1 U21801 ( .C1(n18868), .C2(n18769), .A(n18768), .B(n18767), .ZN(
        n18774) );
  NAND2_X1 U21802 ( .A1(n13108), .A2(n18838), .ZN(n18877) );
  INV_X1 U21803 ( .A(n18877), .ZN(n18771) );
  OAI211_X1 U21804 ( .C1(n18772), .C2(n18775), .A(n18771), .B(n18770), .ZN(
        n18773) );
  OAI211_X1 U21805 ( .C1(n18870), .C2(n18775), .A(n18774), .B(n18773), .ZN(
        P2_U2844) );
  OAI22_X1 U21806 ( .A1(n18777), .A2(n9925), .B1(n18776), .B2(n18865), .ZN(
        n18778) );
  AOI211_X1 U21807 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n18862), .A(n15127), 
        .B(n18778), .ZN(n18786) );
  NAND2_X1 U21808 ( .A1(n13108), .A2(n18779), .ZN(n18780) );
  XNOR2_X1 U21809 ( .A(n18781), .B(n18780), .ZN(n18784) );
  OAI22_X1 U21810 ( .A1(n18841), .A2(n18904), .B1(n18858), .B2(n18782), .ZN(
        n18783) );
  AOI21_X1 U21811 ( .B1(n18838), .B2(n18784), .A(n18783), .ZN(n18785) );
  OAI211_X1 U21812 ( .C1(n18787), .C2(n18871), .A(n18786), .B(n18785), .ZN(
        P2_U2845) );
  NOR2_X1 U21813 ( .A1(n18810), .A2(n18788), .ZN(n18789) );
  XOR2_X1 U21814 ( .A(n18790), .B(n18789), .Z(n18797) );
  INV_X1 U21815 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19620) );
  AOI22_X1 U21816 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18842), .B1(
        n18847), .B2(n18791), .ZN(n18792) );
  OAI211_X1 U21817 ( .C1(n19620), .C2(n18845), .A(n18792), .B(n14056), .ZN(
        n18795) );
  OAI22_X1 U21818 ( .A1(n18841), .A2(n18907), .B1(n18858), .B2(n18793), .ZN(
        n18794) );
  AOI211_X1 U21819 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n18861), .A(n18795), .B(
        n18794), .ZN(n18796) );
  OAI21_X1 U21820 ( .B1(n19582), .B2(n18797), .A(n18796), .ZN(P2_U2846) );
  OAI21_X1 U21821 ( .B1(n19619), .B2(n18845), .A(n14056), .ZN(n18801) );
  OAI22_X1 U21822 ( .A1(n18799), .A2(n18871), .B1(n18798), .B2(n18865), .ZN(
        n18800) );
  AOI211_X1 U21823 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n18861), .A(n18801), .B(
        n18800), .ZN(n18808) );
  NAND2_X1 U21824 ( .A1(n13108), .A2(n18802), .ZN(n18803) );
  XNOR2_X1 U21825 ( .A(n18804), .B(n18803), .ZN(n18806) );
  AOI22_X1 U21826 ( .A1(n18838), .A2(n18806), .B1(n18868), .B2(n18805), .ZN(
        n18807) );
  OAI211_X1 U21827 ( .C1(n18841), .C2(n18910), .A(n18808), .B(n18807), .ZN(
        P2_U2847) );
  NOR2_X1 U21828 ( .A1(n18810), .A2(n18809), .ZN(n18811) );
  XOR2_X1 U21829 ( .A(n18812), .B(n18811), .Z(n18819) );
  AOI22_X1 U21830 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18842), .B1(
        n18813), .B2(n18847), .ZN(n18814) );
  OAI211_X1 U21831 ( .C1(n10750), .C2(n18845), .A(n18814), .B(n14056), .ZN(
        n18817) );
  OAI22_X1 U21832 ( .A1(n18841), .A2(n18911), .B1(n18858), .B2(n18815), .ZN(
        n18816) );
  AOI211_X1 U21833 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n18861), .A(n18817), .B(
        n18816), .ZN(n18818) );
  OAI21_X1 U21834 ( .B1(n19582), .B2(n18819), .A(n18818), .ZN(P2_U2848) );
  OAI21_X1 U21835 ( .B1(n19616), .B2(n18845), .A(n14056), .ZN(n18823) );
  OAI22_X1 U21836 ( .A1(n18821), .A2(n18871), .B1(n18820), .B2(n18865), .ZN(
        n18822) );
  AOI211_X1 U21837 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n18861), .A(n18823), .B(
        n18822), .ZN(n18829) );
  NAND2_X1 U21838 ( .A1(n13108), .A2(n18824), .ZN(n18825) );
  XNOR2_X1 U21839 ( .A(n18826), .B(n18825), .ZN(n18827) );
  AOI22_X1 U21840 ( .A1(n18838), .A2(n18827), .B1(n18868), .B2(n9716), .ZN(
        n18828) );
  OAI211_X1 U21841 ( .C1(n18841), .C2(n18912), .A(n18829), .B(n18828), .ZN(
        P2_U2849) );
  AOI22_X1 U21842 ( .A1(P2_EBX_REG_5__SCAN_IN), .A2(n18861), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18842), .ZN(n18830) );
  OAI21_X1 U21843 ( .B1(n18831), .B2(n18865), .A(n18830), .ZN(n18832) );
  AOI211_X1 U21844 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18862), .A(n15127), .B(
        n18832), .ZN(n18840) );
  NOR2_X1 U21845 ( .A1(n18810), .A2(n18833), .ZN(n18835) );
  XNOR2_X1 U21846 ( .A(n18835), .B(n18834), .ZN(n18837) );
  AOI22_X1 U21847 ( .A1(n18838), .A2(n18837), .B1(n18868), .B2(n18836), .ZN(
        n18839) );
  OAI211_X1 U21848 ( .C1(n18841), .C2(n18919), .A(n18840), .B(n18839), .ZN(
        P2_U2850) );
  AOI22_X1 U21849 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18842), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n18861), .ZN(n18850) );
  NAND2_X1 U21850 ( .A1(n18859), .A2(n18843), .ZN(n18844) );
  OAI211_X1 U21851 ( .C1(n19612), .C2(n18845), .A(n18844), .B(n14056), .ZN(
        n18846) );
  AOI21_X1 U21852 ( .B1(n18848), .B2(n18847), .A(n18846), .ZN(n18849) );
  OAI211_X1 U21853 ( .C1(n18915), .C2(n18851), .A(n18850), .B(n18849), .ZN(
        n18852) );
  INV_X1 U21854 ( .A(n18852), .ZN(n18857) );
  AND2_X1 U21855 ( .A1(n13108), .A2(n18853), .ZN(n18855) );
  AOI21_X1 U21856 ( .B1(n19048), .B2(n18855), .A(n19582), .ZN(n18854) );
  OAI21_X1 U21857 ( .B1(n19048), .B2(n18855), .A(n18854), .ZN(n18856) );
  OAI211_X1 U21858 ( .C1(n19056), .C2(n18858), .A(n18857), .B(n18856), .ZN(
        P2_U2851) );
  NAND2_X1 U21859 ( .A1(n18860), .A2(n18859), .ZN(n18864) );
  AOI22_X1 U21860 ( .A1(n18862), .A2(P2_REIP_REG_0__SCAN_IN), .B1(
        P2_EBX_REG_0__SCAN_IN), .B2(n18861), .ZN(n18863) );
  OAI211_X1 U21861 ( .C1(n18866), .C2(n18865), .A(n18864), .B(n18863), .ZN(
        n18867) );
  AOI21_X1 U21862 ( .B1(n18869), .B2(n18868), .A(n18867), .ZN(n18876) );
  NAND2_X1 U21863 ( .A1(n18871), .A2(n18870), .ZN(n18874) );
  AOI22_X1 U21864 ( .A1(n18874), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18873), .B2(n18872), .ZN(n18875) );
  OAI211_X1 U21865 ( .C1(n18878), .C2(n18877), .A(n18876), .B(n18875), .ZN(
        P2_U2855) );
  AOI22_X1 U21866 ( .A1(n15890), .A2(n18932), .B1(n18883), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n18880) );
  AOI22_X1 U21867 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n18931), .B1(n18884), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n18879) );
  NAND2_X1 U21868 ( .A1(n18880), .A2(n18879), .ZN(P2_U2888) );
  AOI22_X1 U21869 ( .A1(n18882), .A2(n18881), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n18931), .ZN(n18889) );
  AOI22_X1 U21870 ( .A1(n18884), .A2(BUF2_REG_16__SCAN_IN), .B1(n18883), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n18888) );
  AOI22_X1 U21871 ( .A1(n18886), .A2(n18890), .B1(n18932), .B2(n18885), .ZN(
        n18887) );
  NAND3_X1 U21872 ( .A1(n18889), .A2(n18888), .A3(n18887), .ZN(P2_U2903) );
  INV_X1 U21873 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n18980) );
  AOI22_X1 U21874 ( .A1(n18892), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18891), .ZN(n19047) );
  OAI222_X1 U21875 ( .A1(n18893), .A2(n18920), .B1(n18980), .B2(n18922), .C1(
        n19047), .C2(n18940), .ZN(P2_U2904) );
  AOI22_X1 U21876 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n18931), .B1(n18894), 
        .B2(n18913), .ZN(n18895) );
  OAI21_X1 U21877 ( .B1(n18920), .B2(n18896), .A(n18895), .ZN(P2_U2905) );
  INV_X1 U21878 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20715) );
  OAI222_X1 U21879 ( .A1(n18897), .A2(n18920), .B1(n20715), .B2(n18922), .C1(
        n18940), .C2(n19042), .ZN(P2_U2906) );
  AOI22_X1 U21880 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n18931), .B1(n18898), 
        .B2(n18913), .ZN(n18899) );
  OAI21_X1 U21881 ( .B1(n18920), .B2(n18900), .A(n18899), .ZN(P2_U2907) );
  INV_X1 U21882 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18987) );
  OAI222_X1 U21883 ( .A1(n18901), .A2(n18920), .B1(n18987), .B2(n18922), .C1(
        n18940), .C2(n19040), .ZN(P2_U2908) );
  AOI22_X1 U21884 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n18931), .B1(n18902), 
        .B2(n18913), .ZN(n18903) );
  OAI21_X1 U21885 ( .B1(n18920), .B2(n18904), .A(n18903), .ZN(P2_U2909) );
  AOI22_X1 U21886 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n18931), .B1(n18905), .B2(
        n18913), .ZN(n18906) );
  OAI21_X1 U21887 ( .B1(n18920), .B2(n18907), .A(n18906), .ZN(P2_U2910) );
  AOI22_X1 U21888 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n18931), .B1(n18908), .B2(
        n18913), .ZN(n18909) );
  OAI21_X1 U21889 ( .B1(n18920), .B2(n18910), .A(n18909), .ZN(P2_U2911) );
  INV_X1 U21890 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18995) );
  OAI222_X1 U21891 ( .A1(n18911), .A2(n18920), .B1(n18995), .B2(n18922), .C1(
        n18940), .C2(n19038), .ZN(P2_U2912) );
  INV_X1 U21892 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18998) );
  OAI222_X1 U21893 ( .A1(n18912), .A2(n18920), .B1(n18998), .B2(n18922), .C1(
        n18940), .C2(n19036), .ZN(P2_U2913) );
  AOI22_X1 U21894 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n18931), .B1(n18914), .B2(
        n18913), .ZN(n18918) );
  OR3_X1 U21895 ( .A1(n18916), .A2(n18915), .A3(n18936), .ZN(n18917) );
  OAI211_X1 U21896 ( .C1(n18920), .C2(n18919), .A(n18918), .B(n18917), .ZN(
        P2_U2914) );
  INV_X1 U21897 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18921) );
  OAI22_X1 U21898 ( .A1(n19676), .A2(n18923), .B1(n18922), .B2(n18921), .ZN(
        n18924) );
  INV_X1 U21899 ( .A(n18924), .ZN(n18930) );
  AOI21_X1 U21900 ( .B1(n18927), .B2(n18926), .A(n18925), .ZN(n18928) );
  OR2_X1 U21901 ( .A1(n18928), .A2(n18936), .ZN(n18929) );
  OAI211_X1 U21902 ( .C1(n19030), .C2(n18940), .A(n18930), .B(n18929), .ZN(
        P2_U2916) );
  AOI22_X1 U21903 ( .A1(n19694), .A2(n18932), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n18931), .ZN(n18939) );
  AOI21_X1 U21904 ( .B1(n18935), .B2(n18934), .A(n18933), .ZN(n18937) );
  OR2_X1 U21905 ( .A1(n18937), .A2(n18936), .ZN(n18938) );
  OAI211_X1 U21906 ( .C1(n19026), .C2(n18940), .A(n18939), .B(n18938), .ZN(
        P2_U2918) );
  NAND3_X1 U21907 ( .A1(n18942), .A2(n18941), .A3(n19720), .ZN(n18944) );
  NAND2_X1 U21908 ( .A1(n18944), .A2(n18943), .ZN(n18945) );
  NOR2_X4 U21909 ( .A1(n18988), .A2(n18978), .ZN(n18996) );
  AND2_X1 U21910 ( .A1(n18996), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  INV_X1 U21911 ( .A(n18946), .ZN(n18947) );
  AOI22_X1 U21912 ( .A1(n18988), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n18948) );
  OAI21_X1 U21913 ( .B1(n12972), .B2(n18976), .A(n18948), .ZN(P2_U2921) );
  AOI22_X1 U21914 ( .A1(n18988), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n18949) );
  OAI21_X1 U21915 ( .B1(n18950), .B2(n18976), .A(n18949), .ZN(P2_U2922) );
  AOI22_X1 U21916 ( .A1(n18988), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n18951) );
  OAI21_X1 U21917 ( .B1(n18952), .B2(n18976), .A(n18951), .ZN(P2_U2923) );
  AOI22_X1 U21918 ( .A1(n18988), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n18953) );
  OAI21_X1 U21919 ( .B1(n18954), .B2(n18976), .A(n18953), .ZN(P2_U2924) );
  AOI22_X1 U21920 ( .A1(n18988), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n18955) );
  OAI21_X1 U21921 ( .B1(n18956), .B2(n18976), .A(n18955), .ZN(P2_U2925) );
  AOI22_X1 U21922 ( .A1(n18988), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n18957) );
  OAI21_X1 U21923 ( .B1(n18958), .B2(n18976), .A(n18957), .ZN(P2_U2926) );
  AOI22_X1 U21924 ( .A1(n18988), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n18959) );
  OAI21_X1 U21925 ( .B1(n18960), .B2(n18976), .A(n18959), .ZN(P2_U2927) );
  AOI22_X1 U21926 ( .A1(n18988), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n18961) );
  OAI21_X1 U21927 ( .B1(n18962), .B2(n18976), .A(n18961), .ZN(P2_U2928) );
  INV_X1 U21928 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n18964) );
  AOI22_X1 U21929 ( .A1(n18988), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n18963) );
  OAI21_X1 U21930 ( .B1(n18964), .B2(n18976), .A(n18963), .ZN(P2_U2929) );
  AOI22_X1 U21931 ( .A1(n18988), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n18965) );
  OAI21_X1 U21932 ( .B1(n18966), .B2(n18976), .A(n18965), .ZN(P2_U2930) );
  INV_X1 U21933 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n18968) );
  AOI22_X1 U21934 ( .A1(n18988), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n18967) );
  OAI21_X1 U21935 ( .B1(n18968), .B2(n18976), .A(n18967), .ZN(P2_U2931) );
  AOI22_X1 U21936 ( .A1(n18988), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n18969) );
  OAI21_X1 U21937 ( .B1(n18970), .B2(n18976), .A(n18969), .ZN(P2_U2932) );
  INV_X1 U21938 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n18972) );
  AOI22_X1 U21939 ( .A1(n18988), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n18971) );
  OAI21_X1 U21940 ( .B1(n18972), .B2(n18976), .A(n18971), .ZN(P2_U2933) );
  AOI22_X1 U21941 ( .A1(n18988), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n18973) );
  OAI21_X1 U21942 ( .B1(n18974), .B2(n18976), .A(n18973), .ZN(P2_U2934) );
  INV_X1 U21943 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n18977) );
  AOI22_X1 U21944 ( .A1(n18988), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n18975) );
  OAI21_X1 U21945 ( .B1(n18977), .B2(n18976), .A(n18975), .ZN(P2_U2935) );
  AOI22_X1 U21946 ( .A1(n18988), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18979) );
  OAI21_X1 U21947 ( .B1(n18980), .B2(n19010), .A(n18979), .ZN(P2_U2936) );
  AOI22_X1 U21948 ( .A1(n18988), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18981) );
  OAI21_X1 U21949 ( .B1(n18982), .B2(n19010), .A(n18981), .ZN(P2_U2937) );
  AOI22_X1 U21950 ( .A1(n18988), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18983) );
  OAI21_X1 U21951 ( .B1(n20715), .B2(n19010), .A(n18983), .ZN(P2_U2938) );
  AOI22_X1 U21952 ( .A1(n18988), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18984) );
  OAI21_X1 U21953 ( .B1(n18985), .B2(n19010), .A(n18984), .ZN(P2_U2939) );
  AOI22_X1 U21954 ( .A1(n18988), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18986) );
  OAI21_X1 U21955 ( .B1(n18987), .B2(n19010), .A(n18986), .ZN(P2_U2940) );
  AOI22_X1 U21956 ( .A1(n18988), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18989) );
  OAI21_X1 U21957 ( .B1(n20697), .B2(n19010), .A(n18989), .ZN(P2_U2941) );
  AOI22_X1 U21958 ( .A1(n19008), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18990) );
  OAI21_X1 U21959 ( .B1(n18991), .B2(n19010), .A(n18990), .ZN(P2_U2942) );
  AOI22_X1 U21960 ( .A1(n19008), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18992) );
  OAI21_X1 U21961 ( .B1(n18993), .B2(n19010), .A(n18992), .ZN(P2_U2943) );
  AOI22_X1 U21962 ( .A1(n19008), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18994) );
  OAI21_X1 U21963 ( .B1(n18995), .B2(n19010), .A(n18994), .ZN(P2_U2944) );
  AOI22_X1 U21964 ( .A1(n19008), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18997) );
  OAI21_X1 U21965 ( .B1(n18998), .B2(n19010), .A(n18997), .ZN(P2_U2945) );
  INV_X1 U21966 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19000) );
  AOI22_X1 U21967 ( .A1(n19008), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18999) );
  OAI21_X1 U21968 ( .B1(n19000), .B2(n19010), .A(n18999), .ZN(P2_U2946) );
  INV_X1 U21969 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19002) );
  AOI22_X1 U21970 ( .A1(n19008), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19001) );
  OAI21_X1 U21971 ( .B1(n19002), .B2(n19010), .A(n19001), .ZN(P2_U2947) );
  AOI22_X1 U21972 ( .A1(n19008), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19003) );
  OAI21_X1 U21973 ( .B1(n18921), .B2(n19010), .A(n19003), .ZN(P2_U2948) );
  AOI22_X1 U21974 ( .A1(n19008), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19004) );
  OAI21_X1 U21975 ( .B1(n19005), .B2(n19010), .A(n19004), .ZN(P2_U2949) );
  AOI22_X1 U21976 ( .A1(n19008), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19006) );
  OAI21_X1 U21977 ( .B1(n19007), .B2(n19010), .A(n19006), .ZN(P2_U2950) );
  INV_X1 U21978 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19011) );
  AOI22_X1 U21979 ( .A1(n19008), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18996), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19009) );
  OAI21_X1 U21980 ( .B1(n19011), .B2(n19010), .A(n19009), .ZN(P2_U2951) );
  AOI22_X1 U21981 ( .A1(n19016), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19043), .ZN(n19012) );
  OAI21_X1 U21982 ( .B1(n19024), .B2(n19046), .A(n19012), .ZN(P2_U2952) );
  AOI22_X1 U21983 ( .A1(n19016), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19043), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n19013) );
  OAI21_X1 U21984 ( .B1(n19026), .B2(n19046), .A(n19013), .ZN(P2_U2953) );
  AOI22_X1 U21985 ( .A1(n19016), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19043), .ZN(n19014) );
  OAI21_X1 U21986 ( .B1(n19028), .B2(n19046), .A(n19014), .ZN(P2_U2954) );
  AOI22_X1 U21987 ( .A1(n19016), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19043), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n19015) );
  OAI21_X1 U21988 ( .B1(n19030), .B2(n19046), .A(n19015), .ZN(P2_U2955) );
  AOI22_X1 U21989 ( .A1(n19016), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19043), .ZN(n19017) );
  OAI21_X1 U21990 ( .B1(n19032), .B2(n19046), .A(n19017), .ZN(P2_U2956) );
  AOI22_X1 U21991 ( .A1(n19044), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19043), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n19018) );
  OAI21_X1 U21992 ( .B1(n19034), .B2(n19046), .A(n19018), .ZN(P2_U2957) );
  AOI22_X1 U21993 ( .A1(n19044), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19043), .ZN(n19019) );
  OAI21_X1 U21994 ( .B1(n19036), .B2(n19046), .A(n19019), .ZN(P2_U2958) );
  AOI22_X1 U21995 ( .A1(n19044), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19043), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n19020) );
  OAI21_X1 U21996 ( .B1(n19038), .B2(n19046), .A(n19020), .ZN(P2_U2959) );
  AOI22_X1 U21997 ( .A1(n19016), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19043), .ZN(n19021) );
  OAI21_X1 U21998 ( .B1(n19040), .B2(n19046), .A(n19021), .ZN(P2_U2963) );
  AOI22_X1 U21999 ( .A1(n19044), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19043), .ZN(n19022) );
  OAI21_X1 U22000 ( .B1(n19042), .B2(n19046), .A(n19022), .ZN(P2_U2965) );
  AOI22_X1 U22001 ( .A1(n19016), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19043), .ZN(n19023) );
  OAI21_X1 U22002 ( .B1(n19024), .B2(n19046), .A(n19023), .ZN(P2_U2967) );
  AOI22_X1 U22003 ( .A1(n19016), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19043), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n19025) );
  OAI21_X1 U22004 ( .B1(n19026), .B2(n19046), .A(n19025), .ZN(P2_U2968) );
  AOI22_X1 U22005 ( .A1(n19044), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19043), .ZN(n19027) );
  OAI21_X1 U22006 ( .B1(n19028), .B2(n19046), .A(n19027), .ZN(P2_U2969) );
  AOI22_X1 U22007 ( .A1(n19044), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19043), .ZN(n19029) );
  OAI21_X1 U22008 ( .B1(n19030), .B2(n19046), .A(n19029), .ZN(P2_U2970) );
  AOI22_X1 U22009 ( .A1(n19044), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19043), .ZN(n19031) );
  OAI21_X1 U22010 ( .B1(n19032), .B2(n19046), .A(n19031), .ZN(P2_U2971) );
  AOI22_X1 U22011 ( .A1(n19044), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n19043), .ZN(n19033) );
  OAI21_X1 U22012 ( .B1(n19034), .B2(n19046), .A(n19033), .ZN(P2_U2972) );
  AOI22_X1 U22013 ( .A1(n19044), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19043), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n19035) );
  OAI21_X1 U22014 ( .B1(n19036), .B2(n19046), .A(n19035), .ZN(P2_U2973) );
  AOI22_X1 U22015 ( .A1(n19044), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19043), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n19037) );
  OAI21_X1 U22016 ( .B1(n19038), .B2(n19046), .A(n19037), .ZN(P2_U2974) );
  AOI22_X1 U22017 ( .A1(n19044), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n19043), .ZN(n19039) );
  OAI21_X1 U22018 ( .B1(n19040), .B2(n19046), .A(n19039), .ZN(P2_U2978) );
  AOI22_X1 U22019 ( .A1(n19044), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19043), .ZN(n19041) );
  OAI21_X1 U22020 ( .B1(n19042), .B2(n19046), .A(n19041), .ZN(P2_U2980) );
  AOI22_X1 U22021 ( .A1(n19044), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(
        P2_EAX_REG_15__SCAN_IN), .B2(n19043), .ZN(n19045) );
  OAI21_X1 U22022 ( .B1(n19047), .B2(n19046), .A(n19045), .ZN(P2_U2982) );
  AOI22_X1 U22023 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n15127), .B1(n19049), 
        .B2(n19048), .ZN(n19060) );
  NAND2_X1 U22024 ( .A1(n19051), .A2(n19050), .ZN(n19055) );
  NAND2_X1 U22025 ( .A1(n19053), .A2(n19052), .ZN(n19054) );
  OAI211_X1 U22026 ( .C1(n19057), .C2(n19056), .A(n19055), .B(n19054), .ZN(
        n19058) );
  INV_X1 U22027 ( .A(n19058), .ZN(n19059) );
  OAI211_X1 U22028 ( .C1(n19061), .C2(n20762), .A(n19060), .B(n19059), .ZN(
        P2_U3010) );
  AOI22_X1 U22029 ( .A1(n19525), .A2(n19554), .B1(n19074), .B2(n19465), .ZN(
        n19063) );
  AOI22_X1 U22030 ( .A1(n19466), .A2(n19075), .B1(n19104), .B2(n19142), .ZN(
        n19062) );
  OAI211_X1 U22031 ( .C1(n19065), .C2(n19064), .A(n19063), .B(n19062), .ZN(
        P2_U3049) );
  INV_X1 U22032 ( .A(n19478), .ZN(n19539) );
  AOI22_X1 U22033 ( .A1(n19539), .A2(n19554), .B1(n19074), .B2(n19473), .ZN(
        n19067) );
  AOI22_X1 U22034 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19076), .B1(
        n19475), .B2(n19075), .ZN(n19066) );
  OAI211_X1 U22035 ( .C1(n19542), .C2(n19095), .A(n19067), .B(n19066), .ZN(
        P2_U3051) );
  AOI22_X1 U22036 ( .A1(n19546), .A2(n19554), .B1(n19074), .B2(n19479), .ZN(
        n19069) );
  AOI22_X1 U22037 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19076), .B1(
        n19481), .B2(n19075), .ZN(n19068) );
  OAI211_X1 U22038 ( .C1(n19549), .C2(n19095), .A(n19069), .B(n19068), .ZN(
        P2_U3052) );
  INV_X1 U22039 ( .A(n19558), .ZN(n19487) );
  AOI22_X1 U22040 ( .A1(n19487), .A2(n19554), .B1(n19074), .B2(n19486), .ZN(
        n19071) );
  AOI22_X1 U22041 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19076), .B1(
        n19488), .B2(n19075), .ZN(n19070) );
  OAI211_X1 U22042 ( .C1(n19491), .C2(n19095), .A(n19071), .B(n19070), .ZN(
        P2_U3053) );
  AOI22_X1 U22043 ( .A1(n19562), .A2(n19554), .B1(n19074), .B2(n19492), .ZN(
        n19073) );
  AOI22_X1 U22044 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19076), .B1(
        n19493), .B2(n19075), .ZN(n19072) );
  OAI211_X1 U22045 ( .C1(n19565), .C2(n19095), .A(n19073), .B(n19072), .ZN(
        P2_U3054) );
  AOI22_X1 U22046 ( .A1(n19571), .A2(n19554), .B1(n19074), .B2(n19497), .ZN(
        n19078) );
  AOI22_X1 U22047 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19076), .B1(
        n19500), .B2(n19075), .ZN(n19077) );
  OAI211_X1 U22048 ( .C1(n19577), .C2(n19095), .A(n19078), .B(n19077), .ZN(
        P2_U3055) );
  INV_X1 U22049 ( .A(n19079), .ZN(n19080) );
  NOR2_X1 U22050 ( .A1(n19200), .A2(n19131), .ZN(n19102) );
  NOR2_X1 U22051 ( .A1(n19080), .A2(n19102), .ZN(n19085) );
  NOR2_X1 U22052 ( .A1(n19131), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19082) );
  INV_X1 U22053 ( .A(n19082), .ZN(n19081) );
  OAI22_X1 U22054 ( .A1(n19085), .A2(n19504), .B1(n19081), .B2(n19454), .ZN(
        n19103) );
  AOI22_X1 U22055 ( .A1(n19103), .A2(n19462), .B1(n19451), .B2(n19102), .ZN(
        n19088) );
  INV_X1 U22056 ( .A(n19201), .ZN(n19674) );
  AOI21_X1 U22057 ( .B1(n19674), .B2(n19083), .A(n19082), .ZN(n19084) );
  AOI211_X1 U22058 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19085), .A(n19392), 
        .B(n19084), .ZN(n19086) );
  AOI22_X1 U22059 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19105), .B1(
        n19126), .B2(n19518), .ZN(n19087) );
  OAI211_X1 U22060 ( .C1(n19521), .C2(n19095), .A(n19088), .B(n19087), .ZN(
        P2_U3056) );
  AOI22_X1 U22061 ( .A1(n19103), .A2(n19466), .B1(n19465), .B2(n19102), .ZN(
        n19090) );
  AOI22_X1 U22062 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19525), .ZN(n19089) );
  OAI211_X1 U22063 ( .C1(n19528), .C2(n19108), .A(n19090), .B(n19089), .ZN(
        P2_U3057) );
  AOI22_X1 U22064 ( .A1(n19103), .A2(n19470), .B1(n19469), .B2(n19102), .ZN(
        n19092) );
  AOI22_X1 U22065 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19532), .ZN(n19091) );
  OAI211_X1 U22066 ( .C1(n19535), .C2(n19108), .A(n19092), .B(n19091), .ZN(
        P2_U3058) );
  AOI22_X1 U22067 ( .A1(n19103), .A2(n19475), .B1(n19473), .B2(n19102), .ZN(
        n19094) );
  AOI22_X1 U22068 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19105), .B1(
        n19126), .B2(n19474), .ZN(n19093) );
  OAI211_X1 U22069 ( .C1(n19478), .C2(n19095), .A(n19094), .B(n19093), .ZN(
        P2_U3059) );
  AOI22_X1 U22070 ( .A1(n19103), .A2(n19481), .B1(n19479), .B2(n19102), .ZN(
        n19097) );
  AOI22_X1 U22071 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19546), .ZN(n19096) );
  OAI211_X1 U22072 ( .C1(n19549), .C2(n19108), .A(n19097), .B(n19096), .ZN(
        P2_U3060) );
  AOI22_X1 U22073 ( .A1(n19103), .A2(n19488), .B1(n19486), .B2(n19102), .ZN(
        n19099) );
  AOI22_X1 U22074 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19487), .ZN(n19098) );
  OAI211_X1 U22075 ( .C1(n19491), .C2(n19108), .A(n19099), .B(n19098), .ZN(
        P2_U3061) );
  AOI22_X1 U22076 ( .A1(n19103), .A2(n19493), .B1(n19492), .B2(n19102), .ZN(
        n19101) );
  AOI22_X1 U22077 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19562), .ZN(n19100) );
  OAI211_X1 U22078 ( .C1(n19565), .C2(n19108), .A(n19101), .B(n19100), .ZN(
        P2_U3062) );
  AOI22_X1 U22079 ( .A1(n19103), .A2(n19500), .B1(n19497), .B2(n19102), .ZN(
        n19107) );
  AOI22_X1 U22080 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19571), .ZN(n19106) );
  OAI211_X1 U22081 ( .C1(n19577), .C2(n19108), .A(n19107), .B(n19106), .ZN(
        P2_U3063) );
  AOI22_X1 U22082 ( .A1(n19125), .A2(n19466), .B1(n19124), .B2(n19465), .ZN(
        n19110) );
  AOI22_X1 U22083 ( .A1(n19126), .A2(n19525), .B1(n19157), .B2(n19142), .ZN(
        n19109) );
  OAI211_X1 U22084 ( .C1(n19130), .C2(n10228), .A(n19110), .B(n19109), .ZN(
        P2_U3065) );
  INV_X1 U22085 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n19113) );
  AOI22_X1 U22086 ( .A1(n19125), .A2(n19470), .B1(n19124), .B2(n19469), .ZN(
        n19112) );
  AOI22_X1 U22087 ( .A1(n19126), .A2(n19532), .B1(n19157), .B2(n19145), .ZN(
        n19111) );
  OAI211_X1 U22088 ( .C1(n19130), .C2(n19113), .A(n19112), .B(n19111), .ZN(
        P2_U3066) );
  AOI22_X1 U22089 ( .A1(n19125), .A2(n19475), .B1(n19124), .B2(n19473), .ZN(
        n19115) );
  AOI22_X1 U22090 ( .A1(n19126), .A2(n19539), .B1(n19157), .B2(n19474), .ZN(
        n19114) );
  OAI211_X1 U22091 ( .C1(n19130), .C2(n10284), .A(n19115), .B(n19114), .ZN(
        P2_U3067) );
  INV_X1 U22092 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n19118) );
  AOI22_X1 U22093 ( .A1(n19125), .A2(n19481), .B1(n19124), .B2(n19479), .ZN(
        n19117) );
  INV_X1 U22094 ( .A(n19549), .ZN(n19480) );
  AOI22_X1 U22095 ( .A1(n19157), .A2(n19480), .B1(n19126), .B2(n19546), .ZN(
        n19116) );
  OAI211_X1 U22096 ( .C1(n19130), .C2(n19118), .A(n19117), .B(n19116), .ZN(
        P2_U3068) );
  AOI22_X1 U22097 ( .A1(n19125), .A2(n19488), .B1(n19124), .B2(n19486), .ZN(
        n19120) );
  AOI22_X1 U22098 ( .A1(n19157), .A2(n19553), .B1(n19126), .B2(n19487), .ZN(
        n19119) );
  OAI211_X1 U22099 ( .C1(n19130), .C2(n10391), .A(n19120), .B(n19119), .ZN(
        P2_U3069) );
  AOI22_X1 U22100 ( .A1(n19125), .A2(n19493), .B1(n19124), .B2(n19492), .ZN(
        n19122) );
  AOI22_X1 U22101 ( .A1(n19126), .A2(n19562), .B1(n19157), .B2(n19408), .ZN(
        n19121) );
  OAI211_X1 U22102 ( .C1(n19130), .C2(n19123), .A(n19122), .B(n19121), .ZN(
        P2_U3070) );
  INV_X1 U22103 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19129) );
  AOI22_X1 U22104 ( .A1(n19125), .A2(n19500), .B1(n19124), .B2(n19497), .ZN(
        n19128) );
  AOI22_X1 U22105 ( .A1(n19126), .A2(n19571), .B1(n19157), .B2(n19158), .ZN(
        n19127) );
  OAI211_X1 U22106 ( .C1(n19130), .C2(n19129), .A(n19128), .B(n19127), .ZN(
        P2_U3071) );
  AOI21_X1 U22107 ( .B1(n19674), .B2(n19358), .A(n19454), .ZN(n19134) );
  NOR2_X1 U22108 ( .A1(n19696), .A2(n19131), .ZN(n19138) );
  NOR2_X1 U22109 ( .A1(n19347), .A2(n19131), .ZN(n19156) );
  INV_X1 U22110 ( .A(n19156), .ZN(n19135) );
  AOI21_X1 U22111 ( .B1(n19132), .B2(n19135), .A(n19504), .ZN(n19133) );
  AOI22_X1 U22112 ( .A1(n19157), .A2(n19323), .B1(n19451), .B2(n19156), .ZN(
        n19141) );
  INV_X1 U22113 ( .A(n19134), .ZN(n19139) );
  AOI21_X1 U22114 ( .B1(n19136), .B2(n19135), .A(n19392), .ZN(n19137) );
  AOI22_X1 U22115 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19159), .B1(
        n19195), .B2(n19518), .ZN(n19140) );
  OAI211_X1 U22116 ( .C1(n19162), .C2(n19509), .A(n19141), .B(n19140), .ZN(
        P2_U3072) );
  AOI22_X1 U22117 ( .A1(n19142), .A2(n19195), .B1(n19465), .B2(n19156), .ZN(
        n19144) );
  AOI22_X1 U22118 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19159), .B1(
        n19157), .B2(n19525), .ZN(n19143) );
  OAI211_X1 U22119 ( .C1(n19162), .C2(n19523), .A(n19144), .B(n19143), .ZN(
        P2_U3073) );
  AOI22_X1 U22120 ( .A1(n19145), .A2(n19195), .B1(n19469), .B2(n19156), .ZN(
        n19147) );
  AOI22_X1 U22121 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19159), .B1(
        n19157), .B2(n19532), .ZN(n19146) );
  OAI211_X1 U22122 ( .C1(n19162), .C2(n19530), .A(n19147), .B(n19146), .ZN(
        P2_U3074) );
  AOI22_X1 U22123 ( .A1(n19157), .A2(n19539), .B1(n19473), .B2(n19156), .ZN(
        n19149) );
  AOI22_X1 U22124 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19159), .B1(
        n19195), .B2(n19474), .ZN(n19148) );
  OAI211_X1 U22125 ( .C1(n19162), .C2(n19537), .A(n19149), .B(n19148), .ZN(
        P2_U3075) );
  AOI22_X1 U22126 ( .A1(n19480), .A2(n19195), .B1(n19479), .B2(n19156), .ZN(
        n19151) );
  AOI22_X1 U22127 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19159), .B1(
        n19157), .B2(n19546), .ZN(n19150) );
  OAI211_X1 U22128 ( .C1(n19162), .C2(n19544), .A(n19151), .B(n19150), .ZN(
        P2_U3076) );
  AOI22_X1 U22129 ( .A1(n19157), .A2(n19487), .B1(n19486), .B2(n19156), .ZN(
        n19153) );
  AOI22_X1 U22130 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19159), .B1(
        n19195), .B2(n19553), .ZN(n19152) );
  OAI211_X1 U22131 ( .C1(n19162), .C2(n19551), .A(n19153), .B(n19152), .ZN(
        P2_U3077) );
  AOI22_X1 U22132 ( .A1(n19157), .A2(n19562), .B1(n19492), .B2(n19156), .ZN(
        n19155) );
  AOI22_X1 U22133 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19159), .B1(
        n19195), .B2(n19408), .ZN(n19154) );
  OAI211_X1 U22134 ( .C1(n19162), .C2(n19560), .A(n19155), .B(n19154), .ZN(
        P2_U3078) );
  AOI22_X1 U22135 ( .A1(n19571), .A2(n19157), .B1(n19497), .B2(n19156), .ZN(
        n19161) );
  AOI22_X1 U22136 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19159), .B1(
        n19195), .B2(n19158), .ZN(n19160) );
  OAI211_X1 U22137 ( .C1(n19162), .C2(n19568), .A(n19161), .B(n19160), .ZN(
        P2_U3079) );
  INV_X1 U22138 ( .A(n19163), .ZN(n19389) );
  NAND2_X1 U22139 ( .A1(n19680), .A2(n19389), .ZN(n19174) );
  INV_X1 U22140 ( .A(n19164), .ZN(n19168) );
  INV_X1 U22141 ( .A(n19170), .ZN(n19166) );
  NAND2_X1 U22142 ( .A1(n19165), .A2(n19696), .ZN(n19207) );
  NOR2_X1 U22143 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19207), .ZN(
        n19193) );
  OAI21_X1 U22144 ( .B1(n19166), .B2(n19193), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19167) );
  OAI21_X1 U22145 ( .B1(n19174), .B2(n19168), .A(n19167), .ZN(n19194) );
  AOI22_X1 U22146 ( .A1(n19194), .A2(n19462), .B1(n19451), .B2(n19193), .ZN(
        n19179) );
  INV_X1 U22147 ( .A(n19193), .ZN(n19169) );
  OAI211_X1 U22148 ( .C1(n19170), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19169), 
        .B(n19454), .ZN(n19177) );
  INV_X1 U22149 ( .A(n19390), .ZN(n19175) );
  OAI21_X1 U22150 ( .B1(n19195), .B2(n19225), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19173) );
  OAI21_X1 U22151 ( .B1(n19175), .B2(n19174), .A(n19173), .ZN(n19176) );
  NAND3_X1 U22152 ( .A1(n19177), .A2(n19515), .A3(n19176), .ZN(n19196) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19196), .B1(
        n19225), .B2(n19518), .ZN(n19178) );
  OAI211_X1 U22154 ( .C1(n19521), .C2(n19190), .A(n19179), .B(n19178), .ZN(
        P2_U3080) );
  AOI22_X1 U22155 ( .A1(n19194), .A2(n19466), .B1(n19465), .B2(n19193), .ZN(
        n19181) );
  AOI22_X1 U22156 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19196), .B1(
        n19195), .B2(n19525), .ZN(n19180) );
  OAI211_X1 U22157 ( .C1(n19528), .C2(n19223), .A(n19181), .B(n19180), .ZN(
        P2_U3081) );
  AOI22_X1 U22158 ( .A1(n19194), .A2(n19470), .B1(n19469), .B2(n19193), .ZN(
        n19183) );
  AOI22_X1 U22159 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19196), .B1(
        n19195), .B2(n19532), .ZN(n19182) );
  OAI211_X1 U22160 ( .C1(n19535), .C2(n19223), .A(n19183), .B(n19182), .ZN(
        P2_U3082) );
  AOI22_X1 U22161 ( .A1(n19194), .A2(n19475), .B1(n19473), .B2(n19193), .ZN(
        n19185) );
  AOI22_X1 U22162 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19196), .B1(
        n19225), .B2(n19474), .ZN(n19184) );
  OAI211_X1 U22163 ( .C1(n19478), .C2(n19190), .A(n19185), .B(n19184), .ZN(
        P2_U3083) );
  AOI22_X1 U22164 ( .A1(n19194), .A2(n19481), .B1(n19479), .B2(n19193), .ZN(
        n19187) );
  AOI22_X1 U22165 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19196), .B1(
        n19225), .B2(n19480), .ZN(n19186) );
  OAI211_X1 U22166 ( .C1(n19485), .C2(n19190), .A(n19187), .B(n19186), .ZN(
        P2_U3084) );
  AOI22_X1 U22167 ( .A1(n19194), .A2(n19488), .B1(n19486), .B2(n19193), .ZN(
        n19189) );
  AOI22_X1 U22168 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19196), .B1(
        n19225), .B2(n19553), .ZN(n19188) );
  OAI211_X1 U22169 ( .C1(n19558), .C2(n19190), .A(n19189), .B(n19188), .ZN(
        P2_U3085) );
  AOI22_X1 U22170 ( .A1(n19194), .A2(n19493), .B1(n19492), .B2(n19193), .ZN(
        n19192) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19196), .B1(
        n19195), .B2(n19562), .ZN(n19191) );
  OAI211_X1 U22172 ( .C1(n19565), .C2(n19223), .A(n19192), .B(n19191), .ZN(
        P2_U3086) );
  AOI22_X1 U22173 ( .A1(n19194), .A2(n19500), .B1(n19497), .B2(n19193), .ZN(
        n19198) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19196), .B1(
        n19195), .B2(n19571), .ZN(n19197) );
  OAI211_X1 U22175 ( .C1(n19577), .C2(n19223), .A(n19198), .B(n19197), .ZN(
        P2_U3087) );
  NOR2_X1 U22176 ( .A1(n19200), .A2(n19234), .ZN(n19224) );
  AOI22_X1 U22177 ( .A1(n19518), .A2(n19254), .B1(n19451), .B2(n19224), .ZN(
        n19210) );
  OR2_X1 U22178 ( .A1(n19201), .A2(n19422), .ZN(n19202) );
  NAND2_X1 U22179 ( .A1(n19202), .A2(n19681), .ZN(n19208) );
  INV_X1 U22180 ( .A(n19208), .ZN(n19204) );
  NOR2_X1 U22181 ( .A1(n19203), .A2(n19224), .ZN(n19206) );
  AOI22_X1 U22182 ( .A1(n19204), .A2(n19207), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19206), .ZN(n19205) );
  OAI211_X1 U22183 ( .C1(n19224), .C2(n19697), .A(n19205), .B(n19515), .ZN(
        n19227) );
  OAI22_X1 U22184 ( .A1(n19208), .A2(n19207), .B1(n19206), .B2(n19504), .ZN(
        n19226) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19227), .B1(
        n19462), .B2(n19226), .ZN(n19209) );
  OAI211_X1 U22186 ( .C1(n19521), .C2(n19223), .A(n19210), .B(n19209), .ZN(
        P2_U3088) );
  AOI22_X1 U22187 ( .A1(n19525), .A2(n19225), .B1(n19465), .B2(n19224), .ZN(
        n19212) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19227), .B1(
        n19466), .B2(n19226), .ZN(n19211) );
  OAI211_X1 U22189 ( .C1(n19528), .C2(n19249), .A(n19212), .B(n19211), .ZN(
        P2_U3089) );
  AOI22_X1 U22190 ( .A1(n19532), .A2(n19225), .B1(n19469), .B2(n19224), .ZN(
        n19214) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19227), .B1(
        n19470), .B2(n19226), .ZN(n19213) );
  OAI211_X1 U22192 ( .C1(n19535), .C2(n19249), .A(n19214), .B(n19213), .ZN(
        P2_U3090) );
  AOI22_X1 U22193 ( .A1(n19474), .A2(n19254), .B1(n19473), .B2(n19224), .ZN(
        n19216) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19227), .B1(
        n19475), .B2(n19226), .ZN(n19215) );
  OAI211_X1 U22195 ( .C1(n19478), .C2(n19223), .A(n19216), .B(n19215), .ZN(
        P2_U3091) );
  AOI22_X1 U22196 ( .A1(n19225), .A2(n19546), .B1(n19479), .B2(n19224), .ZN(
        n19218) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19227), .B1(
        n19481), .B2(n19226), .ZN(n19217) );
  OAI211_X1 U22198 ( .C1(n19549), .C2(n19249), .A(n19218), .B(n19217), .ZN(
        P2_U3092) );
  AOI22_X1 U22199 ( .A1(n19225), .A2(n19487), .B1(n19486), .B2(n19224), .ZN(
        n19220) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19227), .B1(
        n19488), .B2(n19226), .ZN(n19219) );
  OAI211_X1 U22201 ( .C1(n19491), .C2(n19249), .A(n19220), .B(n19219), .ZN(
        P2_U3093) );
  AOI22_X1 U22202 ( .A1(n19408), .A2(n19254), .B1(n19492), .B2(n19224), .ZN(
        n19222) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19227), .B1(
        n19493), .B2(n19226), .ZN(n19221) );
  OAI211_X1 U22204 ( .C1(n19412), .C2(n19223), .A(n19222), .B(n19221), .ZN(
        P2_U3094) );
  AOI22_X1 U22205 ( .A1(n19571), .A2(n19225), .B1(n19497), .B2(n19224), .ZN(
        n19229) );
  AOI22_X1 U22206 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19227), .B1(
        n19500), .B2(n19226), .ZN(n19228) );
  OAI211_X1 U22207 ( .C1(n19577), .C2(n19249), .A(n19229), .B(n19228), .ZN(
        P2_U3095) );
  NOR2_X1 U22208 ( .A1(n19317), .A2(n19234), .ZN(n19252) );
  OAI21_X1 U22209 ( .B1(n19230), .B2(n19252), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19231) );
  OAI21_X1 U22210 ( .B1(n19234), .B2(n19322), .A(n19231), .ZN(n19253) );
  AOI22_X1 U22211 ( .A1(n19253), .A2(n19462), .B1(n19451), .B2(n19252), .ZN(
        n19238) );
  AOI21_X1 U22212 ( .B1(n19232), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19236) );
  OAI21_X1 U22213 ( .B1(n19254), .B2(n19274), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19233) );
  OAI21_X1 U22214 ( .B1(n19389), .B2(n19234), .A(n19233), .ZN(n19235) );
  OAI211_X1 U22215 ( .C1(n19252), .C2(n19236), .A(n19235), .B(n19515), .ZN(
        n19255) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19255), .B1(
        n19274), .B2(n19518), .ZN(n19237) );
  OAI211_X1 U22217 ( .C1(n19521), .C2(n19249), .A(n19238), .B(n19237), .ZN(
        P2_U3096) );
  AOI22_X1 U22218 ( .A1(n19253), .A2(n19466), .B1(n19465), .B2(n19252), .ZN(
        n19240) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19525), .ZN(n19239) );
  OAI211_X1 U22220 ( .C1(n19528), .C2(n19270), .A(n19240), .B(n19239), .ZN(
        P2_U3097) );
  AOI22_X1 U22221 ( .A1(n19253), .A2(n19470), .B1(n19469), .B2(n19252), .ZN(
        n19242) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19532), .ZN(n19241) );
  OAI211_X1 U22223 ( .C1(n19535), .C2(n19270), .A(n19242), .B(n19241), .ZN(
        P2_U3098) );
  AOI22_X1 U22224 ( .A1(n19253), .A2(n19475), .B1(n19473), .B2(n19252), .ZN(
        n19244) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19255), .B1(
        n19274), .B2(n19474), .ZN(n19243) );
  OAI211_X1 U22226 ( .C1(n19478), .C2(n19249), .A(n19244), .B(n19243), .ZN(
        P2_U3099) );
  AOI22_X1 U22227 ( .A1(n19253), .A2(n19481), .B1(n19479), .B2(n19252), .ZN(
        n19246) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19546), .ZN(n19245) );
  OAI211_X1 U22229 ( .C1(n19549), .C2(n19270), .A(n19246), .B(n19245), .ZN(
        P2_U3100) );
  AOI22_X1 U22230 ( .A1(n19253), .A2(n19488), .B1(n19486), .B2(n19252), .ZN(
        n19248) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19255), .B1(
        n19274), .B2(n19553), .ZN(n19247) );
  OAI211_X1 U22232 ( .C1(n19558), .C2(n19249), .A(n19248), .B(n19247), .ZN(
        P2_U3101) );
  AOI22_X1 U22233 ( .A1(n19253), .A2(n19493), .B1(n19492), .B2(n19252), .ZN(
        n19251) );
  AOI22_X1 U22234 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19562), .ZN(n19250) );
  OAI211_X1 U22235 ( .C1(n19565), .C2(n19270), .A(n19251), .B(n19250), .ZN(
        P2_U3102) );
  AOI22_X1 U22236 ( .A1(n19253), .A2(n19500), .B1(n19497), .B2(n19252), .ZN(
        n19257) );
  AOI22_X1 U22237 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19255), .B1(
        n19254), .B2(n19571), .ZN(n19256) );
  OAI211_X1 U22238 ( .C1(n19577), .C2(n19270), .A(n19257), .B(n19256), .ZN(
        P2_U3103) );
  AOI22_X1 U22239 ( .A1(n19273), .A2(n19462), .B1(n19451), .B2(n19285), .ZN(
        n19259) );
  AOI22_X1 U22240 ( .A1(n19306), .A2(n19518), .B1(n19274), .B2(n19323), .ZN(
        n19258) );
  OAI211_X1 U22241 ( .C1(n19261), .C2(n19260), .A(n19259), .B(n19258), .ZN(
        P2_U3104) );
  AOI22_X1 U22242 ( .A1(n19273), .A2(n19466), .B1(n19465), .B2(n19285), .ZN(
        n19263) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19275), .B1(
        n19274), .B2(n19525), .ZN(n19262) );
  OAI211_X1 U22244 ( .C1(n19528), .C2(n19302), .A(n19263), .B(n19262), .ZN(
        P2_U3105) );
  AOI22_X1 U22245 ( .A1(n19273), .A2(n19475), .B1(n19473), .B2(n19285), .ZN(
        n19265) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19275), .B1(
        n19274), .B2(n19539), .ZN(n19264) );
  OAI211_X1 U22247 ( .C1(n19542), .C2(n19302), .A(n19265), .B(n19264), .ZN(
        P2_U3107) );
  AOI22_X1 U22248 ( .A1(n19273), .A2(n19481), .B1(n19479), .B2(n19285), .ZN(
        n19267) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19275), .B1(
        n19306), .B2(n19480), .ZN(n19266) );
  OAI211_X1 U22250 ( .C1(n19485), .C2(n19270), .A(n19267), .B(n19266), .ZN(
        P2_U3108) );
  AOI22_X1 U22251 ( .A1(n19273), .A2(n19488), .B1(n19486), .B2(n19285), .ZN(
        n19269) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19275), .B1(
        n19306), .B2(n19553), .ZN(n19268) );
  OAI211_X1 U22253 ( .C1(n19558), .C2(n19270), .A(n19269), .B(n19268), .ZN(
        P2_U3109) );
  AOI22_X1 U22254 ( .A1(n19273), .A2(n19493), .B1(n19492), .B2(n19285), .ZN(
        n19272) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19275), .B1(
        n19274), .B2(n19562), .ZN(n19271) );
  OAI211_X1 U22256 ( .C1(n19565), .C2(n19302), .A(n19272), .B(n19271), .ZN(
        P2_U3110) );
  AOI22_X1 U22257 ( .A1(n19273), .A2(n19500), .B1(n19497), .B2(n19285), .ZN(
        n19277) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19275), .B1(
        n19274), .B2(n19571), .ZN(n19276) );
  OAI211_X1 U22259 ( .C1(n19577), .C2(n19302), .A(n19277), .B(n19276), .ZN(
        P2_U3111) );
  NOR2_X1 U22260 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19278), .ZN(
        n19305) );
  AOI22_X1 U22261 ( .A1(n19518), .A2(n19299), .B1(n19451), .B2(n19305), .ZN(
        n19290) );
  AOI21_X1 U22262 ( .B1(n19302), .B2(n19311), .A(n19668), .ZN(n19279) );
  NOR2_X1 U22263 ( .A1(n19279), .A2(n19454), .ZN(n19284) );
  INV_X1 U22264 ( .A(n19280), .ZN(n19286) );
  AOI21_X1 U22265 ( .B1(n19286), .B2(n19697), .A(n19681), .ZN(n19281) );
  AOI21_X1 U22266 ( .B1(n19284), .B2(n19282), .A(n19281), .ZN(n19283) );
  OAI21_X1 U22267 ( .B1(n19285), .B2(n19305), .A(n19284), .ZN(n19288) );
  OAI21_X1 U22268 ( .B1(n19286), .B2(n19305), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19287) );
  NAND2_X1 U22269 ( .A1(n19288), .A2(n19287), .ZN(n19307) );
  AOI22_X1 U22270 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19308), .B1(
        n19462), .B2(n19307), .ZN(n19289) );
  OAI211_X1 U22271 ( .C1(n19521), .C2(n19302), .A(n19290), .B(n19289), .ZN(
        P2_U3112) );
  AOI22_X1 U22272 ( .A1(n19525), .A2(n19306), .B1(n19465), .B2(n19305), .ZN(
        n19292) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19466), .ZN(n19291) );
  OAI211_X1 U22274 ( .C1(n19528), .C2(n19311), .A(n19292), .B(n19291), .ZN(
        P2_U3113) );
  AOI22_X1 U22275 ( .A1(n19532), .A2(n19306), .B1(n19469), .B2(n19305), .ZN(
        n19294) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19470), .ZN(n19293) );
  OAI211_X1 U22277 ( .C1(n19535), .C2(n19311), .A(n19294), .B(n19293), .ZN(
        P2_U3114) );
  AOI22_X1 U22278 ( .A1(n19539), .A2(n19306), .B1(n19473), .B2(n19305), .ZN(
        n19296) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19475), .ZN(n19295) );
  OAI211_X1 U22280 ( .C1(n19542), .C2(n19311), .A(n19296), .B(n19295), .ZN(
        P2_U3115) );
  AOI22_X1 U22281 ( .A1(n19480), .A2(n19299), .B1(n19479), .B2(n19305), .ZN(
        n19298) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19481), .ZN(n19297) );
  OAI211_X1 U22283 ( .C1(n19485), .C2(n19302), .A(n19298), .B(n19297), .ZN(
        P2_U3116) );
  AOI22_X1 U22284 ( .A1(n19553), .A2(n19299), .B1(n19486), .B2(n19305), .ZN(
        n19301) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19488), .ZN(n19300) );
  OAI211_X1 U22286 ( .C1(n19558), .C2(n19302), .A(n19301), .B(n19300), .ZN(
        P2_U3117) );
  AOI22_X1 U22287 ( .A1(n19306), .A2(n19562), .B1(n19492), .B2(n19305), .ZN(
        n19304) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19493), .ZN(n19303) );
  OAI211_X1 U22289 ( .C1(n19565), .C2(n19311), .A(n19304), .B(n19303), .ZN(
        P2_U3118) );
  AOI22_X1 U22290 ( .A1(n19571), .A2(n19306), .B1(n19497), .B2(n19305), .ZN(
        n19310) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19308), .B1(
        n19307), .B2(n19500), .ZN(n19309) );
  OAI211_X1 U22292 ( .C1(n19577), .C2(n19311), .A(n19310), .B(n19309), .ZN(
        P2_U3119) );
  INV_X1 U22293 ( .A(n19449), .ZN(n19313) );
  AOI21_X1 U22294 ( .B1(n19336), .B2(n19376), .A(n19668), .ZN(n19314) );
  OAI21_X1 U22295 ( .B1(n19315), .B2(n19314), .A(n19697), .ZN(n19316) );
  AOI21_X1 U22296 ( .B1(n10392), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19316), 
        .ZN(n19318) );
  NOR2_X1 U22297 ( .A1(n19317), .A2(n19349), .ZN(n19341) );
  OR2_X1 U22298 ( .A1(n19318), .A2(n19341), .ZN(n19319) );
  AND2_X1 U22299 ( .A1(n19319), .A2(n19515), .ZN(n19327) );
  INV_X1 U22300 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19326) );
  INV_X1 U22301 ( .A(n10392), .ZN(n19320) );
  OAI21_X1 U22302 ( .B1(n19320), .B2(n19341), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19321) );
  OAI21_X1 U22303 ( .B1(n19349), .B2(n19322), .A(n19321), .ZN(n19342) );
  AOI22_X1 U22304 ( .A1(n19342), .A2(n19462), .B1(n19451), .B2(n19341), .ZN(
        n19325) );
  AOI22_X1 U22305 ( .A1(n19383), .A2(n19518), .B1(n19343), .B2(n19323), .ZN(
        n19324) );
  OAI211_X1 U22306 ( .C1(n19327), .C2(n19326), .A(n19325), .B(n19324), .ZN(
        P2_U3128) );
  AOI22_X1 U22307 ( .A1(n19342), .A2(n19466), .B1(n19465), .B2(n19341), .ZN(
        n19329) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19344), .B1(
        n19343), .B2(n19525), .ZN(n19328) );
  OAI211_X1 U22309 ( .C1(n19528), .C2(n19376), .A(n19329), .B(n19328), .ZN(
        P2_U3129) );
  AOI22_X1 U22310 ( .A1(n19342), .A2(n19470), .B1(n19469), .B2(n19341), .ZN(
        n19331) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19344), .B1(
        n19343), .B2(n19532), .ZN(n19330) );
  OAI211_X1 U22312 ( .C1(n19535), .C2(n19376), .A(n19331), .B(n19330), .ZN(
        P2_U3130) );
  AOI22_X1 U22313 ( .A1(n19342), .A2(n19475), .B1(n19473), .B2(n19341), .ZN(
        n19333) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19344), .B1(
        n19343), .B2(n19539), .ZN(n19332) );
  OAI211_X1 U22315 ( .C1(n19542), .C2(n19376), .A(n19333), .B(n19332), .ZN(
        P2_U3131) );
  AOI22_X1 U22316 ( .A1(n19342), .A2(n19481), .B1(n19479), .B2(n19341), .ZN(
        n19335) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19344), .B1(
        n19383), .B2(n19480), .ZN(n19334) );
  OAI211_X1 U22318 ( .C1(n19485), .C2(n19336), .A(n19335), .B(n19334), .ZN(
        P2_U3132) );
  AOI22_X1 U22319 ( .A1(n19342), .A2(n19488), .B1(n19486), .B2(n19341), .ZN(
        n19338) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19344), .B1(
        n19343), .B2(n19487), .ZN(n19337) );
  OAI211_X1 U22321 ( .C1(n19491), .C2(n19376), .A(n19338), .B(n19337), .ZN(
        P2_U3133) );
  AOI22_X1 U22322 ( .A1(n19342), .A2(n19493), .B1(n19492), .B2(n19341), .ZN(
        n19340) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19344), .B1(
        n19343), .B2(n19562), .ZN(n19339) );
  OAI211_X1 U22324 ( .C1(n19565), .C2(n19376), .A(n19340), .B(n19339), .ZN(
        P2_U3134) );
  AOI22_X1 U22325 ( .A1(n19342), .A2(n19500), .B1(n19497), .B2(n19341), .ZN(
        n19346) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19344), .B1(
        n19343), .B2(n19571), .ZN(n19345) );
  OAI211_X1 U22327 ( .C1(n19577), .C2(n19376), .A(n19346), .B(n19345), .ZN(
        P2_U3135) );
  NOR2_X1 U22328 ( .A1(n19347), .A2(n19349), .ZN(n19357) );
  NOR2_X1 U22329 ( .A1(n19357), .A2(n19504), .ZN(n19348) );
  OR2_X1 U22330 ( .A1(n19696), .A2(n19349), .ZN(n19354) );
  INV_X1 U22331 ( .A(n19354), .ZN(n19350) );
  AOI21_X1 U22332 ( .B1(n19697), .B2(n19350), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19351) );
  INV_X1 U22333 ( .A(n19357), .ZN(n19380) );
  OAI22_X1 U22334 ( .A1(n19381), .A2(n19509), .B1(n19508), .B2(n19380), .ZN(
        n19352) );
  INV_X1 U22335 ( .A(n19352), .ZN(n19360) );
  NAND2_X1 U22336 ( .A1(n19511), .A2(n19358), .ZN(n19355) );
  AOI21_X1 U22337 ( .B1(n19355), .B2(n19354), .A(n19353), .ZN(n19356) );
  OAI211_X1 U22338 ( .C1(n19357), .C2(n19697), .A(n19356), .B(n19515), .ZN(
        n19384) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19384), .B1(
        n19415), .B2(n19518), .ZN(n19359) );
  OAI211_X1 U22340 ( .C1(n19521), .C2(n19376), .A(n19360), .B(n19359), .ZN(
        P2_U3136) );
  OAI22_X1 U22341 ( .A1(n19381), .A2(n19523), .B1(n19522), .B2(n19380), .ZN(
        n19361) );
  INV_X1 U22342 ( .A(n19361), .ZN(n19363) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19384), .B1(
        n19383), .B2(n19525), .ZN(n19362) );
  OAI211_X1 U22344 ( .C1(n19528), .C2(n19411), .A(n19363), .B(n19362), .ZN(
        P2_U3137) );
  OAI22_X1 U22345 ( .A1(n19381), .A2(n19530), .B1(n19529), .B2(n19380), .ZN(
        n19364) );
  INV_X1 U22346 ( .A(n19364), .ZN(n19366) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19384), .B1(
        n19383), .B2(n19532), .ZN(n19365) );
  OAI211_X1 U22348 ( .C1(n19535), .C2(n19411), .A(n19366), .B(n19365), .ZN(
        P2_U3138) );
  OAI22_X1 U22349 ( .A1(n19381), .A2(n19537), .B1(n19536), .B2(n19380), .ZN(
        n19367) );
  INV_X1 U22350 ( .A(n19367), .ZN(n19369) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19384), .B1(
        n19415), .B2(n19474), .ZN(n19368) );
  OAI211_X1 U22352 ( .C1(n19478), .C2(n19376), .A(n19369), .B(n19368), .ZN(
        P2_U3139) );
  INV_X1 U22353 ( .A(n19479), .ZN(n19543) );
  OAI22_X1 U22354 ( .A1(n19381), .A2(n19544), .B1(n19543), .B2(n19380), .ZN(
        n19370) );
  INV_X1 U22355 ( .A(n19370), .ZN(n19372) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19384), .B1(
        n19383), .B2(n19546), .ZN(n19371) );
  OAI211_X1 U22357 ( .C1(n19549), .C2(n19411), .A(n19372), .B(n19371), .ZN(
        P2_U3140) );
  OAI22_X1 U22358 ( .A1(n19381), .A2(n19551), .B1(n19550), .B2(n19380), .ZN(
        n19373) );
  INV_X1 U22359 ( .A(n19373), .ZN(n19375) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19384), .B1(
        n19415), .B2(n19553), .ZN(n19374) );
  OAI211_X1 U22361 ( .C1(n19558), .C2(n19376), .A(n19375), .B(n19374), .ZN(
        P2_U3141) );
  OAI22_X1 U22362 ( .A1(n19381), .A2(n19560), .B1(n19559), .B2(n19380), .ZN(
        n19377) );
  INV_X1 U22363 ( .A(n19377), .ZN(n19379) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19384), .B1(
        n19383), .B2(n19562), .ZN(n19378) );
  OAI211_X1 U22365 ( .C1(n19565), .C2(n19411), .A(n19379), .B(n19378), .ZN(
        P2_U3142) );
  OAI22_X1 U22366 ( .A1(n19381), .A2(n19568), .B1(n19566), .B2(n19380), .ZN(
        n19382) );
  INV_X1 U22367 ( .A(n19382), .ZN(n19386) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19384), .B1(
        n19383), .B2(n19571), .ZN(n19385) );
  OAI211_X1 U22369 ( .C1(n19577), .C2(n19411), .A(n19386), .B(n19385), .ZN(
        P2_U3143) );
  NAND4_X1 U22370 ( .A1(n19390), .A2(n19389), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A4(n19697), .ZN(n19388) );
  INV_X1 U22371 ( .A(n10402), .ZN(n19387) );
  NAND3_X1 U22372 ( .A1(n19696), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19421) );
  NOR2_X1 U22373 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19421), .ZN(
        n19413) );
  NOR3_X1 U22374 ( .A1(n19387), .A2(n19413), .A3(n19504), .ZN(n19391) );
  AOI21_X1 U22375 ( .B1(n19504), .B2(n19388), .A(n19391), .ZN(n19414) );
  AOI22_X1 U22376 ( .A1(n19414), .A2(n19462), .B1(n19451), .B2(n19413), .ZN(
        n19397) );
  OAI21_X1 U22377 ( .B1(n19415), .B2(n19445), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19394) );
  NAND3_X1 U22378 ( .A1(n19390), .A2(n19389), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19393) );
  AOI211_X1 U22379 ( .C1(n19394), .C2(n19393), .A(n19392), .B(n19391), .ZN(
        n19395) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19416), .B1(
        n19445), .B2(n19518), .ZN(n19396) );
  OAI211_X1 U22381 ( .C1(n19521), .C2(n19411), .A(n19397), .B(n19396), .ZN(
        P2_U3144) );
  AOI22_X1 U22382 ( .A1(n19414), .A2(n19466), .B1(n19465), .B2(n19413), .ZN(
        n19399) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19525), .ZN(n19398) );
  OAI211_X1 U22384 ( .C1(n19528), .C2(n19437), .A(n19399), .B(n19398), .ZN(
        P2_U3145) );
  AOI22_X1 U22385 ( .A1(n19414), .A2(n19470), .B1(n19469), .B2(n19413), .ZN(
        n19401) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19532), .ZN(n19400) );
  OAI211_X1 U22387 ( .C1(n19535), .C2(n19437), .A(n19401), .B(n19400), .ZN(
        P2_U3146) );
  AOI22_X1 U22388 ( .A1(n19414), .A2(n19475), .B1(n19473), .B2(n19413), .ZN(
        n19403) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19416), .B1(
        n19445), .B2(n19474), .ZN(n19402) );
  OAI211_X1 U22390 ( .C1(n19478), .C2(n19411), .A(n19403), .B(n19402), .ZN(
        P2_U3147) );
  AOI22_X1 U22391 ( .A1(n19414), .A2(n19481), .B1(n19479), .B2(n19413), .ZN(
        n19405) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19546), .ZN(n19404) );
  OAI211_X1 U22393 ( .C1(n19549), .C2(n19437), .A(n19405), .B(n19404), .ZN(
        P2_U3148) );
  AOI22_X1 U22394 ( .A1(n19414), .A2(n19488), .B1(n19486), .B2(n19413), .ZN(
        n19407) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19416), .B1(
        n19445), .B2(n19553), .ZN(n19406) );
  OAI211_X1 U22396 ( .C1(n19558), .C2(n19411), .A(n19407), .B(n19406), .ZN(
        P2_U3149) );
  AOI22_X1 U22397 ( .A1(n19414), .A2(n19493), .B1(n19492), .B2(n19413), .ZN(
        n19410) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19416), .B1(
        n19445), .B2(n19408), .ZN(n19409) );
  OAI211_X1 U22399 ( .C1(n19412), .C2(n19411), .A(n19410), .B(n19409), .ZN(
        P2_U3150) );
  AOI22_X1 U22400 ( .A1(n19414), .A2(n19500), .B1(n19497), .B2(n19413), .ZN(
        n19418) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19571), .ZN(n19417) );
  OAI211_X1 U22402 ( .C1(n19577), .C2(n19437), .A(n19418), .B(n19417), .ZN(
        P2_U3151) );
  INV_X1 U22403 ( .A(n10379), .ZN(n19419) );
  NOR2_X1 U22404 ( .A1(n19703), .A2(n19421), .ZN(n19453) );
  OAI21_X1 U22405 ( .B1(n19419), .B2(n19453), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19420) );
  OAI21_X1 U22406 ( .B1(n19421), .B2(n19454), .A(n19420), .ZN(n19444) );
  AOI22_X1 U22407 ( .A1(n19444), .A2(n19462), .B1(n19451), .B2(n19453), .ZN(
        n19430) );
  INV_X1 U22408 ( .A(n19511), .ZN(n19423) );
  OAI21_X1 U22409 ( .B1(n19423), .B2(n19422), .A(n19421), .ZN(n19426) );
  INV_X1 U22410 ( .A(n19453), .ZN(n19424) );
  OAI211_X1 U22411 ( .C1(n10379), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19424), 
        .B(n19454), .ZN(n19425) );
  NAND3_X1 U22412 ( .A1(n19426), .A2(n19515), .A3(n19425), .ZN(n19446) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19446), .B1(
        n19498), .B2(n19518), .ZN(n19429) );
  OAI211_X1 U22414 ( .C1(n19521), .C2(n19437), .A(n19430), .B(n19429), .ZN(
        P2_U3152) );
  AOI22_X1 U22415 ( .A1(n19444), .A2(n19466), .B1(n19465), .B2(n19453), .ZN(
        n19432) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19525), .ZN(n19431) );
  OAI211_X1 U22417 ( .C1(n19528), .C2(n19484), .A(n19432), .B(n19431), .ZN(
        P2_U3153) );
  AOI22_X1 U22418 ( .A1(n19444), .A2(n19470), .B1(n19469), .B2(n19453), .ZN(
        n19434) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19532), .ZN(n19433) );
  OAI211_X1 U22420 ( .C1(n19535), .C2(n19484), .A(n19434), .B(n19433), .ZN(
        P2_U3154) );
  AOI22_X1 U22421 ( .A1(n19444), .A2(n19475), .B1(n19473), .B2(n19453), .ZN(
        n19436) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19446), .B1(
        n19498), .B2(n19474), .ZN(n19435) );
  OAI211_X1 U22423 ( .C1(n19478), .C2(n19437), .A(n19436), .B(n19435), .ZN(
        P2_U3155) );
  AOI22_X1 U22424 ( .A1(n19444), .A2(n19481), .B1(n19479), .B2(n19453), .ZN(
        n19439) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19546), .ZN(n19438) );
  OAI211_X1 U22426 ( .C1(n19549), .C2(n19484), .A(n19439), .B(n19438), .ZN(
        P2_U3156) );
  AOI22_X1 U22427 ( .A1(n19444), .A2(n19488), .B1(n19486), .B2(n19453), .ZN(
        n19441) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19487), .ZN(n19440) );
  OAI211_X1 U22429 ( .C1(n19491), .C2(n19484), .A(n19441), .B(n19440), .ZN(
        P2_U3157) );
  AOI22_X1 U22430 ( .A1(n19444), .A2(n19493), .B1(n19492), .B2(n19453), .ZN(
        n19443) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19562), .ZN(n19442) );
  OAI211_X1 U22432 ( .C1(n19565), .C2(n19484), .A(n19443), .B(n19442), .ZN(
        P2_U3158) );
  AOI22_X1 U22433 ( .A1(n19444), .A2(n19500), .B1(n19497), .B2(n19453), .ZN(
        n19448) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19446), .B1(
        n19445), .B2(n19571), .ZN(n19447) );
  OAI211_X1 U22435 ( .C1(n19577), .C2(n19484), .A(n19448), .B(n19447), .ZN(
        P2_U3159) );
  NAND2_X1 U22436 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19450), .ZN(
        n19513) );
  NOR2_X1 U22437 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19513), .ZN(
        n19496) );
  AOI22_X1 U22438 ( .A1(n19518), .A2(n19572), .B1(n19451), .B2(n19496), .ZN(
        n19464) );
  OAI21_X1 U22439 ( .B1(n19572), .B2(n19498), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19452) );
  NAND2_X1 U22440 ( .A1(n19452), .A2(n19681), .ZN(n19461) );
  NOR2_X1 U22441 ( .A1(n19496), .A2(n19453), .ZN(n19460) );
  INV_X1 U22442 ( .A(n19460), .ZN(n19457) );
  INV_X1 U22443 ( .A(n19496), .ZN(n19455) );
  OAI211_X1 U22444 ( .C1(n10388), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19455), 
        .B(n19454), .ZN(n19456) );
  OAI211_X1 U22445 ( .C1(n19461), .C2(n19457), .A(n19515), .B(n19456), .ZN(
        n19501) );
  INV_X1 U22446 ( .A(n10388), .ZN(n19458) );
  OAI21_X1 U22447 ( .B1(n19458), .B2(n19496), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19459) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19501), .B1(
        n19462), .B2(n19499), .ZN(n19463) );
  OAI211_X1 U22449 ( .C1(n19521), .C2(n19484), .A(n19464), .B(n19463), .ZN(
        P2_U3160) );
  AOI22_X1 U22450 ( .A1(n19525), .A2(n19498), .B1(n19465), .B2(n19496), .ZN(
        n19468) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19501), .B1(
        n19466), .B2(n19499), .ZN(n19467) );
  OAI211_X1 U22452 ( .C1(n19528), .C2(n19557), .A(n19468), .B(n19467), .ZN(
        P2_U3161) );
  AOI22_X1 U22453 ( .A1(n19532), .A2(n19498), .B1(n19469), .B2(n19496), .ZN(
        n19472) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19501), .B1(
        n19470), .B2(n19499), .ZN(n19471) );
  OAI211_X1 U22455 ( .C1(n19535), .C2(n19557), .A(n19472), .B(n19471), .ZN(
        P2_U3162) );
  AOI22_X1 U22456 ( .A1(n19474), .A2(n19572), .B1(n19473), .B2(n19496), .ZN(
        n19477) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19501), .B1(
        n19475), .B2(n19499), .ZN(n19476) );
  OAI211_X1 U22458 ( .C1(n19478), .C2(n19484), .A(n19477), .B(n19476), .ZN(
        P2_U3163) );
  AOI22_X1 U22459 ( .A1(n19480), .A2(n19572), .B1(n19479), .B2(n19496), .ZN(
        n19483) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19501), .B1(
        n19481), .B2(n19499), .ZN(n19482) );
  OAI211_X1 U22461 ( .C1(n19485), .C2(n19484), .A(n19483), .B(n19482), .ZN(
        P2_U3164) );
  AOI22_X1 U22462 ( .A1(n19487), .A2(n19498), .B1(n19486), .B2(n19496), .ZN(
        n19490) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19501), .B1(
        n19488), .B2(n19499), .ZN(n19489) );
  OAI211_X1 U22464 ( .C1(n19491), .C2(n19557), .A(n19490), .B(n19489), .ZN(
        P2_U3165) );
  AOI22_X1 U22465 ( .A1(n19562), .A2(n19498), .B1(n19492), .B2(n19496), .ZN(
        n19495) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19501), .B1(
        n19493), .B2(n19499), .ZN(n19494) );
  OAI211_X1 U22467 ( .C1(n19565), .C2(n19557), .A(n19495), .B(n19494), .ZN(
        P2_U3166) );
  AOI22_X1 U22468 ( .A1(n19571), .A2(n19498), .B1(n19497), .B2(n19496), .ZN(
        n19503) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19501), .B1(
        n19500), .B2(n19499), .ZN(n19502) );
  OAI211_X1 U22470 ( .C1(n19577), .C2(n19557), .A(n19503), .B(n19502), .ZN(
        P2_U3167) );
  NOR2_X1 U22471 ( .A1(n19517), .A2(n19504), .ZN(n19505) );
  INV_X1 U22472 ( .A(n19513), .ZN(n19506) );
  AOI21_X1 U22473 ( .B1(n19697), .B2(n19506), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19507) );
  OR2_X1 U22474 ( .A1(n19512), .A2(n19507), .ZN(n19569) );
  OAI22_X1 U22475 ( .A1(n19569), .A2(n19509), .B1(n19567), .B2(n19508), .ZN(
        n19510) );
  INV_X1 U22476 ( .A(n19510), .ZN(n19520) );
  NAND2_X1 U22477 ( .A1(n19511), .A2(n19673), .ZN(n19514) );
  AOI21_X1 U22478 ( .B1(n19514), .B2(n19513), .A(n19512), .ZN(n19516) );
  OAI211_X1 U22479 ( .C1(n19517), .C2(n19697), .A(n19516), .B(n19515), .ZN(
        n19573) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19573), .B1(
        n19554), .B2(n19518), .ZN(n19519) );
  OAI211_X1 U22481 ( .C1(n19521), .C2(n19557), .A(n19520), .B(n19519), .ZN(
        P2_U3168) );
  OAI22_X1 U22482 ( .A1(n19569), .A2(n19523), .B1(n19567), .B2(n19522), .ZN(
        n19524) );
  INV_X1 U22483 ( .A(n19524), .ZN(n19527) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19525), .ZN(n19526) );
  OAI211_X1 U22485 ( .C1(n19528), .C2(n19576), .A(n19527), .B(n19526), .ZN(
        P2_U3169) );
  OAI22_X1 U22486 ( .A1(n19569), .A2(n19530), .B1(n19567), .B2(n19529), .ZN(
        n19531) );
  INV_X1 U22487 ( .A(n19531), .ZN(n19534) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19532), .ZN(n19533) );
  OAI211_X1 U22489 ( .C1(n19535), .C2(n19576), .A(n19534), .B(n19533), .ZN(
        P2_U3170) );
  OAI22_X1 U22490 ( .A1(n19569), .A2(n19537), .B1(n19567), .B2(n19536), .ZN(
        n19538) );
  INV_X1 U22491 ( .A(n19538), .ZN(n19541) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19539), .ZN(n19540) );
  OAI211_X1 U22493 ( .C1(n19542), .C2(n19576), .A(n19541), .B(n19540), .ZN(
        P2_U3171) );
  OAI22_X1 U22494 ( .A1(n19569), .A2(n19544), .B1(n19567), .B2(n19543), .ZN(
        n19545) );
  INV_X1 U22495 ( .A(n19545), .ZN(n19548) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19546), .ZN(n19547) );
  OAI211_X1 U22497 ( .C1(n19549), .C2(n19576), .A(n19548), .B(n19547), .ZN(
        P2_U3172) );
  OAI22_X1 U22498 ( .A1(n19569), .A2(n19551), .B1(n19567), .B2(n19550), .ZN(
        n19552) );
  INV_X1 U22499 ( .A(n19552), .ZN(n19556) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19573), .B1(
        n19554), .B2(n19553), .ZN(n19555) );
  OAI211_X1 U22501 ( .C1(n19558), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P2_U3173) );
  OAI22_X1 U22502 ( .A1(n19569), .A2(n19560), .B1(n19567), .B2(n19559), .ZN(
        n19561) );
  INV_X1 U22503 ( .A(n19561), .ZN(n19564) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19562), .ZN(n19563) );
  OAI211_X1 U22505 ( .C1(n19565), .C2(n19576), .A(n19564), .B(n19563), .ZN(
        P2_U3174) );
  OAI22_X1 U22506 ( .A1(n19569), .A2(n19568), .B1(n19567), .B2(n19566), .ZN(
        n19570) );
  INV_X1 U22507 ( .A(n19570), .ZN(n19575) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19573), .B1(
        n19572), .B2(n19571), .ZN(n19574) );
  OAI211_X1 U22509 ( .C1(n19577), .C2(n19576), .A(n19575), .B(n19574), .ZN(
        P2_U3175) );
  AOI21_X1 U22510 ( .B1(n19669), .B2(n19578), .A(n19720), .ZN(n19584) );
  NAND2_X1 U22511 ( .A1(n19579), .A2(n19721), .ZN(n19583) );
  OAI211_X1 U22512 ( .C1(n19580), .C2(n19583), .A(n19722), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19581) );
  OAI211_X1 U22513 ( .C1(n19584), .C2(n19583), .A(n19582), .B(n19581), .ZN(
        P2_U3177) );
  AND2_X1 U22514 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19585), .ZN(
        P2_U3179) );
  AND2_X1 U22515 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19585), .ZN(
        P2_U3180) );
  AND2_X1 U22516 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19585), .ZN(
        P2_U3181) );
  AND2_X1 U22517 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19585), .ZN(
        P2_U3182) );
  AND2_X1 U22518 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19585), .ZN(
        P2_U3183) );
  AND2_X1 U22519 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19585), .ZN(
        P2_U3184) );
  AND2_X1 U22520 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19585), .ZN(
        P2_U3185) );
  AND2_X1 U22521 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19585), .ZN(
        P2_U3186) );
  AND2_X1 U22522 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19585), .ZN(
        P2_U3187) );
  AND2_X1 U22523 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19585), .ZN(
        P2_U3188) );
  AND2_X1 U22524 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19585), .ZN(
        P2_U3189) );
  AND2_X1 U22525 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19585), .ZN(
        P2_U3190) );
  AND2_X1 U22526 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19585), .ZN(
        P2_U3191) );
  AND2_X1 U22527 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19585), .ZN(
        P2_U3192) );
  AND2_X1 U22528 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19585), .ZN(
        P2_U3193) );
  AND2_X1 U22529 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19585), .ZN(
        P2_U3194) );
  AND2_X1 U22530 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19585), .ZN(
        P2_U3195) );
  AND2_X1 U22531 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19585), .ZN(
        P2_U3196) );
  AND2_X1 U22532 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19585), .ZN(
        P2_U3197) );
  AND2_X1 U22533 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19585), .ZN(
        P2_U3198) );
  AND2_X1 U22534 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19585), .ZN(
        P2_U3199) );
  AND2_X1 U22535 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19585), .ZN(
        P2_U3200) );
  AND2_X1 U22536 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19585), .ZN(P2_U3201) );
  AND2_X1 U22537 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19585), .ZN(P2_U3202) );
  AND2_X1 U22538 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19585), .ZN(P2_U3203) );
  AND2_X1 U22539 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19585), .ZN(P2_U3204) );
  AND2_X1 U22540 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19585), .ZN(P2_U3205) );
  AND2_X1 U22541 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19585), .ZN(P2_U3206) );
  AND2_X1 U22542 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19585), .ZN(P2_U3207) );
  AND2_X1 U22543 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19585), .ZN(P2_U3208) );
  NOR2_X1 U22544 ( .A1(n19587), .A2(n19586), .ZN(n19598) );
  INV_X1 U22545 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19735) );
  OR3_X1 U22546 ( .A1(n19598), .A2(n19735), .A3(n19602), .ZN(n19589) );
  AOI211_X1 U22547 ( .C1(n19603), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19600), .B(n19736), .ZN(n19588) );
  INV_X1 U22548 ( .A(NA), .ZN(n19599) );
  NOR2_X1 U22549 ( .A1(n19599), .A2(n19591), .ZN(n19607) );
  AOI211_X1 U22550 ( .C1(n19608), .C2(n19589), .A(n19588), .B(n19607), .ZN(
        n19590) );
  INV_X1 U22551 ( .A(n19590), .ZN(P2_U3209) );
  AOI21_X1 U22552 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19603), .A(n19608), 
        .ZN(n19596) );
  NOR2_X1 U22553 ( .A1(n19735), .A2(n19596), .ZN(n19592) );
  AOI21_X1 U22554 ( .B1(n19592), .B2(n19591), .A(n19598), .ZN(n19594) );
  INV_X1 U22555 ( .A(n19730), .ZN(n19593) );
  OAI211_X1 U22556 ( .C1(n19603), .C2(n19595), .A(n19594), .B(n19593), .ZN(
        P2_U3210) );
  AOI21_X1 U22557 ( .B1(n19722), .B2(n19597), .A(n19596), .ZN(n19606) );
  AOI22_X1 U22558 ( .A1(n19735), .A2(n19600), .B1(n19599), .B2(n19598), .ZN(
        n19601) );
  AOI211_X1 U22559 ( .C1(n19735), .C2(n19603), .A(n19602), .B(n19601), .ZN(
        n19604) );
  INV_X1 U22560 ( .A(n19604), .ZN(n19605) );
  OAI21_X1 U22561 ( .B1(n19607), .B2(n19606), .A(n19605), .ZN(P2_U3211) );
  OAI222_X1 U22562 ( .A1(n19655), .A2(n10128), .B1(n19609), .B2(n19736), .C1(
        n10168), .C2(n19656), .ZN(P2_U3212) );
  OAI222_X1 U22563 ( .A1(n19655), .A2(n10180), .B1(n19610), .B2(n19736), .C1(
        n10128), .C2(n19656), .ZN(P2_U3213) );
  OAI222_X1 U22564 ( .A1(n19655), .A2(n19612), .B1(n19611), .B2(n19736), .C1(
        n10180), .C2(n19656), .ZN(P2_U3214) );
  INV_X1 U22565 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19614) );
  OAI222_X1 U22566 ( .A1(n19655), .A2(n19614), .B1(n19613), .B2(n19736), .C1(
        n19612), .C2(n19656), .ZN(P2_U3215) );
  OAI222_X1 U22567 ( .A1(n19655), .A2(n19616), .B1(n19615), .B2(n19736), .C1(
        n19614), .C2(n19656), .ZN(P2_U3216) );
  OAI222_X1 U22568 ( .A1(n19655), .A2(n10750), .B1(n19617), .B2(n19736), .C1(
        n19616), .C2(n19656), .ZN(P2_U3217) );
  OAI222_X1 U22569 ( .A1(n19655), .A2(n19619), .B1(n19618), .B2(n19736), .C1(
        n10750), .C2(n19656), .ZN(P2_U3218) );
  OAI222_X1 U22570 ( .A1(n19655), .A2(n19620), .B1(n20683), .B2(n19736), .C1(
        n19619), .C2(n19656), .ZN(P2_U3219) );
  OAI222_X1 U22571 ( .A1(n19655), .A2(n19622), .B1(n19621), .B2(n19736), .C1(
        n19620), .C2(n19656), .ZN(P2_U3220) );
  OAI222_X1 U22572 ( .A1(n19655), .A2(n10767), .B1(n19623), .B2(n19736), .C1(
        n19622), .C2(n19656), .ZN(P2_U3221) );
  OAI222_X1 U22573 ( .A1(n19655), .A2(n19625), .B1(n19624), .B2(n19736), .C1(
        n10767), .C2(n19656), .ZN(P2_U3222) );
  OAI222_X1 U22574 ( .A1(n19655), .A2(n10776), .B1(n19626), .B2(n19736), .C1(
        n19625), .C2(n19656), .ZN(P2_U3223) );
  OAI222_X1 U22575 ( .A1(n19655), .A2(n19628), .B1(n19627), .B2(n19736), .C1(
        n10776), .C2(n19656), .ZN(P2_U3224) );
  OAI222_X1 U22576 ( .A1(n19655), .A2(n19630), .B1(n19629), .B2(n19736), .C1(
        n19628), .C2(n19656), .ZN(P2_U3225) );
  OAI222_X1 U22577 ( .A1(n19655), .A2(n19632), .B1(n19631), .B2(n19736), .C1(
        n19630), .C2(n19656), .ZN(P2_U3226) );
  OAI222_X1 U22578 ( .A1(n19655), .A2(n19634), .B1(n19633), .B2(n19736), .C1(
        n19632), .C2(n19656), .ZN(P2_U3227) );
  OAI222_X1 U22579 ( .A1(n19655), .A2(n15066), .B1(n19635), .B2(n19736), .C1(
        n19634), .C2(n19656), .ZN(P2_U3228) );
  OAI222_X1 U22580 ( .A1(n19655), .A2(n19637), .B1(n19636), .B2(n19736), .C1(
        n15066), .C2(n19656), .ZN(P2_U3229) );
  INV_X1 U22581 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19639) );
  OAI222_X1 U22582 ( .A1(n19655), .A2(n19639), .B1(n19638), .B2(n19736), .C1(
        n19637), .C2(n19656), .ZN(P2_U3230) );
  OAI222_X1 U22583 ( .A1(n19655), .A2(n19641), .B1(n19640), .B2(n19736), .C1(
        n19639), .C2(n19656), .ZN(P2_U3231) );
  OAI222_X1 U22584 ( .A1(n19655), .A2(n10811), .B1(n19642), .B2(n19736), .C1(
        n19641), .C2(n19656), .ZN(P2_U3232) );
  OAI222_X1 U22585 ( .A1(n19655), .A2(n19644), .B1(n19643), .B2(n19736), .C1(
        n10811), .C2(n19656), .ZN(P2_U3233) );
  OAI222_X1 U22586 ( .A1(n19655), .A2(n15947), .B1(n19645), .B2(n19736), .C1(
        n19644), .C2(n19656), .ZN(P2_U3234) );
  OAI222_X1 U22587 ( .A1(n19655), .A2(n19647), .B1(n19646), .B2(n19736), .C1(
        n15947), .C2(n19656), .ZN(P2_U3235) );
  OAI222_X1 U22588 ( .A1(n19655), .A2(n19649), .B1(n19648), .B2(n19736), .C1(
        n19647), .C2(n19656), .ZN(P2_U3236) );
  OAI222_X1 U22589 ( .A1(n19655), .A2(n19651), .B1(n19650), .B2(n19736), .C1(
        n19649), .C2(n19656), .ZN(P2_U3237) );
  OAI222_X1 U22590 ( .A1(n19656), .A2(n19651), .B1(n20678), .B2(n19736), .C1(
        n14956), .C2(n19655), .ZN(P2_U3238) );
  OAI222_X1 U22591 ( .A1(n19655), .A2(n19653), .B1(n19652), .B2(n19736), .C1(
        n14956), .C2(n19656), .ZN(P2_U3239) );
  INV_X1 U22592 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19657) );
  OAI222_X1 U22593 ( .A1(n19655), .A2(n19657), .B1(n19654), .B2(n19736), .C1(
        n19653), .C2(n19656), .ZN(P2_U3240) );
  OAI222_X1 U22594 ( .A1(n19655), .A2(n19659), .B1(n19658), .B2(n19736), .C1(
        n19657), .C2(n19656), .ZN(P2_U3241) );
  AOI22_X1 U22595 ( .A1(n19736), .A2(n19661), .B1(n19660), .B2(n19737), .ZN(
        P2_U3585) );
  MUX2_X1 U22596 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19737), .Z(P2_U3586) );
  OAI22_X1 U22597 ( .A1(n19737), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19736), .ZN(n19662) );
  INV_X1 U22598 ( .A(n19662), .ZN(P2_U3587) );
  OAI22_X1 U22599 ( .A1(n19737), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19736), .ZN(n19663) );
  INV_X1 U22600 ( .A(n19663), .ZN(P2_U3588) );
  OAI21_X1 U22601 ( .B1(n19667), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19665), 
        .ZN(n19664) );
  INV_X1 U22602 ( .A(n19664), .ZN(P2_U3591) );
  OAI21_X1 U22603 ( .B1(n19667), .B2(n19666), .A(n19665), .ZN(P2_U3592) );
  NOR3_X1 U22604 ( .A1(n19670), .A2(n19669), .A3(n19668), .ZN(n19672) );
  INV_X1 U22605 ( .A(n19671), .ZN(n19719) );
  NOR2_X1 U22606 ( .A1(n19672), .A2(n19719), .ZN(n19684) );
  NAND3_X1 U22607 ( .A1(n19674), .A2(n19681), .A3(n19673), .ZN(n19675) );
  OAI21_X1 U22608 ( .B1(n19676), .B2(n19697), .A(n19675), .ZN(n19677) );
  AOI21_X1 U22609 ( .B1(n19678), .B2(n19684), .A(n19677), .ZN(n19679) );
  AOI22_X1 U22610 ( .A1(n19704), .A2(n19680), .B1(n19679), .B2(n19701), .ZN(
        P2_U3602) );
  NAND2_X1 U22611 ( .A1(n19681), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19691) );
  OAI21_X1 U22612 ( .B1(n19689), .B2(n19691), .A(n19682), .ZN(n19683) );
  AOI22_X1 U22613 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19685), .B1(n19684), 
        .B2(n19683), .ZN(n19686) );
  AOI22_X1 U22614 ( .A1(n19704), .A2(n19687), .B1(n19686), .B2(n19701), .ZN(
        P2_U3603) );
  OR3_X1 U22615 ( .A1(n19689), .A2(n19719), .A3(n19688), .ZN(n19690) );
  OAI21_X1 U22616 ( .B1(n19692), .B2(n19691), .A(n19690), .ZN(n19693) );
  AOI21_X1 U22617 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19694), .A(n19693), 
        .ZN(n19695) );
  AOI22_X1 U22618 ( .A1(n19704), .A2(n19696), .B1(n19695), .B2(n19701), .ZN(
        P2_U3604) );
  OAI22_X1 U22619 ( .A1(n19698), .A2(n19719), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19697), .ZN(n19699) );
  AOI21_X1 U22620 ( .B1(n19700), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19699), 
        .ZN(n19702) );
  AOI22_X1 U22621 ( .A1(n19704), .A2(n19703), .B1(n19702), .B2(n19701), .ZN(
        P2_U3605) );
  AOI22_X1 U22622 ( .A1(n19736), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19705), 
        .B2(n19737), .ZN(P2_U3608) );
  INV_X1 U22623 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19718) );
  INV_X1 U22624 ( .A(n19706), .ZN(n19717) );
  INV_X1 U22625 ( .A(n19707), .ZN(n19711) );
  INV_X1 U22626 ( .A(n19708), .ZN(n19709) );
  OAI22_X1 U22627 ( .A1(n19712), .A2(n19711), .B1(n19710), .B2(n19709), .ZN(
        n19713) );
  INV_X1 U22628 ( .A(n19713), .ZN(n19716) );
  NOR2_X1 U22629 ( .A1(n19717), .A2(n19714), .ZN(n19715) );
  AOI22_X1 U22630 ( .A1(n19718), .A2(n19717), .B1(n19716), .B2(n19715), .ZN(
        P2_U3609) );
  OAI22_X1 U22631 ( .A1(n19722), .A2(n19721), .B1(n19720), .B2(n19719), .ZN(
        n19723) );
  NOR2_X1 U22632 ( .A1(n19724), .A2(n19723), .ZN(n19734) );
  NOR4_X1 U22633 ( .A1(n9627), .A2(n9583), .A3(n19729), .A4(n19730), .ZN(
        n19725) );
  AOI21_X1 U22634 ( .B1(n19727), .B2(n19726), .A(n19725), .ZN(n19733) );
  AOI211_X1 U22635 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19730), .A(n19729), 
        .B(n19728), .ZN(n19731) );
  NOR2_X1 U22636 ( .A1(n19734), .A2(n19731), .ZN(n19732) );
  AOI22_X1 U22637 ( .A1(n19735), .A2(n19734), .B1(n19733), .B2(n19732), .ZN(
        P2_U3610) );
  OAI22_X1 U22638 ( .A1(n19737), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19736), .ZN(n19738) );
  INV_X1 U22639 ( .A(n19738), .ZN(P2_U3611) );
  NOR2_X1 U22640 ( .A1(n20566), .A2(n20570), .ZN(n19745) );
  INV_X1 U22641 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19739) );
  AND2_X1 U22642 ( .A1(n20570), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20637) );
  AOI21_X1 U22643 ( .B1(n19745), .B2(n19739), .A(n20637), .ZN(P1_U2802) );
  OAI21_X1 U22644 ( .B1(n19741), .B2(n19740), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19742) );
  OAI21_X1 U22645 ( .B1(n19743), .B2(n20790), .A(n19742), .ZN(P1_U2803) );
  INV_X2 U22646 ( .A(n20637), .ZN(n20650) );
  NOR2_X1 U22647 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20572) );
  OAI21_X1 U22648 ( .B1(n20572), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20650), .ZN(
        n19744) );
  OAI21_X1 U22649 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20650), .A(n19744), 
        .ZN(P1_U2804) );
  NOR2_X1 U22650 ( .A1(n20637), .A2(n19745), .ZN(n20621) );
  OAI21_X1 U22651 ( .B1(BS16), .B2(n20572), .A(n20621), .ZN(n20619) );
  OAI21_X1 U22652 ( .B1(n20621), .B2(n20641), .A(n20619), .ZN(P1_U2805) );
  OAI21_X1 U22653 ( .B1(n19748), .B2(n19747), .A(n19746), .ZN(P1_U2806) );
  NOR4_X1 U22654 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19752) );
  NOR4_X1 U22655 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19751) );
  NOR4_X1 U22656 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19750) );
  NOR4_X1 U22657 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19749) );
  NAND4_X1 U22658 ( .A1(n19752), .A2(n19751), .A3(n19750), .A4(n19749), .ZN(
        n19758) );
  NOR4_X1 U22659 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19756) );
  AOI211_X1 U22660 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19755) );
  NOR4_X1 U22661 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19754) );
  NOR4_X1 U22662 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19753) );
  NAND4_X1 U22663 ( .A1(n19756), .A2(n19755), .A3(n19754), .A4(n19753), .ZN(
        n19757) );
  NOR2_X1 U22664 ( .A1(n19758), .A2(n19757), .ZN(n20635) );
  INV_X1 U22665 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19760) );
  NOR3_X1 U22666 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A3(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19761) );
  OAI21_X1 U22667 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19761), .A(n20635), .ZN(
        n19759) );
  OAI21_X1 U22668 ( .B1(n20635), .B2(n19760), .A(n19759), .ZN(P1_U2807) );
  INV_X1 U22669 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20620) );
  AOI21_X1 U22670 ( .B1(n13878), .B2(n20620), .A(n19761), .ZN(n19763) );
  INV_X1 U22671 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19762) );
  INV_X1 U22672 ( .A(n20635), .ZN(n20630) );
  AOI22_X1 U22673 ( .A1(n20635), .A2(n19763), .B1(n19762), .B2(n20630), .ZN(
        P1_U2808) );
  INV_X1 U22674 ( .A(n19835), .ZN(n19788) );
  AOI21_X1 U22675 ( .B1(n19789), .B2(n19764), .A(n19788), .ZN(n19787) );
  AOI22_X1 U22676 ( .A1(n19797), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n19766), .B2(
        n19765), .ZN(n19767) );
  OAI211_X1 U22677 ( .C1(n19769), .C2(n19768), .A(n19767), .B(n19820), .ZN(
        n19770) );
  AOI21_X1 U22678 ( .B1(n19828), .B2(n19837), .A(n19770), .ZN(n19773) );
  AOI22_X1 U22679 ( .A1(n19838), .A2(n19809), .B1(n19774), .B2(n19771), .ZN(
        n19772) );
  OAI211_X1 U22680 ( .C1(n19787), .C2(n19774), .A(n19773), .B(n19772), .ZN(
        P1_U2831) );
  NOR4_X1 U22681 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19804), .A3(n19799), .A4(
        n19798), .ZN(n19782) );
  AOI21_X1 U22682 ( .B1(n19823), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19775), .ZN(n19776) );
  OAI21_X1 U22683 ( .B1(n19821), .B2(n19777), .A(n19776), .ZN(n19778) );
  AOI21_X1 U22684 ( .B1(n19797), .B2(P1_EBX_REG_8__SCAN_IN), .A(n19778), .ZN(
        n19779) );
  OAI21_X1 U22685 ( .B1(n19780), .B2(n19793), .A(n19779), .ZN(n19781) );
  OR2_X1 U22686 ( .A1(n19782), .A2(n19781), .ZN(n19783) );
  AOI21_X1 U22687 ( .B1(n19784), .B2(n19809), .A(n19783), .ZN(n19785) );
  OAI21_X1 U22688 ( .B1(n19787), .B2(n19786), .A(n19785), .ZN(P1_U2832) );
  AOI21_X1 U22689 ( .B1(n19789), .B2(n19799), .A(n19788), .ZN(n19806) );
  NAND2_X1 U22690 ( .A1(n19823), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19790) );
  OAI211_X1 U22691 ( .C1(n19821), .C2(n19791), .A(n19790), .B(n19820), .ZN(
        n19796) );
  INV_X1 U22692 ( .A(n19792), .ZN(n19794) );
  NOR2_X1 U22693 ( .A1(n19794), .A2(n19793), .ZN(n19795) );
  AOI211_X1 U22694 ( .C1(n19797), .C2(P1_EBX_REG_7__SCAN_IN), .A(n19796), .B(
        n19795), .ZN(n19803) );
  NOR2_X1 U22695 ( .A1(n19799), .A2(n19798), .ZN(n19800) );
  AOI22_X1 U22696 ( .A1(n19801), .A2(n19809), .B1(n19804), .B2(n19800), .ZN(
        n19802) );
  OAI211_X1 U22697 ( .C1(n19806), .C2(n19804), .A(n19803), .B(n19802), .ZN(
        P1_U2833) );
  AOI22_X1 U22698 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19823), .B1(
        n19828), .B2(n19841), .ZN(n19811) );
  INV_X1 U22699 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19844) );
  OAI22_X1 U22700 ( .A1(n19825), .A2(n19844), .B1(n19805), .B2(n19821), .ZN(
        n19808) );
  INV_X1 U22701 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20581) );
  NAND2_X1 U22702 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19835), .ZN(n19814) );
  AOI21_X1 U22703 ( .B1(n20581), .B2(n19814), .A(n19806), .ZN(n19807) );
  AOI211_X1 U22704 ( .C1(n19842), .C2(n19809), .A(n19808), .B(n19807), .ZN(
        n19810) );
  NAND3_X1 U22705 ( .A1(n19811), .A2(n19810), .A3(n19820), .ZN(P1_U2834) );
  AOI22_X1 U22706 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19823), .B1(
        n19828), .B2(n19845), .ZN(n19818) );
  OAI22_X1 U22707 ( .A1(n19825), .A2(n19850), .B1(n19821), .B2(n19812), .ZN(
        n19813) );
  AOI21_X1 U22708 ( .B1(n19848), .B2(n19833), .A(n19813), .ZN(n19817) );
  OAI21_X1 U22709 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n19815), .A(n19814), .ZN(
        n19816) );
  NAND4_X1 U22710 ( .A1(n19818), .A2(n19817), .A3(n19820), .A4(n19816), .ZN(
        P1_U2835) );
  NAND2_X1 U22711 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n19819), .ZN(n19836) );
  INV_X1 U22712 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20579) );
  OAI21_X1 U22713 ( .B1(n19821), .B2(n19915), .A(n19820), .ZN(n19822) );
  AOI21_X1 U22714 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19823), .A(
        n19822), .ZN(n19824) );
  OAI21_X1 U22715 ( .B1(n19826), .B2(n19825), .A(n19824), .ZN(n19827) );
  AOI21_X1 U22716 ( .B1(n19828), .B2(n19918), .A(n19827), .ZN(n19829) );
  OAI21_X1 U22717 ( .B1(n19831), .B2(n19830), .A(n19829), .ZN(n19832) );
  AOI21_X1 U22718 ( .B1(n19910), .B2(n19833), .A(n19832), .ZN(n19834) );
  OAI221_X1 U22719 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n19836), .C1(n20579), 
        .C2(n19835), .A(n19834), .ZN(P1_U2836) );
  INV_X1 U22720 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19840) );
  AOI22_X1 U22721 ( .A1(n19838), .A2(n19847), .B1(n19846), .B2(n19837), .ZN(
        n19839) );
  OAI21_X1 U22722 ( .B1(n19851), .B2(n19840), .A(n19839), .ZN(P1_U2863) );
  AOI22_X1 U22723 ( .A1(n19842), .A2(n19847), .B1(n19846), .B2(n19841), .ZN(
        n19843) );
  OAI21_X1 U22724 ( .B1(n19851), .B2(n19844), .A(n19843), .ZN(P1_U2866) );
  AOI22_X1 U22725 ( .A1(n19848), .A2(n19847), .B1(n19846), .B2(n19845), .ZN(
        n19849) );
  OAI21_X1 U22726 ( .B1(n19851), .B2(n19850), .A(n19849), .ZN(P1_U2867) );
  AOI22_X1 U22727 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19854), .B1(n19872), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19852) );
  OAI21_X1 U22728 ( .B1(n20791), .B2(n19853), .A(n19852), .ZN(P1_U2921) );
  INV_X1 U22729 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19856) );
  AOI22_X1 U22730 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19855) );
  OAI21_X1 U22731 ( .B1(n19856), .B2(n19875), .A(n19855), .ZN(P1_U2922) );
  AOI22_X1 U22732 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19857) );
  OAI21_X1 U22733 ( .B1(n14135), .B2(n19875), .A(n19857), .ZN(P1_U2923) );
  AOI22_X1 U22734 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19858) );
  OAI21_X1 U22735 ( .B1(n14101), .B2(n19875), .A(n19858), .ZN(P1_U2924) );
  AOI22_X1 U22736 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19859) );
  OAI21_X1 U22737 ( .B1(n14068), .B2(n19875), .A(n19859), .ZN(P1_U2925) );
  AOI22_X1 U22738 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19860) );
  OAI21_X1 U22739 ( .B1(n13986), .B2(n19875), .A(n19860), .ZN(P1_U2926) );
  INV_X1 U22740 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U22741 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19861) );
  OAI21_X1 U22742 ( .B1(n19862), .B2(n19875), .A(n19861), .ZN(P1_U2927) );
  INV_X1 U22743 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U22744 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19863) );
  OAI21_X1 U22745 ( .B1(n19864), .B2(n19875), .A(n19863), .ZN(P1_U2928) );
  AOI22_X1 U22746 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19865) );
  OAI21_X1 U22747 ( .B1(n11662), .B2(n19875), .A(n19865), .ZN(P1_U2929) );
  AOI22_X1 U22748 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19866) );
  OAI21_X1 U22749 ( .B1(n11651), .B2(n19875), .A(n19866), .ZN(P1_U2930) );
  AOI22_X1 U22750 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19867) );
  OAI21_X1 U22751 ( .B1(n13598), .B2(n19875), .A(n19867), .ZN(P1_U2931) );
  AOI22_X1 U22752 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19868) );
  OAI21_X1 U22753 ( .B1(n20749), .B2(n19875), .A(n19868), .ZN(P1_U2932) );
  AOI22_X1 U22754 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19869) );
  OAI21_X1 U22755 ( .B1(n11631), .B2(n19875), .A(n19869), .ZN(P1_U2933) );
  AOI22_X1 U22756 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U22757 ( .B1(n11601), .B2(n19875), .A(n19870), .ZN(P1_U2934) );
  AOI22_X1 U22758 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19871) );
  OAI21_X1 U22759 ( .B1(n11607), .B2(n19875), .A(n19871), .ZN(P1_U2935) );
  AOI22_X1 U22760 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19873), .B1(n19872), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U22761 ( .B1(n19876), .B2(n19875), .A(n19874), .ZN(P1_U2936) );
  AOI22_X1 U22762 ( .A1(n19905), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19904), .ZN(n19878) );
  NAND2_X1 U22763 ( .A1(n19890), .A2(n19877), .ZN(n19892) );
  NAND2_X1 U22764 ( .A1(n19878), .A2(n19892), .ZN(P1_U2945) );
  AOI22_X1 U22765 ( .A1(n19905), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n19880) );
  NAND2_X1 U22766 ( .A1(n19890), .A2(n19879), .ZN(n19894) );
  NAND2_X1 U22767 ( .A1(n19880), .A2(n19894), .ZN(P1_U2946) );
  AOI22_X1 U22768 ( .A1(n19905), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n19882) );
  NAND2_X1 U22769 ( .A1(n19890), .A2(n19881), .ZN(n19896) );
  NAND2_X1 U22770 ( .A1(n19882), .A2(n19896), .ZN(P1_U2947) );
  AOI22_X1 U22771 ( .A1(n19905), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n19884) );
  NAND2_X1 U22772 ( .A1(n19890), .A2(n19883), .ZN(n19898) );
  NAND2_X1 U22773 ( .A1(n19884), .A2(n19898), .ZN(P1_U2948) );
  AOI22_X1 U22774 ( .A1(n19905), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n19886) );
  NAND2_X1 U22775 ( .A1(n19890), .A2(n19885), .ZN(n19900) );
  NAND2_X1 U22776 ( .A1(n19886), .A2(n19900), .ZN(P1_U2949) );
  AOI22_X1 U22777 ( .A1(n19905), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n19888) );
  NAND2_X1 U22778 ( .A1(n19890), .A2(n19887), .ZN(n19902) );
  NAND2_X1 U22779 ( .A1(n19888), .A2(n19902), .ZN(P1_U2950) );
  AOI22_X1 U22780 ( .A1(n19905), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n19891) );
  NAND2_X1 U22781 ( .A1(n19890), .A2(n19889), .ZN(n19906) );
  NAND2_X1 U22782 ( .A1(n19891), .A2(n19906), .ZN(P1_U2951) );
  AOI22_X1 U22783 ( .A1(n19905), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n19893) );
  NAND2_X1 U22784 ( .A1(n19893), .A2(n19892), .ZN(P1_U2960) );
  AOI22_X1 U22785 ( .A1(n19905), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n19895) );
  NAND2_X1 U22786 ( .A1(n19895), .A2(n19894), .ZN(P1_U2961) );
  AOI22_X1 U22787 ( .A1(n19905), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n19897) );
  NAND2_X1 U22788 ( .A1(n19897), .A2(n19896), .ZN(P1_U2962) );
  AOI22_X1 U22789 ( .A1(n19905), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n19899) );
  NAND2_X1 U22790 ( .A1(n19899), .A2(n19898), .ZN(P1_U2963) );
  AOI22_X1 U22791 ( .A1(n19905), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n19901) );
  NAND2_X1 U22792 ( .A1(n19901), .A2(n19900), .ZN(P1_U2964) );
  AOI22_X1 U22793 ( .A1(n19905), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n19903) );
  NAND2_X1 U22794 ( .A1(n19903), .A2(n19902), .ZN(P1_U2965) );
  AOI22_X1 U22795 ( .A1(n19905), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n19907) );
  NAND2_X1 U22796 ( .A1(n19907), .A2(n19906), .ZN(P1_U2966) );
  AOI22_X1 U22797 ( .A1(n19908), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n12105), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U22798 ( .A1(n9582), .A2(n19912), .B1(n19911), .B2(n19910), .ZN(
        n19913) );
  OAI211_X1 U22799 ( .C1(n19916), .C2(n19915), .A(n19914), .B(n19913), .ZN(
        P1_U2995) );
  AOI21_X1 U22800 ( .B1(n19951), .B2(n19950), .A(n19917), .ZN(n19934) );
  AOI222_X1 U22801 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n12105), .B1(n19925), 
        .B2(n19918), .C1(n19929), .C2(n9582), .ZN(n19921) );
  OAI211_X1 U22802 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n19928), .B(n19919), .ZN(n19920) );
  OAI211_X1 U22803 ( .C1(n19934), .C2(n19922), .A(n19921), .B(n19920), .ZN(
        P1_U3027) );
  INV_X1 U22804 ( .A(n19923), .ZN(n19924) );
  AOI21_X1 U22805 ( .B1(n19926), .B2(n19925), .A(n19924), .ZN(n19932) );
  INV_X1 U22806 ( .A(n19927), .ZN(n19930) );
  AOI22_X1 U22807 ( .A1(n19930), .A2(n19929), .B1(n19933), .B2(n19928), .ZN(
        n19931) );
  OAI211_X1 U22808 ( .C1(n19934), .C2(n19933), .A(n19932), .B(n19931), .ZN(
        P1_U3028) );
  NAND2_X1 U22809 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19935), .ZN(
        n19955) );
  NOR3_X1 U22810 ( .A1(n19937), .A2(n19941), .A3(n19936), .ZN(n19939) );
  AOI211_X1 U22811 ( .C1(n19941), .C2(n19940), .A(n19939), .B(n19938), .ZN(
        n19953) );
  OAI22_X1 U22812 ( .A1(n19945), .A2(n19944), .B1(n19943), .B2(n19942), .ZN(
        n19949) );
  NOR2_X1 U22813 ( .A1(n19947), .A2(n19946), .ZN(n19948) );
  AOI211_X1 U22814 ( .C1(n19951), .C2(n19950), .A(n19949), .B(n19948), .ZN(
        n19952) );
  OAI221_X1 U22815 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19955), .C1(
        n19954), .C2(n19953), .A(n19952), .ZN(P1_U3029) );
  NOR2_X1 U22816 ( .A1(n11548), .A2(n19956), .ZN(P1_U3032) );
  NOR2_X2 U22817 ( .A1(n19957), .A2(n19960), .ZN(n19958) );
  AOI22_X1 U22818 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20001), .B1(DATAI_24_), 
        .B2(n19958), .ZN(n20505) );
  INV_X1 U22819 ( .A(n20505), .ZN(n20454) );
  NAND2_X1 U22820 ( .A1(n20002), .A2(n12501), .ZN(n20364) );
  NOR3_X1 U22821 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20013) );
  NAND2_X1 U22822 ( .A1(n20416), .A2(n20013), .ZN(n19969) );
  INV_X1 U22823 ( .A(n19969), .ZN(n20003) );
  AOI22_X1 U22824 ( .A1(n20547), .A2(n20454), .B1(n20495), .B2(n20003), .ZN(
        n19978) );
  AND2_X1 U22825 ( .A1(n20234), .A2(n20287), .ZN(n19974) );
  INV_X1 U22826 ( .A(n19964), .ZN(n19973) );
  NAND2_X1 U22827 ( .A1(n19973), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20445) );
  NAND3_X1 U22828 ( .A1(n20029), .A2(n20418), .A3(n19966), .ZN(n19967) );
  NAND2_X1 U22829 ( .A1(n20418), .A2(n20641), .ZN(n20358) );
  NAND2_X1 U22830 ( .A1(n19967), .A2(n20358), .ZN(n19972) );
  OR2_X1 U22831 ( .A1(n20233), .A2(n19968), .ZN(n20072) );
  OR2_X1 U22832 ( .A1(n20072), .A2(n9648), .ZN(n19975) );
  AOI22_X1 U22833 ( .A1(n19972), .A2(n19975), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n19969), .ZN(n19970) );
  OAI211_X1 U22834 ( .C1(n19974), .C2(n20640), .A(n20294), .B(n19970), .ZN(
        n20006) );
  NOR2_X2 U22835 ( .A1(n19971), .A2(n20119), .ZN(n20496) );
  INV_X1 U22836 ( .A(n19972), .ZN(n19976) );
  NOR2_X1 U22837 ( .A1(n19973), .A2(n20640), .ZN(n20288) );
  INV_X1 U22838 ( .A(n20288), .ZN(n20236) );
  INV_X1 U22839 ( .A(n19974), .ZN(n20115) );
  OAI22_X1 U22840 ( .A1(n19976), .A2(n19975), .B1(n20236), .B2(n20115), .ZN(
        n20005) );
  AOI22_X1 U22841 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20006), .B1(
        n20496), .B2(n20005), .ZN(n19977) );
  OAI211_X1 U22842 ( .C1(n20457), .C2(n20029), .A(n19978), .B(n19977), .ZN(
        P1_U3033) );
  AOI22_X1 U22843 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20001), .B1(DATAI_25_), 
        .B2(n19958), .ZN(n20511) );
  INV_X1 U22844 ( .A(n20511), .ZN(n20458) );
  NAND2_X1 U22845 ( .A1(n20002), .A2(n19979), .ZN(n20377) );
  AOI22_X1 U22846 ( .A1(n20547), .A2(n20458), .B1(n20506), .B2(n20003), .ZN(
        n19982) );
  NOR2_X2 U22847 ( .A1(n19980), .A2(n20119), .ZN(n20507) );
  AOI22_X1 U22848 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20006), .B1(
        n20507), .B2(n20005), .ZN(n19981) );
  OAI211_X1 U22849 ( .C1(n20461), .C2(n20029), .A(n19982), .B(n19981), .ZN(
        P1_U3034) );
  AOI22_X2 U22850 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20001), .B1(DATAI_18_), 
        .B2(n19958), .ZN(n20465) );
  AOI22_X1 U22851 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20001), .B1(DATAI_26_), 
        .B2(n19958), .ZN(n20517) );
  INV_X1 U22852 ( .A(n20517), .ZN(n20462) );
  NAND2_X1 U22853 ( .A1(n20002), .A2(n19983), .ZN(n20382) );
  AOI22_X1 U22854 ( .A1(n20547), .A2(n20462), .B1(n20512), .B2(n20003), .ZN(
        n19986) );
  NOR2_X2 U22855 ( .A1(n19984), .A2(n20119), .ZN(n20513) );
  AOI22_X1 U22856 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20006), .B1(
        n20513), .B2(n20005), .ZN(n19985) );
  OAI211_X1 U22857 ( .C1(n20465), .C2(n20029), .A(n19986), .B(n19985), .ZN(
        P1_U3035) );
  AOI22_X1 U22858 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20001), .B1(DATAI_19_), 
        .B2(n19958), .ZN(n20469) );
  AOI22_X1 U22859 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20001), .B1(DATAI_27_), 
        .B2(n19958), .ZN(n20523) );
  INV_X1 U22860 ( .A(n20523), .ZN(n20466) );
  NAND2_X1 U22861 ( .A1(n20002), .A2(n19987), .ZN(n20387) );
  AOI22_X1 U22862 ( .A1(n20547), .A2(n20466), .B1(n20518), .B2(n20003), .ZN(
        n19990) );
  NOR2_X2 U22863 ( .A1(n19988), .A2(n20119), .ZN(n20519) );
  AOI22_X1 U22864 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20006), .B1(
        n20519), .B2(n20005), .ZN(n19989) );
  OAI211_X1 U22865 ( .C1(n20469), .C2(n20029), .A(n19990), .B(n19989), .ZN(
        P1_U3036) );
  AOI22_X1 U22866 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20001), .B1(DATAI_20_), 
        .B2(n19958), .ZN(n20473) );
  AOI22_X1 U22867 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20001), .B1(DATAI_28_), 
        .B2(n19958), .ZN(n20529) );
  INV_X1 U22868 ( .A(n20529), .ZN(n20470) );
  NAND2_X1 U22869 ( .A1(n20002), .A2(n11180), .ZN(n20392) );
  AOI22_X1 U22870 ( .A1(n20547), .A2(n20470), .B1(n20524), .B2(n20003), .ZN(
        n19993) );
  NOR2_X2 U22871 ( .A1(n19991), .A2(n20119), .ZN(n20525) );
  AOI22_X1 U22872 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20006), .B1(
        n20525), .B2(n20005), .ZN(n19992) );
  OAI211_X1 U22873 ( .C1(n20473), .C2(n20029), .A(n19993), .B(n19992), .ZN(
        P1_U3037) );
  AOI22_X1 U22874 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20001), .B1(DATAI_21_), 
        .B2(n19958), .ZN(n20477) );
  AOI22_X1 U22875 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20001), .B1(DATAI_29_), 
        .B2(n19958), .ZN(n20535) );
  INV_X1 U22876 ( .A(n20535), .ZN(n20474) );
  NAND2_X1 U22877 ( .A1(n20002), .A2(n19994), .ZN(n20397) );
  AOI22_X1 U22878 ( .A1(n20547), .A2(n20474), .B1(n20530), .B2(n20003), .ZN(
        n19997) );
  NOR2_X2 U22879 ( .A1(n19995), .A2(n20119), .ZN(n20531) );
  AOI22_X1 U22880 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20006), .B1(
        n20531), .B2(n20005), .ZN(n19996) );
  OAI211_X1 U22881 ( .C1(n20477), .C2(n20029), .A(n19997), .B(n19996), .ZN(
        P1_U3038) );
  AOI22_X1 U22882 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20001), .B1(DATAI_22_), 
        .B2(n19958), .ZN(n20481) );
  AOI22_X1 U22883 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20001), .B1(DATAI_30_), 
        .B2(n19958), .ZN(n20541) );
  INV_X1 U22884 ( .A(n20541), .ZN(n20478) );
  NAND2_X1 U22885 ( .A1(n20002), .A2(n11270), .ZN(n20402) );
  AOI22_X1 U22886 ( .A1(n20547), .A2(n20478), .B1(n20536), .B2(n20003), .ZN(
        n20000) );
  NOR2_X2 U22887 ( .A1(n19998), .A2(n20119), .ZN(n20537) );
  AOI22_X1 U22888 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20006), .B1(
        n20537), .B2(n20005), .ZN(n19999) );
  OAI211_X1 U22889 ( .C1(n20481), .C2(n20029), .A(n20000), .B(n19999), .ZN(
        P1_U3039) );
  AOI22_X1 U22890 ( .A1(DATAI_23_), .A2(n19958), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20001), .ZN(n20489) );
  AOI22_X1 U22891 ( .A1(DATAI_31_), .A2(n19958), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20001), .ZN(n20552) );
  INV_X1 U22892 ( .A(n20552), .ZN(n20484) );
  NAND2_X1 U22893 ( .A1(n20002), .A2(n11254), .ZN(n20408) );
  AOI22_X1 U22894 ( .A1(n20547), .A2(n20484), .B1(n20542), .B2(n20003), .ZN(
        n20008) );
  NOR2_X2 U22895 ( .A1(n20119), .A2(n20004), .ZN(n20544) );
  AOI22_X1 U22896 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20006), .B1(
        n20544), .B2(n20005), .ZN(n20007) );
  OAI211_X1 U22897 ( .C1(n20489), .C2(n20029), .A(n20008), .B(n20007), .ZN(
        P1_U3040) );
  INV_X1 U22898 ( .A(n20072), .ZN(n20038) );
  INV_X1 U22899 ( .A(n20009), .ZN(n20261) );
  INV_X1 U22900 ( .A(n20013), .ZN(n20010) );
  NOR2_X1 U22901 ( .A1(n20416), .A2(n20010), .ZN(n20030) );
  AOI21_X1 U22902 ( .B1(n20038), .B2(n20261), .A(n20030), .ZN(n20011) );
  OAI22_X1 U22903 ( .A1(n20011), .A2(n20493), .B1(n20010), .B2(n20640), .ZN(
        n20031) );
  AOI22_X1 U22904 ( .A1(n20031), .A2(n20496), .B1(n20495), .B2(n20030), .ZN(
        n20015) );
  OAI21_X1 U22905 ( .B1(n20076), .B2(n20641), .A(n20011), .ZN(n20012) );
  OAI221_X1 U22906 ( .B1(n20418), .B2(n20013), .C1(n20493), .C2(n20012), .A(
        n20499), .ZN(n20033) );
  AOI22_X1 U22907 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n20454), .ZN(n20014) );
  OAI211_X1 U22908 ( .C1(n20457), .C2(n20064), .A(n20015), .B(n20014), .ZN(
        P1_U3041) );
  AOI22_X1 U22909 ( .A1(n20031), .A2(n20507), .B1(n20506), .B2(n20030), .ZN(
        n20017) );
  AOI22_X1 U22910 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n20458), .ZN(n20016) );
  OAI211_X1 U22911 ( .C1(n20461), .C2(n20064), .A(n20017), .B(n20016), .ZN(
        P1_U3042) );
  AOI22_X1 U22912 ( .A1(n20031), .A2(n20513), .B1(n20512), .B2(n20030), .ZN(
        n20019) );
  AOI22_X1 U22913 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n20462), .ZN(n20018) );
  OAI211_X1 U22914 ( .C1(n20465), .C2(n20064), .A(n20019), .B(n20018), .ZN(
        P1_U3043) );
  AOI22_X1 U22915 ( .A1(n20031), .A2(n20519), .B1(n20518), .B2(n20030), .ZN(
        n20021) );
  AOI22_X1 U22916 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n20466), .ZN(n20020) );
  OAI211_X1 U22917 ( .C1(n20469), .C2(n20064), .A(n20021), .B(n20020), .ZN(
        P1_U3044) );
  AOI22_X1 U22918 ( .A1(n20031), .A2(n20525), .B1(n20524), .B2(n20030), .ZN(
        n20023) );
  AOI22_X1 U22919 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n20470), .ZN(n20022) );
  OAI211_X1 U22920 ( .C1(n20473), .C2(n20064), .A(n20023), .B(n20022), .ZN(
        P1_U3045) );
  AOI22_X1 U22921 ( .A1(n20031), .A2(n20531), .B1(n20530), .B2(n20030), .ZN(
        n20025) );
  INV_X1 U22922 ( .A(n20064), .ZN(n20026) );
  INV_X1 U22923 ( .A(n20477), .ZN(n20532) );
  AOI22_X1 U22924 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20033), .B1(
        n20026), .B2(n20532), .ZN(n20024) );
  OAI211_X1 U22925 ( .C1(n20535), .C2(n20029), .A(n20025), .B(n20024), .ZN(
        P1_U3046) );
  AOI22_X1 U22926 ( .A1(n20031), .A2(n20537), .B1(n20536), .B2(n20030), .ZN(
        n20028) );
  INV_X1 U22927 ( .A(n20481), .ZN(n20538) );
  AOI22_X1 U22928 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20033), .B1(
        n20026), .B2(n20538), .ZN(n20027) );
  OAI211_X1 U22929 ( .C1(n20541), .C2(n20029), .A(n20028), .B(n20027), .ZN(
        P1_U3047) );
  AOI22_X1 U22930 ( .A1(n20031), .A2(n20544), .B1(n20542), .B2(n20030), .ZN(
        n20035) );
  AOI22_X1 U22931 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20033), .B1(
        n20032), .B2(n20484), .ZN(n20034) );
  OAI211_X1 U22932 ( .C1(n20489), .C2(n20064), .A(n20035), .B(n20034), .ZN(
        P1_U3048) );
  NOR3_X1 U22933 ( .A1(n11542), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20078) );
  NAND2_X1 U22934 ( .A1(n20416), .A2(n20078), .ZN(n20063) );
  OAI22_X1 U22935 ( .A1(n20064), .A2(n20505), .B1(n20364), .B2(n20063), .ZN(
        n20036) );
  INV_X1 U22936 ( .A(n20036), .ZN(n20044) );
  NAND2_X1 U22937 ( .A1(n20106), .A2(n20064), .ZN(n20037) );
  AOI21_X1 U22938 ( .B1(n20037), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20493), 
        .ZN(n20040) );
  NAND2_X1 U22939 ( .A1(n20038), .A2(n9648), .ZN(n20041) );
  AOI22_X1 U22940 ( .A1(n20040), .A2(n20041), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20063), .ZN(n20039) );
  OR2_X1 U22941 ( .A1(n20287), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20171) );
  NAND2_X1 U22942 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20171), .ZN(n20168) );
  NAND3_X1 U22943 ( .A1(n20294), .A2(n20039), .A3(n20168), .ZN(n20067) );
  INV_X1 U22944 ( .A(n20040), .ZN(n20042) );
  AOI22_X1 U22945 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20067), .B1(
        n20496), .B2(n20066), .ZN(n20043) );
  OAI211_X1 U22946 ( .C1(n20457), .C2(n20106), .A(n20044), .B(n20043), .ZN(
        P1_U3049) );
  OAI22_X1 U22947 ( .A1(n20064), .A2(n20511), .B1(n20063), .B2(n20377), .ZN(
        n20045) );
  INV_X1 U22948 ( .A(n20045), .ZN(n20047) );
  AOI22_X1 U22949 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20067), .B1(
        n20507), .B2(n20066), .ZN(n20046) );
  OAI211_X1 U22950 ( .C1(n20461), .C2(n20106), .A(n20047), .B(n20046), .ZN(
        P1_U3050) );
  OAI22_X1 U22951 ( .A1(n20064), .A2(n20517), .B1(n20063), .B2(n20382), .ZN(
        n20048) );
  INV_X1 U22952 ( .A(n20048), .ZN(n20050) );
  AOI22_X1 U22953 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20067), .B1(
        n20513), .B2(n20066), .ZN(n20049) );
  OAI211_X1 U22954 ( .C1(n20465), .C2(n20106), .A(n20050), .B(n20049), .ZN(
        P1_U3051) );
  OAI22_X1 U22955 ( .A1(n20106), .A2(n20469), .B1(n20063), .B2(n20387), .ZN(
        n20051) );
  INV_X1 U22956 ( .A(n20051), .ZN(n20053) );
  AOI22_X1 U22957 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20067), .B1(
        n20519), .B2(n20066), .ZN(n20052) );
  OAI211_X1 U22958 ( .C1(n20523), .C2(n20064), .A(n20053), .B(n20052), .ZN(
        P1_U3052) );
  OAI22_X1 U22959 ( .A1(n20106), .A2(n20473), .B1(n20063), .B2(n20392), .ZN(
        n20054) );
  INV_X1 U22960 ( .A(n20054), .ZN(n20056) );
  AOI22_X1 U22961 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20067), .B1(
        n20525), .B2(n20066), .ZN(n20055) );
  OAI211_X1 U22962 ( .C1(n20529), .C2(n20064), .A(n20056), .B(n20055), .ZN(
        P1_U3053) );
  OAI22_X1 U22963 ( .A1(n20106), .A2(n20477), .B1(n20063), .B2(n20397), .ZN(
        n20057) );
  INV_X1 U22964 ( .A(n20057), .ZN(n20059) );
  AOI22_X1 U22965 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20067), .B1(
        n20531), .B2(n20066), .ZN(n20058) );
  OAI211_X1 U22966 ( .C1(n20535), .C2(n20064), .A(n20059), .B(n20058), .ZN(
        P1_U3054) );
  OAI22_X1 U22967 ( .A1(n20106), .A2(n20481), .B1(n20063), .B2(n20402), .ZN(
        n20060) );
  INV_X1 U22968 ( .A(n20060), .ZN(n20062) );
  AOI22_X1 U22969 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20067), .B1(
        n20537), .B2(n20066), .ZN(n20061) );
  OAI211_X1 U22970 ( .C1(n20541), .C2(n20064), .A(n20062), .B(n20061), .ZN(
        P1_U3055) );
  OAI22_X1 U22971 ( .A1(n20064), .A2(n20552), .B1(n20063), .B2(n20408), .ZN(
        n20065) );
  INV_X1 U22972 ( .A(n20065), .ZN(n20069) );
  AOI22_X1 U22973 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20067), .B1(
        n20544), .B2(n20066), .ZN(n20068) );
  OAI211_X1 U22974 ( .C1(n20489), .C2(n20106), .A(n20069), .B(n20068), .ZN(
        P1_U3056) );
  INV_X1 U22975 ( .A(n20076), .ZN(n20070) );
  AOI21_X1 U22976 ( .B1(n20070), .B2(n20497), .A(n20493), .ZN(n20081) );
  AND2_X1 U22977 ( .A1(n20071), .A2(n11614), .ZN(n20329) );
  INV_X1 U22978 ( .A(n20329), .ZN(n20491) );
  OR2_X1 U22979 ( .A1(n20072), .A2(n20491), .ZN(n20074) );
  INV_X1 U22980 ( .A(n20328), .ZN(n20073) );
  NAND2_X1 U22981 ( .A1(n20073), .A2(n20363), .ZN(n20105) );
  INV_X1 U22982 ( .A(n20080), .ZN(n20075) );
  INV_X1 U22983 ( .A(n20496), .ZN(n20376) );
  OAI22_X1 U22984 ( .A1(n20100), .A2(n20457), .B1(n20364), .B2(n20105), .ZN(
        n20077) );
  INV_X1 U22985 ( .A(n20077), .ZN(n20084) );
  INV_X1 U22986 ( .A(n20078), .ZN(n20079) );
  AOI22_X1 U22987 ( .A1(n20081), .A2(n20080), .B1(n20493), .B2(n20079), .ZN(
        n20082) );
  NAND2_X1 U22988 ( .A1(n20499), .A2(n20082), .ZN(n20108) );
  INV_X1 U22989 ( .A(n20106), .ZN(n20102) );
  AOI22_X1 U22990 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20108), .B1(
        n20102), .B2(n20454), .ZN(n20083) );
  OAI211_X1 U22991 ( .C1(n20111), .C2(n20376), .A(n20084), .B(n20083), .ZN(
        P1_U3057) );
  INV_X1 U22992 ( .A(n20507), .ZN(n20381) );
  OAI22_X1 U22993 ( .A1(n20100), .A2(n20461), .B1(n20377), .B2(n20105), .ZN(
        n20085) );
  INV_X1 U22994 ( .A(n20085), .ZN(n20087) );
  AOI22_X1 U22995 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20108), .B1(
        n20102), .B2(n20458), .ZN(n20086) );
  OAI211_X1 U22996 ( .C1(n20111), .C2(n20381), .A(n20087), .B(n20086), .ZN(
        P1_U3058) );
  INV_X1 U22997 ( .A(n20513), .ZN(n20386) );
  OAI22_X1 U22998 ( .A1(n20100), .A2(n20465), .B1(n20382), .B2(n20105), .ZN(
        n20088) );
  INV_X1 U22999 ( .A(n20088), .ZN(n20090) );
  AOI22_X1 U23000 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20108), .B1(
        n20102), .B2(n20462), .ZN(n20089) );
  OAI211_X1 U23001 ( .C1(n20111), .C2(n20386), .A(n20090), .B(n20089), .ZN(
        P1_U3059) );
  INV_X1 U23002 ( .A(n20519), .ZN(n20391) );
  OAI22_X1 U23003 ( .A1(n20106), .A2(n20523), .B1(n20105), .B2(n20387), .ZN(
        n20091) );
  INV_X1 U23004 ( .A(n20091), .ZN(n20093) );
  INV_X1 U23005 ( .A(n20469), .ZN(n20520) );
  AOI22_X1 U23006 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20108), .B1(
        n20137), .B2(n20520), .ZN(n20092) );
  OAI211_X1 U23007 ( .C1(n20111), .C2(n20391), .A(n20093), .B(n20092), .ZN(
        P1_U3060) );
  INV_X1 U23008 ( .A(n20525), .ZN(n20396) );
  OAI22_X1 U23009 ( .A1(n20106), .A2(n20529), .B1(n20105), .B2(n20392), .ZN(
        n20094) );
  INV_X1 U23010 ( .A(n20094), .ZN(n20096) );
  INV_X1 U23011 ( .A(n20473), .ZN(n20526) );
  AOI22_X1 U23012 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20108), .B1(
        n20137), .B2(n20526), .ZN(n20095) );
  OAI211_X1 U23013 ( .C1(n20111), .C2(n20396), .A(n20096), .B(n20095), .ZN(
        P1_U3061) );
  INV_X1 U23014 ( .A(n20531), .ZN(n20401) );
  OAI22_X1 U23015 ( .A1(n20100), .A2(n20477), .B1(n20105), .B2(n20397), .ZN(
        n20097) );
  INV_X1 U23016 ( .A(n20097), .ZN(n20099) );
  AOI22_X1 U23017 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20108), .B1(
        n20102), .B2(n20474), .ZN(n20098) );
  OAI211_X1 U23018 ( .C1(n20111), .C2(n20401), .A(n20099), .B(n20098), .ZN(
        P1_U3062) );
  INV_X1 U23019 ( .A(n20537), .ZN(n20406) );
  OAI22_X1 U23020 ( .A1(n20100), .A2(n20481), .B1(n20105), .B2(n20402), .ZN(
        n20101) );
  INV_X1 U23021 ( .A(n20101), .ZN(n20104) );
  AOI22_X1 U23022 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20108), .B1(
        n20102), .B2(n20478), .ZN(n20103) );
  OAI211_X1 U23023 ( .C1(n20111), .C2(n20406), .A(n20104), .B(n20103), .ZN(
        P1_U3063) );
  INV_X1 U23024 ( .A(n20544), .ZN(n20414) );
  OAI22_X1 U23025 ( .A1(n20106), .A2(n20552), .B1(n20408), .B2(n20105), .ZN(
        n20107) );
  INV_X1 U23026 ( .A(n20107), .ZN(n20110) );
  INV_X1 U23027 ( .A(n20489), .ZN(n20546) );
  AOI22_X1 U23028 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20108), .B1(
        n20137), .B2(n20546), .ZN(n20109) );
  OAI211_X1 U23029 ( .C1(n20111), .C2(n20414), .A(n20110), .B(n20109), .ZN(
        P1_U3064) );
  NOR3_X1 U23030 ( .A1(n15558), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20144) );
  INV_X1 U23031 ( .A(n20144), .ZN(n20141) );
  NOR2_X1 U23032 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20141), .ZN(
        n20136) );
  NOR2_X1 U23033 ( .A1(n13417), .A2(n20113), .ZN(n20202) );
  NAND3_X1 U23034 ( .A1(n20202), .A2(n20418), .A3(n13694), .ZN(n20114) );
  OAI21_X1 U23035 ( .B1(n20115), .B2(n20445), .A(n20114), .ZN(n20135) );
  AOI22_X1 U23036 ( .A1(n20495), .A2(n20136), .B1(n20496), .B2(n20135), .ZN(
        n20122) );
  INV_X1 U23037 ( .A(n20202), .ZN(n20118) );
  INV_X1 U23038 ( .A(n20165), .ZN(n20116) );
  OAI21_X1 U23039 ( .B1(n20137), .B2(n20116), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20117) );
  OAI21_X1 U23040 ( .B1(n9648), .B2(n20118), .A(n20117), .ZN(n20120) );
  AOI22_X1 U23041 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20138), .B1(
        n20137), .B2(n20454), .ZN(n20121) );
  OAI211_X1 U23042 ( .C1(n20457), .C2(n20165), .A(n20122), .B(n20121), .ZN(
        P1_U3065) );
  AOI22_X1 U23043 ( .A1(n20506), .A2(n20136), .B1(n20507), .B2(n20135), .ZN(
        n20124) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20138), .B1(
        n20137), .B2(n20458), .ZN(n20123) );
  OAI211_X1 U23045 ( .C1(n20461), .C2(n20165), .A(n20124), .B(n20123), .ZN(
        P1_U3066) );
  AOI22_X1 U23046 ( .A1(n20512), .A2(n20136), .B1(n20513), .B2(n20135), .ZN(
        n20126) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20138), .B1(
        n20137), .B2(n20462), .ZN(n20125) );
  OAI211_X1 U23048 ( .C1(n20465), .C2(n20165), .A(n20126), .B(n20125), .ZN(
        P1_U3067) );
  AOI22_X1 U23049 ( .A1(n20518), .A2(n20136), .B1(n20519), .B2(n20135), .ZN(
        n20128) );
  AOI22_X1 U23050 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20138), .B1(
        n20137), .B2(n20466), .ZN(n20127) );
  OAI211_X1 U23051 ( .C1(n20469), .C2(n20165), .A(n20128), .B(n20127), .ZN(
        P1_U3068) );
  AOI22_X1 U23052 ( .A1(n20524), .A2(n20136), .B1(n20525), .B2(n20135), .ZN(
        n20130) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20138), .B1(
        n20137), .B2(n20470), .ZN(n20129) );
  OAI211_X1 U23054 ( .C1(n20473), .C2(n20165), .A(n20130), .B(n20129), .ZN(
        P1_U3069) );
  AOI22_X1 U23055 ( .A1(n20530), .A2(n20136), .B1(n20531), .B2(n20135), .ZN(
        n20132) );
  AOI22_X1 U23056 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20138), .B1(
        n20137), .B2(n20474), .ZN(n20131) );
  OAI211_X1 U23057 ( .C1(n20477), .C2(n20165), .A(n20132), .B(n20131), .ZN(
        P1_U3070) );
  AOI22_X1 U23058 ( .A1(n20536), .A2(n20136), .B1(n20537), .B2(n20135), .ZN(
        n20134) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20138), .B1(
        n20137), .B2(n20478), .ZN(n20133) );
  OAI211_X1 U23060 ( .C1(n20481), .C2(n20165), .A(n20134), .B(n20133), .ZN(
        P1_U3071) );
  AOI22_X1 U23061 ( .A1(n20542), .A2(n20136), .B1(n20544), .B2(n20135), .ZN(
        n20140) );
  AOI22_X1 U23062 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20138), .B1(
        n20137), .B2(n20484), .ZN(n20139) );
  OAI211_X1 U23063 ( .C1(n20489), .C2(n20165), .A(n20140), .B(n20139), .ZN(
        P1_U3072) );
  NOR2_X1 U23064 ( .A1(n20416), .A2(n20141), .ZN(n20159) );
  AOI21_X1 U23065 ( .B1(n20202), .B2(n20261), .A(n20159), .ZN(n20142) );
  OAI22_X1 U23066 ( .A1(n20142), .A2(n20493), .B1(n20141), .B2(n20640), .ZN(
        n20160) );
  AOI22_X1 U23067 ( .A1(n20160), .A2(n20496), .B1(n20495), .B2(n20159), .ZN(
        n20146) );
  OAI21_X1 U23068 ( .B1(n20207), .B2(n20641), .A(n20142), .ZN(n20143) );
  OAI221_X1 U23069 ( .B1(n20418), .B2(n20144), .C1(n20493), .C2(n20143), .A(
        n20499), .ZN(n20162) );
  INV_X1 U23070 ( .A(n20457), .ZN(n20502) );
  AOI22_X1 U23071 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20162), .B1(
        n20161), .B2(n20502), .ZN(n20145) );
  OAI211_X1 U23072 ( .C1(n20505), .C2(n20165), .A(n20146), .B(n20145), .ZN(
        P1_U3073) );
  AOI22_X1 U23073 ( .A1(n20160), .A2(n20507), .B1(n20506), .B2(n20159), .ZN(
        n20148) );
  INV_X1 U23074 ( .A(n20461), .ZN(n20508) );
  AOI22_X1 U23075 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20162), .B1(
        n20161), .B2(n20508), .ZN(n20147) );
  OAI211_X1 U23076 ( .C1(n20511), .C2(n20165), .A(n20148), .B(n20147), .ZN(
        P1_U3074) );
  AOI22_X1 U23077 ( .A1(n20160), .A2(n20513), .B1(n20512), .B2(n20159), .ZN(
        n20150) );
  INV_X1 U23078 ( .A(n20465), .ZN(n20514) );
  AOI22_X1 U23079 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20162), .B1(
        n20161), .B2(n20514), .ZN(n20149) );
  OAI211_X1 U23080 ( .C1(n20517), .C2(n20165), .A(n20150), .B(n20149), .ZN(
        P1_U3075) );
  AOI22_X1 U23081 ( .A1(n20160), .A2(n20519), .B1(n20518), .B2(n20159), .ZN(
        n20152) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20162), .B1(
        n20161), .B2(n20520), .ZN(n20151) );
  OAI211_X1 U23083 ( .C1(n20523), .C2(n20165), .A(n20152), .B(n20151), .ZN(
        P1_U3076) );
  AOI22_X1 U23084 ( .A1(n20160), .A2(n20525), .B1(n20524), .B2(n20159), .ZN(
        n20154) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20162), .B1(
        n20161), .B2(n20526), .ZN(n20153) );
  OAI211_X1 U23086 ( .C1(n20529), .C2(n20165), .A(n20154), .B(n20153), .ZN(
        P1_U3077) );
  AOI22_X1 U23087 ( .A1(n20160), .A2(n20531), .B1(n20530), .B2(n20159), .ZN(
        n20156) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20162), .B1(
        n20161), .B2(n20532), .ZN(n20155) );
  OAI211_X1 U23089 ( .C1(n20535), .C2(n20165), .A(n20156), .B(n20155), .ZN(
        P1_U3078) );
  AOI22_X1 U23090 ( .A1(n20160), .A2(n20537), .B1(n20536), .B2(n20159), .ZN(
        n20158) );
  AOI22_X1 U23091 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20162), .B1(
        n20161), .B2(n20538), .ZN(n20157) );
  OAI211_X1 U23092 ( .C1(n20541), .C2(n20165), .A(n20158), .B(n20157), .ZN(
        P1_U3079) );
  AOI22_X1 U23093 ( .A1(n20160), .A2(n20544), .B1(n20542), .B2(n20159), .ZN(
        n20164) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20162), .B1(
        n20161), .B2(n20546), .ZN(n20163) );
  OAI211_X1 U23095 ( .C1(n20552), .C2(n20165), .A(n20164), .B(n20163), .ZN(
        P1_U3080) );
  NAND2_X1 U23096 ( .A1(n20416), .A2(n11402), .ZN(n20194) );
  OAI22_X1 U23097 ( .A1(n20200), .A2(n20505), .B1(n20364), .B2(n20194), .ZN(
        n20166) );
  INV_X1 U23098 ( .A(n20166), .ZN(n20175) );
  NAND2_X1 U23099 ( .A1(n20229), .A2(n20200), .ZN(n20167) );
  AOI21_X1 U23100 ( .B1(n20167), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20493), 
        .ZN(n20170) );
  NAND2_X1 U23101 ( .A1(n20202), .A2(n9648), .ZN(n20172) );
  AOI22_X1 U23102 ( .A1(n20170), .A2(n20172), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20194), .ZN(n20169) );
  NAND3_X1 U23103 ( .A1(n20452), .A2(n20169), .A3(n20168), .ZN(n20197) );
  INV_X1 U23104 ( .A(n20170), .ZN(n20173) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20197), .B1(
        n20496), .B2(n20196), .ZN(n20174) );
  OAI211_X1 U23106 ( .C1(n20457), .C2(n20229), .A(n20175), .B(n20174), .ZN(
        P1_U3081) );
  OAI22_X1 U23107 ( .A1(n20200), .A2(n20511), .B1(n20377), .B2(n20194), .ZN(
        n20176) );
  INV_X1 U23108 ( .A(n20176), .ZN(n20178) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20197), .B1(
        n20507), .B2(n20196), .ZN(n20177) );
  OAI211_X1 U23110 ( .C1(n20461), .C2(n20229), .A(n20178), .B(n20177), .ZN(
        P1_U3082) );
  OAI22_X1 U23111 ( .A1(n20200), .A2(n20517), .B1(n20382), .B2(n20194), .ZN(
        n20179) );
  INV_X1 U23112 ( .A(n20179), .ZN(n20181) );
  AOI22_X1 U23113 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20197), .B1(
        n20513), .B2(n20196), .ZN(n20180) );
  OAI211_X1 U23114 ( .C1(n20465), .C2(n20229), .A(n20181), .B(n20180), .ZN(
        P1_U3083) );
  OAI22_X1 U23115 ( .A1(n20200), .A2(n20523), .B1(n20387), .B2(n20194), .ZN(
        n20182) );
  INV_X1 U23116 ( .A(n20182), .ZN(n20184) );
  AOI22_X1 U23117 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20197), .B1(
        n20519), .B2(n20196), .ZN(n20183) );
  OAI211_X1 U23118 ( .C1(n20469), .C2(n20229), .A(n20184), .B(n20183), .ZN(
        P1_U3084) );
  OAI22_X1 U23119 ( .A1(n20229), .A2(n20473), .B1(n20392), .B2(n20194), .ZN(
        n20185) );
  INV_X1 U23120 ( .A(n20185), .ZN(n20187) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20197), .B1(
        n20525), .B2(n20196), .ZN(n20186) );
  OAI211_X1 U23122 ( .C1(n20529), .C2(n20200), .A(n20187), .B(n20186), .ZN(
        P1_U3085) );
  OAI22_X1 U23123 ( .A1(n20229), .A2(n20477), .B1(n20397), .B2(n20194), .ZN(
        n20188) );
  INV_X1 U23124 ( .A(n20188), .ZN(n20190) );
  AOI22_X1 U23125 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20197), .B1(
        n20531), .B2(n20196), .ZN(n20189) );
  OAI211_X1 U23126 ( .C1(n20535), .C2(n20200), .A(n20190), .B(n20189), .ZN(
        P1_U3086) );
  OAI22_X1 U23127 ( .A1(n20200), .A2(n20541), .B1(n20402), .B2(n20194), .ZN(
        n20191) );
  INV_X1 U23128 ( .A(n20191), .ZN(n20193) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20197), .B1(
        n20537), .B2(n20196), .ZN(n20192) );
  OAI211_X1 U23130 ( .C1(n20481), .C2(n20229), .A(n20193), .B(n20192), .ZN(
        P1_U3087) );
  OAI22_X1 U23131 ( .A1(n20229), .A2(n20489), .B1(n20408), .B2(n20194), .ZN(
        n20195) );
  INV_X1 U23132 ( .A(n20195), .ZN(n20199) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20197), .B1(
        n20544), .B2(n20196), .ZN(n20198) );
  OAI211_X1 U23134 ( .C1(n20552), .C2(n20200), .A(n20199), .B(n20198), .ZN(
        P1_U3088) );
  INV_X1 U23135 ( .A(n20201), .ZN(n20224) );
  AOI21_X1 U23136 ( .B1(n20202), .B2(n20329), .A(n20224), .ZN(n20204) );
  OAI22_X1 U23137 ( .A1(n20204), .A2(n20493), .B1(n20203), .B2(n20640), .ZN(
        n20225) );
  AOI22_X1 U23138 ( .A1(n20225), .A2(n20496), .B1(n20495), .B2(n20224), .ZN(
        n20209) );
  NAND2_X1 U23139 ( .A1(n20205), .A2(n20204), .ZN(n20206) );
  OAI221_X1 U23140 ( .B1(n20418), .B2(n11402), .C1(n20493), .C2(n20206), .A(
        n20499), .ZN(n20226) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20226), .B1(
        n20257), .B2(n20502), .ZN(n20208) );
  OAI211_X1 U23142 ( .C1(n20505), .C2(n20229), .A(n20209), .B(n20208), .ZN(
        P1_U3089) );
  AOI22_X1 U23143 ( .A1(n20225), .A2(n20507), .B1(n20506), .B2(n20224), .ZN(
        n20211) );
  INV_X1 U23144 ( .A(n20229), .ZN(n20212) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20226), .B1(
        n20212), .B2(n20458), .ZN(n20210) );
  OAI211_X1 U23146 ( .C1(n20461), .C2(n20215), .A(n20211), .B(n20210), .ZN(
        P1_U3090) );
  AOI22_X1 U23147 ( .A1(n20225), .A2(n20513), .B1(n20512), .B2(n20224), .ZN(
        n20214) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20226), .B1(
        n20212), .B2(n20462), .ZN(n20213) );
  OAI211_X1 U23149 ( .C1(n20465), .C2(n20215), .A(n20214), .B(n20213), .ZN(
        P1_U3091) );
  AOI22_X1 U23150 ( .A1(n20225), .A2(n20519), .B1(n20518), .B2(n20224), .ZN(
        n20217) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20226), .B1(
        n20257), .B2(n20520), .ZN(n20216) );
  OAI211_X1 U23152 ( .C1(n20523), .C2(n20229), .A(n20217), .B(n20216), .ZN(
        P1_U3092) );
  AOI22_X1 U23153 ( .A1(n20225), .A2(n20525), .B1(n20524), .B2(n20224), .ZN(
        n20219) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20226), .B1(
        n20257), .B2(n20526), .ZN(n20218) );
  OAI211_X1 U23155 ( .C1(n20529), .C2(n20229), .A(n20219), .B(n20218), .ZN(
        P1_U3093) );
  AOI22_X1 U23156 ( .A1(n20225), .A2(n20531), .B1(n20530), .B2(n20224), .ZN(
        n20221) );
  AOI22_X1 U23157 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20226), .B1(
        n20257), .B2(n20532), .ZN(n20220) );
  OAI211_X1 U23158 ( .C1(n20535), .C2(n20229), .A(n20221), .B(n20220), .ZN(
        P1_U3094) );
  AOI22_X1 U23159 ( .A1(n20225), .A2(n20537), .B1(n20536), .B2(n20224), .ZN(
        n20223) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20226), .B1(
        n20257), .B2(n20538), .ZN(n20222) );
  OAI211_X1 U23161 ( .C1(n20541), .C2(n20229), .A(n20223), .B(n20222), .ZN(
        P1_U3095) );
  AOI22_X1 U23162 ( .A1(n20225), .A2(n20544), .B1(n20542), .B2(n20224), .ZN(
        n20228) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20226), .B1(
        n20257), .B2(n20546), .ZN(n20227) );
  OAI211_X1 U23164 ( .C1(n20552), .C2(n20229), .A(n20228), .B(n20227), .ZN(
        P1_U3096) );
  INV_X1 U23165 ( .A(n13690), .ZN(n20230) );
  INV_X1 U23166 ( .A(n20334), .ZN(n20232) );
  AND2_X1 U23167 ( .A1(n20233), .A2(n13417), .ZN(n20330) );
  NOR3_X1 U23168 ( .A1(n20363), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20265) );
  INV_X1 U23169 ( .A(n20265), .ZN(n20262) );
  NOR2_X1 U23170 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20262), .ZN(
        n20255) );
  AOI21_X1 U23171 ( .B1(n20330), .B2(n13694), .A(n20255), .ZN(n20238) );
  INV_X1 U23172 ( .A(n20234), .ZN(n20235) );
  AND2_X1 U23173 ( .A1(n20235), .A2(n20287), .ZN(n20361) );
  INV_X1 U23174 ( .A(n20361), .ZN(n20367) );
  OAI22_X1 U23175 ( .A1(n20238), .A2(n20493), .B1(n20236), .B2(n20367), .ZN(
        n20256) );
  AOI22_X1 U23176 ( .A1(n20256), .A2(n20496), .B1(n20495), .B2(n20255), .ZN(
        n20242) );
  INV_X1 U23177 ( .A(n20285), .ZN(n20237) );
  OAI21_X1 U23178 ( .B1(n20237), .B2(n20257), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20239) );
  NAND2_X1 U23179 ( .A1(n20239), .A2(n20238), .ZN(n20240) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20454), .ZN(n20241) );
  OAI211_X1 U23181 ( .C1(n20457), .C2(n20285), .A(n20242), .B(n20241), .ZN(
        P1_U3097) );
  AOI22_X1 U23182 ( .A1(n20256), .A2(n20507), .B1(n20506), .B2(n20255), .ZN(
        n20244) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20458), .ZN(n20243) );
  OAI211_X1 U23184 ( .C1(n20461), .C2(n20285), .A(n20244), .B(n20243), .ZN(
        P1_U3098) );
  AOI22_X1 U23185 ( .A1(n20256), .A2(n20513), .B1(n20512), .B2(n20255), .ZN(
        n20246) );
  AOI22_X1 U23186 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20462), .ZN(n20245) );
  OAI211_X1 U23187 ( .C1(n20465), .C2(n20285), .A(n20246), .B(n20245), .ZN(
        P1_U3099) );
  AOI22_X1 U23188 ( .A1(n20256), .A2(n20519), .B1(n20518), .B2(n20255), .ZN(
        n20248) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20466), .ZN(n20247) );
  OAI211_X1 U23190 ( .C1(n20469), .C2(n20285), .A(n20248), .B(n20247), .ZN(
        P1_U3100) );
  AOI22_X1 U23191 ( .A1(n20256), .A2(n20525), .B1(n20524), .B2(n20255), .ZN(
        n20250) );
  AOI22_X1 U23192 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20470), .ZN(n20249) );
  OAI211_X1 U23193 ( .C1(n20473), .C2(n20285), .A(n20250), .B(n20249), .ZN(
        P1_U3101) );
  AOI22_X1 U23194 ( .A1(n20256), .A2(n20531), .B1(n20530), .B2(n20255), .ZN(
        n20252) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20474), .ZN(n20251) );
  OAI211_X1 U23196 ( .C1(n20477), .C2(n20285), .A(n20252), .B(n20251), .ZN(
        P1_U3102) );
  AOI22_X1 U23197 ( .A1(n20256), .A2(n20537), .B1(n20536), .B2(n20255), .ZN(
        n20254) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20478), .ZN(n20253) );
  OAI211_X1 U23199 ( .C1(n20481), .C2(n20285), .A(n20254), .B(n20253), .ZN(
        P1_U3103) );
  AOI22_X1 U23200 ( .A1(n20256), .A2(n20544), .B1(n20542), .B2(n20255), .ZN(
        n20260) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20258), .B1(
        n20257), .B2(n20484), .ZN(n20259) );
  OAI211_X1 U23202 ( .C1(n20489), .C2(n20285), .A(n20260), .B(n20259), .ZN(
        P1_U3104) );
  NOR2_X1 U23203 ( .A1(n20416), .A2(n20262), .ZN(n20280) );
  AOI21_X1 U23204 ( .B1(n20330), .B2(n20261), .A(n20280), .ZN(n20263) );
  OAI22_X1 U23205 ( .A1(n20263), .A2(n20493), .B1(n20262), .B2(n20640), .ZN(
        n20281) );
  AOI22_X1 U23206 ( .A1(n20281), .A2(n20496), .B1(n20495), .B2(n20280), .ZN(
        n20267) );
  OAI21_X1 U23207 ( .B1(n20334), .B2(n20641), .A(n20263), .ZN(n20264) );
  OAI221_X1 U23208 ( .B1(n20418), .B2(n20265), .C1(n20493), .C2(n20264), .A(
        n20499), .ZN(n20282) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20282), .B1(
        n20322), .B2(n20502), .ZN(n20266) );
  OAI211_X1 U23210 ( .C1(n20505), .C2(n20285), .A(n20267), .B(n20266), .ZN(
        P1_U3105) );
  AOI22_X1 U23211 ( .A1(n20281), .A2(n20507), .B1(n20506), .B2(n20280), .ZN(
        n20269) );
  AOI22_X1 U23212 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20282), .B1(
        n20322), .B2(n20508), .ZN(n20268) );
  OAI211_X1 U23213 ( .C1(n20511), .C2(n20285), .A(n20269), .B(n20268), .ZN(
        P1_U3106) );
  AOI22_X1 U23214 ( .A1(n20281), .A2(n20513), .B1(n20512), .B2(n20280), .ZN(
        n20271) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20282), .B1(
        n20322), .B2(n20514), .ZN(n20270) );
  OAI211_X1 U23216 ( .C1(n20517), .C2(n20285), .A(n20271), .B(n20270), .ZN(
        P1_U3107) );
  AOI22_X1 U23217 ( .A1(n20281), .A2(n20519), .B1(n20518), .B2(n20280), .ZN(
        n20273) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20282), .B1(
        n20322), .B2(n20520), .ZN(n20272) );
  OAI211_X1 U23219 ( .C1(n20523), .C2(n20285), .A(n20273), .B(n20272), .ZN(
        P1_U3108) );
  AOI22_X1 U23220 ( .A1(n20281), .A2(n20525), .B1(n20524), .B2(n20280), .ZN(
        n20275) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20282), .B1(
        n20322), .B2(n20526), .ZN(n20274) );
  OAI211_X1 U23222 ( .C1(n20529), .C2(n20285), .A(n20275), .B(n20274), .ZN(
        P1_U3109) );
  AOI22_X1 U23223 ( .A1(n20281), .A2(n20531), .B1(n20530), .B2(n20280), .ZN(
        n20277) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20282), .B1(
        n20322), .B2(n20532), .ZN(n20276) );
  OAI211_X1 U23225 ( .C1(n20535), .C2(n20285), .A(n20277), .B(n20276), .ZN(
        P1_U3110) );
  AOI22_X1 U23226 ( .A1(n20281), .A2(n20537), .B1(n20536), .B2(n20280), .ZN(
        n20279) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20282), .B1(
        n20322), .B2(n20538), .ZN(n20278) );
  OAI211_X1 U23228 ( .C1(n20541), .C2(n20285), .A(n20279), .B(n20278), .ZN(
        P1_U3111) );
  AOI22_X1 U23229 ( .A1(n20281), .A2(n20544), .B1(n20542), .B2(n20280), .ZN(
        n20284) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20282), .B1(
        n20322), .B2(n20546), .ZN(n20283) );
  OAI211_X1 U23231 ( .C1(n20552), .C2(n20285), .A(n20284), .B(n20283), .ZN(
        P1_U3112) );
  NAND3_X1 U23232 ( .A1(n20320), .A2(n20306), .A3(n20418), .ZN(n20286) );
  NAND2_X1 U23233 ( .A1(n20286), .A2(n20358), .ZN(n20291) );
  OR2_X1 U23234 ( .A1(n20287), .A2(n20363), .ZN(n20446) );
  INV_X1 U23235 ( .A(n20446), .ZN(n20289) );
  NOR3_X1 U23236 ( .A1(n20363), .A2(n11542), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20336) );
  INV_X1 U23237 ( .A(n20336), .ZN(n20331) );
  NOR2_X1 U23238 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20331), .ZN(
        n20292) );
  INV_X1 U23239 ( .A(n20292), .ZN(n20319) );
  OAI22_X1 U23240 ( .A1(n20320), .A2(n20457), .B1(n20364), .B2(n20319), .ZN(
        n20290) );
  INV_X1 U23241 ( .A(n20290), .ZN(n20299) );
  INV_X1 U23242 ( .A(n20291), .ZN(n20297) );
  NAND2_X1 U23243 ( .A1(n20446), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20451) );
  OAI21_X1 U23244 ( .B1(n20371), .B2(n20292), .A(n20451), .ZN(n20293) );
  INV_X1 U23245 ( .A(n20293), .ZN(n20295) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20454), .ZN(n20298) );
  OAI211_X1 U23247 ( .C1(n20326), .C2(n20376), .A(n20299), .B(n20298), .ZN(
        P1_U3113) );
  OAI22_X1 U23248 ( .A1(n20306), .A2(n20511), .B1(n20377), .B2(n20319), .ZN(
        n20300) );
  INV_X1 U23249 ( .A(n20300), .ZN(n20302) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20323), .B1(
        n20353), .B2(n20508), .ZN(n20301) );
  OAI211_X1 U23251 ( .C1(n20326), .C2(n20381), .A(n20302), .B(n20301), .ZN(
        P1_U3114) );
  OAI22_X1 U23252 ( .A1(n20320), .A2(n20465), .B1(n20382), .B2(n20319), .ZN(
        n20303) );
  INV_X1 U23253 ( .A(n20303), .ZN(n20305) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20462), .ZN(n20304) );
  OAI211_X1 U23255 ( .C1(n20326), .C2(n20386), .A(n20305), .B(n20304), .ZN(
        P1_U3115) );
  OAI22_X1 U23256 ( .A1(n20306), .A2(n20523), .B1(n20387), .B2(n20319), .ZN(
        n20307) );
  INV_X1 U23257 ( .A(n20307), .ZN(n20309) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20323), .B1(
        n20353), .B2(n20520), .ZN(n20308) );
  OAI211_X1 U23259 ( .C1(n20326), .C2(n20391), .A(n20309), .B(n20308), .ZN(
        P1_U3116) );
  OAI22_X1 U23260 ( .A1(n20320), .A2(n20473), .B1(n20392), .B2(n20319), .ZN(
        n20310) );
  INV_X1 U23261 ( .A(n20310), .ZN(n20312) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20470), .ZN(n20311) );
  OAI211_X1 U23263 ( .C1(n20326), .C2(n20396), .A(n20312), .B(n20311), .ZN(
        P1_U3117) );
  OAI22_X1 U23264 ( .A1(n20320), .A2(n20477), .B1(n20397), .B2(n20319), .ZN(
        n20313) );
  INV_X1 U23265 ( .A(n20313), .ZN(n20315) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20474), .ZN(n20314) );
  OAI211_X1 U23267 ( .C1(n20326), .C2(n20401), .A(n20315), .B(n20314), .ZN(
        P1_U3118) );
  OAI22_X1 U23268 ( .A1(n20320), .A2(n20481), .B1(n20402), .B2(n20319), .ZN(
        n20316) );
  INV_X1 U23269 ( .A(n20316), .ZN(n20318) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20478), .ZN(n20317) );
  OAI211_X1 U23271 ( .C1(n20326), .C2(n20406), .A(n20318), .B(n20317), .ZN(
        P1_U3119) );
  OAI22_X1 U23272 ( .A1(n20320), .A2(n20489), .B1(n20408), .B2(n20319), .ZN(
        n20321) );
  INV_X1 U23273 ( .A(n20321), .ZN(n20325) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20323), .B1(
        n20322), .B2(n20484), .ZN(n20324) );
  OAI211_X1 U23275 ( .C1(n20326), .C2(n20414), .A(n20325), .B(n20324), .ZN(
        P1_U3120) );
  NOR2_X1 U23276 ( .A1(n20328), .A2(n20363), .ZN(n20351) );
  AOI21_X1 U23277 ( .B1(n20330), .B2(n20329), .A(n20351), .ZN(n20332) );
  OAI22_X1 U23278 ( .A1(n20332), .A2(n20493), .B1(n20331), .B2(n20640), .ZN(
        n20352) );
  AOI22_X1 U23279 ( .A1(n20352), .A2(n20496), .B1(n20495), .B2(n20351), .ZN(
        n20338) );
  OAI21_X1 U23280 ( .B1(n20334), .B2(n20333), .A(n20332), .ZN(n20335) );
  OAI221_X1 U23281 ( .B1(n20418), .B2(n20336), .C1(n20493), .C2(n20335), .A(
        n20499), .ZN(n20354) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20454), .ZN(n20337) );
  OAI211_X1 U23283 ( .C1(n20457), .C2(n20373), .A(n20338), .B(n20337), .ZN(
        P1_U3121) );
  AOI22_X1 U23284 ( .A1(n20352), .A2(n20507), .B1(n20506), .B2(n20351), .ZN(
        n20340) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20458), .ZN(n20339) );
  OAI211_X1 U23286 ( .C1(n20461), .C2(n20373), .A(n20340), .B(n20339), .ZN(
        P1_U3122) );
  AOI22_X1 U23287 ( .A1(n20352), .A2(n20513), .B1(n20512), .B2(n20351), .ZN(
        n20342) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20462), .ZN(n20341) );
  OAI211_X1 U23289 ( .C1(n20465), .C2(n20373), .A(n20342), .B(n20341), .ZN(
        P1_U3123) );
  AOI22_X1 U23290 ( .A1(n20352), .A2(n20519), .B1(n20518), .B2(n20351), .ZN(
        n20344) );
  AOI22_X1 U23291 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20466), .ZN(n20343) );
  OAI211_X1 U23292 ( .C1(n20469), .C2(n20373), .A(n20344), .B(n20343), .ZN(
        P1_U3124) );
  AOI22_X1 U23293 ( .A1(n20352), .A2(n20525), .B1(n20524), .B2(n20351), .ZN(
        n20346) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20470), .ZN(n20345) );
  OAI211_X1 U23295 ( .C1(n20473), .C2(n20373), .A(n20346), .B(n20345), .ZN(
        P1_U3125) );
  AOI22_X1 U23296 ( .A1(n20352), .A2(n20531), .B1(n20530), .B2(n20351), .ZN(
        n20348) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20474), .ZN(n20347) );
  OAI211_X1 U23298 ( .C1(n20477), .C2(n20373), .A(n20348), .B(n20347), .ZN(
        P1_U3126) );
  AOI22_X1 U23299 ( .A1(n20352), .A2(n20537), .B1(n20536), .B2(n20351), .ZN(
        n20350) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20478), .ZN(n20349) );
  OAI211_X1 U23301 ( .C1(n20481), .C2(n20373), .A(n20350), .B(n20349), .ZN(
        P1_U3127) );
  AOI22_X1 U23302 ( .A1(n20352), .A2(n20544), .B1(n20542), .B2(n20351), .ZN(
        n20356) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20484), .ZN(n20355) );
  OAI211_X1 U23304 ( .C1(n20489), .C2(n20373), .A(n20356), .B(n20355), .ZN(
        P1_U3128) );
  NAND3_X1 U23305 ( .A1(n20373), .A2(n20418), .A3(n20442), .ZN(n20359) );
  NAND2_X1 U23306 ( .A1(n20359), .A2(n20358), .ZN(n20369) );
  OR2_X1 U23307 ( .A1(n13417), .A2(n20360), .ZN(n20417) );
  NOR2_X1 U23308 ( .A1(n20417), .A2(n9648), .ZN(n20366) );
  INV_X1 U23309 ( .A(n20445), .ZN(n20362) );
  NOR3_X1 U23310 ( .A1(n15558), .A2(n20363), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20421) );
  INV_X1 U23311 ( .A(n20421), .ZN(n20419) );
  NOR2_X1 U23312 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20419), .ZN(
        n20372) );
  INV_X1 U23313 ( .A(n20372), .ZN(n20407) );
  OAI22_X1 U23314 ( .A1(n20442), .A2(n20457), .B1(n20364), .B2(n20407), .ZN(
        n20365) );
  INV_X1 U23315 ( .A(n20365), .ZN(n20375) );
  INV_X1 U23316 ( .A(n20366), .ZN(n20368) );
  AOI22_X1 U23317 ( .A1(n20369), .A2(n20368), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20367), .ZN(n20370) );
  OAI211_X1 U23318 ( .C1(n20372), .C2(n20371), .A(n20452), .B(n20370), .ZN(
        n20411) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20454), .ZN(n20374) );
  OAI211_X1 U23320 ( .C1(n20415), .C2(n20376), .A(n20375), .B(n20374), .ZN(
        P1_U3129) );
  OAI22_X1 U23321 ( .A1(n20442), .A2(n20461), .B1(n20377), .B2(n20407), .ZN(
        n20378) );
  INV_X1 U23322 ( .A(n20378), .ZN(n20380) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20458), .ZN(n20379) );
  OAI211_X1 U23324 ( .C1(n20415), .C2(n20381), .A(n20380), .B(n20379), .ZN(
        P1_U3130) );
  OAI22_X1 U23325 ( .A1(n20442), .A2(n20465), .B1(n20382), .B2(n20407), .ZN(
        n20383) );
  INV_X1 U23326 ( .A(n20383), .ZN(n20385) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20462), .ZN(n20384) );
  OAI211_X1 U23328 ( .C1(n20415), .C2(n20386), .A(n20385), .B(n20384), .ZN(
        P1_U3131) );
  OAI22_X1 U23329 ( .A1(n20442), .A2(n20469), .B1(n20387), .B2(n20407), .ZN(
        n20388) );
  INV_X1 U23330 ( .A(n20388), .ZN(n20390) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20466), .ZN(n20389) );
  OAI211_X1 U23332 ( .C1(n20415), .C2(n20391), .A(n20390), .B(n20389), .ZN(
        P1_U3132) );
  OAI22_X1 U23333 ( .A1(n20442), .A2(n20473), .B1(n20392), .B2(n20407), .ZN(
        n20393) );
  INV_X1 U23334 ( .A(n20393), .ZN(n20395) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20470), .ZN(n20394) );
  OAI211_X1 U23336 ( .C1(n20415), .C2(n20396), .A(n20395), .B(n20394), .ZN(
        P1_U3133) );
  OAI22_X1 U23337 ( .A1(n20442), .A2(n20477), .B1(n20397), .B2(n20407), .ZN(
        n20398) );
  INV_X1 U23338 ( .A(n20398), .ZN(n20400) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20474), .ZN(n20399) );
  OAI211_X1 U23340 ( .C1(n20415), .C2(n20401), .A(n20400), .B(n20399), .ZN(
        P1_U3134) );
  OAI22_X1 U23341 ( .A1(n20442), .A2(n20481), .B1(n20402), .B2(n20407), .ZN(
        n20403) );
  INV_X1 U23342 ( .A(n20403), .ZN(n20405) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20478), .ZN(n20404) );
  OAI211_X1 U23344 ( .C1(n20415), .C2(n20406), .A(n20405), .B(n20404), .ZN(
        P1_U3135) );
  OAI22_X1 U23345 ( .A1(n20442), .A2(n20489), .B1(n20408), .B2(n20407), .ZN(
        n20409) );
  INV_X1 U23346 ( .A(n20409), .ZN(n20413) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20411), .B1(
        n20410), .B2(n20484), .ZN(n20412) );
  OAI211_X1 U23348 ( .C1(n20415), .C2(n20414), .A(n20413), .B(n20412), .ZN(
        P1_U3136) );
  NOR2_X1 U23349 ( .A1(n20416), .A2(n20419), .ZN(n20437) );
  INV_X1 U23350 ( .A(n20437), .ZN(n20420) );
  INV_X1 U23351 ( .A(n20417), .ZN(n20449) );
  NAND2_X1 U23352 ( .A1(n20449), .A2(n20418), .ZN(n20490) );
  OAI222_X1 U23353 ( .A1(n20420), .A2(n20493), .B1(n20640), .B2(n20419), .C1(
        n20009), .C2(n20490), .ZN(n20438) );
  AOI22_X1 U23354 ( .A1(n20438), .A2(n20496), .B1(n20495), .B2(n20437), .ZN(
        n20424) );
  NOR2_X1 U23355 ( .A1(n20444), .A2(n20493), .ZN(n20498) );
  OAI221_X1 U23356 ( .B1(n20421), .B2(P1_STATEBS16_REG_SCAN_IN), .C1(n20421), 
        .C2(n20498), .A(n20499), .ZN(n20439) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20439), .B1(
        n20485), .B2(n20502), .ZN(n20423) );
  OAI211_X1 U23358 ( .C1(n20505), .C2(n20442), .A(n20424), .B(n20423), .ZN(
        P1_U3137) );
  AOI22_X1 U23359 ( .A1(n20438), .A2(n20507), .B1(n20506), .B2(n20437), .ZN(
        n20426) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20439), .B1(
        n20485), .B2(n20508), .ZN(n20425) );
  OAI211_X1 U23361 ( .C1(n20511), .C2(n20442), .A(n20426), .B(n20425), .ZN(
        P1_U3138) );
  AOI22_X1 U23362 ( .A1(n20438), .A2(n20513), .B1(n20512), .B2(n20437), .ZN(
        n20428) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20439), .B1(
        n20485), .B2(n20514), .ZN(n20427) );
  OAI211_X1 U23364 ( .C1(n20517), .C2(n20442), .A(n20428), .B(n20427), .ZN(
        P1_U3139) );
  AOI22_X1 U23365 ( .A1(n20438), .A2(n20519), .B1(n20518), .B2(n20437), .ZN(
        n20430) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20439), .B1(
        n20485), .B2(n20520), .ZN(n20429) );
  OAI211_X1 U23367 ( .C1(n20523), .C2(n20442), .A(n20430), .B(n20429), .ZN(
        P1_U3140) );
  AOI22_X1 U23368 ( .A1(n20438), .A2(n20525), .B1(n20524), .B2(n20437), .ZN(
        n20432) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20439), .B1(
        n20485), .B2(n20526), .ZN(n20431) );
  OAI211_X1 U23370 ( .C1(n20529), .C2(n20442), .A(n20432), .B(n20431), .ZN(
        P1_U3141) );
  AOI22_X1 U23371 ( .A1(n20438), .A2(n20531), .B1(n20530), .B2(n20437), .ZN(
        n20434) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20439), .B1(
        n20485), .B2(n20532), .ZN(n20433) );
  OAI211_X1 U23373 ( .C1(n20535), .C2(n20442), .A(n20434), .B(n20433), .ZN(
        P1_U3142) );
  AOI22_X1 U23374 ( .A1(n20438), .A2(n20537), .B1(n20536), .B2(n20437), .ZN(
        n20436) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20439), .B1(
        n20485), .B2(n20538), .ZN(n20435) );
  OAI211_X1 U23376 ( .C1(n20541), .C2(n20442), .A(n20436), .B(n20435), .ZN(
        P1_U3143) );
  AOI22_X1 U23377 ( .A1(n20438), .A2(n20544), .B1(n20542), .B2(n20437), .ZN(
        n20441) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20439), .B1(
        n20485), .B2(n20546), .ZN(n20440) );
  OAI211_X1 U23379 ( .C1(n20552), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P1_U3144) );
  INV_X1 U23380 ( .A(n20500), .ZN(n20492) );
  NOR2_X1 U23381 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20492), .ZN(
        n20483) );
  OAI22_X1 U23382 ( .A1(n20490), .A2(n13694), .B1(n20446), .B2(n20445), .ZN(
        n20482) );
  AOI22_X1 U23383 ( .A1(n20495), .A2(n20483), .B1(n20482), .B2(n20496), .ZN(
        n20456) );
  INV_X1 U23384 ( .A(n20485), .ZN(n20447) );
  AOI21_X1 U23385 ( .B1(n20447), .B2(n20551), .A(n20641), .ZN(n20448) );
  AOI21_X1 U23386 ( .B1(n20449), .B2(n9648), .A(n20448), .ZN(n20450) );
  NOR2_X1 U23387 ( .A1(n20450), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20453) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20486), .B1(
        n20485), .B2(n20454), .ZN(n20455) );
  OAI211_X1 U23389 ( .C1(n20457), .C2(n20551), .A(n20456), .B(n20455), .ZN(
        P1_U3145) );
  AOI22_X1 U23390 ( .A1(n20506), .A2(n20483), .B1(n20482), .B2(n20507), .ZN(
        n20460) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20486), .B1(
        n20485), .B2(n20458), .ZN(n20459) );
  OAI211_X1 U23392 ( .C1(n20461), .C2(n20551), .A(n20460), .B(n20459), .ZN(
        P1_U3146) );
  AOI22_X1 U23393 ( .A1(n20512), .A2(n20483), .B1(n20482), .B2(n20513), .ZN(
        n20464) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20486), .B1(
        n20485), .B2(n20462), .ZN(n20463) );
  OAI211_X1 U23395 ( .C1(n20465), .C2(n20551), .A(n20464), .B(n20463), .ZN(
        P1_U3147) );
  AOI22_X1 U23396 ( .A1(n20518), .A2(n20483), .B1(n20482), .B2(n20519), .ZN(
        n20468) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20486), .B1(
        n20485), .B2(n20466), .ZN(n20467) );
  OAI211_X1 U23398 ( .C1(n20469), .C2(n20551), .A(n20468), .B(n20467), .ZN(
        P1_U3148) );
  AOI22_X1 U23399 ( .A1(n20524), .A2(n20483), .B1(n20482), .B2(n20525), .ZN(
        n20472) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20486), .B1(
        n20485), .B2(n20470), .ZN(n20471) );
  OAI211_X1 U23401 ( .C1(n20473), .C2(n20551), .A(n20472), .B(n20471), .ZN(
        P1_U3149) );
  AOI22_X1 U23402 ( .A1(n20530), .A2(n20483), .B1(n20482), .B2(n20531), .ZN(
        n20476) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20486), .B1(
        n20485), .B2(n20474), .ZN(n20475) );
  OAI211_X1 U23404 ( .C1(n20477), .C2(n20551), .A(n20476), .B(n20475), .ZN(
        P1_U3150) );
  AOI22_X1 U23405 ( .A1(n20536), .A2(n20483), .B1(n20482), .B2(n20537), .ZN(
        n20480) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20486), .B1(
        n20485), .B2(n20478), .ZN(n20479) );
  OAI211_X1 U23407 ( .C1(n20481), .C2(n20551), .A(n20480), .B(n20479), .ZN(
        P1_U3151) );
  AOI22_X1 U23408 ( .A1(n20542), .A2(n20483), .B1(n20544), .B2(n20482), .ZN(
        n20488) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20486), .B1(
        n20485), .B2(n20484), .ZN(n20487) );
  OAI211_X1 U23410 ( .C1(n20489), .C2(n20551), .A(n20488), .B(n20487), .ZN(
        P1_U3152) );
  OAI222_X1 U23411 ( .A1(n20493), .A2(n20494), .B1(n20640), .B2(n20492), .C1(
        n20491), .C2(n20490), .ZN(n20545) );
  INV_X1 U23412 ( .A(n20494), .ZN(n20543) );
  AOI22_X1 U23413 ( .A1(n20545), .A2(n20496), .B1(n20543), .B2(n20495), .ZN(
        n20504) );
  AND2_X1 U23414 ( .A1(n20498), .A2(n20497), .ZN(n20501) );
  OAI21_X1 U23415 ( .B1(n20501), .B2(n20500), .A(n20499), .ZN(n20548) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20502), .ZN(n20503) );
  OAI211_X1 U23417 ( .C1(n20505), .C2(n20551), .A(n20504), .B(n20503), .ZN(
        P1_U3153) );
  AOI22_X1 U23418 ( .A1(n20545), .A2(n20507), .B1(n20543), .B2(n20506), .ZN(
        n20510) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20508), .ZN(n20509) );
  OAI211_X1 U23420 ( .C1(n20511), .C2(n20551), .A(n20510), .B(n20509), .ZN(
        P1_U3154) );
  AOI22_X1 U23421 ( .A1(n20545), .A2(n20513), .B1(n20543), .B2(n20512), .ZN(
        n20516) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20514), .ZN(n20515) );
  OAI211_X1 U23423 ( .C1(n20517), .C2(n20551), .A(n20516), .B(n20515), .ZN(
        P1_U3155) );
  AOI22_X1 U23424 ( .A1(n20545), .A2(n20519), .B1(n20543), .B2(n20518), .ZN(
        n20522) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20520), .ZN(n20521) );
  OAI211_X1 U23426 ( .C1(n20523), .C2(n20551), .A(n20522), .B(n20521), .ZN(
        P1_U3156) );
  AOI22_X1 U23427 ( .A1(n20545), .A2(n20525), .B1(n20543), .B2(n20524), .ZN(
        n20528) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20526), .ZN(n20527) );
  OAI211_X1 U23429 ( .C1(n20529), .C2(n20551), .A(n20528), .B(n20527), .ZN(
        P1_U3157) );
  AOI22_X1 U23430 ( .A1(n20545), .A2(n20531), .B1(n20543), .B2(n20530), .ZN(
        n20534) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20532), .ZN(n20533) );
  OAI211_X1 U23432 ( .C1(n20535), .C2(n20551), .A(n20534), .B(n20533), .ZN(
        P1_U3158) );
  AOI22_X1 U23433 ( .A1(n20545), .A2(n20537), .B1(n20543), .B2(n20536), .ZN(
        n20540) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20538), .ZN(n20539) );
  OAI211_X1 U23435 ( .C1(n20541), .C2(n20551), .A(n20540), .B(n20539), .ZN(
        P1_U3159) );
  AOI22_X1 U23436 ( .A1(n20545), .A2(n20544), .B1(n20543), .B2(n20542), .ZN(
        n20550) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20548), .B1(
        n20547), .B2(n20546), .ZN(n20549) );
  OAI211_X1 U23438 ( .C1(n20552), .C2(n20551), .A(n20550), .B(n20549), .ZN(
        P1_U3160) );
  NOR2_X1 U23439 ( .A1(n20790), .A2(n20553), .ZN(n20555) );
  OAI21_X1 U23440 ( .B1(n20555), .B2(n20640), .A(n20554), .ZN(P1_U3163) );
  AND2_X1 U23441 ( .A1(n20556), .A2(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(
        P1_U3164) );
  AND2_X1 U23442 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20556), .ZN(
        P1_U3165) );
  AND2_X1 U23443 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20556), .ZN(
        P1_U3166) );
  AND2_X1 U23444 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20556), .ZN(
        P1_U3167) );
  AND2_X1 U23445 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20556), .ZN(
        P1_U3168) );
  AND2_X1 U23446 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20556), .ZN(
        P1_U3169) );
  AND2_X1 U23447 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20556), .ZN(
        P1_U3170) );
  AND2_X1 U23448 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20556), .ZN(
        P1_U3171) );
  AND2_X1 U23449 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20556), .ZN(
        P1_U3172) );
  AND2_X1 U23450 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20556), .ZN(
        P1_U3173) );
  AND2_X1 U23451 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20556), .ZN(
        P1_U3174) );
  AND2_X1 U23452 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20556), .ZN(
        P1_U3175) );
  AND2_X1 U23453 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20556), .ZN(
        P1_U3176) );
  AND2_X1 U23454 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20556), .ZN(
        P1_U3177) );
  AND2_X1 U23455 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20556), .ZN(
        P1_U3178) );
  AND2_X1 U23456 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20556), .ZN(
        P1_U3179) );
  AND2_X1 U23457 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20556), .ZN(
        P1_U3180) );
  AND2_X1 U23458 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20556), .ZN(
        P1_U3181) );
  AND2_X1 U23459 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20556), .ZN(
        P1_U3182) );
  AND2_X1 U23460 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20556), .ZN(
        P1_U3183) );
  AND2_X1 U23461 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20556), .ZN(
        P1_U3184) );
  AND2_X1 U23462 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20556), .ZN(
        P1_U3185) );
  AND2_X1 U23463 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20556), .ZN(P1_U3186) );
  AND2_X1 U23464 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20556), .ZN(P1_U3187) );
  AND2_X1 U23465 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20556), .ZN(P1_U3188) );
  AND2_X1 U23466 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20556), .ZN(P1_U3189) );
  AND2_X1 U23467 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20556), .ZN(P1_U3190) );
  AND2_X1 U23468 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20556), .ZN(P1_U3191) );
  AND2_X1 U23469 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20556), .ZN(P1_U3192) );
  AND2_X1 U23470 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20556), .ZN(P1_U3193) );
  NOR2_X1 U23471 ( .A1(n20564), .A2(n20570), .ZN(n20561) );
  INV_X1 U23472 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20573) );
  NAND2_X1 U23473 ( .A1(n20562), .A2(n20573), .ZN(n20559) );
  INV_X1 U23474 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20568) );
  NOR2_X1 U23475 ( .A1(n20568), .A2(NA), .ZN(n20565) );
  INV_X1 U23476 ( .A(n20565), .ZN(n20557) );
  AOI22_X1 U23477 ( .A1(HOLD), .A2(n20559), .B1(n20558), .B2(n20557), .ZN(
        n20560) );
  OAI22_X1 U23478 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20561), .B1(n20637), 
        .B2(n20560), .ZN(P1_U3194) );
  AOI21_X1 U23479 ( .B1(NA), .B2(n20562), .A(P1_STATE_REG_0__SCAN_IN), .ZN(
        n20563) );
  OAI22_X1 U23480 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20565), .B1(n20564), 
        .B2(n20563), .ZN(n20571) );
  OAI21_X1 U23481 ( .B1(NA), .B2(n20647), .A(n20566), .ZN(n20567) );
  OAI211_X1 U23482 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20568), .A(HOLD), .B(
        n20567), .ZN(n20569) );
  OAI22_X1 U23483 ( .A1(n20572), .A2(n20571), .B1(n20570), .B2(n20569), .ZN(
        P1_U3196) );
  INV_X1 U23484 ( .A(n20603), .ZN(n20611) );
  NOR2_X1 U23485 ( .A1(n20573), .A2(n20650), .ZN(n20612) );
  INV_X1 U23486 ( .A(n20612), .ZN(n20606) );
  AOI222_X1 U23487 ( .A1(n20611), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20609), .ZN(n20574) );
  INV_X1 U23488 ( .A(n20574), .ZN(P1_U3197) );
  AOI222_X1 U23489 ( .A1(n20609), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20611), .ZN(n20575) );
  INV_X1 U23490 ( .A(n20575), .ZN(P1_U3198) );
  OAI222_X1 U23491 ( .A1(n20606), .A2(n20577), .B1(n20576), .B2(n20637), .C1(
        n20579), .C2(n20603), .ZN(P1_U3199) );
  AOI22_X1 U23492 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20650), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20611), .ZN(n20578) );
  OAI21_X1 U23493 ( .B1(n20579), .B2(n20606), .A(n20578), .ZN(P1_U3200) );
  AOI22_X1 U23494 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20650), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20612), .ZN(n20580) );
  OAI21_X1 U23495 ( .B1(n20581), .B2(n20603), .A(n20580), .ZN(P1_U3201) );
  AOI222_X1 U23496 ( .A1(n20609), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20611), .ZN(n20582) );
  INV_X1 U23497 ( .A(n20582), .ZN(P1_U3202) );
  AOI222_X1 U23498 ( .A1(n20609), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20611), .ZN(n20583) );
  INV_X1 U23499 ( .A(n20583), .ZN(P1_U3203) );
  AOI222_X1 U23500 ( .A1(n20611), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20609), .ZN(n20584) );
  INV_X1 U23501 ( .A(n20584), .ZN(P1_U3204) );
  AOI222_X1 U23502 ( .A1(n20609), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20611), .ZN(n20585) );
  INV_X1 U23503 ( .A(n20585), .ZN(P1_U3205) );
  AOI22_X1 U23504 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20650), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20611), .ZN(n20586) );
  OAI21_X1 U23505 ( .B1(n14651), .B2(n20606), .A(n20586), .ZN(P1_U3206) );
  INV_X1 U23506 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20588) );
  AOI22_X1 U23507 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20650), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20611), .ZN(n20587) );
  OAI21_X1 U23508 ( .B1(n20588), .B2(n20606), .A(n20587), .ZN(P1_U3207) );
  AOI22_X1 U23509 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20650), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20609), .ZN(n20589) );
  OAI21_X1 U23510 ( .B1(n14642), .B2(n20603), .A(n20589), .ZN(P1_U3208) );
  AOI222_X1 U23511 ( .A1(n20609), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20611), .ZN(n20590) );
  INV_X1 U23512 ( .A(n20590), .ZN(P1_U3209) );
  AOI222_X1 U23513 ( .A1(n20611), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20609), .ZN(n20591) );
  INV_X1 U23514 ( .A(n20591), .ZN(P1_U3210) );
  AOI222_X1 U23515 ( .A1(n20609), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20611), .ZN(n20592) );
  INV_X1 U23516 ( .A(n20592), .ZN(P1_U3211) );
  AOI222_X1 U23517 ( .A1(n20612), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20611), .ZN(n20593) );
  INV_X1 U23518 ( .A(n20593), .ZN(P1_U3212) );
  AOI22_X1 U23519 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20650), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20611), .ZN(n20594) );
  OAI21_X1 U23520 ( .B1(n15778), .B2(n20606), .A(n20594), .ZN(P1_U3213) );
  AOI22_X1 U23521 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20650), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20609), .ZN(n20595) );
  OAI21_X1 U23522 ( .B1(n20722), .B2(n20603), .A(n20595), .ZN(P1_U3214) );
  AOI222_X1 U23523 ( .A1(n20611), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20609), .ZN(n20596) );
  INV_X1 U23524 ( .A(n20596), .ZN(P1_U3215) );
  AOI222_X1 U23525 ( .A1(n20612), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20611), .ZN(n20597) );
  INV_X1 U23526 ( .A(n20597), .ZN(P1_U3216) );
  AOI222_X1 U23527 ( .A1(n20612), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20611), .ZN(n20598) );
  INV_X1 U23528 ( .A(n20598), .ZN(P1_U3217) );
  AOI222_X1 U23529 ( .A1(n20611), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20609), .ZN(n20599) );
  INV_X1 U23530 ( .A(n20599), .ZN(P1_U3218) );
  AOI222_X1 U23531 ( .A1(n20612), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20611), .ZN(n20600) );
  INV_X1 U23532 ( .A(n20600), .ZN(P1_U3219) );
  AOI222_X1 U23533 ( .A1(n20612), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20611), .ZN(n20601) );
  INV_X1 U23534 ( .A(n20601), .ZN(P1_U3220) );
  AOI222_X1 U23535 ( .A1(n20612), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20611), .ZN(n20602) );
  INV_X1 U23536 ( .A(n20602), .ZN(P1_U3221) );
  INV_X1 U23537 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20605) );
  INV_X1 U23538 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20705) );
  OAI222_X1 U23539 ( .A1(n20606), .A2(n20605), .B1(n20705), .B2(n20637), .C1(
        n20604), .C2(n20603), .ZN(P1_U3222) );
  AOI222_X1 U23540 ( .A1(n20609), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20611), .ZN(n20607) );
  INV_X1 U23541 ( .A(n20607), .ZN(P1_U3223) );
  AOI222_X1 U23542 ( .A1(n20609), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20611), .ZN(n20608) );
  INV_X1 U23543 ( .A(n20608), .ZN(P1_U3224) );
  AOI222_X1 U23544 ( .A1(n20611), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20609), .ZN(n20610) );
  INV_X1 U23545 ( .A(n20610), .ZN(P1_U3225) );
  AOI222_X1 U23546 ( .A1(n20612), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20650), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20611), .ZN(n20613) );
  INV_X1 U23547 ( .A(n20613), .ZN(P1_U3226) );
  OAI22_X1 U23548 ( .A1(n20650), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20637), .ZN(n20614) );
  INV_X1 U23549 ( .A(n20614), .ZN(P1_U3458) );
  OAI22_X1 U23550 ( .A1(n20650), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20637), .ZN(n20615) );
  INV_X1 U23551 ( .A(n20615), .ZN(P1_U3459) );
  OAI22_X1 U23552 ( .A1(n20650), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20637), .ZN(n20616) );
  INV_X1 U23553 ( .A(n20616), .ZN(P1_U3460) );
  OAI22_X1 U23554 ( .A1(n20650), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20637), .ZN(n20617) );
  INV_X1 U23555 ( .A(n20617), .ZN(P1_U3461) );
  OAI21_X1 U23556 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20621), .A(n20619), 
        .ZN(n20618) );
  INV_X1 U23557 ( .A(n20618), .ZN(P1_U3464) );
  OAI21_X1 U23558 ( .B1(n20621), .B2(n20620), .A(n20619), .ZN(P1_U3465) );
  INV_X1 U23559 ( .A(n20622), .ZN(n20626) );
  OAI22_X1 U23560 ( .A1(n20626), .A2(n20625), .B1(n20624), .B2(n20623), .ZN(
        n20628) );
  MUX2_X1 U23561 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20628), .S(
        n20627), .Z(P1_U3469) );
  AOI21_X1 U23562 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20629) );
  AOI22_X1 U23563 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20629), .B2(n13878), .ZN(n20632) );
  INV_X1 U23564 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20631) );
  AOI22_X1 U23565 ( .A1(n20635), .A2(n20632), .B1(n20631), .B2(n20630), .ZN(
        P1_U3481) );
  INV_X1 U23566 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20634) );
  OAI21_X1 U23567 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20635), .ZN(n20633) );
  OAI21_X1 U23568 ( .B1(n20635), .B2(n20634), .A(n20633), .ZN(P1_U3482) );
  AOI22_X1 U23569 ( .A1(n20637), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20636), 
        .B2(n20650), .ZN(P1_U3483) );
  INV_X1 U23570 ( .A(n20638), .ZN(n20639) );
  AOI211_X1 U23571 ( .C1(n20642), .C2(n20641), .A(n20640), .B(n20639), .ZN(
        n20644) );
  OAI21_X1 U23572 ( .B1(n20644), .B2(n20790), .A(n20643), .ZN(n20649) );
  AOI211_X1 U23573 ( .C1(n19873), .C2(n20647), .A(n20646), .B(n20645), .ZN(
        n20648) );
  MUX2_X1 U23574 ( .A(n20649), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20648), 
        .Z(P1_U3485) );
  MUX2_X1 U23575 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20650), .Z(P1_U3486) );
  NOR2_X1 U23576 ( .A1(keyinput29), .A2(keyinput47), .ZN(n20651) );
  NAND3_X1 U23577 ( .A1(keyinput50), .A2(keyinput22), .A3(n20651), .ZN(n20656)
         );
  NAND3_X1 U23578 ( .A1(keyinput11), .A2(keyinput55), .A3(keyinput60), .ZN(
        n20655) );
  NOR3_X1 U23579 ( .A1(keyinput41), .A2(keyinput35), .A3(keyinput6), .ZN(
        n20653) );
  NOR3_X1 U23580 ( .A1(keyinput9), .A2(keyinput24), .A3(keyinput23), .ZN(
        n20652) );
  NAND4_X1 U23581 ( .A1(keyinput34), .A2(n20653), .A3(keyinput49), .A4(n20652), 
        .ZN(n20654) );
  NOR4_X1 U23582 ( .A1(keyinput44), .A2(n20656), .A3(n20655), .A4(n20654), 
        .ZN(n20805) );
  NOR3_X1 U23583 ( .A1(keyinput18), .A2(keyinput54), .A3(keyinput53), .ZN(
        n20661) );
  INV_X1 U23584 ( .A(keyinput32), .ZN(n20727) );
  NOR4_X1 U23585 ( .A1(keyinput31), .A2(keyinput28), .A3(keyinput63), .A4(
        n20727), .ZN(n20660) );
  NAND4_X1 U23586 ( .A1(keyinput62), .A2(keyinput27), .A3(keyinput13), .A4(
        keyinput16), .ZN(n20658) );
  NAND2_X1 U23587 ( .A1(keyinput43), .A2(keyinput40), .ZN(n20657) );
  NOR4_X1 U23588 ( .A1(keyinput14), .A2(keyinput8), .A3(n20658), .A4(n20657), 
        .ZN(n20659) );
  NAND4_X1 U23589 ( .A1(keyinput51), .A2(n20661), .A3(n20660), .A4(n20659), 
        .ZN(n20672) );
  NOR4_X1 U23590 ( .A1(keyinput1), .A2(keyinput5), .A3(keyinput17), .A4(
        keyinput37), .ZN(n20665) );
  NOR4_X1 U23591 ( .A1(keyinput57), .A2(keyinput12), .A3(keyinput4), .A4(
        keyinput20), .ZN(n20664) );
  NOR4_X1 U23592 ( .A1(keyinput36), .A2(keyinput48), .A3(keyinput56), .A4(
        keyinput0), .ZN(n20663) );
  NOR4_X1 U23593 ( .A1(keyinput39), .A2(keyinput58), .A3(keyinput59), .A4(
        keyinput15), .ZN(n20662) );
  NAND4_X1 U23594 ( .A1(n20665), .A2(n20664), .A3(n20663), .A4(n20662), .ZN(
        n20671) );
  NAND4_X1 U23595 ( .A1(keyinput45), .A2(keyinput33), .A3(keyinput61), .A4(
        keyinput52), .ZN(n20670) );
  NAND3_X1 U23596 ( .A1(keyinput7), .A2(keyinput25), .A3(keyinput21), .ZN(
        n20668) );
  NAND4_X1 U23597 ( .A1(keyinput42), .A2(keyinput46), .A3(keyinput38), .A4(
        keyinput2), .ZN(n20667) );
  NAND4_X1 U23598 ( .A1(keyinput10), .A2(keyinput30), .A3(keyinput26), .A4(
        keyinput19), .ZN(n20666) );
  OR4_X1 U23599 ( .A1(keyinput3), .A2(n20668), .A3(n20667), .A4(n20666), .ZN(
        n20669) );
  NOR4_X1 U23600 ( .A1(n20672), .A2(n20671), .A3(n20670), .A4(n20669), .ZN(
        n20804) );
  INV_X1 U23601 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n20675) );
  INV_X1 U23602 ( .A(keyinput41), .ZN(n20674) );
  AOI22_X1 U23603 ( .A1(n20675), .A2(keyinput34), .B1(P3_M_IO_N_REG_SCAN_IN), 
        .B2(n20674), .ZN(n20673) );
  OAI221_X1 U23604 ( .B1(n20675), .B2(keyinput34), .C1(n20674), .C2(
        P3_M_IO_N_REG_SCAN_IN), .A(n20673), .ZN(n20688) );
  INV_X1 U23605 ( .A(keyinput35), .ZN(n20677) );
  AOI22_X1 U23606 ( .A1(n20678), .A2(keyinput6), .B1(
        P3_DATAWIDTH_REG_28__SCAN_IN), .B2(n20677), .ZN(n20676) );
  OAI221_X1 U23607 ( .B1(n20678), .B2(keyinput6), .C1(n20677), .C2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A(n20676), .ZN(n20687) );
  INV_X1 U23608 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20680) );
  AOI22_X1 U23609 ( .A1(n20681), .A2(keyinput29), .B1(n20680), .B2(keyinput50), 
        .ZN(n20679) );
  OAI221_X1 U23610 ( .B1(n20681), .B2(keyinput29), .C1(n20680), .C2(keyinput50), .A(n20679), .ZN(n20686) );
  AOI22_X1 U23611 ( .A1(n20684), .A2(keyinput22), .B1(n20683), .B2(keyinput47), 
        .ZN(n20682) );
  OAI221_X1 U23612 ( .B1(n20684), .B2(keyinput22), .C1(n20683), .C2(keyinput47), .A(n20682), .ZN(n20685) );
  NOR4_X1 U23613 ( .A1(n20688), .A2(n20687), .A3(n20686), .A4(n20685), .ZN(
        n20739) );
  AOI22_X1 U23614 ( .A1(n20691), .A2(keyinput9), .B1(keyinput49), .B2(n20690), 
        .ZN(n20689) );
  OAI221_X1 U23615 ( .B1(n20691), .B2(keyinput9), .C1(n20690), .C2(keyinput49), 
        .A(n20689), .ZN(n20703) );
  INV_X1 U23616 ( .A(DATAI_19_), .ZN(n20694) );
  INV_X1 U23617 ( .A(keyinput24), .ZN(n20693) );
  AOI22_X1 U23618 ( .A1(n20694), .A2(keyinput23), .B1(
        P2_DATAWIDTH_REG_3__SCAN_IN), .B2(n20693), .ZN(n20692) );
  OAI221_X1 U23619 ( .B1(n20694), .B2(keyinput23), .C1(n20693), .C2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A(n20692), .ZN(n20702) );
  AOI22_X1 U23620 ( .A1(n20697), .A2(keyinput11), .B1(keyinput44), .B2(n20696), 
        .ZN(n20695) );
  OAI221_X1 U23621 ( .B1(n20697), .B2(keyinput11), .C1(n20696), .C2(keyinput44), .A(n20695), .ZN(n20701) );
  AOI22_X1 U23622 ( .A1(n20699), .A2(keyinput55), .B1(keyinput60), .B2(n11876), 
        .ZN(n20698) );
  OAI221_X1 U23623 ( .B1(n20699), .B2(keyinput55), .C1(n11876), .C2(keyinput60), .A(n20698), .ZN(n20700) );
  NOR4_X1 U23624 ( .A1(n20703), .A2(n20702), .A3(n20701), .A4(n20700), .ZN(
        n20738) );
  INV_X1 U23625 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n20706) );
  AOI22_X1 U23626 ( .A1(n20706), .A2(keyinput18), .B1(keyinput54), .B2(n20705), 
        .ZN(n20704) );
  OAI221_X1 U23627 ( .B1(n20706), .B2(keyinput18), .C1(n20705), .C2(keyinput54), .A(n20704), .ZN(n20719) );
  INV_X1 U23628 ( .A(P3_UWORD_REG_12__SCAN_IN), .ZN(n20709) );
  INV_X1 U23629 ( .A(keyinput51), .ZN(n20708) );
  AOI22_X1 U23630 ( .A1(n20709), .A2(keyinput53), .B1(
        P3_DATAWIDTH_REG_9__SCAN_IN), .B2(n20708), .ZN(n20707) );
  OAI221_X1 U23631 ( .B1(n20709), .B2(keyinput53), .C1(n20708), .C2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A(n20707), .ZN(n20718) );
  INV_X1 U23632 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n20712) );
  INV_X1 U23633 ( .A(P1_LWORD_REG_11__SCAN_IN), .ZN(n20711) );
  AOI22_X1 U23634 ( .A1(n20712), .A2(keyinput62), .B1(keyinput27), .B2(n20711), 
        .ZN(n20710) );
  OAI221_X1 U23635 ( .B1(n20712), .B2(keyinput62), .C1(n20711), .C2(keyinput27), .A(n20710), .ZN(n20717) );
  INV_X1 U23636 ( .A(keyinput16), .ZN(n20714) );
  AOI22_X1 U23637 ( .A1(n20715), .A2(keyinput13), .B1(
        P2_DATAWIDTH_REG_11__SCAN_IN), .B2(n20714), .ZN(n20713) );
  OAI221_X1 U23638 ( .B1(n20715), .B2(keyinput13), .C1(n20714), .C2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A(n20713), .ZN(n20716) );
  NOR4_X1 U23639 ( .A1(n20719), .A2(n20718), .A3(n20717), .A4(n20716), .ZN(
        n20737) );
  INV_X1 U23640 ( .A(keyinput8), .ZN(n20721) );
  AOI22_X1 U23641 ( .A1(n20722), .A2(keyinput14), .B1(
        P2_DATAWIDTH_REG_15__SCAN_IN), .B2(n20721), .ZN(n20720) );
  OAI221_X1 U23642 ( .B1(n20722), .B2(keyinput14), .C1(n20721), .C2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A(n20720), .ZN(n20735) );
  INV_X1 U23643 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20725) );
  AOI22_X1 U23644 ( .A1(n20725), .A2(keyinput43), .B1(keyinput40), .B2(n20724), 
        .ZN(n20723) );
  OAI221_X1 U23645 ( .B1(n20725), .B2(keyinput43), .C1(n20724), .C2(keyinput40), .A(n20723), .ZN(n20734) );
  INV_X1 U23646 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n20728) );
  AOI22_X1 U23647 ( .A1(n20728), .A2(keyinput28), .B1(
        P1_DATAWIDTH_REG_31__SCAN_IN), .B2(n20727), .ZN(n20726) );
  OAI221_X1 U23648 ( .B1(n20728), .B2(keyinput28), .C1(n20727), .C2(
        P1_DATAWIDTH_REG_31__SCAN_IN), .A(n20726), .ZN(n20733) );
  INV_X1 U23649 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20731) );
  INV_X1 U23650 ( .A(keyinput63), .ZN(n20730) );
  AOI22_X1 U23651 ( .A1(n20731), .A2(keyinput31), .B1(
        P3_DATAWIDTH_REG_3__SCAN_IN), .B2(n20730), .ZN(n20729) );
  OAI221_X1 U23652 ( .B1(n20731), .B2(keyinput31), .C1(n20730), .C2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A(n20729), .ZN(n20732) );
  NOR4_X1 U23653 ( .A1(n20735), .A2(n20734), .A3(n20733), .A4(n20732), .ZN(
        n20736) );
  NAND4_X1 U23654 ( .A1(n20739), .A2(n20738), .A3(n20737), .A4(n20736), .ZN(
        n20803) );
  INV_X1 U23655 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20741) );
  AOI22_X1 U23656 ( .A1(n20741), .A2(keyinput1), .B1(n12799), .B2(keyinput37), 
        .ZN(n20740) );
  OAI221_X1 U23657 ( .B1(n20741), .B2(keyinput1), .C1(n12799), .C2(keyinput37), 
        .A(n20740), .ZN(n20753) );
  AOI22_X1 U23658 ( .A1(n20744), .A2(keyinput38), .B1(keyinput26), .B2(n20743), 
        .ZN(n20742) );
  OAI221_X1 U23659 ( .B1(n20744), .B2(keyinput38), .C1(n20743), .C2(keyinput26), .A(n20742), .ZN(n20752) );
  INV_X1 U23660 ( .A(keyinput39), .ZN(n20746) );
  AOI22_X1 U23661 ( .A1(n20747), .A2(keyinput48), .B1(
        P3_BYTEENABLE_REG_1__SCAN_IN), .B2(n20746), .ZN(n20745) );
  OAI221_X1 U23662 ( .B1(n20747), .B2(keyinput48), .C1(n20746), .C2(
        P3_BYTEENABLE_REG_1__SCAN_IN), .A(n20745), .ZN(n20751) );
  AOI22_X1 U23663 ( .A1(n20749), .A2(keyinput56), .B1(n12853), .B2(keyinput59), 
        .ZN(n20748) );
  OAI221_X1 U23664 ( .B1(n20749), .B2(keyinput56), .C1(n12853), .C2(keyinput59), .A(n20748), .ZN(n20750) );
  NOR4_X1 U23665 ( .A1(n20753), .A2(n20752), .A3(n20751), .A4(n20750), .ZN(
        n20801) );
  AOI22_X1 U23666 ( .A1(n20756), .A2(keyinput7), .B1(keyinput25), .B2(n20755), 
        .ZN(n20754) );
  OAI221_X1 U23667 ( .B1(n20756), .B2(keyinput7), .C1(n20755), .C2(keyinput25), 
        .A(n20754), .ZN(n20768) );
  INV_X1 U23668 ( .A(keyinput2), .ZN(n20758) );
  AOI22_X1 U23669 ( .A1(n20759), .A2(keyinput58), .B1(P2_BE_N_REG_3__SCAN_IN), 
        .B2(n20758), .ZN(n20757) );
  OAI221_X1 U23670 ( .B1(n20759), .B2(keyinput58), .C1(n20758), .C2(
        P2_BE_N_REG_3__SCAN_IN), .A(n20757), .ZN(n20767) );
  INV_X1 U23671 ( .A(P3_LWORD_REG_1__SCAN_IN), .ZN(n20761) );
  AOI22_X1 U23672 ( .A1(n20762), .A2(keyinput33), .B1(keyinput19), .B2(n20761), 
        .ZN(n20760) );
  OAI221_X1 U23673 ( .B1(n20762), .B2(keyinput33), .C1(n20761), .C2(keyinput19), .A(n20760), .ZN(n20766) );
  INV_X1 U23674 ( .A(keyinput15), .ZN(n20764) );
  AOI22_X1 U23675 ( .A1(n10204), .A2(keyinput52), .B1(
        P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20764), .ZN(n20763) );
  OAI221_X1 U23676 ( .B1(n10204), .B2(keyinput52), .C1(n20764), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(n20763), .ZN(n20765) );
  NOR4_X1 U23677 ( .A1(n20768), .A2(n20767), .A3(n20766), .A4(n20765), .ZN(
        n20800) );
  INV_X1 U23678 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20771) );
  INV_X1 U23679 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n20770) );
  AOI22_X1 U23680 ( .A1(n20771), .A2(keyinput42), .B1(keyinput10), .B2(n20770), 
        .ZN(n20769) );
  OAI221_X1 U23681 ( .B1(n20771), .B2(keyinput42), .C1(n20770), .C2(keyinput10), .A(n20769), .ZN(n20783) );
  INV_X1 U23682 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n20773) );
  AOI22_X1 U23683 ( .A1(n20774), .A2(keyinput12), .B1(n20773), .B2(keyinput3), 
        .ZN(n20772) );
  OAI221_X1 U23684 ( .B1(n20774), .B2(keyinput12), .C1(n20773), .C2(keyinput3), 
        .A(n20772), .ZN(n20782) );
  INV_X1 U23685 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n20776) );
  AOI22_X1 U23686 ( .A1(n20777), .A2(keyinput5), .B1(n20776), .B2(keyinput0), 
        .ZN(n20775) );
  OAI221_X1 U23687 ( .B1(n20777), .B2(keyinput5), .C1(n20776), .C2(keyinput0), 
        .A(n20775), .ZN(n20781) );
  INV_X1 U23688 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20779) );
  AOI22_X1 U23689 ( .A1(n11548), .A2(keyinput17), .B1(keyinput21), .B2(n20779), 
        .ZN(n20778) );
  OAI221_X1 U23690 ( .B1(n11548), .B2(keyinput17), .C1(n20779), .C2(keyinput21), .A(n20778), .ZN(n20780) );
  NOR4_X1 U23691 ( .A1(n20783), .A2(n20782), .A3(n20781), .A4(n20780), .ZN(
        n20799) );
  AOI22_X1 U23692 ( .A1(n20786), .A2(keyinput57), .B1(n20785), .B2(keyinput36), 
        .ZN(n20784) );
  OAI221_X1 U23693 ( .B1(n20786), .B2(keyinput57), .C1(n20785), .C2(keyinput36), .A(n20784), .ZN(n20797) );
  INV_X1 U23694 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20788) );
  AOI22_X1 U23695 ( .A1(n20788), .A2(keyinput20), .B1(n12773), .B2(keyinput61), 
        .ZN(n20787) );
  OAI221_X1 U23696 ( .B1(n20788), .B2(keyinput20), .C1(n12773), .C2(keyinput61), .A(n20787), .ZN(n20796) );
  AOI22_X1 U23697 ( .A1(n20791), .A2(keyinput4), .B1(n20790), .B2(keyinput30), 
        .ZN(n20789) );
  OAI221_X1 U23698 ( .B1(n20791), .B2(keyinput4), .C1(n20790), .C2(keyinput30), 
        .A(n20789), .ZN(n20795) );
  AOI22_X1 U23699 ( .A1(n10385), .A2(keyinput45), .B1(keyinput46), .B2(n20793), 
        .ZN(n20792) );
  OAI221_X1 U23700 ( .B1(n10385), .B2(keyinput45), .C1(n20793), .C2(keyinput46), .A(n20792), .ZN(n20794) );
  NOR4_X1 U23701 ( .A1(n20797), .A2(n20796), .A3(n20795), .A4(n20794), .ZN(
        n20798) );
  NAND4_X1 U23702 ( .A1(n20801), .A2(n20800), .A3(n20799), .A4(n20798), .ZN(
        n20802) );
  AOI211_X1 U23703 ( .C1(n20805), .C2(n20804), .A(n20803), .B(n20802), .ZN(
        n20819) );
  AOI22_X1 U23704 ( .A1(n20809), .A2(n20808), .B1(n20807), .B2(n20806), .ZN(
        n20810) );
  INV_X1 U23705 ( .A(n20810), .ZN(n20816) );
  OAI22_X1 U23706 ( .A1(n20814), .A2(n20813), .B1(n20812), .B2(n20811), .ZN(
        n20815) );
  AOI211_X1 U23707 ( .C1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .C2(n20817), .A(
        n20816), .B(n20815), .ZN(n20818) );
  XNOR2_X1 U23708 ( .A(n20819), .B(n20818), .ZN(P3_U2936) );
  INV_X1 U11069 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11104) );
  INV_X2 U11035 ( .A(n12280), .ZN(n16945) );
  CLKBUF_X2 U11028 ( .A(n10198), .Z(n13533) );
  BUF_X2 U11037 ( .A(n10179), .Z(n9651) );
  BUF_X2 U11064 ( .A(n10854), .Z(n9584) );
  BUF_X1 U11080 ( .A(n10854), .Z(n9583) );
  CLKBUF_X1 U11108 ( .A(n11326), .Z(n11299) );
  CLKBUF_X1 U11127 ( .A(n10120), .Z(n10855) );
  CLKBUF_X1 U11132 ( .A(n10155), .Z(n10842) );
  INV_X1 U11170 ( .A(n16872), .ZN(n12280) );
  INV_X1 U11180 ( .A(n10478), .ZN(n10894) );
  CLKBUF_X1 U11452 ( .A(n10165), .Z(n13450) );
  INV_X1 U11469 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19697) );
  CLKBUF_X1 U11508 ( .A(n10136), .Z(n12954) );
  CLKBUF_X1 U11562 ( .A(n10184), .Z(n10196) );
  CLKBUF_X1 U12284 ( .A(n17252), .Z(n17245) );
  CLKBUF_X1 U12285 ( .A(n16990), .Z(n9588) );
  CLKBUF_X1 U12316 ( .A(n16249), .Z(n16262) );
  CLKBUF_X1 U12649 ( .A(n13021), .Z(n20820) );
  CLKBUF_X1 U12782 ( .A(n11409), .Z(n11284) );
  CLKBUF_X1 U13199 ( .A(n18600), .Z(n17203) );
endmodule

