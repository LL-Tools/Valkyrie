

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530;

  AOI211_X1 U4893 ( .C1(n9342), .C2(n7698), .A(n9768), .B(n7788), .ZN(n7707)
         );
  NAND2_X1 U4894 ( .A1(n8601), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8639) );
  INV_X1 U4895 ( .A(n8160), .ZN(n8978) );
  CLKBUF_X2 U4896 ( .A(n6083), .Z(n6827) );
  NAND2_X1 U4897 ( .A1(n6910), .A2(n6724), .ZN(n4402) );
  BUF_X2 U4898 ( .A(n5488), .Z(n4716) );
  INV_X1 U4899 ( .A(n10013), .ZN(n9281) );
  INV_X1 U4900 ( .A(n7320), .ZN(n5716) );
  CLKBUF_X2 U4901 ( .A(n7584), .Z(n4395) );
  CLKBUF_X2 U4902 ( .A(n7297), .Z(n4725) );
  INV_X1 U4903 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5364) );
  NOR2_X1 U4904 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5358) );
  NOR2_X1 U4905 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5361) );
  NOR2_X1 U4906 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5357) );
  NAND4_X1 U4907 ( .A1(n10478), .A2(n5365), .A3(n5619), .A4(n5364), .ZN(n5665)
         );
  INV_X1 U4908 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4567) );
  INV_X1 U4909 ( .A(n7174), .ZN(n7249) );
  INV_X1 U4910 ( .A(n6565), .ZN(n5488) );
  NAND2_X1 U4912 ( .A1(n9610), .A2(n8273), .ZN(n6634) );
  NAND3_X1 U4913 ( .A1(n4567), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4568) );
  INV_X2 U4914 ( .A(n4402), .ZN(n7293) );
  INV_X1 U4915 ( .A(n8704), .ZN(n7164) );
  BUF_X1 U4916 ( .A(n6043), .Z(n6227) );
  XNOR2_X1 U4917 ( .A(n5993), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9114) );
  INV_X1 U4918 ( .A(n9183), .ZN(n7092) );
  NAND2_X1 U4919 ( .A1(n5519), .A2(n5269), .ZN(n5526) );
  INV_X1 U4920 ( .A(n5243), .ZN(n4396) );
  INV_X1 U4921 ( .A(n9507), .ZN(n9772) );
  INV_X1 U4922 ( .A(n4396), .ZN(n4397) );
  AOI211_X1 U4923 ( .C1(n8701), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8688), .B(
        n8687), .ZN(n8689) );
  CLKBUF_X3 U4925 ( .A(n4705), .Z(n4387) );
  OAI21_X1 U4926 ( .B1(n7888), .B2(n6953), .A(n6952), .ZN(n7958) );
  AOI21_X2 U4927 ( .B1(n9519), .B2(n10087), .A(n5880), .ZN(n4937) );
  NAND4_X2 U4928 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n8550)
         );
  INV_X2 U4929 ( .A(n8999), .ZN(n4392) );
  AND3_X4 U4930 ( .A1(n4462), .A2(n6037), .A3(n6038), .ZN(n8999) );
  NAND2_X4 U4931 ( .A1(n4569), .A2(n4568), .ZN(n7297) );
  BUF_X4 U4932 ( .A(n5555), .Z(n4388) );
  BUF_X4 U4933 ( .A(n5555), .Z(n4389) );
  AND2_X2 U4934 ( .A1(n5384), .A2(n9932), .ZN(n5555) );
  BUF_X1 U4935 ( .A(n6034), .Z(n7392) );
  INV_X4 U4936 ( .A(n4397), .ZN(n4815) );
  BUF_X4 U4937 ( .A(n9114), .Z(n4393) );
  NOR2_X2 U4938 ( .A1(n8646), .A2(n4682), .ZN(n8648) );
  NAND2_X1 U4939 ( .A1(n7320), .A2(n4397), .ZN(n4390) );
  NAND2_X2 U4940 ( .A1(n7320), .A2(n4758), .ZN(n6565) );
  AOI21_X2 U4941 ( .B1(n8596), .B2(n8595), .A(n4638), .ZN(n8617) );
  OR2_X1 U4942 ( .A1(n7698), .A2(n9342), .ZN(n7697) );
  NAND3_X2 U4943 ( .A1(n4840), .A2(n4839), .A3(n6772), .ZN(n8896) );
  AOI21_X2 U4944 ( .B1(n8639), .B2(n8637), .A(n8638), .ZN(n8646) );
  INV_X2 U4945 ( .A(n6048), .ZN(n6398) );
  INV_X1 U4946 ( .A(n6397), .ZN(n7530) );
  NAND4_X4 U4947 ( .A1(n6017), .A2(n5058), .A3(n5057), .A4(n5056), .ZN(n6397)
         );
  NOR2_X2 U4948 ( .A1(n4448), .A2(n8914), .ZN(n7484) );
  AND2_X2 U4949 ( .A1(n4835), .A2(n10136), .ZN(n8914) );
  OAI211_X2 U4950 ( .C1(n8987), .C2(n6400), .A(n6399), .B(n6731), .ZN(n10113)
         );
  AOI21_X2 U4951 ( .B1(n8053), .B2(n5479), .A(n5478), .ZN(n7997) );
  INV_X1 U4952 ( .A(n5775), .ZN(n4391) );
  BUF_X4 U4953 ( .A(n6934), .Z(n7040) );
  NOR4_X1 U4954 ( .A1(n8832), .A2(n8846), .A3(n8858), .A4(n6876), .ZN(n6877)
         );
  OR2_X1 U4955 ( .A1(n8871), .A2(n6875), .ZN(n6876) );
  NAND2_X2 U4956 ( .A1(n8190), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8260) );
  AOI21_X2 U4957 ( .B1(n9307), .B2(n9306), .A(n5223), .ZN(n9242) );
  XNOR2_X2 U4958 ( .A(n6226), .B(n6331), .ZN(n8704) );
  AOI22_X2 U4959 ( .A1(n8183), .A2(n8182), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n8181), .ZN(n8242) );
  AND2_X1 U4960 ( .A1(n4791), .A2(n4430), .ZN(n8745) );
  OAI21_X1 U4961 ( .B1(n6539), .B2(n6599), .A(n6617), .ZN(n6540) );
  NAND2_X1 U4962 ( .A1(n6409), .A2(n4837), .ZN(n8843) );
  NAND2_X1 U4963 ( .A1(n8856), .A2(n6785), .ZN(n6409) );
  AND2_X1 U4964 ( .A1(n5111), .A2(n9224), .ZN(n5114) );
  NAND2_X1 U4965 ( .A1(n8025), .A2(n8026), .ZN(n8000) );
  NAND2_X2 U4966 ( .A1(n8108), .A2(n8006), .ZN(n8026) );
  NAND2_X2 U4967 ( .A1(n4394), .A2(n6936), .ZN(n6459) );
  NAND2_X1 U4968 ( .A1(n7873), .A2(n10021), .ZN(n6653) );
  INV_X1 U4969 ( .A(n7170), .ZN(n7174) );
  INV_X1 U4970 ( .A(n6634), .ZN(n6630) );
  INV_X1 U4971 ( .A(n8551), .ZN(n7772) );
  OAI21_X1 U4972 ( .B1(n8332), .B2(n5563), .A(n5451), .ZN(n4672) );
  NAND2_X1 U4973 ( .A1(n5846), .A2(n6914), .ZN(n6917) );
  INV_X1 U4974 ( .A(n8549), .ZN(n8221) );
  INV_X1 U4975 ( .A(n8547), .ZN(n8504) );
  OR2_X1 U4976 ( .A1(n5603), .A2(n5602), .ZN(n5625) );
  OAI211_X1 U4977 ( .C1(n7320), .C2(n9422), .A(n5444), .B(n5443), .ZN(n7894)
         );
  NAND2_X1 U4978 ( .A1(n6060), .A2(n6059), .ZN(n8458) );
  CLKBUF_X2 U4979 ( .A(n6035), .Z(n6083) );
  NAND2_X1 U4980 ( .A1(n5516), .A2(n5268), .ZN(n5519) );
  CLKBUF_X1 U4981 ( .A(n6084), .Z(n4398) );
  INV_X1 U4982 ( .A(n5384), .ZN(n8340) );
  XNOR2_X1 U4983 ( .A(n5383), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U4984 ( .A1(n5842), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5906) );
  INV_X1 U4985 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4572) );
  NOR2_X1 U4986 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5981) );
  INV_X1 U4987 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5905) );
  AOI211_X1 U4988 ( .C1(n8660), .C2(n8670), .A(n8659), .B(n8658), .ZN(n8661)
         );
  OAI21_X1 U4989 ( .B1(n4822), .B2(n4819), .A(n4820), .ZN(n4818) );
  NAND2_X1 U4990 ( .A1(n4658), .A2(n5833), .ZN(n5187) );
  OR2_X1 U4991 ( .A1(n9806), .A2(n4726), .ZN(n9910) );
  NOR2_X1 U4992 ( .A1(n6626), .A2(n9610), .ZN(n6627) );
  CLKBUF_X1 U4993 ( .A(n6417), .Z(n4637) );
  CLKBUF_X1 U4994 ( .A(n9604), .Z(n9605) );
  OAI21_X1 U4995 ( .B1(n9620), .B2(n5754), .A(n5753), .ZN(n9604) );
  AND2_X1 U4996 ( .A1(n9785), .A2(n9784), .ZN(n4660) );
  INV_X1 U4997 ( .A(n6637), .ZN(n6689) );
  NAND2_X1 U4998 ( .A1(n6846), .A2(n6845), .ZN(n6894) );
  NAND2_X1 U4999 ( .A1(n6567), .A2(n6566), .ZN(n9766) );
  NAND2_X1 U5000 ( .A1(n6554), .A2(n6553), .ZN(n9507) );
  XNOR2_X1 U5001 ( .A(n6563), .B(n6562), .ZN(n9109) );
  OAI21_X1 U5002 ( .B1(n6560), .B2(n6559), .A(n6558), .ZN(n6563) );
  INV_X1 U5003 ( .A(n6593), .ZN(n5833) );
  XNOR2_X1 U5004 ( .A(n6560), .B(n6559), .ZN(n8339) );
  CLKBUF_X1 U5005 ( .A(n9164), .Z(n4720) );
  OAI21_X1 U5006 ( .B1(n6548), .B2(n6547), .A(n6546), .ZN(n6560) );
  OR2_X1 U5007 ( .A1(n5391), .A2(n9777), .ZN(n6617) );
  AND2_X1 U5008 ( .A1(n4890), .A2(n9954), .ZN(n9464) );
  XNOR2_X1 U5009 ( .A(n6548), .B(SI_29_), .ZN(n9117) );
  OR2_X1 U5010 ( .A1(n9540), .A2(n9798), .ZN(n6599) );
  INV_X1 U5011 ( .A(n4981), .ZN(n4980) );
  XNOR2_X1 U5012 ( .A(n6545), .B(n6544), .ZN(n6548) );
  NAND2_X1 U5013 ( .A1(n5375), .A2(n5374), .ZN(n5391) );
  NAND2_X1 U5014 ( .A1(n6598), .A2(n6612), .ZN(n9553) );
  AND2_X1 U5015 ( .A1(n5231), .A2(n4683), .ZN(n8190) );
  OAI21_X1 U5016 ( .B1(n5231), .B2(n8259), .A(n4986), .ZN(n4981) );
  NAND2_X1 U5017 ( .A1(n4847), .A2(n5921), .ZN(n6545) );
  NAND2_X1 U5018 ( .A1(n8863), .A2(n4423), .ZN(n8847) );
  NAND2_X1 U5019 ( .A1(n6309), .A2(n6308), .ZN(n9021) );
  OAI211_X1 U5020 ( .C1(n5867), .C2(n4589), .A(n4587), .B(n6640), .ZN(n9645)
         );
  NAND2_X1 U5021 ( .A1(n8188), .A2(n8202), .ZN(n5231) );
  AND2_X1 U5022 ( .A1(n5196), .A2(n5709), .ZN(n5195) );
  NAND2_X1 U5023 ( .A1(n4614), .A2(n9954), .ZN(n4613) );
  OR2_X1 U5024 ( .A1(n9056), .A2(n8468), .ZN(n6789) );
  NAND2_X1 U5025 ( .A1(n5744), .A2(n5743), .ZN(n9837) );
  AND2_X1 U5026 ( .A1(n6720), .A2(n6795), .ZN(n8810) );
  NAND2_X1 U5027 ( .A1(n6248), .A2(n6247), .ZN(n9056) );
  OAI21_X1 U5028 ( .B1(n8017), .B2(n4468), .A(n4770), .ZN(n8902) );
  NAND2_X1 U5029 ( .A1(n4585), .A2(n5725), .ZN(n9845) );
  NAND2_X1 U5030 ( .A1(n6240), .A2(n6239), .ZN(n9062) );
  XNOR2_X1 U5031 ( .A(n5742), .B(n5741), .ZN(n8265) );
  INV_X1 U5032 ( .A(n7219), .ZN(n8954) );
  NOR2_X1 U5033 ( .A1(n7982), .A2(n4539), .ZN(n7986) );
  NAND2_X1 U5034 ( .A1(n5700), .A2(n5699), .ZN(n9863) );
  XNOR2_X1 U5035 ( .A(n5737), .B(n5724), .ZN(n8210) );
  NAND2_X1 U5036 ( .A1(n6011), .A2(n6010), .ZN(n9077) );
  NAND2_X1 U5037 ( .A1(n4578), .A2(n5309), .ZN(n5712) );
  XNOR2_X1 U5038 ( .A(n5693), .B(n5692), .ZN(n7934) );
  XNOR2_X1 U5039 ( .A(n5682), .B(n5681), .ZN(n7864) );
  NAND2_X1 U5040 ( .A1(n4575), .A2(n5305), .ZN(n5693) );
  NAND2_X1 U5041 ( .A1(n5637), .A2(n5636), .ZN(n9746) );
  NAND3_X1 U5042 ( .A1(n4974), .A2(n4973), .A3(n4972), .ZN(n7655) );
  NAND2_X1 U5043 ( .A1(n4975), .A2(n7640), .ZN(n7653) );
  NAND2_X1 U5044 ( .A1(n6168), .A2(n6167), .ZN(n8900) );
  NAND2_X1 U5045 ( .A1(n6159), .A2(n6158), .ZN(n8160) );
  OR2_X1 U5046 ( .A1(n7550), .A2(n7549), .ZN(n7619) );
  CLKBUF_X1 U5047 ( .A(n8880), .Z(n8925) );
  NAND2_X1 U5048 ( .A1(n5566), .A2(n5565), .ZN(n10062) );
  NOR2_X2 U5049 ( .A1(n5673), .A2(n5672), .ZN(n9258) );
  AND2_X1 U5050 ( .A1(n4554), .A2(n4553), .ZN(n7518) );
  AND2_X1 U5051 ( .A1(n6743), .A2(n6749), .ZN(n7729) );
  NAND2_X1 U5052 ( .A1(n6459), .A2(n6653), .ZN(n8053) );
  NAND2_X1 U5053 ( .A1(n6133), .A2(n6132), .ZN(n8983) );
  AND2_X1 U5054 ( .A1(n5612), .A2(n5595), .ZN(n7416) );
  NOR2_X2 U5055 ( .A1(n7697), .A2(n7894), .ZN(n7874) );
  INV_X1 U5056 ( .A(n10027), .ZN(n8006) );
  NAND2_X1 U5057 ( .A1(n9183), .A2(n6934), .ZN(n4650) );
  INV_X1 U5058 ( .A(n6934), .ZN(n9179) );
  NAND2_X1 U5059 ( .A1(n5551), .A2(n5550), .ZN(n10054) );
  NAND2_X1 U5060 ( .A1(n6080), .A2(n6079), .ZN(n7732) );
  AND2_X1 U5061 ( .A1(n6069), .A2(n6068), .ZN(n10152) );
  BUF_X2 U5062 ( .A(n4672), .Z(n4394) );
  NAND3_X2 U5063 ( .A1(n6917), .A2(n7291), .A3(n6916), .ZN(n6934) );
  NAND4_X2 U5064 ( .A1(n5465), .A2(n5464), .A3(n5463), .A4(n5462), .ZN(n9389)
         );
  INV_X1 U5065 ( .A(n7894), .ZN(n10006) );
  INV_X1 U5066 ( .A(n9176), .ZN(n6941) );
  OAI211_X2 U5067 ( .C1(n7120), .C2(n6914), .A(n7291), .B(n8036), .ZN(n9183)
         );
  OR2_X1 U5069 ( .A1(n5168), .A2(n5167), .ZN(n5162) );
  AND4_X1 U5070 ( .A1(n5458), .A2(n5457), .A3(n5456), .A4(n5455), .ZN(n6936)
         );
  INV_X1 U5071 ( .A(n5934), .ZN(n5846) );
  NAND2_X1 U5072 ( .A1(n5483), .A2(n5450), .ZN(n8332) );
  BUF_X2 U5073 ( .A(n5527), .Z(n5923) );
  NAND2_X1 U5074 ( .A1(n4987), .A2(n7444), .ZN(n7557) );
  AND2_X1 U5075 ( .A1(n5291), .A2(n5169), .ZN(n5168) );
  OR2_X1 U5076 ( .A1(n5449), .A2(SI_5_), .ZN(n5450) );
  NAND2_X1 U5077 ( .A1(n8340), .A2(n5385), .ZN(n5775) );
  NAND2_X1 U5078 ( .A1(n6036), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5057) );
  NOR2_X1 U5079 ( .A1(n8315), .A2(n9939), .ZN(n4710) );
  NAND2_X1 U5080 ( .A1(n5714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5715) );
  CLKBUF_X3 U5081 ( .A(n4415), .Z(n6246) );
  NAND2_X1 U5082 ( .A1(n4738), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U5083 ( .A1(n5885), .A2(n5886), .ZN(n8315) );
  INV_X1 U5084 ( .A(n5385), .ZN(n9932) );
  NAND2_X1 U5085 ( .A1(n5093), .A2(n5256), .ZN(n5481) );
  INV_X1 U5086 ( .A(n6039), .ZN(n6127) );
  NAND2_X1 U5087 ( .A1(n5142), .A2(n4425), .ZN(n5141) );
  AND2_X1 U5088 ( .A1(n8212), .A2(n6645), .ZN(n6915) );
  OAI211_X1 U5089 ( .C1(n5906), .C2(n5150), .A(n5147), .B(n5145), .ZN(n9944)
         );
  INV_X1 U5090 ( .A(n8273), .ZN(n6914) );
  NAND2_X1 U5091 ( .A1(n4654), .A2(n4454), .ZN(n9939) );
  XNOR2_X1 U5092 ( .A(n4593), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5384) );
  AND2_X1 U5093 ( .A1(n9114), .A2(n5994), .ZN(n6084) );
  NAND2_X1 U5094 ( .A1(n7440), .A2(n7506), .ZN(n7445) );
  XNOR2_X1 U5095 ( .A(n5906), .B(n5905), .ZN(n8273) );
  NAND2_X1 U5096 ( .A1(n5889), .A2(n4719), .ZN(n5083) );
  NAND3_X1 U5097 ( .A1(n4671), .A2(n4848), .A3(n5401), .ZN(n5441) );
  NAND2_X1 U5098 ( .A1(n4594), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4593) );
  NAND2_X1 U5099 ( .A1(n5255), .A2(n5472), .ZN(n5092) );
  NAND2_X1 U5100 ( .A1(n6353), .A2(n4618), .ZN(n8266) );
  NAND2_X1 U5101 ( .A1(n6365), .A2(n6366), .ZN(n8312) );
  XNOR2_X1 U5102 ( .A(n5845), .B(n5844), .ZN(n8269) );
  NAND2_X1 U5103 ( .A1(n6004), .A2(n4464), .ZN(n4816) );
  CLKBUF_X1 U5104 ( .A(n5841), .Z(n5842) );
  NAND2_X2 U5105 ( .A1(n4397), .A2(P2_U3151), .ZN(n9132) );
  OR2_X1 U5106 ( .A1(n4849), .A2(n5246), .ZN(n5401) );
  XNOR2_X1 U5107 ( .A(n5270), .B(SI_8_), .ZN(n5525) );
  CLKBUF_X1 U5108 ( .A(n6000), .Z(n6005) );
  XNOR2_X1 U5109 ( .A(n5274), .B(SI_9_), .ZN(n5546) );
  NOR2_X1 U5110 ( .A1(n5367), .A2(n5214), .ZN(n5213) );
  AND2_X1 U5111 ( .A1(n5259), .A2(n5258), .ZN(n5480) );
  XNOR2_X1 U5112 ( .A(n6012), .B(P2_IR_REG_2__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U5113 ( .A1(n6041), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6012) );
  AND2_X1 U5114 ( .A1(n6090), .A2(n6008), .ZN(n4628) );
  NAND2_X2 U5115 ( .A1(n6042), .A2(n6041), .ZN(n7599) );
  NAND3_X1 U5116 ( .A1(n4572), .A2(n4571), .A3(n4570), .ZN(n4569) );
  MUX2_X1 U5117 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6040), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6042) );
  INV_X1 U5118 ( .A(n7433), .ZN(n6041) );
  NOR2_X1 U5119 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5363) );
  INV_X1 U5120 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6185) );
  INV_X1 U5121 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6128) );
  NOR2_X1 U5122 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5972) );
  NOR2_X1 U5123 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5971) );
  INV_X1 U5124 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n10243) );
  INV_X1 U5125 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6008) );
  INV_X4 U5126 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5127 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5578) );
  NOR2_X1 U5128 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5371) );
  INV_X1 U5129 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5365) );
  NOR2_X1 U5130 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5359) );
  NOR2_X2 U5131 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5835) );
  INV_X1 U5132 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5844) );
  NOR3_X1 U5133 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .A3(
        P2_IR_REG_2__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U5134 ( .A1(n7958), .A2(n6958), .ZN(n6961) );
  INV_X1 U5135 ( .A(n5848), .ZN(n7692) );
  OAI21_X2 U5136 ( .B1(n7936), .B2(n6757), .A(n4706), .ZN(n6405) );
  NAND2_X2 U5137 ( .A1(n6402), .A2(n6864), .ZN(n7936) );
  BUF_X4 U5138 ( .A(n6084), .Z(n4399) );
  NOR2_X2 U5139 ( .A1(n6920), .A2(n9338), .ZN(n9209) );
  OAI21_X2 U5140 ( .B1(n9210), .B2(n9338), .A(n9337), .ZN(n9336) );
  AND2_X2 U5141 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  OAI21_X2 U5142 ( .B1(n8896), .B2(n6407), .A(n6776), .ZN(n8868) );
  OR2_X2 U5143 ( .A1(n5934), .A2(n4530), .ZN(n7120) );
  NOR2_X2 U5144 ( .A1(n8054), .A2(n4394), .ZN(n8002) );
  INV_X1 U5145 ( .A(n7320), .ZN(n4400) );
  NOR2_X2 U5146 ( .A1(n7890), .A2(n7889), .ZN(n7888) );
  INV_X1 U5147 ( .A(n5576), .ZN(n4558) );
  AND2_X1 U5148 ( .A1(n4951), .A2(n9591), .ZN(n4955) );
  NAND2_X1 U5149 ( .A1(n9845), .A2(n9833), .ZN(n6507) );
  OAI21_X1 U5150 ( .B1(n6584), .B2(n8139), .A(n6481), .ZN(n5855) );
  NAND2_X1 U5151 ( .A1(n5794), .A2(n5795), .ZN(n4844) );
  AOI22_X1 U5152 ( .A1(n8729), .A2(n6320), .B1(n6319), .B2(n7280), .ZN(n7144)
         );
  OR2_X1 U5153 ( .A1(n9812), .A2(n9598), .ZN(n6602) );
  AND2_X1 U5154 ( .A1(n9573), .A2(n4595), .ZN(n9558) );
  NOR2_X1 U5155 ( .A1(n9560), .A2(n4596), .ZN(n4595) );
  INV_X1 U5156 ( .A(n6602), .ZN(n4596) );
  OR2_X1 U5157 ( .A1(n6663), .A2(n4475), .ZN(n4752) );
  AND2_X1 U5158 ( .A1(n6469), .A2(n6657), .ZN(n4754) );
  OAI21_X1 U5159 ( .B1(n6509), .B2(n6506), .A(n6508), .ZN(n6521) );
  NAND2_X1 U5160 ( .A1(n8049), .A2(n10013), .ZN(n6452) );
  AND3_X1 U5161 ( .A1(n4551), .A2(n6718), .A3(n4550), .ZN(n6824) );
  NAND2_X1 U5162 ( .A1(n6837), .A2(n4402), .ZN(n6718) );
  OAI21_X1 U5163 ( .B1(n9117), .B2(n4548), .A(n4545), .ZN(n4550) );
  INV_X1 U5164 ( .A(n9665), .ZN(n5199) );
  NAND2_X1 U5165 ( .A1(n5312), .A2(n5311), .ZN(n5315) );
  XNOR2_X1 U5166 ( .A(n7761), .B(n7249), .ZN(n7181) );
  INV_X1 U5167 ( .A(n4393), .ZN(n5043) );
  OR2_X1 U5168 ( .A1(n6838), .A2(n6837), .ZN(n7141) );
  OR2_X1 U5169 ( .A1(n6323), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8334) );
  INV_X1 U5170 ( .A(n8730), .ZN(n7148) );
  AND2_X1 U5171 ( .A1(n9027), .A2(n8422), .ZN(n6818) );
  AND2_X1 U5172 ( .A1(n9044), .A2(n8790), .ZN(n8773) );
  AND2_X1 U5173 ( .A1(n5032), .A2(n5033), .ZN(n5031) );
  INV_X1 U5174 ( .A(n8823), .ZN(n5032) );
  OR2_X1 U5175 ( .A1(n9068), .A2(n8835), .ZN(n6788) );
  NAND2_X1 U5176 ( .A1(n8875), .A2(n4424), .ZN(n8857) );
  OR2_X1 U5177 ( .A1(n8963), .A2(n8889), .ZN(n6779) );
  NAND2_X1 U5178 ( .A1(n4401), .A2(n5026), .ZN(n5025) );
  INV_X1 U5179 ( .A(n6155), .ZN(n5026) );
  INV_X1 U5180 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5181 ( .A1(n4650), .A2(n8325), .ZN(n6926) );
  NAND2_X1 U5182 ( .A1(n4892), .A2(n4891), .ZN(n4890) );
  NAND2_X1 U5183 ( .A1(n9466), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4891) );
  OR2_X1 U5184 ( .A1(n9779), .A2(n9521), .ZN(n6618) );
  NOR2_X1 U5185 ( .A1(n5182), .A2(n5793), .ZN(n5180) );
  NOR2_X1 U5186 ( .A1(n9600), .A2(n9825), .ZN(n5780) );
  INV_X1 U5187 ( .A(n9606), .ZN(n4961) );
  OR2_X1 U5188 ( .A1(n9845), .A2(n9851), .ZN(n5733) );
  NOR2_X1 U5189 ( .A1(n9845), .A2(n9657), .ZN(n5076) );
  OR2_X1 U5190 ( .A1(n9863), .A2(n9261), .ZN(n6515) );
  OR2_X1 U5191 ( .A1(n9877), .A2(n9725), .ZN(n6671) );
  NAND2_X1 U5192 ( .A1(n4737), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5603) );
  INV_X1 U5193 ( .A(n5584), .ZN(n4737) );
  OR2_X1 U5194 ( .A1(n10054), .A2(n10039), .ZN(n6470) );
  INV_X1 U5195 ( .A(n5563), .ZN(n5527) );
  NAND2_X1 U5196 ( .A1(n5355), .A2(n5354), .ZN(n5917) );
  NAND4_X1 U5197 ( .A1(n4656), .A2(n5596), .A3(n4655), .A4(n5844), .ZN(n5841)
         );
  AOI21_X1 U5198 ( .B1(n5782), .B2(n4562), .A(n4561), .ZN(n4560) );
  INV_X1 U5199 ( .A(n5782), .ZN(n4563) );
  INV_X1 U5200 ( .A(n5333), .ZN(n4562) );
  AND2_X1 U5201 ( .A1(n5344), .A2(n5343), .ZN(n5795) );
  OAI21_X1 U5202 ( .B1(n5712), .B2(n5713), .A(n5315), .ZN(n5737) );
  NAND2_X1 U5203 ( .A1(n5305), .A2(n5304), .ZN(n5681) );
  NOR2_X1 U5204 ( .A1(n4466), .A2(n4556), .ZN(n4555) );
  INV_X1 U5205 ( .A(n5283), .ZN(n4556) );
  NAND2_X1 U5206 ( .A1(n4557), .A2(n5283), .ZN(n5594) );
  OR2_X1 U5207 ( .A1(n5594), .A2(n5593), .ZN(n5612) );
  NAND2_X1 U5208 ( .A1(n4629), .A2(n4441), .ZN(n7968) );
  AND2_X1 U5209 ( .A1(n7835), .A2(n7182), .ZN(n5014) );
  AND2_X1 U5210 ( .A1(n6222), .A2(n6221), .ZN(n7222) );
  NAND2_X1 U5211 ( .A1(n4398), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U5212 ( .A1(n7559), .A2(n7560), .ZN(n7606) );
  NAND2_X1 U5213 ( .A1(n7141), .A2(n7140), .ZN(n7151) );
  NAND2_X1 U5214 ( .A1(n6311), .A2(n6310), .ZN(n6323) );
  INV_X1 U5215 ( .A(n6312), .ZN(n6311) );
  NAND2_X1 U5216 ( .A1(n4774), .A2(n6141), .ZN(n8151) );
  NAND2_X1 U5217 ( .A1(n8017), .A2(n6140), .ZN(n4774) );
  INV_X1 U5218 ( .A(n8266), .ZN(n6724) );
  INV_X1 U5219 ( .A(n8740), .ZN(n7280) );
  XNOR2_X1 U5220 ( .A(n7285), .B(n7148), .ZN(n6883) );
  INV_X1 U5221 ( .A(n4776), .ZN(n8729) );
  OAI21_X1 U5222 ( .B1(n8774), .B2(n4470), .A(n4777), .ZN(n4776) );
  AOI21_X1 U5223 ( .B1(n4778), .B2(n6307), .A(n4789), .ZN(n4777) );
  OR2_X1 U5224 ( .A1(n9039), .A2(n8778), .ZN(n8759) );
  NOR2_X1 U5225 ( .A1(n6276), .A2(n4453), .ZN(n4788) );
  NAND2_X1 U5226 ( .A1(n8774), .A2(n6277), .ZN(n4784) );
  AND2_X1 U5227 ( .A1(n6264), .A2(n6263), .ZN(n8777) );
  INV_X1 U5228 ( .A(n8832), .ZN(n6410) );
  XNOR2_X1 U5229 ( .A(n9077), .B(n8861), .ZN(n8846) );
  OR2_X1 U5230 ( .A1(n9083), .A2(n8878), .ZN(n6784) );
  OR2_X1 U5231 ( .A1(n4842), .A2(n6767), .ZN(n4839) );
  NAND2_X1 U5232 ( .A1(n5992), .A2(n5991), .ZN(n5994) );
  NOR2_X1 U5233 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5989) );
  AND2_X1 U5234 ( .A1(n9169), .A2(n7047), .ZN(n7048) );
  INV_X1 U5235 ( .A(n9194), .ZN(n5105) );
  AND2_X1 U5236 ( .A1(n9218), .A2(n5134), .ZN(n5124) );
  NAND2_X1 U5237 ( .A1(n5110), .A2(n5109), .ZN(n5115) );
  INV_X1 U5238 ( .A(n4507), .ZN(n5109) );
  INV_X1 U5239 ( .A(n5812), .ZN(n5872) );
  AND2_X1 U5240 ( .A1(n8122), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8123) );
  INV_X1 U5241 ( .A(n9481), .ZN(n4686) );
  INV_X1 U5242 ( .A(n9480), .ZN(n4687) );
  NAND2_X1 U5243 ( .A1(n4886), .A2(n4510), .ZN(n9958) );
  INV_X1 U5244 ( .A(n9961), .ZN(n4885) );
  XNOR2_X1 U5245 ( .A(n4598), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U5246 ( .A1(n9962), .A2(n9495), .ZN(n4598) );
  NAND2_X1 U5247 ( .A1(n5948), .A2(n4418), .ZN(n9785) );
  NAND2_X1 U5248 ( .A1(n5391), .A2(n9777), .ZN(n6440) );
  INV_X1 U5249 ( .A(n5154), .ZN(n5153) );
  NAND2_X1 U5250 ( .A1(n9558), .A2(n5157), .ZN(n5156) );
  OAI21_X1 U5251 ( .B1(n5155), .B2(n5833), .A(n6439), .ZN(n5154) );
  AND2_X1 U5252 ( .A1(n5175), .A2(n5805), .ZN(n5174) );
  NOR2_X1 U5253 ( .A1(n9808), .A2(n5078), .ZN(n5077) );
  INV_X1 U5254 ( .A(n5079), .ZN(n5078) );
  AND2_X1 U5255 ( .A1(n5818), .A2(n5817), .ZN(n9562) );
  NAND2_X1 U5256 ( .A1(n4950), .A2(n4947), .ZN(n9573) );
  AND2_X1 U5257 ( .A1(n4493), .A2(n4948), .ZN(n4947) );
  NAND2_X1 U5258 ( .A1(n4955), .A2(n9629), .ZN(n4950) );
  INV_X1 U5259 ( .A(n9816), .ZN(n9598) );
  AOI21_X1 U5260 ( .B1(n6443), .B2(n4961), .A(n4959), .ZN(n4958) );
  INV_X1 U5261 ( .A(n6526), .ZN(n4959) );
  AND2_X1 U5262 ( .A1(n9837), .A2(n9842), .ZN(n6443) );
  XNOR2_X1 U5263 ( .A(n9837), .B(n9824), .ZN(n9628) );
  NAND2_X1 U5264 ( .A1(n6515), .A2(n6517), .ZN(n9667) );
  OR2_X1 U5265 ( .A1(n9869), .A2(n9874), .ZN(n6673) );
  AND2_X1 U5266 ( .A1(n6658), .A2(n5856), .ZN(n4938) );
  INV_X1 U5267 ( .A(n8230), .ZN(n5856) );
  AND2_X1 U5268 ( .A1(n9405), .A2(n7318), .ZN(n10053) );
  INV_X1 U5269 ( .A(n9986), .ZN(n10065) );
  NAND2_X1 U5270 ( .A1(n4471), .A2(n5370), .ZN(n5214) );
  XNOR2_X1 U5271 ( .A(n5917), .B(n5918), .ZN(n8316) );
  XNOR2_X1 U5272 ( .A(n8712), .B(n4643), .ZN(n4642) );
  INV_X1 U5273 ( .A(n8713), .ZN(n4643) );
  OAI22_X1 U5274 ( .A1(n8711), .A2(n8710), .B1(n8709), .B2(n10231), .ZN(n8712)
         );
  OR2_X1 U5275 ( .A1(n9193), .A2(n5108), .ZN(n5107) );
  OR2_X1 U5276 ( .A1(n9192), .A2(n9380), .ZN(n5108) );
  NOR2_X1 U5277 ( .A1(n4433), .A2(n4603), .ZN(n7359) );
  NAND2_X1 U5278 ( .A1(n4920), .A2(n4402), .ZN(n6727) );
  MUX2_X1 U5279 ( .A(n6753), .B(n6752), .S(n7293), .Z(n6755) );
  NAND2_X1 U5280 ( .A1(n4805), .A2(n7293), .ZN(n4804) );
  INV_X1 U5281 ( .A(n6757), .ZN(n4805) );
  NOR2_X1 U5282 ( .A1(n6755), .A2(n7821), .ZN(n4926) );
  AOI21_X1 U5283 ( .B1(n4798), .B2(n4797), .A(n4467), .ZN(n6750) );
  NOR2_X1 U5284 ( .A1(n6744), .A2(n6745), .ZN(n4797) );
  NAND2_X1 U5285 ( .A1(n6747), .A2(n6746), .ZN(n4798) );
  INV_X1 U5286 ( .A(n6787), .ZN(n4793) );
  NAND2_X1 U5287 ( .A1(n6485), .A2(n6630), .ZN(n4664) );
  OAI21_X1 U5288 ( .B1(n6809), .B2(n8773), .A(n6880), .ZN(n4936) );
  AND2_X1 U5289 ( .A1(n8759), .A2(n7293), .ZN(n4935) );
  NOR2_X1 U5290 ( .A1(n4932), .A2(n7293), .ZN(n4931) );
  INV_X1 U5291 ( .A(n8758), .ZN(n4932) );
  NAND2_X1 U5292 ( .A1(n4429), .A2(n6519), .ZN(n4544) );
  AND2_X1 U5293 ( .A1(n7871), .A2(n8025), .ZN(n4668) );
  INV_X1 U5294 ( .A(n6584), .ZN(n4669) );
  INV_X1 U5295 ( .A(n4625), .ZN(n4624) );
  OAI21_X1 U5296 ( .B1(n8377), .B2(n4626), .A(n5224), .ZN(n4625) );
  MUX2_X1 U5297 ( .A(n7148), .B(n7147), .S(n4402), .Z(n6834) );
  NAND2_X1 U5298 ( .A1(n4810), .A2(n4811), .ZN(n4559) );
  AND2_X1 U5299 ( .A1(n8758), .A2(n8771), .ZN(n6880) );
  INV_X1 U5300 ( .A(n5662), .ZN(n5298) );
  AOI21_X1 U5301 ( .B1(n5168), .B2(n5292), .A(n5165), .ZN(n5164) );
  OR2_X1 U5302 ( .A1(n5167), .A2(n5293), .ZN(n5165) );
  INV_X1 U5303 ( .A(n8385), .ZN(n5004) );
  AND2_X1 U5304 ( .A1(n5001), .A2(n4623), .ZN(n4622) );
  NAND2_X1 U5305 ( .A1(n4624), .A2(n4626), .ZN(n4623) );
  AND2_X1 U5306 ( .A1(n5002), .A2(n8399), .ZN(n5001) );
  NAND2_X1 U5307 ( .A1(n8467), .A2(n5224), .ZN(n5002) );
  NAND2_X1 U5308 ( .A1(n7215), .A2(n8878), .ZN(n5023) );
  NAND2_X1 U5309 ( .A1(n9018), .A2(n8542), .ZN(n6839) );
  AOI21_X1 U5310 ( .B1(n7577), .B2(n7578), .A(n4899), .ZN(n7425) );
  NAND2_X1 U5311 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  NOR2_X1 U5312 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n4869) );
  INV_X1 U5313 ( .A(n6282), .ZN(n6281) );
  AND2_X1 U5314 ( .A1(n6230), .A2(n4875), .ZN(n4874) );
  INV_X1 U5315 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n4875) );
  INV_X1 U5316 ( .A(n6232), .ZN(n6231) );
  AND2_X1 U5317 ( .A1(n5968), .A2(n4872), .ZN(n4871) );
  INV_X1 U5318 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4872) );
  INV_X1 U5319 ( .A(n6193), .ZN(n5969) );
  INV_X1 U5320 ( .A(n6861), .ZN(n8012) );
  AND2_X1 U5321 ( .A1(n5962), .A2(n4879), .ZN(n4878) );
  INV_X1 U5322 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n4879) );
  AND2_X1 U5323 ( .A1(n8218), .A2(n8548), .ZN(n6861) );
  NAND2_X1 U5324 ( .A1(n6112), .A2(n4768), .ZN(n4767) );
  INV_X1 U5325 ( .A(n6102), .ZN(n4768) );
  INV_X1 U5326 ( .A(n6119), .ZN(n5963) );
  AND2_X1 U5327 ( .A1(n4474), .A2(n6868), .ZN(n5046) );
  NOR2_X1 U5328 ( .A1(n10109), .A2(n10147), .ZN(n6745) );
  AND2_X1 U5329 ( .A1(n7163), .A2(n7334), .ZN(n6702) );
  AND2_X1 U5330 ( .A1(n6378), .A2(n7336), .ZN(n6430) );
  INV_X1 U5331 ( .A(n4780), .ZN(n4778) );
  AND2_X1 U5332 ( .A1(n9027), .A2(n8747), .ZN(n4789) );
  INV_X1 U5333 ( .A(n6277), .ZN(n4782) );
  NOR2_X1 U5334 ( .A1(n6812), .A2(n4787), .ZN(n4786) );
  INV_X1 U5335 ( .A(n4788), .ZN(n4787) );
  INV_X1 U5336 ( .A(n4422), .ZN(n5030) );
  NAND2_X1 U5337 ( .A1(n8494), .A2(n8412), .ZN(n6764) );
  OR2_X1 U5338 ( .A1(n9093), .A2(n8536), .ZN(n6775) );
  NAND2_X1 U5339 ( .A1(n4769), .A2(n4407), .ZN(n4771) );
  INV_X1 U5340 ( .A(n5025), .ZN(n4769) );
  INV_X1 U5341 ( .A(n6140), .ZN(n4772) );
  OR2_X1 U5342 ( .A1(n6057), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6064) );
  AOI22_X1 U5343 ( .A1(n4412), .A2(n8106), .B1(n6963), .B2(n5120), .ZN(n5119)
         );
  XNOR2_X1 U5344 ( .A(n4692), .B(n7040), .ZN(n6919) );
  NAND2_X1 U5345 ( .A1(n4581), .A2(n4580), .ZN(n4744) );
  NOR2_X1 U5346 ( .A1(n6540), .A2(n6630), .ZN(n4580) );
  NAND2_X1 U5347 ( .A1(n4582), .A2(n6612), .ZN(n4581) );
  NAND2_X1 U5348 ( .A1(n4745), .A2(n4746), .ZN(n4582) );
  NOR2_X1 U5349 ( .A1(n4613), .A2(n9468), .ZN(n4616) );
  NOR2_X1 U5350 ( .A1(n5810), .A2(n9363), .ZN(n4742) );
  INV_X1 U5351 ( .A(n4742), .ZN(n5825) );
  OR2_X1 U5352 ( .A1(n9801), .A2(n9562), .ZN(n6598) );
  NOR2_X1 U5353 ( .A1(n9812), .A2(n9600), .ZN(n5079) );
  NAND2_X1 U5354 ( .A1(n4417), .A2(n5723), .ZN(n5209) );
  NOR2_X1 U5355 ( .A1(n5734), .A2(n5211), .ZN(n5210) );
  INV_X1 U5356 ( .A(n5723), .ZN(n5211) );
  INV_X1 U5357 ( .A(n4965), .ZN(n4588) );
  NOR2_X1 U5358 ( .A1(n5072), .A2(n5860), .ZN(n5071) );
  NAND2_X1 U5359 ( .A1(n9895), .A2(n5073), .ZN(n5072) );
  NOR2_X1 U5360 ( .A1(n10043), .A2(n10054), .ZN(n5065) );
  INV_X1 U5361 ( .A(n5193), .ZN(n5192) );
  OAI21_X1 U5362 ( .B1(n8171), .B2(n5194), .A(n8142), .ZN(n5193) );
  INV_X1 U5363 ( .A(n5544), .ZN(n5194) );
  NAND2_X1 U5364 ( .A1(n5377), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5538) );
  INV_X1 U5365 ( .A(n5505), .ZN(n5377) );
  NAND2_X1 U5366 ( .A1(n9294), .A2(n10043), .ZN(n6465) );
  INV_X1 U5367 ( .A(n6447), .ZN(n4718) );
  INV_X1 U5368 ( .A(n9342), .ZN(n6929) );
  INV_X1 U5369 ( .A(n7665), .ZN(n7663) );
  NAND2_X1 U5370 ( .A1(n8228), .A2(n5858), .ZN(n9983) );
  AND2_X1 U5371 ( .A1(n5354), .A2(n5353), .ZN(n5822) );
  AND2_X1 U5372 ( .A1(n5349), .A2(n5348), .ZN(n5807) );
  AND2_X1 U5373 ( .A1(n5339), .A2(n5338), .ZN(n5782) );
  AOI21_X1 U5374 ( .B1(n4853), .B2(n4856), .A(n4852), .ZN(n4851) );
  INV_X1 U5375 ( .A(n5768), .ZN(n4852) );
  NOR2_X1 U5376 ( .A1(n5310), .A2(n4574), .ZN(n4573) );
  INV_X1 U5377 ( .A(n5305), .ZN(n4574) );
  INV_X1 U5378 ( .A(n5692), .ZN(n5310) );
  INV_X1 U5379 ( .A(n4861), .ZN(n4860) );
  OAI21_X1 U5380 ( .B1(n5322), .B2(n4862), .A(n5321), .ZN(n4861) );
  NAND2_X1 U5381 ( .A1(n5713), .A2(n5315), .ZN(n4862) );
  XNOR2_X1 U5382 ( .A(n5307), .B(SI_18_), .ZN(n5692) );
  NAND2_X1 U5383 ( .A1(n4579), .A2(n4576), .ZN(n4575) );
  NOR2_X1 U5384 ( .A1(n4577), .A2(n5681), .ZN(n4576) );
  INV_X1 U5385 ( .A(n5299), .ZN(n4577) );
  NAND2_X1 U5386 ( .A1(n5298), .A2(SI_16_), .ZN(n5299) );
  NAND2_X1 U5387 ( .A1(n5288), .A2(n10342), .ZN(n5614) );
  NAND2_X1 U5388 ( .A1(n5267), .A2(SI_7_), .ZN(n5269) );
  INV_X1 U5389 ( .A(n5092), .ZN(n5256) );
  OR2_X1 U5390 ( .A1(n7297), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U5391 ( .A1(n5251), .A2(SI_3_), .ZN(n5470) );
  INV_X1 U5392 ( .A(SI_13_), .ZN(n10342) );
  INV_X1 U5393 ( .A(n8312), .ZN(n6371) );
  XNOR2_X1 U5394 ( .A(n7170), .B(n10114), .ZN(n7175) );
  NAND2_X1 U5395 ( .A1(n4998), .A2(n8999), .ZN(n7169) );
  INV_X1 U5396 ( .A(n7240), .ZN(n5008) );
  AND2_X1 U5397 ( .A1(n8217), .A2(n7191), .ZN(n5006) );
  AND2_X1 U5398 ( .A1(n5994), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5042) );
  AND2_X1 U5399 ( .A1(n6852), .A2(n6348), .ZN(n6837) );
  NAND2_X1 U5400 ( .A1(n4917), .A2(n9118), .ZN(n4916) );
  AND2_X1 U5401 ( .A1(n4393), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4917) );
  OAI21_X1 U5402 ( .B1(n9125), .B2(n4712), .A(n4711), .ZN(n7451) );
  NAND2_X1 U5403 ( .A1(n9125), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4711) );
  OR2_X1 U5404 ( .A1(n7555), .A2(n7419), .ZN(n4907) );
  NAND2_X1 U5405 ( .A1(n4977), .A2(n7640), .ZN(n4976) );
  INV_X1 U5406 ( .A(n7605), .ZN(n4977) );
  NAND2_X1 U5407 ( .A1(n7606), .A2(n4443), .ZN(n4972) );
  NAND2_X1 U5408 ( .A1(n7616), .A2(n7615), .ZN(n7649) );
  NAND2_X1 U5409 ( .A1(n8189), .A2(n8243), .ZN(n4683) );
  NAND2_X1 U5410 ( .A1(n8196), .A2(n8195), .ZN(n8253) );
  OR2_X1 U5411 ( .A1(n8243), .A2(n10343), .ZN(n4913) );
  NAND2_X1 U5412 ( .A1(n8604), .A2(n8605), .ZN(n8630) );
  NAND2_X1 U5413 ( .A1(n4996), .A2(n4993), .ZN(n4991) );
  INV_X1 U5414 ( .A(n8669), .ZN(n4993) );
  AOI22_X1 U5415 ( .A1(n8665), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n4895), .B2(
        n8664), .ZN(n8711) );
  NAND2_X1 U5416 ( .A1(n6281), .A2(n4869), .ZN(n6300) );
  OR2_X1 U5417 ( .A1(n6268), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6282) );
  OR2_X1 U5418 ( .A1(n6258), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6268) );
  OR2_X1 U5419 ( .A1(n6216), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U5420 ( .A1(n5969), .A2(n4871), .ZN(n6206) );
  NAND2_X1 U5421 ( .A1(n5969), .A2(n5968), .ZN(n6204) );
  NAND2_X1 U5422 ( .A1(n5965), .A2(n5964), .ZN(n6169) );
  INV_X1 U5423 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5964) );
  INV_X1 U5424 ( .A(n6160), .ZN(n5965) );
  NAND2_X1 U5425 ( .A1(n5024), .A2(n6126), .ZN(n8017) );
  AND2_X1 U5426 ( .A1(n7824), .A2(n6749), .ZN(n5061) );
  NAND2_X1 U5427 ( .A1(n4405), .A2(n5047), .ZN(n7827) );
  INV_X1 U5428 ( .A(n6723), .ZN(n4835) );
  AND2_X1 U5429 ( .A1(n6389), .A2(n4402), .ZN(n6703) );
  NAND2_X1 U5430 ( .A1(n4549), .A2(n6717), .ZN(n6838) );
  AND2_X1 U5431 ( .A1(n7155), .A2(n7154), .ZN(n4823) );
  OAI21_X1 U5432 ( .B1(n7151), .B2(n4427), .A(n5227), .ZN(n7152) );
  NOR2_X1 U5433 ( .A1(n8888), .A2(n6837), .ZN(n6350) );
  INV_X1 U5434 ( .A(n8728), .ZN(n8726) );
  AOI21_X1 U5435 ( .B1(n4828), .B2(n4830), .A(n6816), .ZN(n4827) );
  INV_X1 U5436 ( .A(n4833), .ZN(n4828) );
  AND2_X1 U5437 ( .A1(n8747), .A2(n10107), .ZN(n5055) );
  NAND2_X1 U5438 ( .A1(n6817), .A2(n4449), .ZN(n8728) );
  NOR2_X1 U5439 ( .A1(n4834), .A2(n6814), .ZN(n4833) );
  INV_X1 U5440 ( .A(n8759), .ZN(n4834) );
  OR2_X1 U5441 ( .A1(n6816), .A2(n6818), .ZN(n8736) );
  AND2_X1 U5442 ( .A1(n6415), .A2(n6805), .ZN(n5063) );
  NAND2_X1 U5443 ( .A1(n8789), .A2(n6265), .ZN(n8774) );
  OR2_X1 U5444 ( .A1(n9050), .A2(n8777), .ZN(n6805) );
  OAI21_X1 U5445 ( .B1(n8801), .B2(n4763), .A(n4761), .ZN(n8789) );
  INV_X1 U5446 ( .A(n4762), .ZN(n4761) );
  OAI21_X1 U5447 ( .B1(n8800), .B2(n4763), .A(n8785), .ZN(n4762) );
  INV_X1 U5448 ( .A(n8786), .ZN(n4763) );
  OAI22_X1 U5449 ( .A1(n8809), .A2(n8810), .B1(n9062), .B2(n8824), .ZN(n8801)
         );
  INV_X1 U5450 ( .A(n8847), .ZN(n5035) );
  OR2_X1 U5451 ( .A1(n5036), .A2(n6223), .ZN(n5033) );
  AND2_X1 U5452 ( .A1(n5037), .A2(n6224), .ZN(n5036) );
  NAND2_X1 U5453 ( .A1(n5038), .A2(n5040), .ZN(n5037) );
  OR2_X1 U5454 ( .A1(n8954), .A2(n7222), .ZN(n8820) );
  NAND2_X1 U5455 ( .A1(n8847), .A2(n8846), .ZN(n8845) );
  NOR2_X1 U5456 ( .A1(n8846), .A2(n4838), .ZN(n4837) );
  INV_X1 U5457 ( .A(n6784), .ZN(n4838) );
  NAND2_X1 U5458 ( .A1(n6198), .A2(n8872), .ZN(n6199) );
  NAND2_X1 U5459 ( .A1(n7293), .A2(n7262), .ZN(n8998) );
  NAND2_X1 U5460 ( .A1(n7293), .A2(n7263), .ZN(n8888) );
  INV_X1 U5461 ( .A(n8998), .ZN(n10107) );
  INV_X1 U5462 ( .A(n8888), .ZN(n10108) );
  NAND2_X1 U5463 ( .A1(n6424), .A2(n6896), .ZN(n10111) );
  INV_X1 U5464 ( .A(n10111), .ZN(n10132) );
  NAND2_X2 U5465 ( .A1(n4816), .A2(n6005), .ZN(n9125) );
  OAI21_X1 U5466 ( .B1(n6363), .B2(n6362), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4641) );
  NAND2_X1 U5467 ( .A1(n4620), .A2(n6335), .ZN(n6353) );
  INV_X1 U5468 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6335) );
  INV_X1 U5469 ( .A(n6337), .ZN(n4620) );
  NOR2_X1 U5470 ( .A1(n6334), .A2(n6333), .ZN(n6338) );
  OAI21_X1 U5471 ( .B1(n7100), .B2(n4436), .A(n7113), .ZN(n4520) );
  INV_X1 U5472 ( .A(n5568), .ZN(n4738) );
  NAND2_X1 U5473 ( .A1(n5128), .A2(n5127), .ZN(n5125) );
  AOI21_X1 U5474 ( .B1(n5130), .B2(n5132), .A(n4497), .ZN(n5127) );
  OR2_X1 U5475 ( .A1(n5798), .A2(n10310), .ZN(n5810) );
  AOI21_X1 U5476 ( .B1(n9269), .B2(n5088), .A(n7088), .ZN(n5087) );
  INV_X1 U5477 ( .A(n9144), .ZN(n5088) );
  INV_X1 U5478 ( .A(n9258), .ZN(n9260) );
  NAND2_X1 U5479 ( .A1(n6926), .A2(n4649), .ZN(n7508) );
  AND2_X1 U5480 ( .A1(n6922), .A2(n6921), .ZN(n4649) );
  OR2_X1 U5481 ( .A1(n5115), .A2(n6991), .ZN(n5111) );
  INV_X1 U5482 ( .A(n6981), .ZN(n4527) );
  AND2_X1 U5483 ( .A1(n7126), .A2(n9923), .ZN(n7122) );
  AND2_X1 U5484 ( .A1(n9509), .A2(n9511), .ZN(n6637) );
  AND2_X1 U5485 ( .A1(n7317), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7289) );
  NAND2_X1 U5486 ( .A1(n9429), .A2(n7365), .ZN(n9438) );
  AND2_X1 U5487 ( .A1(n9438), .A2(n9439), .ZN(n9436) );
  OR2_X1 U5488 ( .A1(n7403), .A2(n4434), .ZN(n4554) );
  NOR2_X1 U5489 ( .A1(n7679), .A2(n4501), .ZN(n7684) );
  NOR2_X1 U5490 ( .A1(n8117), .A2(n4882), .ZN(n8120) );
  AND2_X1 U5491 ( .A1(n8122), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U5492 ( .A1(n4674), .A2(n4673), .ZN(n4892) );
  INV_X1 U5493 ( .A(n9454), .ZN(n4673) );
  OR2_X1 U5494 ( .A1(n9451), .A2(n9450), .ZN(n4730) );
  NAND2_X1 U5495 ( .A1(n4730), .A2(n4729), .ZN(n4614) );
  NAND2_X1 U5496 ( .A1(n9466), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U5497 ( .A1(n9483), .A2(n9484), .ZN(n9487) );
  NAND2_X1 U5498 ( .A1(n4742), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U5499 ( .A1(n6612), .A2(n9553), .ZN(n5159) );
  NAND2_X1 U5500 ( .A1(n6612), .A2(n6611), .ZN(n5160) );
  AOI21_X1 U5501 ( .B1(n5180), .B2(n5177), .A(n4460), .ZN(n5176) );
  INV_X1 U5502 ( .A(n5184), .ZN(n5177) );
  NAND2_X1 U5503 ( .A1(n4741), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5798) );
  AND2_X1 U5504 ( .A1(n6602), .A2(n6607), .ZN(n9575) );
  NAND2_X1 U5505 ( .A1(n9593), .A2(n5079), .ZN(n9581) );
  NOR2_X1 U5506 ( .A1(n5780), .A2(n5185), .ZN(n5184) );
  INV_X1 U5507 ( .A(n5186), .ZN(n5185) );
  OAI21_X1 U5508 ( .B1(n5780), .B2(n5183), .A(n5779), .ZN(n5182) );
  NAND2_X1 U5509 ( .A1(n5766), .A2(n5186), .ZN(n5183) );
  OAI21_X1 U5510 ( .B1(n9628), .B2(n6443), .A(n4961), .ZN(n4952) );
  NAND2_X1 U5511 ( .A1(n4953), .A2(n4955), .ZN(n9574) );
  OR2_X1 U5512 ( .A1(n9629), .A2(n4957), .ZN(n4953) );
  NAND2_X1 U5513 ( .A1(n6524), .A2(n6526), .ZN(n9606) );
  NAND2_X1 U5514 ( .A1(n9645), .A2(n9644), .ZN(n9643) );
  CLKBUF_X1 U5515 ( .A(n9648), .Z(n9649) );
  INV_X1 U5516 ( .A(n6673), .ZN(n4968) );
  OAI21_X1 U5517 ( .B1(n9751), .B2(n5865), .A(n5864), .ZN(n9692) );
  NAND2_X1 U5518 ( .A1(n5867), .A2(n9681), .ZN(n9691) );
  NAND2_X1 U5519 ( .A1(n5202), .A2(n4421), .ZN(n5201) );
  INV_X1 U5520 ( .A(n9716), .ZN(n5202) );
  NAND2_X1 U5521 ( .A1(n4945), .A2(n4943), .ZN(n9751) );
  NOR2_X1 U5522 ( .A1(n9754), .A2(n4944), .ZN(n4943) );
  INV_X1 U5523 ( .A(n6474), .ZN(n4944) );
  NAND2_X1 U5524 ( .A1(n8279), .A2(n8278), .ZN(n4945) );
  AND2_X1 U5525 ( .A1(n5601), .A2(n5600), .ZN(n8282) );
  NAND2_X1 U5526 ( .A1(n9983), .A2(n6473), .ZN(n8279) );
  NAND2_X1 U5527 ( .A1(n4939), .A2(n5851), .ZN(n4941) );
  NOR2_X1 U5528 ( .A1(n6656), .A2(n4940), .ZN(n4939) );
  INV_X1 U5529 ( .A(n6459), .ZN(n4940) );
  OR2_X1 U5530 ( .A1(n5854), .A2(n5855), .ZN(n6658) );
  NAND2_X1 U5531 ( .A1(n6657), .A2(n9980), .ZN(n8230) );
  AND2_X1 U5532 ( .A1(n6465), .A2(n8169), .ZN(n8139) );
  CLKBUF_X1 U5533 ( .A(n8166), .Z(n8167) );
  AND4_X1 U5534 ( .A1(n5559), .A2(n5558), .A3(n5557), .A4(n5556), .ZN(n10039)
         );
  AND2_X1 U5535 ( .A1(n7478), .A2(n8212), .ZN(n9975) );
  NAND2_X1 U5536 ( .A1(n5934), .A2(n6915), .ZN(n8036) );
  NAND2_X1 U5537 ( .A1(n6578), .A2(n8325), .ZN(n7665) );
  INV_X1 U5538 ( .A(n9783), .ZN(n9784) );
  NAND2_X1 U5539 ( .A1(n9775), .A2(n9786), .ZN(n5067) );
  NAND2_X1 U5540 ( .A1(n9782), .A2(n4447), .ZN(n5188) );
  INV_X1 U5541 ( .A(n9577), .ZN(n9797) );
  NAND2_X1 U5542 ( .A1(n5797), .A2(n5796), .ZN(n9808) );
  NAND2_X1 U5543 ( .A1(n5686), .A2(n5685), .ZN(n9869) );
  NAND2_X1 U5544 ( .A1(n7864), .A2(n5923), .ZN(n5686) );
  INV_X1 U5545 ( .A(n10071), .ZN(n10078) );
  NAND2_X1 U5546 ( .A1(n9979), .A2(n10045), .ZN(n10087) );
  INV_X1 U5547 ( .A(n10087), .ZN(n10057) );
  NAND2_X1 U5548 ( .A1(n5891), .A2(n5890), .ZN(n9924) );
  NAND2_X1 U5549 ( .A1(n5212), .A2(n5213), .ZN(n5382) );
  OR2_X2 U5550 ( .A1(n5372), .A2(n5369), .ZN(n5082) );
  NAND2_X1 U5551 ( .A1(n5368), .A2(n5369), .ZN(n4653) );
  NAND2_X1 U5552 ( .A1(n5212), .A2(n4946), .ZN(n5889) );
  NOR2_X1 U5553 ( .A1(n5367), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n4946) );
  XNOR2_X1 U5554 ( .A(n5806), .B(n5807), .ZN(n9126) );
  NAND2_X1 U5555 ( .A1(n5883), .A2(n5369), .ZN(n5149) );
  NAND2_X1 U5556 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5150) );
  AND2_X1 U5557 ( .A1(n5151), .A2(n5883), .ZN(n5146) );
  AND2_X1 U5558 ( .A1(n5882), .A2(n5152), .ZN(n5151) );
  NAND2_X1 U5559 ( .A1(n4865), .A2(n5162), .ZN(n5647) );
  NAND2_X1 U5560 ( .A1(n5170), .A2(n5291), .ZN(n5634) );
  NAND2_X1 U5561 ( .A1(n5166), .A2(n5171), .ZN(n5170) );
  NAND2_X1 U5562 ( .A1(n5135), .A2(n5137), .ZN(n5577) );
  OR2_X1 U5563 ( .A1(n5548), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5564) );
  XNOR2_X1 U5564 ( .A(n5545), .B(n5546), .ZN(n7345) );
  OAI21_X1 U5565 ( .B1(n5526), .B2(n5525), .A(n5273), .ZN(n5545) );
  OR2_X1 U5566 ( .A1(n5532), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5548) );
  AOI21_X1 U5567 ( .B1(n5014), .B2(n5013), .A(n4452), .ZN(n5012) );
  INV_X1 U5568 ( .A(n7767), .ZN(n5013) );
  AND2_X1 U5569 ( .A1(n5014), .A2(n7766), .ZN(n4630) );
  AND4_X1 U5570 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n8887)
         );
  AND2_X1 U5571 ( .A1(n6288), .A2(n6287), .ZN(n8778) );
  NAND2_X1 U5572 ( .A1(n7470), .A2(n7472), .ZN(n7471) );
  NAND2_X1 U5573 ( .A1(n6322), .A2(n6321), .ZN(n7285) );
  AOI21_X1 U5574 ( .B1(n8815), .B2(n6246), .A(n6245), .ZN(n8402) );
  AND2_X1 U5575 ( .A1(n6306), .A2(n6305), .ZN(n8422) );
  AND2_X1 U5576 ( .A1(n7264), .A2(n7263), .ZN(n8533) );
  AND2_X1 U5577 ( .A1(n6238), .A2(n6237), .ZN(n8835) );
  NAND2_X1 U5578 ( .A1(n7254), .A2(n7253), .ZN(n8500) );
  INV_X1 U5579 ( .A(n8739), .ZN(n8762) );
  NAND2_X1 U5580 ( .A1(n7259), .A2(n10122), .ZN(n8524) );
  OR2_X1 U5581 ( .A1(n6858), .A2(n6856), .ZN(n6908) );
  NAND2_X1 U5582 ( .A1(n6330), .A2(n6329), .ZN(n8730) );
  NAND2_X1 U5583 ( .A1(n6318), .A2(n6317), .ZN(n8740) );
  INV_X1 U5584 ( .A(n8422), .ZN(n8747) );
  INV_X1 U5585 ( .A(n8778), .ZN(n8746) );
  INV_X1 U5586 ( .A(n8402), .ZN(n8824) );
  INV_X1 U5587 ( .A(n7222), .ZN(n8849) );
  NAND2_X1 U5588 ( .A1(n6035), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5058) );
  NOR2_X1 U5589 ( .A1(n6711), .A2(n10121), .ZN(n8880) );
  NOR2_X1 U5590 ( .A1(n7158), .A2(n10164), .ZN(n4821) );
  NAND2_X1 U5591 ( .A1(n4823), .A2(n7156), .ZN(n4822) );
  NAND2_X1 U5592 ( .A1(n10157), .A2(n10141), .ZN(n9100) );
  OR2_X1 U5593 ( .A1(n6428), .A2(n7258), .ZN(n6434) );
  NAND2_X1 U5594 ( .A1(n6225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6226) );
  AND4_X1 U5595 ( .A1(n5630), .A2(n5629), .A3(n5628), .A4(n5627), .ZN(n9139)
         );
  NOR2_X1 U5596 ( .A1(n9232), .A2(n5099), .ZN(n5098) );
  INV_X1 U5597 ( .A(n5102), .ZN(n5099) );
  NAND2_X1 U5598 ( .A1(n4472), .A2(n5096), .ZN(n5095) );
  NAND2_X1 U5599 ( .A1(n5102), .A2(n5097), .ZN(n5096) );
  NOR2_X1 U5600 ( .A1(n4432), .A2(n5105), .ZN(n5104) );
  NAND2_X1 U5601 ( .A1(n8265), .A2(n5923), .ZN(n5744) );
  INV_X1 U5602 ( .A(n9825), .ZN(n9613) );
  NAND2_X1 U5603 ( .A1(n8210), .A2(n5923), .ZN(n4585) );
  NAND2_X1 U5604 ( .A1(n5623), .A2(n5622), .ZN(n9902) );
  OAI21_X1 U5605 ( .B1(n6632), .B2(n9507), .A(n4695), .ZN(n6633) );
  NAND2_X1 U5606 ( .A1(n5765), .A2(n5764), .ZN(n9815) );
  OR2_X1 U5607 ( .A1(n9612), .A2(n5872), .ZN(n5765) );
  NOR2_X1 U5608 ( .A1(n7379), .A2(n4431), .ZN(n7382) );
  NOR2_X1 U5609 ( .A1(n4518), .A2(n4403), .ZN(n7378) );
  OR2_X1 U5610 ( .A1(n7674), .A2(n4609), .ZN(n7843) );
  NAND2_X1 U5611 ( .A1(n7675), .A2(n4610), .ZN(n4609) );
  INV_X1 U5612 ( .A(n5219), .ZN(n4610) );
  NOR2_X1 U5613 ( .A1(n7849), .A2(n7850), .ZN(n7982) );
  NAND2_X1 U5614 ( .A1(n7847), .A2(n4552), .ZN(n7849) );
  NAND2_X1 U5615 ( .A1(n7681), .A2(n7682), .ZN(n4552) );
  NOR2_X1 U5616 ( .A1(n7986), .A2(n7985), .ZN(n8117) );
  INV_X1 U5617 ( .A(n4606), .ZN(n4605) );
  NOR2_X1 U5618 ( .A1(n9949), .A2(n9464), .ZN(n9483) );
  NOR2_X1 U5619 ( .A1(n9964), .A2(n4735), .ZN(n4734) );
  NAND2_X1 U5620 ( .A1(n4736), .A2(n9496), .ZN(n4735) );
  NOR2_X1 U5621 ( .A1(n4733), .A2(n4732), .ZN(n4731) );
  INV_X1 U5622 ( .A(n9967), .ZN(n4732) );
  NAND2_X1 U5623 ( .A1(n9960), .A2(n9961), .ZN(n4584) );
  NAND2_X1 U5624 ( .A1(n4886), .A2(n4887), .ZN(n9960) );
  NOR2_X1 U5625 ( .A1(n4406), .A2(n9968), .ZN(n4535) );
  XNOR2_X1 U5626 ( .A(n5955), .B(n6595), .ZN(n9787) );
  NAND2_X1 U5627 ( .A1(n5187), .A2(n4420), .ZN(n5834) );
  NAND2_X1 U5628 ( .A1(n9573), .A2(n6602), .ZN(n9559) );
  NAND2_X2 U5630 ( .A1(n5949), .A2(n9671), .ZN(n9997) );
  AND2_X1 U5631 ( .A1(n4799), .A2(n6866), .ZN(n6747) );
  NAND2_X1 U5632 ( .A1(n4800), .A2(n6736), .ZN(n4799) );
  OR2_X1 U5633 ( .A1(n6759), .A2(n7293), .ZN(n4802) );
  OR2_X1 U5634 ( .A1(n6758), .A2(n4804), .ZN(n4803) );
  NAND2_X1 U5635 ( .A1(n6751), .A2(n7293), .ZN(n4925) );
  AND2_X1 U5636 ( .A1(n4928), .A2(n4926), .ZN(n4924) );
  INV_X1 U5637 ( .A(n6481), .ZN(n4753) );
  AOI21_X1 U5638 ( .B1(n6480), .B2(n6479), .A(n6478), .ZN(n6485) );
  AND2_X1 U5639 ( .A1(n6788), .A2(n4402), .ZN(n4922) );
  AOI21_X1 U5640 ( .B1(n4794), .B2(n4792), .A(n4438), .ZN(n6792) );
  NOR2_X1 U5641 ( .A1(n4793), .A2(n8846), .ZN(n4792) );
  NAND2_X1 U5642 ( .A1(n6796), .A2(n6791), .ZN(n4923) );
  OAI21_X1 U5643 ( .B1(n6490), .B2(n6634), .A(n4680), .ZN(n4662) );
  NOR2_X1 U5644 ( .A1(n4435), .A2(n4681), .ZN(n4680) );
  NOR2_X1 U5645 ( .A1(n6491), .A2(n6630), .ZN(n4681) );
  NAND2_X1 U5646 ( .A1(n6504), .A2(n6512), .ZN(n6509) );
  AND2_X1 U5647 ( .A1(n6515), .A2(n6673), .ZN(n4717) );
  NOR2_X1 U5648 ( .A1(n4548), .A2(n4402), .ZN(n4547) );
  AND2_X1 U5649 ( .A1(n8543), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U5650 ( .A1(n6717), .A2(n6127), .ZN(n4546) );
  AOI21_X1 U5651 ( .B1(n4933), .B2(n4931), .A(n4930), .ZN(n4929) );
  NAND2_X1 U5652 ( .A1(n4936), .A2(n4935), .ZN(n4934) );
  AND2_X1 U5653 ( .A1(n6527), .A2(n6634), .ZN(n4704) );
  OAI21_X1 U5654 ( .B1(n4426), .B2(n4543), .A(n6525), .ZN(n4542) );
  NOR2_X1 U5655 ( .A1(n6532), .A2(n4751), .ZN(n4750) );
  INV_X1 U5656 ( .A(n6531), .ZN(n4751) );
  OR2_X1 U5657 ( .A1(n6443), .A2(n6441), .ZN(n6442) );
  INV_X1 U5658 ( .A(n7224), .ZN(n4626) );
  NAND2_X1 U5659 ( .A1(n8554), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4914) );
  INV_X1 U5660 ( .A(n6817), .ZN(n4826) );
  NAND2_X1 U5661 ( .A1(n10152), .A2(n8552), .ZN(n6742) );
  AND2_X1 U5662 ( .A1(n5978), .A2(n6090), .ZN(n6357) );
  NOR2_X1 U5663 ( .A1(n8230), .A2(n4667), .ZN(n4666) );
  OAI21_X1 U5664 ( .B1(n6530), .B2(n6529), .A(n6531), .ZN(n6535) );
  INV_X1 U5665 ( .A(n4747), .ZN(n4746) );
  OAI21_X1 U5666 ( .B1(n4749), .B2(n4748), .A(n6533), .ZN(n4747) );
  INV_X1 U5667 ( .A(n6529), .ZN(n4748) );
  INV_X1 U5668 ( .A(n4750), .ZN(n4749) );
  NOR2_X1 U5669 ( .A1(n9837), .A2(n9842), .ZN(n6608) );
  INV_X1 U5670 ( .A(n6442), .ZN(n6609) );
  NAND2_X1 U5671 ( .A1(n5200), .A2(n5198), .ZN(n5196) );
  NOR2_X1 U5672 ( .A1(n9665), .A2(n4421), .ZN(n5198) );
  AND3_X1 U5673 ( .A1(n6452), .A2(n6646), .A3(n7869), .ZN(n4962) );
  INV_X1 U5674 ( .A(n5339), .ZN(n4561) );
  INV_X1 U5675 ( .A(n5735), .ZN(n5318) );
  OAI22_X1 U5676 ( .A1(SI_20_), .A2(n5318), .B1(n5319), .B2(SI_21_), .ZN(n5322) );
  NOR2_X1 U5677 ( .A1(n5632), .A2(SI_14_), .ZN(n5167) );
  NAND2_X1 U5678 ( .A1(n5632), .A2(SI_14_), .ZN(n5169) );
  INV_X1 U5679 ( .A(n5167), .ZN(n5163) );
  OAI21_X1 U5680 ( .B1(n7297), .B2(n4635), .A(n4634), .ZN(n5270) );
  NAND2_X1 U5681 ( .A1(n7297), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n4634) );
  OAI21_X1 U5682 ( .B1(n4396), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4709), .ZN(
        n5253) );
  NAND2_X1 U5683 ( .A1(n7297), .A2(n7301), .ZN(n4709) );
  NAND2_X1 U5684 ( .A1(n7297), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4702) );
  OR2_X1 U5685 ( .A1(n7297), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U5686 ( .A1(n8753), .A2(n6881), .ZN(n4876) );
  NAND2_X1 U5687 ( .A1(n4809), .A2(n4808), .ZN(n4807) );
  INV_X1 U5688 ( .A(n6834), .ZN(n4808) );
  INV_X1 U5689 ( .A(n6824), .ZN(n4809) );
  NAND2_X1 U5690 ( .A1(n8554), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4986) );
  OAI22_X1 U5691 ( .A1(n4980), .A2(n8572), .B1(n8260), .B2(n4978), .ZN(n8585)
         );
  OR2_X1 U5692 ( .A1(n8259), .A2(n8572), .ZN(n4978) );
  INV_X1 U5693 ( .A(n4914), .ZN(n4909) );
  NOR2_X1 U5694 ( .A1(n8636), .A2(n10210), .ZN(n4682) );
  INV_X1 U5695 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5959) );
  INV_X1 U5696 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U5697 ( .A1(n9117), .A2(n6844), .ZN(n4549) );
  INV_X1 U5698 ( .A(n6307), .ZN(n4779) );
  INV_X1 U5699 ( .A(n8773), .ZN(n6415) );
  INV_X1 U5700 ( .A(n9056), .ZN(n7227) );
  OR2_X1 U5701 ( .A1(n9062), .A2(n8402), .ZN(n6720) );
  AOI21_X1 U5702 ( .B1(n8163), .B2(n6767), .A(n5060), .ZN(n5059) );
  INV_X1 U5703 ( .A(n6771), .ZN(n5060) );
  AND2_X1 U5704 ( .A1(n6404), .A2(n8148), .ZN(n4706) );
  OR2_X1 U5705 ( .A1(n8900), .A2(n8887), .ZN(n6772) );
  OAI21_X1 U5706 ( .B1(n6342), .B2(n4396), .A(n4812), .ZN(n6039) );
  NOR2_X1 U5707 ( .A1(n4814), .A2(n7297), .ZN(n4813) );
  INV_X1 U5708 ( .A(n6005), .ZN(n4814) );
  INV_X1 U5709 ( .A(n6745), .ZN(n4707) );
  NAND2_X1 U5710 ( .A1(n6723), .A2(n4836), .ZN(n6862) );
  INV_X1 U5711 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5980) );
  INV_X1 U5712 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5979) );
  INV_X1 U5713 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5982) );
  NOR2_X1 U5714 ( .A1(n6000), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5986) );
  INV_X1 U5715 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6332) );
  OR2_X1 U5716 ( .A1(n6092), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6114) );
  NOR2_X1 U5717 ( .A1(n5089), .A2(n5086), .ZN(n5085) );
  INV_X1 U5718 ( .A(n9145), .ZN(n5086) );
  INV_X1 U5719 ( .A(n9269), .ZN(n5089) );
  AOI21_X1 U5720 ( .B1(n5119), .B2(n5121), .A(n4458), .ZN(n5118) );
  AND2_X1 U5721 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5452) );
  NAND2_X1 U5722 ( .A1(n5160), .A2(n5159), .ZN(n5155) );
  NOR2_X1 U5723 ( .A1(n5158), .A2(n5833), .ZN(n5157) );
  INV_X1 U5724 ( .A(n5159), .ZN(n5158) );
  AND2_X1 U5725 ( .A1(n5176), .A2(n4439), .ZN(n5173) );
  OR2_X1 U5726 ( .A1(n9808), .A2(n9797), .ZN(n6605) );
  NOR2_X1 U5727 ( .A1(n5771), .A2(n9147), .ZN(n4741) );
  NAND2_X1 U5728 ( .A1(n4951), .A2(n4949), .ZN(n4948) );
  NOR2_X1 U5729 ( .A1(n4958), .A2(n4956), .ZN(n4949) );
  NAND2_X1 U5730 ( .A1(n5071), .A2(n5070), .ZN(n5069) );
  OR2_X1 U5731 ( .A1(n5860), .A2(n9873), .ZN(n6575) );
  NAND2_X1 U5732 ( .A1(n4740), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5655) );
  AND2_X1 U5733 ( .A1(n6586), .A2(n9731), .ZN(n9698) );
  NOR2_X2 U5734 ( .A1(n5625), .A2(n5624), .ZN(n4740) );
  INV_X1 U5735 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5602) );
  INV_X1 U5736 ( .A(n8175), .ZN(n5066) );
  NAND2_X1 U5737 ( .A1(n9390), .A2(n10006), .ZN(n6447) );
  NAND2_X1 U5738 ( .A1(n9212), .A2(n9342), .ZN(n6646) );
  NAND2_X1 U5739 ( .A1(n5407), .A2(n6929), .ZN(n6648) );
  OR2_X1 U5740 ( .A1(n5929), .A2(n5928), .ZN(n7116) );
  INV_X1 U5741 ( .A(n9924), .ZN(n5902) );
  NOR2_X1 U5742 ( .A1(n9759), .A2(n9902), .ZN(n9758) );
  OR2_X1 U5743 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  NAND2_X1 U5744 ( .A1(n5324), .A2(n5323), .ZN(n5327) );
  AND2_X1 U5745 ( .A1(n4860), .A2(n4858), .ZN(n4857) );
  INV_X1 U5746 ( .A(n5755), .ZN(n4858) );
  NOR2_X1 U5747 ( .A1(n5322), .A2(n4864), .ZN(n4863) );
  INV_X1 U5748 ( .A(n5315), .ZN(n4864) );
  NAND2_X1 U5749 ( .A1(n5315), .A2(n5314), .ZN(n5713) );
  INV_X1 U5750 ( .A(n5280), .ZN(n5136) );
  NAND2_X1 U5751 ( .A1(n5253), .A2(n10211), .ZN(n5473) );
  NAND2_X1 U5752 ( .A1(n4600), .A2(n4721), .ZN(n5397) );
  NAND2_X1 U5753 ( .A1(n4849), .A2(n5246), .ZN(n5402) );
  INV_X1 U5754 ( .A(SI_11_), .ZN(n10414) );
  INV_X1 U5755 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5537) );
  OAI21_X1 U5756 ( .B1(n8518), .B2(n8747), .A(n8516), .ZN(n7245) );
  AOI22_X1 U5757 ( .A1(n8476), .A2(n7207), .B1(n7206), .B2(n8545), .ZN(n8353)
         );
  XNOR2_X1 U5758 ( .A(n7170), .B(n6398), .ZN(n7171) );
  INV_X1 U5759 ( .A(n10136), .ZN(n4836) );
  OR2_X1 U5760 ( .A1(n7226), .A2(n8824), .ZN(n5224) );
  INV_X1 U5761 ( .A(n7236), .ZN(n5011) );
  AND2_X1 U5762 ( .A1(n5023), .A2(n7210), .ZN(n5022) );
  XNOR2_X1 U5763 ( .A(n6416), .B(n7174), .ZN(n8443) );
  OR2_X1 U5764 ( .A1(n7223), .A2(n8835), .ZN(n7224) );
  OR2_X1 U5765 ( .A1(n8466), .A2(n8467), .ZN(n8464) );
  AOI21_X1 U5766 ( .B1(n5006), .B2(n5004), .A(n4446), .ZN(n5003) );
  INV_X1 U5767 ( .A(n5006), .ZN(n5005) );
  NOR2_X1 U5768 ( .A1(n5022), .A2(n8434), .ZN(n5018) );
  NOR2_X1 U5769 ( .A1(n7218), .A2(n5041), .ZN(n5017) );
  NAND2_X1 U5770 ( .A1(n4473), .A2(n5023), .ZN(n5021) );
  XNOR2_X1 U5771 ( .A(n7732), .B(n7249), .ZN(n7183) );
  NAND2_X1 U5772 ( .A1(n7765), .A2(n7766), .ZN(n7180) );
  NAND2_X1 U5773 ( .A1(n8418), .A2(n8419), .ZN(n8517) );
  NAND2_X1 U5774 ( .A1(n7211), .A2(n7210), .ZN(n8527) );
  AND2_X1 U5775 ( .A1(n6432), .A2(n6431), .ZN(n7274) );
  NAND2_X1 U5776 ( .A1(n6343), .A2(n6246), .ZN(n6852) );
  INV_X1 U5777 ( .A(n6847), .ZN(n6830) );
  INV_X1 U5778 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6018) );
  XNOR2_X1 U5779 ( .A(n4395), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n7578) );
  NAND2_X1 U5780 ( .A1(n7424), .A2(n7423), .ZN(n7577) );
  XNOR2_X1 U5781 ( .A(n7425), .B(n4644), .ZN(n7496) );
  CLKBUF_X1 U5782 ( .A(n7442), .Z(n7443) );
  OAI22_X1 U5783 ( .A1(n7496), .A2(n7426), .B1(n4644), .B2(n7425), .ZN(n7427)
         );
  AND2_X1 U5784 ( .A1(n4970), .A2(n7561), .ZN(n5233) );
  NAND2_X1 U5785 ( .A1(n7558), .A2(n7633), .ZN(n7561) );
  NAND3_X1 U5786 ( .A1(n4970), .A2(P2_REG2_REG_5__SCAN_IN), .A3(n7561), .ZN(
        n7629) );
  OAI21_X1 U5787 ( .B1(n7628), .B2(n7554), .A(n4906), .ZN(n7602) );
  NAND2_X1 U5788 ( .A1(n7552), .A2(n7633), .ZN(n4906) );
  AOI21_X1 U5789 ( .B1(n7602), .B2(n7601), .A(n4905), .ZN(n7638) );
  NOR2_X1 U5790 ( .A1(n7604), .A2(n7727), .ZN(n4905) );
  NAND2_X1 U5791 ( .A1(n7606), .A2(n7605), .ZN(n4975) );
  NAND2_X1 U5792 ( .A1(n7646), .A2(n7645), .ZN(n7813) );
  OAI21_X1 U5793 ( .B1(n7796), .B2(n7795), .A(n4645), .ZN(n7909) );
  OR2_X1 U5794 ( .A1(n7794), .A2(n10293), .ZN(n4645) );
  NAND2_X1 U5795 ( .A1(n7925), .A2(n7924), .ZN(n8199) );
  OR2_X1 U5796 ( .A1(n6156), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U5797 ( .A1(n8250), .A2(n8249), .ZN(n8562) );
  NAND2_X1 U5798 ( .A1(n4910), .A2(n4908), .ZN(n8571) );
  OR2_X1 U5799 ( .A1(n4911), .A2(n4909), .ZN(n4908) );
  NAND2_X1 U5800 ( .A1(n8242), .A2(n4500), .ZN(n4910) );
  AND2_X1 U5801 ( .A1(n8553), .A2(n4496), .ZN(n4911) );
  NAND2_X1 U5802 ( .A1(n8578), .A2(n8577), .ZN(n8608) );
  NOR2_X1 U5803 ( .A1(n8587), .A2(n8966), .ZN(n4638) );
  AOI21_X1 U5804 ( .B1(n8645), .B2(n8644), .A(n4513), .ZN(n8663) );
  NAND2_X1 U5805 ( .A1(n8627), .A2(n8626), .ZN(n8654) );
  NAND2_X1 U5806 ( .A1(n6281), .A2(n4499), .ZN(n6312) );
  AND2_X1 U5807 ( .A1(n4784), .A2(n6275), .ZN(n8760) );
  INV_X1 U5808 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U5809 ( .A1(n6231), .A2(n4874), .ZN(n6249) );
  NAND2_X1 U5810 ( .A1(n6231), .A2(n6230), .ZN(n6241) );
  AND2_X1 U5811 ( .A1(n6215), .A2(n6214), .ZN(n7219) );
  NAND2_X1 U5812 ( .A1(n5969), .A2(n4414), .ZN(n6216) );
  INV_X1 U5813 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4870) );
  OR2_X1 U5814 ( .A1(n6179), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U5815 ( .A1(n5967), .A2(n5966), .ZN(n6179) );
  INV_X1 U5816 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5966) );
  INV_X1 U5817 ( .A(n6169), .ZN(n5967) );
  AND2_X1 U5818 ( .A1(n6763), .A2(n6764), .ZN(n8148) );
  NAND2_X1 U5819 ( .A1(n5963), .A2(n4455), .ZN(n6160) );
  NAND2_X1 U5820 ( .A1(n5963), .A2(n4878), .ZN(n6148) );
  INV_X1 U5821 ( .A(n8546), .ZN(n8412) );
  AND2_X1 U5822 ( .A1(n4767), .A2(n6113), .ZN(n4766) );
  NAND2_X1 U5823 ( .A1(n5963), .A2(n5962), .ZN(n6134) );
  OR2_X1 U5824 ( .A1(n6106), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6119) );
  NAND4_X1 U5825 ( .A1(n6018), .A2(n5959), .A3(n5958), .A4(n4880), .ZN(n6096)
         );
  INV_X1 U5826 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U5827 ( .A1(n5961), .A2(n5960), .ZN(n6106) );
  INV_X1 U5828 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5960) );
  INV_X1 U5829 ( .A(n6096), .ZN(n5961) );
  NAND2_X1 U5830 ( .A1(n5047), .A2(n6089), .ZN(n7825) );
  NAND2_X1 U5831 ( .A1(n6018), .A2(n5958), .ZN(n6070) );
  AOI22_X1 U5832 ( .A1(n8996), .A2(n10140), .B1(n6397), .B2(n9004), .ZN(n6049)
         );
  NAND2_X1 U5833 ( .A1(n8999), .A2(n9007), .ZN(n8987) );
  AND2_X1 U5834 ( .A1(n7736), .A2(n6420), .ZN(n8990) );
  OR2_X1 U5835 ( .A1(n6705), .A2(n6704), .ZN(n6711) );
  INV_X1 U5836 ( .A(n7285), .ZN(n7147) );
  AND2_X1 U5837 ( .A1(n4781), .A2(n4785), .ZN(n4780) );
  NAND2_X1 U5838 ( .A1(n4790), .A2(n4410), .ZN(n4785) );
  NAND2_X1 U5839 ( .A1(n4786), .A2(n4782), .ZN(n4781) );
  INV_X1 U5840 ( .A(n8736), .ZN(n8738) );
  INV_X1 U5841 ( .A(n4786), .ZN(n4783) );
  NAND2_X1 U5842 ( .A1(n8801), .A2(n8800), .ZN(n8799) );
  AOI21_X1 U5843 ( .B1(n5031), .B2(n5030), .A(n4461), .ZN(n5029) );
  NAND2_X1 U5844 ( .A1(n5031), .A2(n8847), .ZN(n5028) );
  NAND2_X1 U5845 ( .A1(n8857), .A2(n8858), .ZN(n8863) );
  AND3_X1 U5846 ( .A1(n6197), .A2(n6196), .A3(n6195), .ZN(n8889) );
  AND2_X1 U5847 ( .A1(n4775), .A2(n4771), .ZN(n4770) );
  NAND2_X1 U5848 ( .A1(n4401), .A2(n4404), .ZN(n4775) );
  NAND2_X1 U5849 ( .A1(n7827), .A2(n6102), .ZN(n7884) );
  AND2_X1 U5850 ( .A1(n7274), .A2(n7333), .ZN(n7261) );
  NAND2_X1 U5851 ( .A1(n7945), .A2(n10153), .ZN(n10149) );
  XNOR2_X1 U5852 ( .A(n6336), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6910) );
  INV_X1 U5853 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6331) );
  XNOR2_X1 U5854 ( .A(n6058), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7555) );
  INV_X1 U5855 ( .A(n6930), .ZN(n4675) );
  NAND2_X1 U5856 ( .A1(n9258), .A2(n5380), .ZN(n5719) );
  INV_X1 U5857 ( .A(n4677), .ZN(n5726) );
  AND2_X1 U5858 ( .A1(n7109), .A2(n7108), .ZN(n9192) );
  OR2_X1 U5859 ( .A1(n5107), .A2(n7114), .ZN(n5101) );
  AND2_X1 U5860 ( .A1(n7114), .A2(n5106), .ZN(n5102) );
  AND2_X1 U5861 ( .A1(n9193), .A2(n9359), .ZN(n5106) );
  NAND2_X1 U5862 ( .A1(n5117), .A2(n5119), .ZN(n9196) );
  OR2_X1 U5863 ( .A1(n6961), .A2(n5121), .ZN(n5117) );
  AND2_X1 U5864 ( .A1(n6919), .A2(n6918), .ZN(n6920) );
  INV_X1 U5865 ( .A(n9388), .ZN(n8108) );
  NAND2_X1 U5866 ( .A1(n5379), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5673) );
  INV_X1 U5867 ( .A(n5655), .ZN(n5379) );
  OR2_X1 U5868 ( .A1(n5538), .A2(n5537), .ZN(n5553) );
  NAND2_X1 U5869 ( .A1(n5378), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5568) );
  INV_X1 U5870 ( .A(n5553), .ZN(n5378) );
  NAND2_X1 U5871 ( .A1(n5133), .A2(n7053), .ZN(n5132) );
  INV_X1 U5872 ( .A(n7049), .ZN(n5133) );
  OR2_X1 U5873 ( .A1(n5746), .A2(n5745), .ZN(n5759) );
  NAND2_X1 U5874 ( .A1(n5381), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5771) );
  INV_X1 U5875 ( .A(n5759), .ZN(n5381) );
  NAND2_X1 U5876 ( .A1(n5452), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U5877 ( .A1(n5376), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5505) );
  INV_X1 U5878 ( .A(n5493), .ZN(n5376) );
  AND2_X1 U5879 ( .A1(n9766), .A2(n6574), .ZN(n6629) );
  OR3_X1 U5880 ( .A1(n9772), .A2(n6574), .A3(n9382), .ZN(n5222) );
  NAND2_X1 U5881 ( .A1(n6568), .A2(n9766), .ZN(n6572) );
  AND2_X1 U5882 ( .A1(n6689), .A2(n4696), .ZN(n4695) );
  AOI21_X1 U5883 ( .B1(n9507), .B2(n6634), .A(n4697), .ZN(n4696) );
  INV_X1 U5884 ( .A(n6631), .ZN(n4697) );
  AND2_X1 U5885 ( .A1(n9766), .A2(n9382), .ZN(n4698) );
  NAND2_X1 U5886 ( .A1(n9772), .A2(n6634), .ZN(n4845) );
  INV_X1 U5887 ( .A(n6629), .ZN(n6686) );
  NAND2_X1 U5888 ( .A1(n9441), .A2(n9442), .ZN(n9440) );
  NAND2_X1 U5889 ( .A1(n7684), .A2(n7683), .ZN(n7847) );
  NAND2_X1 U5890 ( .A1(n8120), .A2(n8119), .ZN(n8296) );
  NAND2_X1 U5891 ( .A1(n4608), .A2(n4607), .ZN(n4606) );
  INV_X1 U5892 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n4607) );
  NOR2_X1 U5893 ( .A1(n4890), .A2(n9954), .ZN(n4889) );
  NAND2_X1 U5894 ( .A1(n4617), .A2(n4615), .ZN(n9480) );
  NOR2_X1 U5895 ( .A1(n4616), .A2(n9478), .ZN(n4615) );
  OR2_X1 U5896 ( .A1(n4685), .A2(n9468), .ZN(n4617) );
  NAND2_X1 U5897 ( .A1(n9494), .A2(n4511), .ZN(n9962) );
  INV_X1 U5898 ( .A(n9966), .ZN(n4599) );
  NAND2_X1 U5899 ( .A1(n9494), .A2(n9493), .ZN(n9965) );
  AOI21_X1 U5900 ( .B1(n9497), .B2(n4888), .A(n4512), .ZN(n4887) );
  INV_X1 U5901 ( .A(n9486), .ZN(n4888) );
  NAND2_X1 U5902 ( .A1(n4532), .A2(n9497), .ZN(n4886) );
  INV_X1 U5903 ( .A(n9487), .ZN(n4532) );
  INV_X1 U5904 ( .A(n9766), .ZN(n9509) );
  INV_X1 U5905 ( .A(n5869), .ZN(n6594) );
  NAND2_X1 U5906 ( .A1(n6617), .A2(n6440), .ZN(n5869) );
  AND2_X1 U5907 ( .A1(n5390), .A2(n5389), .ZN(n9777) );
  AND2_X1 U5908 ( .A1(n5825), .A2(n5811), .ZN(n9548) );
  INV_X1 U5909 ( .A(n5180), .ZN(n5178) );
  NAND2_X1 U5910 ( .A1(n9593), .A2(n9819), .ZN(n9594) );
  NOR2_X1 U5911 ( .A1(n5075), .A2(n9837), .ZN(n5074) );
  INV_X1 U5912 ( .A(n5076), .ZN(n5075) );
  INV_X1 U5913 ( .A(n5208), .ZN(n5207) );
  OAI21_X1 U5914 ( .B1(n5734), .B2(n5209), .A(n5733), .ZN(n5208) );
  NAND2_X1 U5915 ( .A1(n9670), .A2(n5076), .ZN(n9621) );
  NAND2_X1 U5916 ( .A1(n4967), .A2(n4590), .ZN(n4589) );
  NAND2_X1 U5917 ( .A1(n4588), .A2(n4590), .ZN(n4587) );
  INV_X1 U5918 ( .A(n9650), .ZN(n4590) );
  NAND2_X1 U5919 ( .A1(n9670), .A2(n9854), .ZN(n9633) );
  AND2_X1 U5920 ( .A1(n9663), .A2(n9664), .ZN(n9682) );
  AND2_X1 U5921 ( .A1(n5680), .A2(n5661), .ZN(n5200) );
  AND2_X1 U5922 ( .A1(n6671), .A2(n6487), .ZN(n9702) );
  INV_X1 U5923 ( .A(n9702), .ZN(n5680) );
  INV_X1 U5924 ( .A(n9759), .ZN(n5068) );
  OR2_X1 U5925 ( .A1(n9746), .A2(n9756), .ZN(n9717) );
  NAND2_X1 U5926 ( .A1(n5646), .A2(n5645), .ZN(n9716) );
  AND2_X1 U5927 ( .A1(n5631), .A2(n4492), .ZN(n5203) );
  AND2_X1 U5928 ( .A1(n6575), .A2(n9700), .ZN(n9719) );
  NAND2_X1 U5929 ( .A1(n9750), .A2(n9754), .ZN(n5204) );
  INV_X1 U5930 ( .A(n4740), .ZN(n5639) );
  NAND2_X1 U5931 ( .A1(n8235), .A2(n5065), .ZN(n5064) );
  AOI21_X1 U5932 ( .B1(n5192), .B2(n5194), .A(n4459), .ZN(n5190) );
  AND4_X1 U5933 ( .A1(n5510), .A2(n5509), .A3(n5508), .A4(n5507), .ZN(n10040)
         );
  CLKBUF_X1 U5934 ( .A(n7866), .Z(n7867) );
  INV_X1 U5935 ( .A(n4725), .ZN(n4758) );
  OR2_X1 U5936 ( .A1(n9536), .A2(n5872), .ZN(n5832) );
  NAND2_X1 U5937 ( .A1(n5809), .A2(n5808), .ZN(n9801) );
  NAND2_X1 U5938 ( .A1(n5784), .A2(n5783), .ZN(n9812) );
  OR2_X1 U5939 ( .A1(n6634), .A2(n4530), .ZN(n10045) );
  INV_X1 U5940 ( .A(n8113), .ZN(n10033) );
  AND4_X2 U5941 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n10011)
         );
  OR2_X1 U5942 ( .A1(n6565), .A2(n7301), .ZN(n5476) );
  AND2_X1 U5943 ( .A1(n7115), .A2(n5912), .ZN(n5930) );
  AND3_X1 U5944 ( .A1(n5928), .A2(n5927), .A3(n5932), .ZN(n5913) );
  AND2_X1 U5945 ( .A1(n8273), .A2(n8269), .ZN(n7478) );
  NOR2_X1 U5946 ( .A1(n5215), .A2(n5369), .ZN(n4719) );
  INV_X1 U5947 ( .A(n5843), .ZN(n4597) );
  NAND2_X1 U5948 ( .A1(n4471), .A2(n5844), .ZN(n4760) );
  AND2_X1 U5949 ( .A1(n5333), .A2(n5332), .ZN(n5768) );
  AOI21_X1 U5950 ( .B1(n4857), .B2(n4855), .A(n4854), .ZN(n4853) );
  INV_X1 U5951 ( .A(n5327), .ZN(n4854) );
  INV_X1 U5952 ( .A(n4863), .ZN(n4855) );
  INV_X1 U5953 ( .A(n4857), .ZN(n4856) );
  NAND2_X1 U5954 ( .A1(n4575), .A2(n4573), .ZN(n4578) );
  INV_X1 U5955 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U5956 ( .A1(n5838), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U5957 ( .A1(n4579), .A2(n5299), .ZN(n5682) );
  XNOR2_X1 U5958 ( .A(n5616), .B(n5615), .ZN(n7512) );
  AOI21_X1 U5959 ( .B1(n5141), .B2(n5144), .A(n5560), .ZN(n5139) );
  INV_X1 U5960 ( .A(n5141), .ZN(n5140) );
  NAND2_X1 U5961 ( .A1(n5526), .A2(n5143), .ZN(n5138) );
  XNOR2_X1 U5962 ( .A(n5487), .B(n5486), .ZN(n7312) );
  XNOR2_X1 U5963 ( .A(n5481), .B(n5448), .ZN(n5449) );
  INV_X1 U5964 ( .A(n5480), .ZN(n5448) );
  NAND2_X1 U5965 ( .A1(n5396), .A2(n5363), .ZN(n5466) );
  INV_X1 U5966 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U5967 ( .A1(n5397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5434) );
  INV_X1 U5968 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10344) );
  INV_X1 U5969 ( .A(n8983), .ZN(n8370) );
  AND2_X1 U5970 ( .A1(n7535), .A2(n7173), .ZN(n5000) );
  NAND2_X1 U5971 ( .A1(n8378), .A2(n8377), .ZN(n8376) );
  NAND2_X1 U5972 ( .A1(n4678), .A2(n7168), .ZN(n7481) );
  NAND2_X1 U5973 ( .A1(n8464), .A2(n5224), .ZN(n8398) );
  OAI21_X1 U5974 ( .B1(n7233), .B2(n5009), .A(n5007), .ZN(n8418) );
  INV_X1 U5975 ( .A(n5010), .ZN(n5009) );
  AOI21_X1 U5976 ( .B1(n5010), .B2(n8483), .A(n5008), .ZN(n5007) );
  NOR2_X1 U5977 ( .A1(n7241), .A2(n5011), .ZN(n5010) );
  AND3_X1 U5978 ( .A1(n6209), .A2(n6208), .A3(n6207), .ZN(n8878) );
  NAND2_X1 U5979 ( .A1(n5015), .A2(n5021), .ZN(n8435) );
  NAND2_X1 U5980 ( .A1(n7211), .A2(n5022), .ZN(n5015) );
  NAND2_X1 U5981 ( .A1(n8388), .A2(n5006), .ZN(n8216) );
  INV_X1 U5982 ( .A(n8533), .ZN(n8489) );
  NAND2_X1 U5983 ( .A1(n8376), .A2(n7224), .ZN(n8466) );
  OAI21_X1 U5984 ( .B1(n7211), .B2(n5019), .A(n5016), .ZN(n8510) );
  NAND2_X1 U5985 ( .A1(n5021), .A2(n5020), .ZN(n5019) );
  AOI21_X1 U5986 ( .B1(n5018), .B2(n5021), .A(n5017), .ZN(n5016) );
  INV_X1 U5987 ( .A(n8434), .ZN(n5020) );
  NAND2_X1 U5988 ( .A1(n5014), .A2(n7769), .ZN(n7834) );
  INV_X1 U5989 ( .A(n8524), .ZN(n8541) );
  NAND2_X1 U5990 ( .A1(n6297), .A2(n6296), .ZN(n8739) );
  NAND2_X1 U5991 ( .A1(n6274), .A2(n6273), .ZN(n8790) );
  INV_X1 U5992 ( .A(n8777), .ZN(n8802) );
  OAI21_X1 U5993 ( .B1(n7588), .B2(n7587), .A(n7452), .ZN(n7572) );
  XNOR2_X1 U5994 ( .A(n7552), .B(n7633), .ZN(n7628) );
  XNOR2_X1 U5995 ( .A(n7638), .B(n7640), .ZN(n7641) );
  AND2_X1 U5996 ( .A1(n4976), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U5997 ( .A1(n4988), .A2(n7914), .ZN(n7916) );
  INV_X1 U5998 ( .A(n4989), .ZN(n4988) );
  AND2_X1 U5999 ( .A1(n7802), .A2(n7914), .ZN(n5232) );
  XNOR2_X1 U6000 ( .A(n7909), .B(n7806), .ZN(n7912) );
  NAND2_X1 U6001 ( .A1(n8260), .A2(n5231), .ZN(n4979) );
  NAND2_X1 U6002 ( .A1(n8242), .A2(n4913), .ZN(n4912) );
  XNOR2_X1 U6003 ( .A(n8571), .B(n8572), .ZN(n8574) );
  OAI22_X1 U6004 ( .A1(n8574), .A2(n8573), .B1(n8572), .B2(n8571), .ZN(n8596)
         );
  XNOR2_X1 U6005 ( .A(n8617), .B(n8618), .ZN(n8619) );
  OAI21_X1 U6006 ( .B1(n8619), .B2(n8961), .A(n4896), .ZN(n8645) );
  NAND2_X1 U6007 ( .A1(n4898), .A2(n4897), .ZN(n4896) );
  INV_X1 U6008 ( .A(n8617), .ZN(n4898) );
  XNOR2_X1 U6009 ( .A(n8663), .B(n4895), .ZN(n8665) );
  OR2_X1 U6010 ( .A1(n6710), .A2(n8883), .ZN(n6715) );
  AND2_X1 U6011 ( .A1(n6279), .A2(n6278), .ZN(n8757) );
  OAI21_X1 U6012 ( .B1(n4691), .B2(n10132), .A(n4689), .ZN(n8939) );
  INV_X1 U6013 ( .A(n4690), .ZN(n4689) );
  XNOR2_X1 U6014 ( .A(n8760), .B(n8767), .ZN(n4691) );
  OAI22_X1 U6015 ( .A1(n8762), .A2(n8888), .B1(n8998), .B2(n8761), .ZN(n4690)
         );
  NAND2_X1 U6016 ( .A1(n8845), .A2(n5040), .ZN(n8833) );
  OR2_X1 U6017 ( .A1(n8151), .A2(n6155), .ZN(n5027) );
  NAND2_X1 U6018 ( .A1(n6147), .A2(n6146), .ZN(n8494) );
  NAND2_X1 U6019 ( .A1(n6118), .A2(n6117), .ZN(n8044) );
  NAND2_X1 U6020 ( .A1(n5062), .A2(n6749), .ZN(n7822) );
  NAND2_X1 U6021 ( .A1(n7333), .A2(n6707), .ZN(n10122) );
  INV_X1 U6022 ( .A(n10122), .ZN(n8924) );
  NOR2_X1 U6023 ( .A1(n10166), .A2(n8933), .ZN(n5053) );
  NAND2_X1 U6024 ( .A1(n6192), .A2(n6191), .ZN(n8963) );
  INV_X1 U6025 ( .A(n6894), .ZN(n9015) );
  INV_X1 U6026 ( .A(n6890), .ZN(n9018) );
  NOR2_X1 U6027 ( .A1(n6350), .A2(n6349), .ZN(n6351) );
  NOR2_X1 U6028 ( .A1(n7280), .A2(n8998), .ZN(n6349) );
  OAI21_X1 U6029 ( .B1(n4637), .B2(n4829), .A(n4827), .ZN(n8727) );
  AOI21_X1 U6030 ( .B1(n5049), .B2(n10111), .A(n5048), .ZN(n9019) );
  INV_X1 U6031 ( .A(n5054), .ZN(n5048) );
  AOI21_X1 U6032 ( .B1(n8730), .B2(n10108), .A(n5055), .ZN(n5054) );
  NAND2_X1 U6033 ( .A1(n6299), .A2(n6298), .ZN(n9027) );
  NAND2_X1 U6034 ( .A1(n4832), .A2(n6813), .ZN(n8735) );
  NAND2_X1 U6035 ( .A1(n4637), .A2(n4833), .ZN(n4832) );
  NAND2_X1 U6036 ( .A1(n6290), .A2(n6289), .ZN(n9033) );
  NAND2_X1 U6037 ( .A1(n4637), .A2(n8759), .ZN(n8752) );
  NAND2_X1 U6038 ( .A1(n4784), .A2(n4788), .ZN(n4791) );
  INV_X1 U6039 ( .A(n8757), .ZN(n9039) );
  INV_X1 U6040 ( .A(n6416), .ZN(n9044) );
  NAND2_X1 U6041 ( .A1(n6414), .A2(n6805), .ZN(n8770) );
  NAND2_X1 U6042 ( .A1(n6257), .A2(n6256), .ZN(n9050) );
  NAND2_X1 U6043 ( .A1(n5034), .A2(n5033), .ZN(n8822) );
  NAND2_X1 U6044 ( .A1(n5035), .A2(n4422), .ZN(n5034) );
  NAND2_X1 U6045 ( .A1(n8843), .A2(n6790), .ZN(n8830) );
  NAND2_X1 U6046 ( .A1(n6203), .A2(n6202), .ZN(n9083) );
  NAND2_X1 U6047 ( .A1(n6178), .A2(n6177), .ZN(n9093) );
  NAND2_X1 U6048 ( .A1(n8161), .A2(n6767), .ZN(n8910) );
  INV_X1 U6049 ( .A(n9100), .ZN(n9094) );
  NAND2_X1 U6050 ( .A1(n6076), .A2(n6868), .ZN(n7725) );
  NAND2_X1 U6051 ( .A1(n9110), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5993) );
  INV_X2 U6052 ( .A(n5994), .ZN(n9118) );
  NAND2_X1 U6053 ( .A1(n4640), .A2(n4639), .ZN(n6365) );
  NAND2_X1 U6054 ( .A1(n5974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4639) );
  NOR2_X1 U6055 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4619) );
  INV_X1 U6056 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10438) );
  XNOR2_X1 U6057 ( .A(n6341), .B(n6340), .ZN(n8215) );
  NAND2_X1 U6058 ( .A1(n6339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6341) );
  INV_X1 U6059 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8208) );
  INV_X1 U6060 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7956) );
  INV_X1 U6061 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7907) );
  INV_X1 U6062 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7780) );
  INV_X1 U6063 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10440) );
  INV_X1 U6064 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6024) );
  INV_X1 U6065 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5239) );
  OAI21_X1 U6066 ( .B1(n9232), .B2(n4436), .A(n4519), .ZN(n4524) );
  INV_X1 U6067 ( .A(n4520), .ZN(n4519) );
  OR2_X1 U6068 ( .A1(n4720), .A2(n7049), .ZN(n5129) );
  NOR2_X1 U6069 ( .A1(n5123), .A2(n9299), .ZN(n9217) );
  INV_X1 U6070 ( .A(n5125), .ZN(n5123) );
  AND4_X1 U6071 ( .A1(n5589), .A2(n5588), .A3(n5587), .A4(n5586), .ZN(n10083)
         );
  NAND2_X1 U6072 ( .A1(n5113), .A2(n5116), .ZN(n9225) );
  INV_X1 U6073 ( .A(n5115), .ZN(n5116) );
  INV_X1 U6074 ( .A(n8282), .ZN(n10079) );
  INV_X1 U6075 ( .A(n9869), .ZN(n5866) );
  NAND2_X1 U6076 ( .A1(n9268), .A2(n9269), .ZN(n9267) );
  NAND2_X1 U6077 ( .A1(n5090), .A2(n9144), .ZN(n9268) );
  NAND2_X1 U6078 ( .A1(n5126), .A2(n5130), .ZN(n9301) );
  OR2_X1 U6079 ( .A1(n4720), .A2(n5132), .ZN(n5126) );
  AOI21_X1 U6080 ( .B1(n5114), .B2(n4527), .A(n4444), .ZN(n4526) );
  INV_X1 U6081 ( .A(n5114), .ZN(n4525) );
  AND4_X1 U6082 ( .A1(n5573), .A2(n5572), .A3(n5571), .A4(n5570), .ZN(n9331)
         );
  OR2_X1 U6083 ( .A1(n7125), .A2(n7124), .ZN(n9349) );
  AND2_X1 U6084 ( .A1(n6951), .A2(n6950), .ZN(n6952) );
  INV_X1 U6085 ( .A(n9350), .ZN(n9373) );
  AND2_X1 U6086 ( .A1(n7122), .A2(n7121), .ZN(n9365) );
  NAND2_X1 U6087 ( .A1(n9232), .A2(n7100), .ZN(n9358) );
  AND2_X1 U6088 ( .A1(n7122), .A2(n7127), .ZN(n9359) );
  AND3_X1 U6089 ( .A1(n5679), .A2(n5678), .A3(n5677), .ZN(n9725) );
  INV_X1 U6090 ( .A(n9359), .ZN(n9380) );
  OR3_X1 U6091 ( .A1(n5943), .A2(n5872), .A3(n9186), .ZN(n5878) );
  INV_X1 U6092 ( .A(n9798), .ZN(n9384) );
  INV_X1 U6093 ( .A(n9562), .ZN(n9788) );
  NAND2_X1 U6094 ( .A1(n5804), .A2(n5803), .ZN(n9577) );
  OR2_X1 U6095 ( .A1(n9564), .A2(n5872), .ZN(n5804) );
  NAND2_X1 U6096 ( .A1(n5792), .A2(n5791), .ZN(n9816) );
  OR2_X1 U6097 ( .A1(n9585), .A2(n5872), .ZN(n5792) );
  NAND2_X1 U6098 ( .A1(n5778), .A2(n5777), .ZN(n9825) );
  INV_X1 U6099 ( .A(n10040), .ZN(n9387) );
  NAND2_X1 U6100 ( .A1(n5937), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5465) );
  INV_X1 U6101 ( .A(n9212), .ZN(n5407) );
  XNOR2_X1 U6102 ( .A(n7360), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9399) );
  NAND2_X1 U6103 ( .A1(n4893), .A2(n4631), .ZN(n9397) );
  NAND2_X1 U6104 ( .A1(n7360), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U6105 ( .A1(n4632), .A2(n10375), .ZN(n4631) );
  NAND2_X1 U6106 ( .A1(n4723), .A2(n4722), .ZN(n9415) );
  NAND2_X1 U6107 ( .A1(n4728), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4722) );
  OR2_X1 U6108 ( .A1(n4728), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4723) );
  NAND2_X1 U6109 ( .A1(n9418), .A2(n9417), .ZN(n9416) );
  NAND2_X1 U6110 ( .A1(n4541), .A2(n7362), .ZN(n9418) );
  NAND2_X1 U6111 ( .A1(n4728), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7362) );
  OR2_X1 U6112 ( .A1(n4728), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4541) );
  NOR2_X1 U6113 ( .A1(n7366), .A2(n4884), .ZN(n4883) );
  AOI21_X1 U6114 ( .B1(n7356), .B2(n9440), .A(n7359), .ZN(n7379) );
  AND2_X1 U6115 ( .A1(n9440), .A2(n7356), .ZN(n5237) );
  INV_X1 U6116 ( .A(n7404), .ZN(n4553) );
  INV_X1 U6117 ( .A(n4554), .ZN(n7405) );
  NOR2_X1 U6118 ( .A1(n7520), .A2(n7519), .ZN(n7679) );
  AOI21_X1 U6119 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7522), .A(n7521), .ZN(
        n7524) );
  NAND2_X1 U6120 ( .A1(n7681), .A2(n4612), .ZN(n4611) );
  INV_X1 U6121 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n4612) );
  NOR2_X1 U6122 ( .A1(n7844), .A2(n7845), .ZN(n7979) );
  AND2_X1 U6123 ( .A1(n7983), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4539) );
  NAND2_X1 U6124 ( .A1(n8296), .A2(n4881), .ZN(n8298) );
  NAND2_X1 U6125 ( .A1(n4608), .A2(n8118), .ZN(n4881) );
  INV_X1 U6126 ( .A(n4892), .ZN(n9463) );
  NOR2_X1 U6127 ( .A1(n4416), .A2(n5226), .ZN(n9451) );
  INV_X1 U6128 ( .A(n4730), .ZN(n9465) );
  AND2_X1 U6129 ( .A1(n9948), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9949) );
  OAI21_X1 U6130 ( .B1(n9954), .B2(n4614), .A(n4613), .ZN(n9947) );
  AND2_X1 U6131 ( .A1(n4685), .A2(n4613), .ZN(n9469) );
  NAND2_X1 U6132 ( .A1(n9487), .A2(n9486), .ZN(n9498) );
  NAND2_X1 U6133 ( .A1(n8316), .A2(n5923), .ZN(n5375) );
  XNOR2_X1 U6134 ( .A(n5954), .B(n5869), .ZN(n9531) );
  NAND2_X1 U6135 ( .A1(n5824), .A2(n5823), .ZN(n9540) );
  OAI21_X1 U6136 ( .B1(n9558), .B2(n5160), .A(n5159), .ZN(n9533) );
  NOR2_X1 U6137 ( .A1(n9558), .A2(n6532), .ZN(n9544) );
  NAND2_X1 U6138 ( .A1(n5181), .A2(n5179), .ZN(n9572) );
  INV_X1 U6139 ( .A(n5182), .ZN(n5179) );
  NAND2_X1 U6140 ( .A1(n9605), .A2(n5184), .ZN(n5181) );
  INV_X1 U6141 ( .A(n4952), .ZN(n4960) );
  OAI21_X1 U6142 ( .B1(n9605), .B2(n5766), .A(n5186), .ZN(n9590) );
  INV_X1 U6143 ( .A(n9320), .ZN(n9828) );
  AOI21_X1 U6144 ( .B1(n9629), .B2(n9628), .A(n6443), .ZN(n9607) );
  INV_X1 U6145 ( .A(n9815), .ZN(n9834) );
  NAND2_X1 U6146 ( .A1(n5206), .A2(n5723), .ZN(n9632) );
  OR2_X1 U6147 ( .A1(n9649), .A2(n4417), .ZN(n5206) );
  INV_X1 U6148 ( .A(n4586), .ZN(n9651) );
  OAI21_X1 U6149 ( .B1(n5867), .B2(n4966), .A(n4965), .ZN(n4586) );
  NAND2_X1 U6150 ( .A1(n9691), .A2(n6673), .ZN(n9662) );
  AND2_X1 U6151 ( .A1(n9691), .A2(n4967), .ZN(n9661) );
  NAND2_X1 U6152 ( .A1(n4945), .A2(n6474), .ZN(n9753) );
  NAND2_X1 U6153 ( .A1(n4941), .A2(n6658), .ZN(n8231) );
  NAND2_X1 U6154 ( .A1(n8167), .A2(n8171), .ZN(n5191) );
  INV_X1 U6155 ( .A(n9747), .ZN(n9995) );
  AND2_X1 U6156 ( .A1(n9997), .A2(n5935), .ZN(n9704) );
  NAND2_X2 U6157 ( .A1(n4942), .A2(n4757), .ZN(n5848) );
  NAND2_X1 U6158 ( .A1(n7320), .A2(n4756), .ZN(n4757) );
  NAND2_X1 U6159 ( .A1(n4400), .A2(n4632), .ZN(n4942) );
  OAI22_X1 U6160 ( .A1(n7307), .A2(n4758), .B1(n4815), .B2(n10311), .ZN(n4756)
         );
  NAND2_X1 U6161 ( .A1(n4389), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6162 ( .A1(n9923), .A2(n5933), .ZN(n9671) );
  NAND2_X1 U6163 ( .A1(n7320), .A2(n7295), .ZN(n5080) );
  OR2_X1 U6164 ( .A1(n7320), .A2(n4600), .ZN(n5081) );
  AND2_X1 U6165 ( .A1(n9997), .A2(n7128), .ZN(n9747) );
  NAND2_X1 U6166 ( .A1(n5067), .A2(n4660), .ZN(n4659) );
  OAI21_X1 U6167 ( .B1(n9809), .B2(n10057), .A(n4457), .ZN(n4726) );
  AND2_X1 U6168 ( .A1(n9808), .A2(n10078), .ZN(n4727) );
  AND2_X1 U6169 ( .A1(n9924), .A2(n9923), .ZN(n10001) );
  AND2_X1 U6170 ( .A1(n5213), .A2(n4592), .ZN(n4591) );
  INV_X1 U6171 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4592) );
  OR2_X1 U6172 ( .A1(n5888), .A2(n5368), .ZN(n4654) );
  OAI21_X1 U6173 ( .B1(n5842), .B2(n5367), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5888) );
  INV_X1 U6174 ( .A(n5148), .ZN(n5147) );
  OAI21_X1 U6175 ( .B1(n5151), .B2(n5150), .A(n5149), .ZN(n5148) );
  INV_X1 U6176 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8309) );
  XNOR2_X1 U6177 ( .A(n5767), .B(n5768), .ZN(n8306) );
  OAI21_X1 U6178 ( .B1(n5712), .B2(n4856), .A(n4853), .ZN(n5767) );
  INV_X1 U6179 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8275) );
  INV_X1 U6180 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10371) );
  INV_X1 U6181 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7516) );
  XNOR2_X1 U6182 ( .A(n5581), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8122) );
  AND2_X1 U6183 ( .A1(n5533), .A2(n5548), .ZN(n7680) );
  INV_X1 U6184 ( .A(n5516), .ZN(n5518) );
  XNOR2_X1 U6185 ( .A(n5447), .B(P1_IR_REG_5__SCAN_IN), .ZN(n8330) );
  INV_X1 U6186 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7301) );
  INV_X1 U6187 ( .A(n5441), .ZN(n5438) );
  INV_X1 U6188 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U6189 ( .A1(n4629), .A2(n5012), .ZN(n7970) );
  XNOR2_X1 U6190 ( .A(n8242), .B(n8243), .ZN(n8244) );
  NAND2_X1 U6191 ( .A1(n4714), .A2(n8714), .ZN(n4713) );
  NAND2_X1 U6192 ( .A1(n4642), .A2(n8714), .ZN(n8715) );
  NAND2_X1 U6193 ( .A1(n4764), .A2(n8338), .ZN(P2_U3204) );
  NAND2_X1 U6194 ( .A1(n4822), .A2(n10128), .ZN(n4764) );
  NAND2_X1 U6195 ( .A1(n7159), .A2(n4498), .ZN(n4820) );
  OAI21_X1 U6196 ( .B1(n9019), .B2(n10164), .A(n5050), .ZN(P2_U3486) );
  INV_X1 U6197 ( .A(n5051), .ZN(n5050) );
  OAI21_X1 U6198 ( .B1(n9024), .B2(n8972), .A(n5052), .ZN(n5051) );
  NOR2_X1 U6199 ( .A1(n4437), .A2(n5053), .ZN(n5052) );
  NAND2_X1 U6200 ( .A1(n4636), .A2(n7160), .ZN(n7161) );
  OAI21_X1 U6201 ( .B1(n7306), .B2(n9132), .A(n4900), .ZN(P2_U3293) );
  NOR2_X1 U6202 ( .A1(n4903), .A2(n4901), .ZN(n4900) );
  NOR2_X1 U6203 ( .A1(P2_U3151), .A2(n4902), .ZN(n4901) );
  NOR2_X1 U6204 ( .A1(n9130), .A2(n7305), .ZN(n4903) );
  NOR2_X1 U6205 ( .A1(n5107), .A2(n5097), .ZN(n5100) );
  AND2_X1 U6206 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  AND2_X1 U6207 ( .A1(n4583), .A2(n4481), .ZN(n9970) );
  AOI21_X1 U6208 ( .B1(n9506), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9505), .ZN(
        n4894) );
  NAND2_X1 U6209 ( .A1(n4538), .A2(n5846), .ZN(n4537) );
  NAND2_X1 U6210 ( .A1(n8978), .A2(n8478), .ZN(n4401) );
  NAND2_X1 U6211 ( .A1(n5653), .A2(n5652), .ZN(n5860) );
  CLKBUF_X3 U6212 ( .A(n6014), .Z(n6213) );
  INV_X1 U6213 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9111) );
  OAI211_X1 U6214 ( .C1(P1_IR_REG_31__SCAN_IN), .C2(P1_IR_REG_1__SCAN_IN), .A(
        n4602), .B(n4601), .ZN(n7360) );
  AND2_X1 U6215 ( .A1(n8330), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4403) );
  INV_X1 U6216 ( .A(n6275), .ZN(n6276) );
  NAND2_X1 U6217 ( .A1(n9801), .A2(n9562), .ZN(n6612) );
  NAND2_X1 U6218 ( .A1(n4428), .A2(n6154), .ZN(n4404) );
  NOR2_X1 U6219 ( .A1(n9667), .A2(n4968), .ZN(n4967) );
  AND2_X1 U6220 ( .A1(n7821), .A2(n6089), .ZN(n4405) );
  NAND2_X1 U6221 ( .A1(n5068), .A2(n5071), .ZN(n9705) );
  AND2_X1 U6222 ( .A1(n9504), .A2(n9496), .ZN(n4406) );
  AND2_X1 U6223 ( .A1(n6141), .A2(n4772), .ZN(n4407) );
  AND2_X1 U6224 ( .A1(n6410), .A2(n6790), .ZN(n4408) );
  INV_X1 U6225 ( .A(n5144), .ZN(n5143) );
  NAND2_X1 U6226 ( .A1(n4425), .A2(n5273), .ZN(n5144) );
  NAND2_X1 U6227 ( .A1(n5988), .A2(n6001), .ZN(n4409) );
  INV_X1 U6228 ( .A(n7611), .ZN(n7640) );
  NAND2_X1 U6229 ( .A1(n4430), .A2(n6810), .ZN(n4410) );
  AND2_X1 U6230 ( .A1(n4830), .A2(n6817), .ZN(n4411) );
  NAND2_X1 U6231 ( .A1(n7959), .A2(n5122), .ZN(n4412) );
  NOR2_X1 U6232 ( .A1(n4409), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4413) );
  NAND2_X1 U6233 ( .A1(n9077), .A2(n5041), .ZN(n5040) );
  NAND2_X1 U6234 ( .A1(n5066), .A2(n9204), .ZN(n8135) );
  INV_X1 U6235 ( .A(n8163), .ZN(n6406) );
  NAND2_X1 U6236 ( .A1(n7180), .A2(n7767), .ZN(n7769) );
  AND2_X1 U6237 ( .A1(n4871), .A2(n4870), .ZN(n4414) );
  INV_X1 U6238 ( .A(n9968), .ZN(n4733) );
  INV_X1 U6239 ( .A(n7506), .ZN(n4644) );
  AND2_X1 U6240 ( .A1(n9118), .A2(n4393), .ZN(n4415) );
  INV_X1 U6241 ( .A(n7100), .ZN(n5097) );
  AND2_X1 U6242 ( .A1(n8293), .A2(n4604), .ZN(n4416) );
  NOR2_X1 U6243 ( .A1(n9657), .A2(n9638), .ZN(n4417) );
  INV_X1 U6244 ( .A(n4672), .ZN(n10021) );
  NAND2_X1 U6245 ( .A1(n5925), .A2(n5924), .ZN(n9779) );
  NAND2_X1 U6246 ( .A1(n5758), .A2(n5757), .ZN(n9320) );
  AND2_X1 U6247 ( .A1(n5535), .A2(n5534), .ZN(n9204) );
  NAND2_X1 U6248 ( .A1(n7167), .A2(n7166), .ZN(n7170) );
  NAND2_X1 U6249 ( .A1(n6229), .A2(n6228), .ZN(n9068) );
  OR2_X1 U6250 ( .A1(n5947), .A2(n9779), .ZN(n4418) );
  XNOR2_X1 U6251 ( .A(n8329), .B(n7692), .ZN(n6580) );
  AND2_X1 U6252 ( .A1(n8600), .A2(n8618), .ZN(n4419) );
  NAND2_X1 U6253 ( .A1(n6826), .A2(n6825), .ZN(n6890) );
  XNOR2_X1 U6254 ( .A(n5436), .B(n10227), .ZN(n9422) );
  AND2_X1 U6255 ( .A1(n9670), .A2(n5074), .ZN(n9608) );
  OR2_X1 U6256 ( .A1(n9540), .A2(n9384), .ZN(n4420) );
  NAND2_X1 U6257 ( .A1(n5860), .A2(n9891), .ZN(n4421) );
  AND2_X1 U6258 ( .A1(n5039), .A2(n5040), .ZN(n4422) );
  OR2_X1 U6259 ( .A1(n8429), .A2(n8878), .ZN(n4423) );
  OR2_X1 U6260 ( .A1(n9088), .A2(n8889), .ZN(n4424) );
  INV_X1 U6261 ( .A(n6963), .ZN(n5122) );
  OR2_X1 U6262 ( .A1(n5275), .A2(SI_9_), .ZN(n4425) );
  AND4_X1 U6263 ( .A1(n6511), .A2(n6514), .A3(n6521), .A4(n6510), .ZN(n4426)
         );
  OR3_X1 U6264 ( .A1(n7147), .A2(n7148), .A3(n10132), .ZN(n4427) );
  NAND2_X1 U6265 ( .A1(n8160), .A2(n8904), .ZN(n4428) );
  AND2_X1 U6266 ( .A1(n6520), .A2(n6521), .ZN(n4429) );
  OAI21_X1 U6267 ( .B1(n5334), .B2(n4563), .A(n4560), .ZN(n5794) );
  OAI21_X1 U6268 ( .B1(n8774), .B2(n4783), .A(n4780), .ZN(n8737) );
  NAND2_X1 U6269 ( .A1(n9039), .A2(n8746), .ZN(n4430) );
  INV_X1 U6270 ( .A(n9902), .ZN(n5073) );
  AND2_X1 U6271 ( .A1(n8330), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4431) );
  AND3_X1 U6272 ( .A1(n9193), .A2(n9359), .A3(n9192), .ZN(n4432) );
  INV_X1 U6273 ( .A(n7297), .ZN(n5243) );
  AND2_X1 U6274 ( .A1(n8330), .A2(n7357), .ZN(n4433) );
  INV_X1 U6275 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6023) );
  AND2_X1 U6276 ( .A1(n7407), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4434) );
  NAND4_X1 U6277 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5578), .ZN(n5666)
         );
  XNOR2_X1 U6278 ( .A(n6078), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7604) );
  NOR3_X1 U6279 ( .A1(n6641), .A2(n6497), .A3(n6634), .ZN(n4435) );
  AND2_X1 U6280 ( .A1(n7103), .A2(n7102), .ZN(n4436) );
  NAND2_X1 U6281 ( .A1(n5770), .A2(n5769), .ZN(n9600) );
  NAND2_X1 U6282 ( .A1(n5201), .A2(n5200), .ZN(n9663) );
  AND2_X1 U6283 ( .A1(n9021), .A2(n8967), .ZN(n4437) );
  INV_X1 U6284 ( .A(n8846), .ZN(n5038) );
  AND2_X1 U6285 ( .A1(n6786), .A2(n4402), .ZN(n4438) );
  OR2_X1 U6286 ( .A1(n9808), .A2(n9577), .ZN(n4439) );
  AND2_X1 U6287 ( .A1(n5491), .A2(n5490), .ZN(n10027) );
  AND3_X1 U6288 ( .A1(n8810), .A2(n6789), .A3(n4922), .ZN(n4440) );
  AND2_X1 U6289 ( .A1(n5012), .A2(n7188), .ZN(n4441) );
  NAND2_X1 U6290 ( .A1(n5081), .A2(n5080), .ZN(n8325) );
  AND2_X1 U6291 ( .A1(n6523), .A2(n6522), .ZN(n4442) );
  AND2_X1 U6292 ( .A1(n7605), .A2(n7611), .ZN(n4443) );
  AND2_X1 U6293 ( .A1(n6996), .A2(n6998), .ZN(n4444) );
  AND2_X1 U6294 ( .A1(n6452), .A2(n7869), .ZN(n4445) );
  INV_X2 U6295 ( .A(n5775), .ZN(n5937) );
  AND2_X1 U6296 ( .A1(n7193), .A2(n8548), .ZN(n4446) );
  NOR2_X1 U6297 ( .A1(n9773), .A2(n10057), .ZN(n4447) );
  INV_X1 U6298 ( .A(n5292), .ZN(n5171) );
  AND2_X1 U6299 ( .A1(n7174), .A2(n4836), .ZN(n4448) );
  INV_X1 U6300 ( .A(n9657), .ZN(n9854) );
  NAND2_X1 U6301 ( .A1(n5718), .A2(n5717), .ZN(n9657) );
  INV_X1 U6302 ( .A(n6813), .ZN(n4831) );
  OR2_X1 U6303 ( .A1(n7280), .A2(n9021), .ZN(n4449) );
  OR2_X1 U6304 ( .A1(n6894), .A2(n6891), .ZN(n4450) );
  AND2_X1 U6305 ( .A1(n5222), .A2(n6571), .ZN(n4451) );
  AND2_X1 U6306 ( .A1(n6599), .A2(n6439), .ZN(n6593) );
  AND2_X1 U6307 ( .A1(n7184), .A2(n8551), .ZN(n4452) );
  AND2_X1 U6308 ( .A1(n8757), .A2(n8778), .ZN(n4453) );
  AND2_X1 U6309 ( .A1(n5889), .A2(n4653), .ZN(n4454) );
  AND2_X1 U6310 ( .A1(n4878), .A2(n4877), .ZN(n4455) );
  INV_X1 U6311 ( .A(n9204), .ZN(n10043) );
  INV_X1 U6312 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5370) );
  INV_X1 U6313 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5215) );
  OR2_X1 U6314 ( .A1(n7148), .A2(n7285), .ZN(n4456) );
  NOR2_X1 U6315 ( .A1(n9807), .A2(n4727), .ZN(n4457) );
  NOR2_X1 U6316 ( .A1(n9195), .A2(n6974), .ZN(n4458) );
  NOR2_X1 U6317 ( .A1(n10054), .A2(n9386), .ZN(n4459) );
  NOR2_X1 U6318 ( .A1(n9812), .A2(n9816), .ZN(n4460) );
  NOR2_X1 U6319 ( .A1(n8383), .A2(n8835), .ZN(n4461) );
  OR2_X1 U6320 ( .A1(n9027), .A2(n8422), .ZN(n6820) );
  AND2_X1 U6321 ( .A1(n5045), .A2(n5044), .ZN(n4462) );
  AND2_X1 U6322 ( .A1(n5141), .A2(n5138), .ZN(n4463) );
  INV_X1 U6323 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5369) );
  NAND2_X1 U6324 ( .A1(n10214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4464) );
  AND2_X1 U6325 ( .A1(n6487), .A2(n6488), .ZN(n4465) );
  NAND2_X1 U6326 ( .A1(n5171), .A2(n5163), .ZN(n4466) );
  AND2_X1 U6327 ( .A1(n6748), .A2(n6749), .ZN(n4467) );
  INV_X1 U6328 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5368) );
  INV_X1 U6329 ( .A(n4830), .ZN(n4829) );
  NOR2_X1 U6330 ( .A1(n6818), .A2(n4831), .ZN(n4830) );
  OR2_X1 U6331 ( .A1(n5025), .A2(n4773), .ZN(n4468) );
  AND2_X1 U6332 ( .A1(n5129), .A2(n7048), .ZN(n4469) );
  INV_X1 U6333 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7303) );
  OR2_X1 U6334 ( .A1(n4783), .A2(n4779), .ZN(n4470) );
  INV_X1 U6335 ( .A(n4967), .ZN(n4966) );
  AND2_X1 U6336 ( .A1(n5368), .A2(n5215), .ZN(n4471) );
  AND2_X1 U6337 ( .A1(n5104), .A2(n5101), .ZN(n4472) );
  INV_X1 U6338 ( .A(n6141), .ZN(n4773) );
  INV_X1 U6339 ( .A(n7821), .ZN(n7824) );
  NAND2_X1 U6340 ( .A1(n6756), .A2(n7881), .ZN(n7821) );
  OR2_X1 U6341 ( .A1(n6812), .A2(n6811), .ZN(n8753) );
  INV_X1 U6342 ( .A(n8753), .ZN(n4930) );
  NAND2_X1 U6343 ( .A1(n7551), .A2(n4907), .ZN(n7552) );
  INV_X1 U6344 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10214) );
  INV_X1 U6345 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5883) );
  INV_X1 U6346 ( .A(n6812), .ZN(n4790) );
  NAND2_X1 U6347 ( .A1(n7216), .A2(n7214), .ZN(n4473) );
  OR2_X1 U6348 ( .A1(n7732), .A2(n8551), .ZN(n4474) );
  AND2_X1 U6349 ( .A1(n6657), .A2(n4753), .ZN(n4475) );
  NAND2_X1 U6350 ( .A1(n6618), .A2(n6620), .ZN(n9782) );
  OR2_X1 U6351 ( .A1(n9787), .A2(n9715), .ZN(n4476) );
  OR2_X1 U6352 ( .A1(n6745), .A2(n6735), .ZN(n7742) );
  AND2_X1 U6353 ( .A1(n8527), .A2(n7214), .ZN(n4477) );
  OR2_X1 U6354 ( .A1(n5298), .A2(SI_16_), .ZN(n4478) );
  INV_X1 U6355 ( .A(n9874), .ZN(n9675) );
  AND2_X1 U6356 ( .A1(n5691), .A2(n5690), .ZN(n9874) );
  AND2_X1 U6357 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4479) );
  AND2_X1 U6358 ( .A1(n6415), .A2(n8759), .ZN(n4480) );
  NOR2_X1 U6359 ( .A1(n4734), .A2(n4731), .ZN(n4481) );
  OR2_X1 U6360 ( .A1(n6686), .A2(n6634), .ZN(n4482) );
  AND2_X1 U6361 ( .A1(n5869), .A2(n4420), .ZN(n4483) );
  NOR2_X1 U6362 ( .A1(n9544), .A2(n9553), .ZN(n4484) );
  NOR2_X1 U6363 ( .A1(n9469), .A2(n9468), .ZN(n4485) );
  NAND2_X1 U6364 ( .A1(n7145), .A2(n10111), .ZN(n4486) );
  AND2_X1 U6365 ( .A1(n6198), .A2(n6773), .ZN(n4487) );
  AND2_X1 U6366 ( .A1(n5200), .A2(n5199), .ZN(n4488) );
  INV_X1 U6367 ( .A(n9591), .ZN(n4956) );
  AND2_X1 U6368 ( .A1(n6528), .A2(n9576), .ZN(n9591) );
  INV_X1 U6369 ( .A(n6499), .ZN(n9681) );
  NAND2_X1 U6370 ( .A1(n6501), .A2(n6673), .ZN(n6499) );
  AND2_X1 U6371 ( .A1(n6884), .A2(n7141), .ZN(n4489) );
  AND2_X1 U6372 ( .A1(n5162), .A2(n5293), .ZN(n4490) );
  AND2_X1 U6373 ( .A1(n8726), .A2(n6821), .ZN(n4491) );
  OAI21_X1 U6374 ( .B1(n4827), .B2(n4826), .A(n4449), .ZN(n4825) );
  OR2_X1 U6375 ( .A1(n9746), .A2(n9882), .ZN(n4492) );
  INV_X1 U6376 ( .A(n6223), .ZN(n5039) );
  AND2_X1 U6377 ( .A1(n8954), .A2(n8849), .ZN(n6223) );
  NAND2_X1 U6378 ( .A1(n6396), .A2(n4392), .ZN(n6726) );
  INV_X1 U6379 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5446) );
  INV_X1 U6380 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4721) );
  AND2_X1 U6381 ( .A1(n9575), .A2(n9576), .ZN(n4493) );
  INV_X1 U6382 ( .A(n6766), .ZN(n4928) );
  INV_X1 U6383 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5152) );
  XNOR2_X1 U6384 ( .A(n5281), .B(SI_11_), .ZN(n5576) );
  AND2_X1 U6385 ( .A1(n6406), .A2(n6765), .ZN(n4494) );
  AND2_X1 U6386 ( .A1(n5999), .A2(n5998), .ZN(n8861) );
  XNOR2_X1 U6387 ( .A(n5840), .B(n5839), .ZN(n8212) );
  INV_X1 U6388 ( .A(n8212), .ZN(n4530) );
  INV_X1 U6389 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U6390 ( .A1(n5851), .A2(n6459), .ZN(n7995) );
  AND2_X1 U6391 ( .A1(n8002), .A2(n10027), .ZN(n8003) );
  OR2_X1 U6392 ( .A1(n7048), .A2(n5131), .ZN(n5130) );
  OR2_X1 U6393 ( .A1(n8162), .A2(n8163), .ZN(n8161) );
  INV_X1 U6394 ( .A(n8259), .ZN(n4982) );
  AND2_X1 U6395 ( .A1(n5066), .A2(n5065), .ZN(n4495) );
  NAND2_X1 U6396 ( .A1(n9288), .A2(n6981), .ZN(n9155) );
  NAND2_X1 U6397 ( .A1(n8243), .A2(n10343), .ZN(n4496) );
  NAND2_X1 U6398 ( .A1(n5027), .A2(n6154), .ZN(n8156) );
  NAND2_X1 U6399 ( .A1(n5204), .A2(n5631), .ZN(n9735) );
  NAND2_X1 U6400 ( .A1(n5191), .A2(n5544), .ZN(n8133) );
  NAND2_X1 U6401 ( .A1(n6409), .A2(n6784), .ZN(n8842) );
  OR2_X1 U6402 ( .A1(n5855), .A2(n5852), .ZN(n6656) );
  INV_X1 U6403 ( .A(n6656), .ZN(n4670) );
  AND2_X1 U6404 ( .A1(n7060), .A2(n7059), .ZN(n4497) );
  NOR2_X1 U6405 ( .A1(P2_REG1_REG_29__SCAN_IN), .A2(n10166), .ZN(n4498) );
  AND2_X1 U6406 ( .A1(n4869), .A2(n4868), .ZN(n4499) );
  AND2_X1 U6407 ( .A1(n4914), .A2(n4913), .ZN(n4500) );
  AND2_X1 U6408 ( .A1(n7680), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4501) );
  NOR2_X1 U6409 ( .A1(n9759), .A2(n5072), .ZN(n9721) );
  INV_X1 U6410 ( .A(n9299), .ZN(n5134) );
  NAND2_X1 U6411 ( .A1(n7189), .A2(n8385), .ZN(n8388) );
  NAND2_X1 U6412 ( .A1(n6356), .A2(n6090), .ZN(n4502) );
  AND2_X1 U6413 ( .A1(n4912), .A2(n4496), .ZN(n4503) );
  INV_X1 U6414 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4600) );
  NOR2_X1 U6415 ( .A1(n9452), .A2(n4509), .ZN(n4540) );
  AND2_X1 U6416 ( .A1(n8388), .A2(n7191), .ZN(n4504) );
  AND2_X1 U6417 ( .A1(n4874), .A2(n4873), .ZN(n4505) );
  AND2_X1 U6418 ( .A1(n4979), .A2(n4982), .ZN(n4506) );
  INV_X2 U6419 ( .A(n10159), .ZN(n10157) );
  AND2_X1 U6420 ( .A1(n6434), .A2(n6433), .ZN(n10159) );
  INV_X1 U6421 ( .A(n8572), .ZN(n4984) );
  INV_X1 U6422 ( .A(n8618), .ZN(n4897) );
  XNOR2_X1 U6424 ( .A(n7181), .B(n8552), .ZN(n7767) );
  INV_X1 U6425 ( .A(n7959), .ZN(n5120) );
  AND2_X1 U6426 ( .A1(n6711), .A2(n10122), .ZN(n10130) );
  INV_X1 U6427 ( .A(n8714), .ZN(n8690) );
  NAND2_X1 U6428 ( .A1(n5671), .A2(n5670), .ZN(n9877) );
  INV_X1 U6429 ( .A(n9877), .ZN(n5070) );
  AND2_X1 U6430 ( .A1(n6994), .A2(n6993), .ZN(n4507) );
  AND3_X1 U6431 ( .A1(n4974), .A2(n4976), .A3(n4972), .ZN(n4508) );
  AND2_X1 U6432 ( .A1(n9453), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4509) );
  AND2_X1 U6433 ( .A1(n4885), .A2(n4887), .ZN(n4510) );
  AND2_X1 U6434 ( .A1(n4599), .A2(n9493), .ZN(n4511) );
  NOR2_X1 U6435 ( .A1(n9499), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n4512) );
  AND2_X1 U6436 ( .A1(n8647), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4513) );
  AND2_X1 U6437 ( .A1(n5599), .A2(n5618), .ZN(n8297) );
  INV_X1 U6438 ( .A(n8297), .ZN(n4608) );
  NOR2_X1 U6439 ( .A1(n7674), .A2(n5219), .ZN(n4514) );
  AND2_X1 U6440 ( .A1(n7769), .A2(n7182), .ZN(n4515) );
  AND2_X1 U6441 ( .A1(n7471), .A2(n7173), .ZN(n4516) );
  NAND2_X1 U6442 ( .A1(n9610), .A2(n8269), .ZN(n4517) );
  INV_X1 U6443 ( .A(n8674), .ZN(n4895) );
  INV_X1 U6444 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4868) );
  INV_X1 U6445 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U6446 ( .A1(n5212), .A2(n4591), .ZN(n4594) );
  NOR2_X1 U6447 ( .A1(n7370), .A2(n7369), .ZN(n4518) );
  INV_X1 U6448 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4635) );
  INV_X1 U6449 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n4884) );
  INV_X1 U6450 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n4712) );
  NAND2_X1 U6451 ( .A1(n4521), .A2(n7139), .ZN(P1_U3214) );
  NAND2_X1 U6452 ( .A1(n4522), .A2(n9359), .ZN(n4521) );
  NAND2_X1 U6453 ( .A1(n4524), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U6454 ( .A1(n9358), .A2(n7114), .ZN(n4523) );
  OAI211_X2 U6455 ( .C1(n9288), .C2(n4525), .A(n4526), .B(n5112), .ZN(n9307)
         );
  NAND2_X1 U6456 ( .A1(n4528), .A2(n5118), .ZN(n6977) );
  NAND2_X1 U6457 ( .A1(n6961), .A2(n5119), .ZN(n4528) );
  NAND2_X1 U6458 ( .A1(n4529), .A2(n5085), .ZN(n5084) );
  NAND2_X1 U6459 ( .A1(n4529), .A2(n9145), .ZN(n5090) );
  XNOR2_X1 U6460 ( .A(n4529), .B(n9146), .ZN(n9152) );
  NAND2_X1 U6461 ( .A1(n7075), .A2(n9313), .ZN(n4529) );
  NAND2_X1 U6462 ( .A1(n5667), .A2(n5668), .ZN(n5683) );
  AND3_X2 U6463 ( .A1(n5396), .A2(n5363), .A3(n5446), .ZN(n5668) );
  INV_X1 U6464 ( .A(n5683), .ZN(n5684) );
  AND2_X1 U6465 ( .A1(n4531), .A2(n6932), .ZN(n9337) );
  AND2_X2 U6466 ( .A1(n9336), .A2(n4531), .ZN(n7890) );
  NAND2_X1 U6467 ( .A1(n4676), .A2(n4675), .ZN(n4531) );
  NAND3_X1 U6468 ( .A1(n4537), .A2(n4894), .A3(n4533), .ZN(P1_U3262) );
  NAND2_X1 U6469 ( .A1(n4534), .A2(n5934), .ZN(n4533) );
  NAND2_X1 U6470 ( .A1(n4536), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U6471 ( .A1(n9503), .A2(n9502), .ZN(n4536) );
  OAI22_X1 U6472 ( .A1(n9503), .A2(n9959), .B1(n9504), .B2(n9963), .ZN(n4538)
         );
  INV_X1 U6473 ( .A(n4540), .ZN(n4674) );
  NOR2_X1 U6474 ( .A1(n8298), .A2(n8299), .ZN(n9452) );
  NOR2_X1 U6475 ( .A1(n7378), .A2(n7377), .ZN(n7403) );
  NAND2_X1 U6476 ( .A1(n9416), .A2(n7363), .ZN(n9430) );
  AOI21_X1 U6477 ( .B1(n4542), .B2(n9576), .A(n4704), .ZN(n6530) );
  NAND2_X1 U6478 ( .A1(n4544), .A2(n4442), .ZN(n4543) );
  NAND2_X1 U6479 ( .A1(n4549), .A2(n4547), .ZN(n4551) );
  INV_X1 U6480 ( .A(n6717), .ZN(n4548) );
  INV_X1 U6481 ( .A(n5594), .ZN(n5166) );
  NAND2_X1 U6482 ( .A1(n4555), .A2(n4557), .ZN(n4865) );
  NAND3_X1 U6483 ( .A1(n5135), .A2(n5137), .A3(n4558), .ZN(n4557) );
  NOR2_X1 U6484 ( .A1(n4559), .A2(n6834), .ZN(n6840) );
  NAND2_X1 U6485 ( .A1(n4559), .A2(n4807), .ZN(n6842) );
  NAND2_X1 U6486 ( .A1(n5334), .A2(n5333), .ZN(n5781) );
  NAND2_X1 U6487 ( .A1(n4564), .A2(n4482), .ZN(n6639) );
  NAND3_X1 U6488 ( .A1(n4565), .A2(n6633), .A3(n6686), .ZN(n4564) );
  NAND2_X1 U6489 ( .A1(n4566), .A2(n4698), .ZN(n4565) );
  NAND2_X1 U6490 ( .A1(n4846), .A2(n4845), .ZN(n4566) );
  INV_X1 U6491 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4570) );
  INV_X1 U6492 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4571) );
  NAND3_X1 U6493 ( .A1(n5297), .A2(n5296), .A3(n4478), .ZN(n4579) );
  NAND3_X1 U6494 ( .A1(n4584), .A2(n9958), .A3(n9502), .ZN(n4583) );
  NOR2_X1 U6495 ( .A1(n9464), .A2(n4889), .ZN(n9948) );
  NOR2_X1 U6496 ( .A1(n9436), .A2(n4883), .ZN(n7370) );
  NAND2_X1 U6497 ( .A1(n9430), .A2(n9431), .ZN(n9429) );
  XNOR2_X2 U6498 ( .A(n5434), .B(n5433), .ZN(n4728) );
  AND2_X2 U6499 ( .A1(n4759), .A2(n4597), .ZN(n5372) );
  NAND3_X1 U6500 ( .A1(n4656), .A2(n4655), .A3(n5596), .ZN(n5843) );
  NAND3_X1 U6501 ( .A1(n4476), .A2(n5956), .A3(n5957), .ZN(P1_U3356) );
  NAND2_X1 U6502 ( .A1(n4600), .A2(n4721), .ZN(n4602) );
  NAND3_X1 U6503 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4601) );
  NOR2_X1 U6504 ( .A1(n8330), .A2(n7357), .ZN(n4603) );
  NAND2_X1 U6505 ( .A1(n8293), .A2(n4606), .ZN(n8294) );
  NOR2_X1 U6506 ( .A1(n8295), .A2(n4605), .ZN(n4604) );
  NAND2_X1 U6507 ( .A1(n8125), .A2(n8126), .ZN(n8293) );
  NAND2_X1 U6508 ( .A1(n7843), .A2(n4611), .ZN(n7844) );
  NOR2_X4 U6509 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7433) );
  NAND2_X1 U6510 ( .A1(n7164), .A2(n8266), .ZN(n7165) );
  AOI21_X1 U6511 ( .B1(n6337), .B2(n4479), .A(n4619), .ZN(n4618) );
  NAND2_X1 U6512 ( .A1(n4621), .A2(n4622), .ZN(n7231) );
  NAND2_X1 U6513 ( .A1(n8378), .A2(n4624), .ZN(n4621) );
  NAND3_X1 U6514 ( .A1(n4628), .A2(n4627), .A3(n6356), .ZN(n6334) );
  NAND2_X1 U6515 ( .A1(n4628), .A2(n6356), .ZN(n6363) );
  NAND2_X1 U6516 ( .A1(n5000), .A2(n7471), .ZN(n7534) );
  NAND2_X1 U6517 ( .A1(n7481), .A2(n7169), .ZN(n7470) );
  NAND2_X1 U6518 ( .A1(n4630), .A2(n7765), .ZN(n4629) );
  OAI21_X1 U6519 ( .B1(n7189), .B2(n5005), .A(n5003), .ZN(n8364) );
  INV_X1 U6520 ( .A(n8484), .ZN(n7233) );
  XNOR2_X1 U6521 ( .A(n7170), .B(n6396), .ZN(n4999) );
  XNOR2_X1 U6522 ( .A(n8442), .B(n8443), .ZN(n8444) );
  AOI22_X1 U6523 ( .A1(n8510), .A2(n8509), .B1(n7222), .B2(n7221), .ZN(n8378)
         );
  INV_X1 U6524 ( .A(n8530), .ZN(n7211) );
  INV_X1 U6525 ( .A(n9532), .ZN(n4658) );
  NOR2_X2 U6526 ( .A1(n4659), .A2(n9774), .ZN(n4633) );
  NAND2_X1 U6527 ( .A1(n9397), .A2(n9396), .ZN(n9395) );
  INV_X1 U6528 ( .A(n7360), .ZN(n4632) );
  OAI21_X1 U6529 ( .B1(n9787), .B2(n9881), .A(n4633), .ZN(n9907) );
  NAND2_X1 U6530 ( .A1(n4677), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U6531 ( .A1(n4952), .A2(n4958), .ZN(n4951) );
  NAND3_X1 U6532 ( .A1(n4715), .A2(n4713), .A3(n8689), .ZN(P2_U3200) );
  OAI21_X1 U6533 ( .B1(SI_5_), .B2(n5480), .A(n5485), .ZN(n5262) );
  NAND3_X1 U6534 ( .A1(n6908), .A2(n6907), .A3(n6905), .ZN(n4652) );
  NAND3_X1 U6535 ( .A1(n5263), .A2(n5220), .A3(n5441), .ZN(n4699) );
  NAND2_X1 U6536 ( .A1(n4843), .A2(n5349), .ZN(n5821) );
  OAI22_X1 U6537 ( .A1(n6929), .A2(n6965), .B1(n9212), .B2(n9176), .ZN(n6928)
         );
  OR2_X1 U6538 ( .A1(n5563), .A2(n7306), .ZN(n5406) );
  AOI21_X2 U6539 ( .B1(n9242), .B2(n7028), .A(n7027), .ZN(n9255) );
  NAND2_X1 U6540 ( .A1(n5525), .A2(n5273), .ZN(n4700) );
  NAND2_X1 U6541 ( .A1(n4701), .A2(n4451), .ZN(n4665) );
  INV_X1 U6542 ( .A(n8329), .ZN(n4646) );
  NAND2_X1 U6543 ( .A1(n4646), .A2(n6941), .ZN(n4694) );
  NAND2_X1 U6544 ( .A1(n6357), .A2(n5225), .ZN(n6361) );
  NAND2_X1 U6545 ( .A1(n8765), .A2(n6880), .ZN(n6417) );
  AOI21_X1 U6546 ( .B1(n4824), .B2(n4411), .A(n4825), .ZN(n6888) );
  INV_X1 U6547 ( .A(n8458), .ZN(n10147) );
  AOI21_X2 U6548 ( .B1(n8808), .B2(n6720), .A(n6412), .ZN(n8797) );
  NAND4_X1 U6549 ( .A1(n7156), .A2(n7157), .A3(n4823), .A4(n10157), .ZN(n4636)
         );
  NAND2_X1 U6550 ( .A1(n7728), .A2(n7729), .ZN(n5062) );
  AND3_X2 U6551 ( .A1(n5985), .A2(n5984), .A3(n5983), .ZN(n5225) );
  INV_X1 U6552 ( .A(n7741), .ZN(n4708) );
  NAND2_X1 U6553 ( .A1(n5247), .A2(SI_1_), .ZN(n5398) );
  OAI22_X1 U6554 ( .A1(n8444), .A2(n8790), .B1(n8443), .B2(n8442), .ZN(n8447)
         );
  NAND2_X1 U6555 ( .A1(n4641), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U6556 ( .A1(n7968), .A2(n8384), .ZN(n7189) );
  NAND2_X1 U6557 ( .A1(n6375), .A2(n6374), .ZN(n7163) );
  INV_X1 U6558 ( .A(n5397), .ZN(n5396) );
  AND4_X2 U6559 ( .A1(n5418), .A2(n5416), .A3(n5417), .A4(n5415), .ZN(n8329)
         );
  NAND2_X1 U6560 ( .A1(n5125), .A2(n5124), .ZN(n9216) );
  NAND2_X1 U6561 ( .A1(n4650), .A2(n5848), .ZN(n4693) );
  NAND2_X1 U6562 ( .A1(n6977), .A2(n6976), .ZN(n9288) );
  INV_X2 U6563 ( .A(n4650), .ZN(n6965) );
  NOR2_X2 U6564 ( .A1(n8635), .A2(n4419), .ZN(n8601) );
  NOR2_X2 U6565 ( .A1(n8648), .A2(n8674), .ZN(n8669) );
  NAND2_X1 U6566 ( .A1(n4971), .A2(n7640), .ZN(n4974) );
  NAND2_X1 U6567 ( .A1(n8187), .A2(n8186), .ZN(n8188) );
  NOR2_X2 U6568 ( .A1(n4983), .A2(n8585), .ZN(n8555) );
  NOR2_X1 U6569 ( .A1(n8667), .A2(n4657), .ZN(n8671) );
  NAND2_X1 U6570 ( .A1(n8649), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4994) );
  OAI21_X1 U6571 ( .B1(n4652), .B2(n4651), .A(n6913), .ZN(P2_U3296) );
  INV_X1 U6572 ( .A(n6906), .ZN(n4651) );
  NAND3_X1 U6573 ( .A1(n4699), .A2(n5234), .A3(n5091), .ZN(n5516) );
  NOR2_X2 U6574 ( .A1(n5362), .A2(n5665), .ZN(n4655) );
  INV_X1 U6575 ( .A(n5466), .ZN(n4656) );
  NAND2_X1 U6576 ( .A1(n6414), .A2(n5063), .ZN(n8765) );
  NAND2_X1 U6577 ( .A1(n7802), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U6578 ( .A1(n7651), .A2(n7652), .ZN(n7799) );
  OAI21_X1 U6579 ( .B1(n8260), .B2(n8259), .A(n4980), .ZN(n4985) );
  NOR2_X1 U6580 ( .A1(n4996), .A2(n8669), .ZN(n8649) );
  AOI21_X1 U6581 ( .B1(n8590), .B2(n8588), .A(n8589), .ZN(n8599) );
  OR2_X1 U6582 ( .A1(n8669), .A2(n8668), .ZN(n4657) );
  NAND2_X1 U6583 ( .A1(n9604), .A2(n5173), .ZN(n5172) );
  AND2_X2 U6584 ( .A1(n5187), .A2(n4483), .ZN(n9786) );
  NAND2_X1 U6585 ( .A1(n9413), .A2(n7354), .ZN(n9427) );
  NAND2_X1 U6586 ( .A1(n9398), .A2(n7352), .ZN(n9414) );
  NOR2_X1 U6587 ( .A1(n7981), .A2(n7980), .ZN(n8124) );
  NAND2_X1 U6588 ( .A1(n9427), .A2(n9428), .ZN(n9426) );
  NAND2_X1 U6589 ( .A1(n4724), .A2(n6542), .ZN(n6632) );
  AOI21_X1 U6590 ( .B1(n4754), .B2(n4755), .A(n4752), .ZN(n6483) );
  NAND2_X1 U6591 ( .A1(n6498), .A2(n4661), .ZN(n6500) );
  INV_X1 U6592 ( .A(n4662), .ZN(n4661) );
  AOI21_X1 U6593 ( .B1(n4665), .B2(n4517), .A(n6623), .ZN(n6628) );
  NAND2_X1 U6594 ( .A1(n6484), .A2(n6634), .ZN(n4663) );
  NAND2_X1 U6595 ( .A1(n6580), .A2(n6577), .ZN(n7670) );
  NAND2_X1 U6596 ( .A1(n6458), .A2(n6457), .ZN(n4755) );
  AOI21_X1 U6597 ( .B1(n6492), .B2(n6489), .A(n4465), .ZN(n6490) );
  NAND2_X1 U6598 ( .A1(n4664), .A2(n4663), .ZN(n6492) );
  NOR4_X1 U6599 ( .A1(n9553), .A2(n9560), .A3(n9571), .A4(n6591), .ZN(n6592)
         );
  NOR4_X1 U6600 ( .A1(n9754), .A2(n6587), .A3(n9736), .A4(n9981), .ZN(n6588)
         );
  AND3_X1 U6601 ( .A1(n4670), .A2(n6583), .A3(n4666), .ZN(n6585) );
  NAND3_X1 U6602 ( .A1(n4669), .A2(n8059), .A3(n4668), .ZN(n4667) );
  NAND3_X1 U6603 ( .A1(n5399), .A2(n5402), .A3(n5419), .ZN(n4671) );
  NAND2_X1 U6604 ( .A1(n5546), .A2(n4700), .ZN(n5142) );
  INV_X1 U6605 ( .A(n6931), .ZN(n4676) );
  NAND2_X1 U6606 ( .A1(n4866), .A2(n8266), .ZN(n6902) );
  NAND2_X1 U6607 ( .A1(n5114), .A2(n5115), .ZN(n5112) );
  NAND2_X1 U6608 ( .A1(n5820), .A2(n5819), .ZN(n9532) );
  INV_X1 U6609 ( .A(n4741), .ZN(n5786) );
  NAND2_X1 U6610 ( .A1(n6991), .A2(n6992), .ZN(n5110) );
  NOR2_X2 U6611 ( .A1(n5719), .A2(n9171), .ZN(n4677) );
  AOI21_X1 U6612 ( .B1(n5139), .B2(n5140), .A(n5136), .ZN(n5135) );
  NAND2_X1 U6613 ( .A1(n6809), .A2(n4480), .ZN(n4933) );
  INV_X1 U6614 ( .A(n7483), .ZN(n4678) );
  NAND2_X1 U6615 ( .A1(n7169), .A2(n4997), .ZN(n7483) );
  AOI21_X1 U6616 ( .B1(n4929), .B2(n4934), .A(n6815), .ZN(n6822) );
  OAI21_X1 U6617 ( .B1(n6792), .B2(n4923), .A(n4440), .ZN(n6798) );
  OAI21_X1 U6618 ( .B1(n6446), .B2(n6449), .A(n4679), .ZN(n6450) );
  AND2_X1 U6619 ( .A1(n6650), .A2(n6634), .ZN(n4679) );
  NAND2_X1 U6620 ( .A1(n6573), .A2(n6572), .ZN(n4701) );
  NAND2_X1 U6621 ( .A1(n4684), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4685) );
  XNOR2_X2 U6622 ( .A(n5715), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5934) );
  INV_X1 U6623 ( .A(n9947), .ZN(n4684) );
  NAND2_X1 U6624 ( .A1(n4687), .A2(n4686), .ZN(n9494) );
  NOR2_X1 U6625 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  AOI21_X1 U6626 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7983), .A(n7979), .ZN(
        n7981) );
  NAND3_X1 U6627 ( .A1(n4964), .A2(n4963), .A3(n6448), .ZN(n6445) );
  NAND2_X1 U6628 ( .A1(n7573), .A2(n7439), .ZN(n7440) );
  NAND2_X1 U6629 ( .A1(n4989), .A2(n7914), .ZN(n4990) );
  NAND2_X1 U6630 ( .A1(n8692), .A2(n8691), .ZN(n8693) );
  AOI21_X1 U6631 ( .B1(n7508), .B2(n7507), .A(n6927), .ZN(n9208) );
  NAND2_X1 U6632 ( .A1(n6808), .A2(n6807), .ZN(n6809) );
  NAND2_X1 U6633 ( .A1(n5248), .A2(n5402), .ZN(n4848) );
  OAI21_X1 U6634 ( .B1(n6822), .B2(n8736), .A(n4491), .ZN(n4811) );
  NAND2_X1 U6635 ( .A1(n5263), .A2(n5092), .ZN(n5091) );
  NAND2_X1 U6636 ( .A1(n9426), .A2(n7355), .ZN(n9441) );
  NOR2_X1 U6637 ( .A1(n7524), .A2(n7523), .ZN(n7674) );
  NAND2_X1 U6638 ( .A1(n9414), .A2(n9415), .ZN(n9413) );
  INV_X1 U6639 ( .A(n4685), .ZN(n9945) );
  NAND2_X1 U6640 ( .A1(n6338), .A2(n6340), .ZN(n6337) );
  NAND3_X1 U6641 ( .A1(n4688), .A2(n6799), .A3(n6798), .ZN(n6803) );
  NAND4_X1 U6642 ( .A1(n6797), .A2(n6795), .A3(n6796), .A4(n7293), .ZN(n4688)
         );
  OR2_X1 U6643 ( .A1(n5247), .A2(SI_1_), .ZN(n5399) );
  NOR2_X2 U6644 ( .A1(n6919), .A2(n6918), .ZN(n9338) );
  NAND2_X1 U6645 ( .A1(n4694), .A2(n4693), .ZN(n4692) );
  OR2_X1 U6646 ( .A1(n6538), .A2(n6537), .ZN(n4743) );
  NAND2_X1 U6647 ( .A1(n7670), .A2(n5849), .ZN(n6643) );
  XNOR2_X1 U6648 ( .A(n9501), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U6649 ( .A1(n6643), .A2(n6648), .ZN(n5850) );
  NAND2_X1 U6650 ( .A1(n5156), .A2(n5153), .ZN(n5954) );
  NAND2_X1 U6651 ( .A1(n5917), .A2(n5918), .ZN(n4847) );
  NAND2_X1 U6652 ( .A1(n4844), .A2(n5344), .ZN(n5806) );
  OAI21_X1 U6653 ( .B1(n7297), .B2(n4703), .A(n4702), .ZN(n5251) );
  AND2_X1 U6654 ( .A1(n6448), .A2(n6447), .ZN(n6650) );
  AND3_X2 U6655 ( .A1(n5977), .A2(n7433), .A3(n5976), .ZN(n6090) );
  NAND2_X1 U6656 ( .A1(n4708), .A2(n4707), .ZN(n7749) );
  NAND2_X1 U6657 ( .A1(n4817), .A2(n6740), .ZN(n7728) );
  NAND3_X1 U6658 ( .A1(n6726), .A2(n6730), .A3(n8914), .ZN(n6399) );
  NAND4_X1 U6659 ( .A1(n6090), .A2(n5225), .A3(n10214), .A4(n5978), .ZN(n6000)
         );
  OAI21_X2 U6660 ( .B1(n6888), .B2(n6887), .A(n4456), .ZN(n7142) );
  XNOR2_X1 U6661 ( .A(n8711), .B(n8710), .ZN(n4714) );
  NAND2_X1 U6662 ( .A1(n7749), .A2(n6737), .ZN(n4817) );
  NOR2_X1 U6663 ( .A1(n6824), .A2(n6823), .ZN(n4810) );
  NAND2_X2 U6664 ( .A1(n4710), .A2(n5904), .ZN(n7291) );
  NAND2_X1 U6665 ( .A1(n9164), .A2(n5130), .ZN(n5128) );
  NAND2_X1 U6666 ( .A1(n9254), .A2(n7038), .ZN(n9164) );
  NAND2_X1 U6667 ( .A1(n5084), .A2(n5087), .ZN(n9233) );
  NAND2_X1 U6668 ( .A1(n8485), .A2(n7236), .ZN(n8442) );
  AOI21_X1 U6669 ( .B1(n4967), .B2(n6499), .A(n5868), .ZN(n4965) );
  OAI21_X1 U6670 ( .B1(n8671), .B2(n8672), .A(n8670), .ZN(n4715) );
  NAND2_X1 U6671 ( .A1(n4969), .A2(n7553), .ZN(n4970) );
  OR2_X1 U6672 ( .A1(n7440), .A2(n7506), .ZN(n7441) );
  NAND2_X1 U6673 ( .A1(n9399), .A2(n9404), .ZN(n9398) );
  INV_X1 U6674 ( .A(n4994), .ZN(n8667) );
  NAND2_X1 U6675 ( .A1(n5197), .A2(n5195), .ZN(n5711) );
  NAND2_X1 U6676 ( .A1(n6361), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6003) );
  NOR2_X2 U6677 ( .A1(n6362), .A2(n5975), .ZN(n5978) );
  INV_X1 U6678 ( .A(n6377), .ZN(n6375) );
  OAI21_X1 U6679 ( .B1(n8364), .B2(n7202), .A(n7201), .ZN(n7205) );
  NAND2_X1 U6680 ( .A1(n5435), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6681 ( .A1(n6632), .A2(n9507), .ZN(n4846) );
  NAND2_X1 U6682 ( .A1(n6516), .A2(n4717), .ZN(n6518) );
  NAND2_X1 U6683 ( .A1(n6500), .A2(n9681), .ZN(n6516) );
  NAND2_X1 U6684 ( .A1(n4718), .A2(n4445), .ZN(n4963) );
  NAND2_X2 U6685 ( .A1(n7320), .A2(n4815), .ZN(n5563) );
  NAND2_X2 U6686 ( .A1(n9233), .A2(n9234), .ZN(n9232) );
  XNOR2_X1 U6687 ( .A(n6944), .B(n9179), .ZN(n8070) );
  INV_X4 U6688 ( .A(n6965), .ZN(n9175) );
  NAND2_X1 U6689 ( .A1(n5684), .A2(n5360), .ZN(n5838) );
  NOR2_X1 U6690 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  NAND4_X1 U6691 ( .A1(n4744), .A2(n4743), .A3(n6595), .A4(n4739), .ZN(n4724)
         );
  NAND2_X1 U6692 ( .A1(n4859), .A2(n4860), .ZN(n5756) );
  NAND2_X1 U6693 ( .A1(n9965), .A2(n9966), .ZN(n4736) );
  NAND2_X1 U6694 ( .A1(n7655), .A2(n7653), .ZN(n7651) );
  NOR2_X1 U6695 ( .A1(n8600), .A2(n8618), .ZN(n8635) );
  NAND2_X1 U6696 ( .A1(n7799), .A2(n7798), .ZN(n7800) );
  NAND3_X1 U6697 ( .A1(n6698), .A2(n6699), .A3(n6697), .ZN(P1_U3242) );
  INV_X1 U6698 ( .A(n6543), .ZN(n4739) );
  OAI21_X1 U6699 ( .B1(n9531), .B2(n9881), .A(n4937), .ZN(n5914) );
  NAND2_X1 U6700 ( .A1(n6530), .A2(n4750), .ZN(n4745) );
  NAND2_X1 U6701 ( .A1(n4755), .A2(n6469), .ZN(n6482) );
  NOR2_X1 U6702 ( .A1(n4760), .A2(n5367), .ZN(n4759) );
  NAND3_X1 U6703 ( .A1(n9118), .A2(P2_REG3_REG_1__SCAN_IN), .A3(n4393), .ZN(
        n5044) );
  NOR2_X2 U6704 ( .A1(n9118), .A2(n4393), .ZN(n6035) );
  NAND4_X1 U6705 ( .A1(n6090), .A2(n4413), .A3(n5225), .A4(n5978), .ZN(n9110)
         );
  NAND2_X1 U6706 ( .A1(n4765), .A2(n4766), .ZN(n7941) );
  NAND3_X1 U6707 ( .A1(n4405), .A2(n6112), .A3(n5047), .ZN(n4765) );
  NAND2_X1 U6708 ( .A1(n8902), .A2(n8901), .ZN(n8869) );
  NAND2_X1 U6709 ( .A1(n4795), .A2(n6783), .ZN(n4794) );
  NAND2_X1 U6710 ( .A1(n4796), .A2(n6778), .ZN(n4795) );
  NAND2_X1 U6711 ( .A1(n6774), .A2(n4487), .ZN(n4796) );
  NAND3_X1 U6712 ( .A1(n6729), .A2(n6728), .A3(n8992), .ZN(n4800) );
  NAND3_X1 U6713 ( .A1(n4806), .A2(n4494), .A3(n4801), .ZN(n6770) );
  NAND3_X1 U6714 ( .A1(n4803), .A2(n4928), .A3(n4802), .ZN(n4801) );
  NAND3_X1 U6715 ( .A1(n4924), .A2(n4927), .A3(n4925), .ZN(n4806) );
  NAND2_X1 U6716 ( .A1(n4816), .A2(n4813), .ZN(n4812) );
  NAND2_X2 U6717 ( .A1(n9125), .A2(n6342), .ZN(n6034) );
  NAND2_X1 U6718 ( .A1(n7157), .A2(n4821), .ZN(n4819) );
  INV_X1 U6719 ( .A(n4818), .ZN(P2_U3488) );
  INV_X1 U6720 ( .A(n6417), .ZN(n4824) );
  NAND2_X2 U6721 ( .A1(n8843), .A2(n4408), .ZN(n8819) );
  NAND2_X1 U6722 ( .A1(n6405), .A2(n6764), .ZN(n8162) );
  NAND3_X1 U6723 ( .A1(n4841), .A2(n6405), .A3(n6764), .ZN(n4840) );
  INV_X1 U6724 ( .A(n4842), .ZN(n4841) );
  INV_X1 U6725 ( .A(n5059), .ZN(n4842) );
  NAND2_X1 U6726 ( .A1(n5806), .A2(n5807), .ZN(n4843) );
  NAND2_X1 U6727 ( .A1(n5244), .A2(n5245), .ZN(n4849) );
  NAND2_X1 U6728 ( .A1(n5712), .A2(n4853), .ZN(n4850) );
  NAND2_X1 U6729 ( .A1(n4850), .A2(n4851), .ZN(n5334) );
  NAND2_X1 U6730 ( .A1(n5712), .A2(n4863), .ZN(n4859) );
  NAND2_X1 U6731 ( .A1(n4865), .A2(n4490), .ZN(n5297) );
  NAND4_X1 U6732 ( .A1(n4450), .A2(n6886), .A3(n6885), .A4(n4867), .ZN(n4866)
         );
  AND2_X1 U6733 ( .A1(n6839), .A2(n4489), .ZN(n4867) );
  NAND2_X1 U6734 ( .A1(n6281), .A2(n6280), .ZN(n6291) );
  NAND2_X1 U6735 ( .A1(n6231), .A2(n4505), .ZN(n6258) );
  NOR2_X1 U6736 ( .A1(n8728), .A2(n4876), .ZN(n6882) );
  NAND3_X1 U6737 ( .A1(n6018), .A2(n5959), .A3(n5958), .ZN(n6081) );
  OR2_X1 U6738 ( .A1(n4395), .A2(n7438), .ZN(n7439) );
  XNOR2_X1 U6739 ( .A(n7584), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7575) );
  NOR2_X1 U6740 ( .A1(n4395), .A2(n7420), .ZN(n4899) );
  INV_X1 U6741 ( .A(n4395), .ZN(n4902) );
  NAND3_X1 U6742 ( .A1(n6015), .A2(n6016), .A3(n4904), .ZN(n6048) );
  NAND2_X1 U6743 ( .A1(n6043), .A2(n4395), .ZN(n4904) );
  NAND3_X2 U6744 ( .A1(n6032), .A2(n6031), .A3(n4915), .ZN(n6723) );
  AND2_X1 U6745 ( .A1(n6030), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U6746 ( .A1(n6862), .A2(n6724), .ZN(n4918) );
  NAND2_X1 U6747 ( .A1(n4921), .A2(n4918), .ZN(n4920) );
  NAND3_X1 U6748 ( .A1(n4920), .A2(n6726), .A3(n4402), .ZN(n4919) );
  NAND2_X1 U6749 ( .A1(n4919), .A2(n8987), .ZN(n6725) );
  INV_X1 U6750 ( .A(n8914), .ZN(n4921) );
  NAND2_X1 U6751 ( .A1(n6750), .A2(n4402), .ZN(n4927) );
  INV_X1 U6752 ( .A(n9110), .ZN(n5990) );
  NAND2_X1 U6753 ( .A1(n4941), .A2(n4938), .ZN(n8228) );
  NAND2_X1 U6754 ( .A1(n4954), .A2(n4958), .ZN(n9592) );
  NAND2_X1 U6755 ( .A1(n9629), .A2(n4960), .ZN(n4954) );
  INV_X1 U6756 ( .A(n4958), .ZN(n4957) );
  NAND2_X1 U6757 ( .A1(n5850), .A2(n4962), .ZN(n4964) );
  NAND2_X1 U6758 ( .A1(n5850), .A2(n6646), .ZN(n6446) );
  INV_X1 U6759 ( .A(n7558), .ZN(n4969) );
  INV_X1 U6760 ( .A(n7606), .ZN(n4971) );
  NOR2_X1 U6761 ( .A1(n4985), .A2(n4984), .ZN(n4983) );
  NAND3_X1 U6762 ( .A1(n7441), .A2(n7445), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n7442) );
  NAND2_X1 U6763 ( .A1(n7441), .A2(n7445), .ZN(n7493) );
  NAND2_X1 U6764 ( .A1(n7442), .A2(n7445), .ZN(n4987) );
  NAND2_X1 U6765 ( .A1(n4990), .A2(n7913), .ZN(n8187) );
  NAND2_X1 U6766 ( .A1(n4992), .A2(n4991), .ZN(n8692) );
  INV_X1 U6767 ( .A(n4995), .ZN(n4992) );
  OAI21_X1 U6768 ( .B1(n8669), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8668), .ZN(
        n4995) );
  AND2_X1 U6769 ( .A1(n8648), .A2(n8674), .ZN(n4996) );
  OAI22_X1 U6770 ( .A1(n7912), .A2(n10264), .B1(n7911), .B2(n7910), .ZN(n8183)
         );
  AOI22_X1 U6771 ( .A1(n7641), .A2(P2_REG1_REG_7__SCAN_IN), .B1(n7640), .B2(
        n7639), .ZN(n7796) );
  NAND2_X4 U6772 ( .A1(n9935), .A2(n5871), .ZN(n7320) );
  INV_X1 U6773 ( .A(n4999), .ZN(n4998) );
  NAND2_X1 U6774 ( .A1(n4999), .A2(n4392), .ZN(n4997) );
  INV_X1 U6775 ( .A(n6396), .ZN(n9007) );
  OAI211_X1 U6776 ( .C1(n4516), .C2(n7535), .A(n7534), .B(n8500), .ZN(n7536)
         );
  NAND2_X1 U6777 ( .A1(n7233), .A2(n7232), .ZN(n8485) );
  NAND2_X1 U6778 ( .A1(n7941), .A2(n6125), .ZN(n5024) );
  NAND2_X1 U6779 ( .A1(n5028), .A2(n5029), .ZN(n8809) );
  INV_X1 U6780 ( .A(n8861), .ZN(n5041) );
  NAND2_X1 U6781 ( .A1(n5043), .A2(n5042), .ZN(n5045) );
  NAND2_X1 U6782 ( .A1(n6076), .A2(n5046), .ZN(n5047) );
  XNOR2_X1 U6783 ( .A(n8729), .B(n8728), .ZN(n5049) );
  NAND2_X1 U6784 ( .A1(n5062), .A2(n5061), .ZN(n7820) );
  NAND2_X1 U6785 ( .A1(n8819), .A2(n6793), .ZN(n6411) );
  NOR2_X2 U6786 ( .A1(n8175), .A2(n5064), .ZN(n8233) );
  OAI21_X2 U6787 ( .B1(n8868), .B2(n6782), .A(n6779), .ZN(n8856) );
  XNOR2_X2 U6788 ( .A(n7142), .B(n7151), .ZN(n8333) );
  NOR2_X2 U6789 ( .A1(n9759), .A2(n5069), .ZN(n9683) );
  AND2_X2 U6790 ( .A1(n9593), .A2(n5077), .ZN(n9563) );
  XNOR2_X2 U6791 ( .A(n5082), .B(n5370), .ZN(n5871) );
  NAND2_X2 U6792 ( .A1(n5083), .A2(n5373), .ZN(n9935) );
  NAND2_X1 U6793 ( .A1(n5296), .A2(n5297), .ZN(n5664) );
  NAND2_X1 U6794 ( .A1(n5441), .A2(n5220), .ZN(n5093) );
  NAND2_X1 U6795 ( .A1(n5103), .A2(n5094), .ZN(P1_U3220) );
  NOR2_X1 U6796 ( .A1(n5098), .A2(n5095), .ZN(n5094) );
  NAND2_X1 U6797 ( .A1(n9232), .A2(n5100), .ZN(n5103) );
  NAND2_X1 U6798 ( .A1(n9155), .A2(n6991), .ZN(n5113) );
  NAND2_X1 U6799 ( .A1(n6961), .A2(n7959), .ZN(n8105) );
  NOR2_X1 U6800 ( .A1(n8106), .A2(n6963), .ZN(n5121) );
  INV_X1 U6801 ( .A(n7053), .ZN(n5131) );
  NAND2_X1 U6802 ( .A1(n5526), .A2(n5139), .ZN(n5137) );
  OAI21_X1 U6803 ( .B1(n5526), .B2(n5140), .A(n5139), .ZN(n5562) );
  NAND2_X1 U6804 ( .A1(n5906), .A2(n5151), .ZN(n5886) );
  NAND2_X1 U6805 ( .A1(n5906), .A2(n5146), .ZN(n5145) );
  NAND2_X1 U6806 ( .A1(n5906), .A2(n5882), .ZN(n5884) );
  NAND2_X1 U6807 ( .A1(n5161), .A2(n5164), .ZN(n5295) );
  NAND2_X1 U6808 ( .A1(n5594), .A2(n5168), .ZN(n5161) );
  NAND2_X1 U6809 ( .A1(n5174), .A2(n5172), .ZN(n9554) );
  NAND3_X1 U6810 ( .A1(n5176), .A2(n5178), .A3(n4439), .ZN(n5175) );
  OAI21_X1 U6811 ( .B1(n9605), .B2(n5178), .A(n5176), .ZN(n9557) );
  OR2_X1 U6812 ( .A1(n9320), .A2(n9815), .ZN(n5186) );
  NAND2_X1 U6813 ( .A1(n6648), .A2(n6646), .ZN(n6581) );
  AND4_X2 U6814 ( .A1(n5392), .A2(n5393), .A3(n5395), .A4(n5394), .ZN(n9212)
         );
  NOR2_X1 U6815 ( .A1(n9786), .A2(n5188), .ZN(n9774) );
  NAND2_X1 U6816 ( .A1(n8166), .A2(n5192), .ZN(n5189) );
  NAND2_X1 U6817 ( .A1(n5189), .A2(n5190), .ZN(n8227) );
  NAND2_X1 U6818 ( .A1(n9716), .A2(n4488), .ZN(n5197) );
  NAND2_X1 U6819 ( .A1(n5201), .A2(n5661), .ZN(n9703) );
  NAND2_X1 U6820 ( .A1(n5204), .A2(n5203), .ZN(n5646) );
  NAND2_X1 U6821 ( .A1(n9648), .A2(n5210), .ZN(n5205) );
  NAND2_X1 U6822 ( .A1(n5205), .A2(n5207), .ZN(n9620) );
  INV_X1 U6823 ( .A(n5841), .ZN(n5212) );
  INV_X1 U6824 ( .A(n8527), .ZN(n8528) );
  INV_X1 U6825 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6340) );
  AND2_X2 U6826 ( .A1(n5043), .A2(n9118), .ZN(n6036) );
  OAI21_X1 U6827 ( .B1(n9782), .B2(n9781), .A(n9780), .ZN(n9783) );
  NOR4_X2 U6828 ( .A1(n6637), .A2(n6597), .A3(n6596), .A4(n6629), .ZN(n6623)
         );
  INV_X1 U6829 ( .A(n6632), .ZN(n6573) );
  NAND2_X1 U6830 ( .A1(n8517), .A2(n7246), .ZN(n7248) );
  AOI21_X1 U6831 ( .B1(n7153), .B2(n5217), .A(n7152), .ZN(n7154) );
  OR2_X1 U6832 ( .A1(n7153), .A2(n4486), .ZN(n7155) );
  INV_X1 U6833 ( .A(n6838), .ZN(n8336) );
  NAND2_X1 U6834 ( .A1(n9545), .A2(n9792), .ZN(n9534) );
  XNOR2_X1 U6835 ( .A(n5821), .B(n5822), .ZN(n9124) );
  NAND2_X1 U6836 ( .A1(n6398), .A2(n7530), .ZN(n10104) );
  CLKBUF_X1 U6837 ( .A(n8281), .Z(n9974) );
  NAND2_X1 U6838 ( .A1(n9117), .A2(n5923), .ZN(n5925) );
  BUF_X4 U6839 ( .A(n6036), .Z(n6847) );
  AND2_X1 U6840 ( .A1(n7418), .A2(n4387), .ZN(n8714) );
  OAI211_X1 U6841 ( .C1(n7866), .C2(n5501), .A(n8000), .B(n5500), .ZN(n5503)
         );
  OR2_X2 U6842 ( .A1(n6027), .A2(n6026), .ZN(n10140) );
  INV_X1 U6843 ( .A(n9683), .ZN(n9706) );
  NAND2_X1 U6844 ( .A1(n9683), .A2(n5866), .ZN(n9685) );
  CLKBUF_X1 U6845 ( .A(n5871), .Z(n8317) );
  NAND2_X1 U6846 ( .A1(n7297), .A2(n7298), .ZN(n5245) );
  OAI21_X1 U6847 ( .B1(n7297), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n5241), .ZN(
        n5242) );
  NAND2_X1 U6848 ( .A1(n7297), .A2(n5413), .ZN(n5241) );
  OAI21_X1 U6849 ( .B1(n7297), .B2(n5239), .A(n5238), .ZN(n5247) );
  NAND2_X1 U6850 ( .A1(n5536), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5409) );
  INV_X1 U6851 ( .A(n5536), .ZN(n5875) );
  AND2_X1 U6852 ( .A1(n7321), .A2(n4530), .ZN(n5216) );
  AND2_X1 U6853 ( .A1(n7151), .A2(n5229), .ZN(n5217) );
  OR2_X1 U6854 ( .A1(n10128), .A2(n6712), .ZN(n5218) );
  AND2_X1 U6855 ( .A1(n7680), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5219) );
  AND2_X1 U6856 ( .A1(n5437), .A2(n5473), .ZN(n5220) );
  OR2_X1 U6857 ( .A1(n8336), .A2(n9100), .ZN(n5221) );
  AND2_X1 U6858 ( .A1(n7005), .A2(n7004), .ZN(n5223) );
  AND2_X1 U6859 ( .A1(n9453), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5226) );
  INV_X1 U6860 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6374) );
  CLKBUF_X3 U6861 ( .A(n6941), .Z(n9181) );
  NOR2_X1 U6862 ( .A1(n7150), .A2(n7149), .ZN(n5227) );
  INV_X1 U6863 ( .A(n6889), .ZN(n6886) );
  AND3_X1 U6864 ( .A1(n7257), .A2(n7282), .A3(n8500), .ZN(n5228) );
  AND2_X1 U6865 ( .A1(n7146), .A2(n10111), .ZN(n5229) );
  AND2_X1 U6866 ( .A1(n6715), .A2(n6714), .ZN(n5230) );
  AND2_X2 U6867 ( .A1(n5913), .A2(n5930), .ZN(n10090) );
  AND2_X1 U6868 ( .A1(n5266), .A2(n5484), .ZN(n5234) );
  AND2_X1 U6869 ( .A1(n8871), .A2(n6199), .ZN(n5235) );
  AND2_X1 U6870 ( .A1(n8870), .A2(n8872), .ZN(n5236) );
  INV_X2 U6871 ( .A(n10164), .ZN(n10166) );
  OAI21_X1 U6872 ( .B1(n6800), .B2(n4402), .A(n8787), .ZN(n6801) );
  INV_X1 U6873 ( .A(n6801), .ZN(n6802) );
  MUX2_X1 U6874 ( .A(n6806), .B(n6805), .S(n7293), .Z(n6807) );
  INV_X1 U6875 ( .A(n8897), .ZN(n6198) );
  INV_X1 U6876 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5360) );
  INV_X1 U6877 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5974) );
  INV_X1 U6878 ( .A(n8454), .ZN(n7178) );
  INV_X1 U6879 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6712) );
  OR2_X1 U6880 ( .A1(n7285), .A2(n8730), .ZN(n7143) );
  OR2_X1 U6881 ( .A1(n9050), .A2(n8802), .ZN(n6265) );
  NOR2_X1 U6882 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5976) );
  NOR2_X1 U6883 ( .A1(n6570), .A2(n6569), .ZN(n6571) );
  NAND2_X1 U6884 ( .A1(n7297), .A2(n5257), .ZN(n5258) );
  NAND2_X1 U6885 ( .A1(n8366), .A2(n8547), .ZN(n7194) );
  INV_X1 U6886 ( .A(n6839), .ZN(n6895) );
  NAND2_X1 U6887 ( .A1(n7801), .A2(n7911), .ZN(n7802) );
  NOR2_X1 U6888 ( .A1(n8587), .A2(n8586), .ZN(n8598) );
  NAND2_X1 U6889 ( .A1(n6398), .A2(n6397), .ZN(n6730) );
  NAND2_X1 U6890 ( .A1(n6063), .A2(n6062), .ZN(n7754) );
  INV_X1 U6891 ( .A(n6979), .ZN(n6980) );
  NAND2_X1 U6892 ( .A1(n9195), .A2(n6974), .ZN(n6975) );
  INV_X1 U6893 ( .A(n9383), .ZN(n9521) );
  INV_X1 U6894 ( .A(n5740), .ZN(n5319) );
  NAND2_X1 U6895 ( .A1(n5308), .A2(SI_18_), .ZN(n5309) );
  INV_X1 U6896 ( .A(n5648), .ZN(n5294) );
  NAND2_X1 U6897 ( .A1(n5282), .A2(n10414), .ZN(n5283) );
  INV_X1 U6898 ( .A(n8531), .ZN(n7210) );
  INV_X1 U6899 ( .A(n7200), .ZN(n7201) );
  INV_X1 U6900 ( .A(n9027), .ZN(n7243) );
  INV_X1 U6901 ( .A(n4399), .ZN(n6327) );
  INV_X1 U6902 ( .A(n8188), .ZN(n8189) );
  INV_X1 U6903 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5962) );
  INV_X1 U6904 ( .A(n6034), .ZN(n6043) );
  INV_X1 U6905 ( .A(n8014), .ZN(n8018) );
  OR2_X1 U6906 ( .A1(n6425), .A2(n6424), .ZN(n7271) );
  NOR2_X1 U6907 ( .A1(n6007), .A2(n6006), .ZN(n6356) );
  INV_X1 U6908 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U6909 ( .A1(n6978), .A2(n6980), .ZN(n6981) );
  INV_X1 U6910 ( .A(n4389), .ZN(n5829) );
  INV_X1 U6911 ( .A(n9600), .ZN(n9819) );
  NOR2_X1 U6912 ( .A1(n6578), .A2(n6579), .ZN(n6577) );
  NAND2_X1 U6913 ( .A1(n5302), .A2(n5301), .ZN(n5305) );
  AND2_X1 U6914 ( .A1(n5290), .A2(n5613), .ZN(n5291) );
  NAND2_X1 U6915 ( .A1(n5276), .A2(SI_10_), .ZN(n5280) );
  NAND2_X1 U6916 ( .A1(n7213), .A2(n8544), .ZN(n7214) );
  INV_X1 U6917 ( .A(n8904), .ZN(n8478) );
  OR2_X1 U6918 ( .A1(P2_U3150), .A2(n7400), .ZN(n8622) );
  NAND2_X1 U6919 ( .A1(n6267), .A2(n6266), .ZN(n6416) );
  OR2_X1 U6920 ( .A1(n6861), .A2(n6860), .ZN(n7940) );
  OR2_X1 U6921 ( .A1(n10151), .A2(n6857), .ZN(n10121) );
  OR2_X1 U6922 ( .A1(n6377), .A2(n6388), .ZN(n6426) );
  INV_X1 U6923 ( .A(n8550), .ZN(n7886) );
  AND2_X1 U6924 ( .A1(n7164), .A2(n8215), .ZN(n6857) );
  INV_X1 U6925 ( .A(n8990), .ZN(n7945) );
  NAND2_X1 U6926 ( .A1(n6373), .A2(n6376), .ZN(n6377) );
  INV_X1 U6927 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6354) );
  INV_X1 U6928 ( .A(n9540), .ZN(n9792) );
  INV_X1 U6929 ( .A(n9365), .ZN(n9376) );
  OR2_X1 U6930 ( .A1(n5775), .A2(n7703), .ZN(n5393) );
  INV_X1 U6931 ( .A(n7514), .ZN(n9453) );
  INV_X1 U6932 ( .A(n9985), .ZN(n9757) );
  AOI21_X1 U6933 ( .B1(n5954), .B2(n6594), .A(n5953), .ZN(n5955) );
  INV_X1 U6934 ( .A(n10053), .ZN(n10082) );
  AND2_X1 U6935 ( .A1(n6914), .A2(n6645), .ZN(n7318) );
  OR2_X1 U6936 ( .A1(n5598), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5618) );
  INV_X1 U6937 ( .A(n8790), .ZN(n8761) );
  INV_X1 U6938 ( .A(n8535), .ZN(n8487) );
  AND2_X1 U6939 ( .A1(n6852), .A2(n6851), .ZN(n6891) );
  AND2_X1 U6940 ( .A1(n6255), .A2(n6254), .ZN(n8468) );
  INV_X1 U6941 ( .A(n8705), .ZN(n8634) );
  INV_X1 U6942 ( .A(n8717), .ZN(n8670) );
  INV_X1 U6943 ( .A(n8971), .ZN(n8967) );
  AND2_X1 U6944 ( .A1(n6788), .A2(n6796), .ZN(n8823) );
  NAND2_X1 U6945 ( .A1(n8272), .A2(n8266), .ZN(n10151) );
  AND2_X1 U6946 ( .A1(n8272), .A2(n6857), .ZN(n9008) );
  INV_X1 U6947 ( .A(n10151), .ZN(n10141) );
  AND2_X1 U6948 ( .A1(n7338), .A2(n7292), .ZN(n7333) );
  AND2_X1 U6949 ( .A1(n6093), .A2(n6114), .ZN(n7611) );
  INV_X1 U6950 ( .A(n9349), .ZN(n9372) );
  INV_X1 U6951 ( .A(n9368), .ZN(n9378) );
  AOI21_X1 U6952 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n7407), .A(n7406), .ZN(
        n7410) );
  NAND2_X1 U6953 ( .A1(n6605), .A2(n6611), .ZN(n9560) );
  INV_X1 U6954 ( .A(n9743), .ZN(n9977) );
  INV_X1 U6955 ( .A(n9715), .ZN(n9729) );
  NAND2_X1 U6956 ( .A1(n7120), .A2(n7478), .ZN(n10071) );
  AND2_X1 U6957 ( .A1(n6569), .A2(n6635), .ZN(n9881) );
  INV_X1 U6958 ( .A(n9881), .ZN(n10061) );
  AND2_X1 U6959 ( .A1(n8317), .A2(n7318), .ZN(n9986) );
  AND2_X1 U6960 ( .A1(n7291), .A2(n7289), .ZN(n9923) );
  NAND2_X1 U6961 ( .A1(n5438), .A2(n5439), .ZN(n5442) );
  INV_X1 U6962 ( .A(n8500), .ZN(n8529) );
  INV_X1 U6963 ( .A(n8468), .ZN(n8812) );
  INV_X1 U6964 ( .A(n8887), .ZN(n8545) );
  INV_X1 U6965 ( .A(n8707), .ZN(n8683) );
  NAND2_X1 U6966 ( .A1(n10128), .A2(n6709), .ZN(n8883) );
  INV_X2 U6967 ( .A(n10130), .ZN(n10128) );
  NAND2_X1 U6968 ( .A1(n10166), .A2(n10149), .ZN(n8972) );
  NAND2_X1 U6969 ( .A1(n10166), .A2(n10141), .ZN(n8971) );
  OR2_X1 U6970 ( .A1(n6705), .A2(n6394), .ZN(n10164) );
  NAND2_X1 U6971 ( .A1(n10157), .A2(n10149), .ZN(n9102) );
  AND2_X1 U6972 ( .A1(n7399), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7338) );
  NAND2_X1 U6973 ( .A1(n6377), .A2(n7333), .ZN(n7341) );
  INV_X1 U6974 ( .A(n6910), .ZN(n8272) );
  INV_X1 U6975 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7513) );
  INV_X1 U6976 ( .A(n9746), .ZN(n9895) );
  AND2_X1 U6977 ( .A1(n7119), .A2(n9671), .ZN(n9368) );
  INV_X1 U6978 ( .A(n9777), .ZN(n9789) );
  INV_X1 U6979 ( .A(n9725), .ZN(n9883) );
  NAND2_X1 U6980 ( .A1(n5950), .A2(n5846), .ZN(n9743) );
  INV_X1 U6981 ( .A(n9704), .ZN(n9765) );
  AND2_X2 U6982 ( .A1(n5913), .A2(n5910), .ZN(n10103) );
  INV_X1 U6983 ( .A(n10103), .ZN(n10101) );
  INV_X1 U6984 ( .A(n10090), .ZN(n10088) );
  INV_X1 U6985 ( .A(n10001), .ZN(n10002) );
  INV_X1 U6986 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8211) );
  INV_X1 U6987 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10386) );
  INV_X1 U6988 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7347) );
  INV_X1 U6989 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10212) );
  NAND2_X1 U6990 ( .A1(n6423), .A2(n6422), .ZN(P2_U3487) );
  NAND2_X1 U6991 ( .A1(n6438), .A2(n6437), .ZN(P2_U3455) );
  INV_X1 U6992 ( .A(n9391), .ZN(P1_U3973) );
  MUX2_X1 U6993 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n5914), .S(n10103), .Z(
        P1_U3550) );
  NAND2_X1 U6994 ( .A1(n7297), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5238) );
  INV_X1 U6995 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5240) );
  INV_X1 U6996 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5413) );
  NOR2_X1 U6997 ( .A1(n5242), .A2(n10345), .ZN(n5419) );
  INV_X1 U6998 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7305) );
  INV_X1 U6999 ( .A(SI_2_), .ZN(n5246) );
  INV_X1 U7000 ( .A(n5398), .ZN(n5248) );
  INV_X1 U7001 ( .A(n5251), .ZN(n5250) );
  INV_X1 U7002 ( .A(SI_3_), .ZN(n5249) );
  NAND2_X1 U7003 ( .A1(n5250), .A2(n5249), .ZN(n5437) );
  INV_X1 U7004 ( .A(SI_4_), .ZN(n10211) );
  INV_X1 U7005 ( .A(n5470), .ZN(n5252) );
  NAND2_X1 U7006 ( .A1(n5252), .A2(n5473), .ZN(n5255) );
  INV_X1 U7007 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U7008 ( .A1(n5254), .A2(SI_4_), .ZN(n5472) );
  INV_X1 U7009 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7309) );
  INV_X1 U7010 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5257) );
  INV_X1 U7011 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7323) );
  INV_X1 U7012 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5260) );
  MUX2_X1 U7013 ( .A(n7323), .B(n5260), .S(n7297), .Z(n5264) );
  INV_X1 U7014 ( .A(SI_6_), .ZN(n5261) );
  NAND2_X1 U7015 ( .A1(n5264), .A2(n5261), .ZN(n5485) );
  INV_X1 U7016 ( .A(n5262), .ZN(n5263) );
  NAND3_X1 U7017 ( .A1(n5485), .A2(n5480), .A3(SI_5_), .ZN(n5266) );
  INV_X1 U7018 ( .A(n5264), .ZN(n5265) );
  NAND2_X1 U7019 ( .A1(n5265), .A2(SI_6_), .ZN(n5484) );
  MUX2_X1 U7020 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4725), .Z(n5267) );
  OAI21_X1 U7021 ( .B1(n5267), .B2(SI_7_), .A(n5269), .ZN(n5517) );
  INV_X1 U7022 ( .A(n5517), .ZN(n5268) );
  INV_X1 U7023 ( .A(n5270), .ZN(n5272) );
  INV_X1 U7024 ( .A(SI_8_), .ZN(n5271) );
  NAND2_X1 U7025 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  MUX2_X1 U7026 ( .A(n10440), .B(n7347), .S(n7297), .Z(n5274) );
  INV_X1 U7027 ( .A(n5274), .ZN(n5275) );
  MUX2_X1 U7028 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4725), .Z(n5276) );
  INV_X1 U7029 ( .A(n5276), .ZN(n5278) );
  INV_X1 U7030 ( .A(SI_10_), .ZN(n5277) );
  NAND2_X1 U7031 ( .A1(n5278), .A2(n5277), .ZN(n5279) );
  NAND2_X1 U7032 ( .A1(n5280), .A2(n5279), .ZN(n5560) );
  MUX2_X1 U7033 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4725), .Z(n5281) );
  INV_X1 U7034 ( .A(n5281), .ZN(n5282) );
  MUX2_X1 U7035 ( .A(n7513), .B(n7516), .S(n4725), .Z(n5288) );
  MUX2_X1 U7036 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4725), .Z(n5286) );
  INV_X1 U7037 ( .A(n5286), .ZN(n5285) );
  INV_X1 U7038 ( .A(SI_12_), .ZN(n5284) );
  NAND2_X1 U7039 ( .A1(n5285), .A2(n5284), .ZN(n5592) );
  NAND2_X1 U7040 ( .A1(n5614), .A2(n5592), .ZN(n5292) );
  NAND2_X1 U7041 ( .A1(n5286), .A2(SI_12_), .ZN(n5611) );
  INV_X1 U7042 ( .A(n5611), .ZN(n5287) );
  NAND2_X1 U7043 ( .A1(n5287), .A2(n5614), .ZN(n5290) );
  INV_X1 U7044 ( .A(n5288), .ZN(n5289) );
  NAND2_X1 U7045 ( .A1(n5289), .A2(SI_13_), .ZN(n5613) );
  MUX2_X1 U7046 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4815), .Z(n5632) );
  INV_X1 U7047 ( .A(SI_15_), .ZN(n5293) );
  MUX2_X1 U7048 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4815), .Z(n5648) );
  NAND2_X1 U7049 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  MUX2_X1 U7050 ( .A(n7780), .B(n10386), .S(n4815), .Z(n5662) );
  INV_X1 U7051 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5300) );
  MUX2_X1 U7052 ( .A(n7907), .B(n5300), .S(n4815), .Z(n5302) );
  INV_X1 U7053 ( .A(SI_17_), .ZN(n5301) );
  INV_X1 U7054 ( .A(n5302), .ZN(n5303) );
  NAND2_X1 U7055 ( .A1(n5303), .A2(SI_17_), .ZN(n5304) );
  INV_X1 U7056 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5306) );
  MUX2_X1 U7057 ( .A(n7956), .B(n5306), .S(n4815), .Z(n5307) );
  INV_X1 U7058 ( .A(n5307), .ZN(n5308) );
  MUX2_X1 U7059 ( .A(n8208), .B(n10371), .S(n4815), .Z(n5312) );
  INV_X1 U7060 ( .A(SI_19_), .ZN(n5311) );
  INV_X1 U7061 ( .A(n5312), .ZN(n5313) );
  NAND2_X1 U7062 ( .A1(n5313), .A2(SI_19_), .ZN(n5314) );
  INV_X1 U7063 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8213) );
  MUX2_X1 U7064 ( .A(n8213), .B(n8211), .S(n4815), .Z(n5735) );
  INV_X1 U7065 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8267) );
  MUX2_X1 U7066 ( .A(n10438), .B(n8267), .S(n4815), .Z(n5740) );
  INV_X1 U7067 ( .A(SI_20_), .ZN(n5736) );
  INV_X1 U7068 ( .A(SI_21_), .ZN(n5316) );
  OAI21_X1 U7069 ( .B1(n5735), .B2(n5736), .A(n5316), .ZN(n5320) );
  AND2_X1 U7070 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5317) );
  AOI22_X1 U7071 ( .A1(n5320), .A2(n5319), .B1(n5318), .B2(n5317), .ZN(n5321)
         );
  INV_X1 U7072 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8271) );
  MUX2_X1 U7073 ( .A(n8271), .B(n8275), .S(n4815), .Z(n5324) );
  INV_X1 U7074 ( .A(SI_22_), .ZN(n5323) );
  INV_X1 U7075 ( .A(n5324), .ZN(n5325) );
  NAND2_X1 U7076 ( .A1(n5325), .A2(SI_22_), .ZN(n5326) );
  NAND2_X1 U7077 ( .A1(n5327), .A2(n5326), .ZN(n5755) );
  INV_X1 U7078 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5328) );
  MUX2_X1 U7079 ( .A(n5328), .B(n8309), .S(n4815), .Z(n5330) );
  INV_X1 U7080 ( .A(SI_23_), .ZN(n5329) );
  NAND2_X1 U7081 ( .A1(n5330), .A2(n5329), .ZN(n5333) );
  INV_X1 U7082 ( .A(n5330), .ZN(n5331) );
  NAND2_X1 U7083 ( .A1(n5331), .A2(SI_23_), .ZN(n5332) );
  INV_X1 U7084 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8311) );
  INV_X1 U7085 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8313) );
  MUX2_X1 U7086 ( .A(n8311), .B(n8313), .S(n4815), .Z(n5336) );
  INV_X1 U7087 ( .A(SI_24_), .ZN(n5335) );
  NAND2_X1 U7088 ( .A1(n5336), .A2(n5335), .ZN(n5339) );
  INV_X1 U7089 ( .A(n5336), .ZN(n5337) );
  NAND2_X1 U7090 ( .A1(n5337), .A2(SI_24_), .ZN(n5338) );
  INV_X1 U7091 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9131) );
  INV_X1 U7092 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9941) );
  MUX2_X1 U7093 ( .A(n9131), .B(n9941), .S(n4815), .Z(n5341) );
  INV_X1 U7094 ( .A(SI_25_), .ZN(n5340) );
  NAND2_X1 U7095 ( .A1(n5341), .A2(n5340), .ZN(n5344) );
  INV_X1 U7096 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U7097 ( .A1(n5342), .A2(SI_25_), .ZN(n5343) );
  INV_X1 U7098 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9127) );
  INV_X1 U7099 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9937) );
  MUX2_X1 U7100 ( .A(n9127), .B(n9937), .S(n4815), .Z(n5346) );
  INV_X1 U7101 ( .A(SI_26_), .ZN(n5345) );
  NAND2_X1 U7102 ( .A1(n5346), .A2(n5345), .ZN(n5349) );
  INV_X1 U7103 ( .A(n5346), .ZN(n5347) );
  NAND2_X1 U7104 ( .A1(n5347), .A2(SI_26_), .ZN(n5348) );
  INV_X1 U7105 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10431) );
  INV_X1 U7106 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9936) );
  MUX2_X1 U7107 ( .A(n10431), .B(n9936), .S(n4815), .Z(n5351) );
  INV_X1 U7108 ( .A(SI_27_), .ZN(n5350) );
  NAND2_X1 U7109 ( .A1(n5351), .A2(n5350), .ZN(n5354) );
  INV_X1 U7110 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U7111 ( .A1(n5352), .A2(SI_27_), .ZN(n5353) );
  NAND2_X1 U7112 ( .A1(n5821), .A2(n5822), .ZN(n5355) );
  INV_X1 U7113 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5356) );
  INV_X1 U7114 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8318) );
  MUX2_X1 U7115 ( .A(n5356), .B(n8318), .S(n4815), .Z(n5920) );
  XNOR2_X1 U7116 ( .A(n5920), .B(SI_28_), .ZN(n5918) );
  NAND4_X1 U7117 ( .A1(n5835), .A2(n5361), .A3(n5360), .A4(n5446), .ZN(n5362)
         );
  INV_X2 U7118 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10478) );
  INV_X2 U7119 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5619) );
  INV_X2 U7120 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7121 ( .A1(n5908), .A2(n5905), .ZN(n5881) );
  INV_X1 U7122 ( .A(n5881), .ZN(n5366) );
  NAND3_X1 U7123 ( .A1(n5366), .A2(n5883), .A3(n5152), .ZN(n5367) );
  NOR2_X1 U7124 ( .A1(n5372), .A2(n5371), .ZN(n5373) );
  OR2_X1 U7125 ( .A1(n6565), .A2(n8318), .ZN(n5374) );
  INV_X1 U7126 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5624) );
  INV_X1 U7127 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5672) );
  AND2_X1 U7128 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_18__SCAN_IN), 
        .ZN(n5380) );
  INV_X1 U7129 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9171) );
  INV_X1 U7130 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5745) );
  INV_X1 U7131 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9147) );
  INV_X1 U7132 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10310) );
  INV_X1 U7133 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9363) );
  XNOR2_X1 U7134 ( .A(n5943), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U7135 ( .A1(n5382), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5383) );
  AND2_X4 U7136 ( .A1(n5384), .A2(n5385), .ZN(n5812) );
  NAND2_X1 U7137 ( .A1(n9525), .A2(n5812), .ZN(n5390) );
  INV_X1 U7138 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9520) );
  AND2_X4 U7139 ( .A1(n8340), .A2(n9932), .ZN(n5536) );
  NAND2_X1 U7140 ( .A1(n5536), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U7141 ( .A1(n5937), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5386) );
  OAI211_X1 U7142 ( .C1(n9520), .C2(n5829), .A(n5387), .B(n5386), .ZN(n5388)
         );
  INV_X1 U7143 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U7144 ( .A1(n4388), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U7145 ( .A1(n5812), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U7146 ( .A1(n5536), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5392) );
  INV_X1 U7147 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U7148 ( .A1(n5398), .A2(n5399), .ZN(n5421) );
  INV_X1 U7149 ( .A(n5421), .ZN(n5400) );
  NAND2_X1 U7150 ( .A1(n5400), .A2(n5419), .ZN(n5423) );
  NAND2_X1 U7151 ( .A1(n5423), .A2(n5398), .ZN(n5404) );
  NAND2_X1 U7152 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  XNOR2_X1 U7153 ( .A(n5404), .B(n5403), .ZN(n6013) );
  INV_X1 U7154 ( .A(n6013), .ZN(n7306) );
  OR2_X1 U7155 ( .A1(n4390), .A2(n7298), .ZN(n5405) );
  OAI211_X2 U7156 ( .C1(n7320), .C2(n4728), .A(n5406), .B(n5405), .ZN(n9342)
         );
  INV_X1 U7157 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5408) );
  OR2_X1 U7158 ( .A1(n5775), .A2(n5408), .ZN(n5412) );
  NAND2_X1 U7159 ( .A1(n5812), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5411) );
  NAND4_X2 U7160 ( .A1(n5412), .A2(n5411), .A3(n5410), .A4(n5409), .ZN(n6578)
         );
  NOR2_X1 U7161 ( .A1(n5243), .A2(n10345), .ZN(n5414) );
  XNOR2_X1 U7162 ( .A(n5414), .B(n5413), .ZN(n7295) );
  NAND2_X1 U7163 ( .A1(n4391), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U7164 ( .A1(n5536), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U7165 ( .A1(n5812), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U7166 ( .A1(n4389), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U7167 ( .A1(n7665), .A2(n4648), .ZN(n5424) );
  INV_X1 U7168 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10311) );
  INV_X1 U7169 ( .A(n5419), .ZN(n5420) );
  NAND2_X1 U7170 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  NAND2_X1 U7171 ( .A1(n5423), .A2(n5422), .ZN(n7307) );
  NAND2_X1 U7172 ( .A1(n5424), .A2(n5848), .ZN(n5426) );
  NAND2_X1 U7173 ( .A1(n7663), .A2(n4646), .ZN(n5425) );
  NAND3_X1 U7174 ( .A1(n6581), .A2(n5426), .A3(n5425), .ZN(n5428) );
  NAND2_X1 U7175 ( .A1(n9212), .A2(n6929), .ZN(n5427) );
  NAND2_X1 U7176 ( .A1(n5428), .A2(n5427), .ZN(n7782) );
  INV_X1 U7177 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U7178 ( .A1(n5812), .A2(n7891), .ZN(n5432) );
  NAND2_X1 U7179 ( .A1(n5937), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U7180 ( .A1(n4389), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7181 ( .A1(n5536), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U7182 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  INV_X1 U7183 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7299) );
  OR2_X1 U7184 ( .A1(n6565), .A2(n7299), .ZN(n5444) );
  NAND2_X1 U7185 ( .A1(n5470), .A2(n5437), .ZN(n5439) );
  INV_X1 U7186 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U7187 ( .A1(n5441), .A2(n5440), .ZN(n5471) );
  NAND2_X1 U7188 ( .A1(n5442), .A2(n5471), .ZN(n7302) );
  OR2_X1 U7189 ( .A1(n5563), .A2(n7302), .ZN(n5443) );
  NAND2_X1 U7190 ( .A1(n10011), .A2(n7894), .ZN(n7869) );
  INV_X1 U7191 ( .A(n10011), .ZN(n9390) );
  NAND2_X1 U7192 ( .A1(n7869), .A2(n6447), .ZN(n7784) );
  NAND2_X1 U7193 ( .A1(n7782), .A2(n7784), .ZN(n7783) );
  NAND2_X1 U7194 ( .A1(n10011), .A2(n10006), .ZN(n5445) );
  NAND2_X1 U7195 ( .A1(n7783), .A2(n5445), .ZN(n7866) );
  INV_X1 U7196 ( .A(n5668), .ZN(n5468) );
  NAND2_X1 U7197 ( .A1(n5468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5447) );
  AOI22_X1 U7198 ( .A1(n5488), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5716), .B2(
        n8330), .ZN(n5451) );
  NAND2_X1 U7199 ( .A1(n5449), .A2(SI_5_), .ZN(n5483) );
  NAND2_X1 U7200 ( .A1(n5536), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7201 ( .A1(n4391), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5457) );
  INV_X1 U7202 ( .A(n5452), .ZN(n5460) );
  INV_X1 U7203 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U7204 ( .A1(n5460), .A2(n5453), .ZN(n5454) );
  AND2_X1 U7205 ( .A1(n5493), .A2(n5454), .ZN(n8076) );
  NAND2_X1 U7206 ( .A1(n5812), .A2(n8076), .ZN(n5456) );
  NAND2_X1 U7207 ( .A1(n4388), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5455) );
  NAND4_X1 U7208 ( .A1(n5458), .A2(n5457), .A3(n5456), .A4(n5455), .ZN(n7873)
         );
  NAND2_X1 U7209 ( .A1(n4388), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5464) );
  INV_X1 U7210 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7211 ( .A1(n7891), .A2(n5459), .ZN(n5461) );
  AND2_X1 U7212 ( .A1(n5461), .A2(n5460), .ZN(n9280) );
  NAND2_X1 U7213 ( .A1(n5812), .A2(n9280), .ZN(n5463) );
  NAND2_X1 U7214 ( .A1(n5536), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7215 ( .A1(n5466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5467) );
  MUX2_X1 U7216 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5467), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5469) );
  NAND2_X1 U7217 ( .A1(n5469), .A2(n5468), .ZN(n7366) );
  NAND2_X1 U7218 ( .A1(n5471), .A2(n5470), .ZN(n5475) );
  NAND2_X1 U7219 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  XNOR2_X1 U7220 ( .A(n5475), .B(n5474), .ZN(n7300) );
  NAND2_X1 U7221 ( .A1(n5527), .A2(n7300), .ZN(n5477) );
  OAI211_X1 U7222 ( .C1(n7320), .C2(n7366), .A(n5477), .B(n5476), .ZN(n10013)
         );
  NOR2_X1 U7223 ( .A1(n9389), .A2(n10013), .ZN(n5479) );
  NOR2_X1 U7224 ( .A1(n7873), .A2(n4394), .ZN(n5478) );
  INV_X1 U7225 ( .A(n7997), .ZN(n5501) );
  NAND2_X1 U7226 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  NAND2_X1 U7227 ( .A1(n5483), .A2(n5482), .ZN(n5487) );
  NAND2_X1 U7228 ( .A1(n5485), .A2(n5484), .ZN(n5486) );
  NAND2_X1 U7229 ( .A1(n7312), .A2(n5527), .ZN(n5491) );
  INV_X1 U7230 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7231 ( .A1(n5668), .A2(n5489), .ZN(n5528) );
  NAND2_X1 U7232 ( .A1(n5528), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5512) );
  XNOR2_X1 U7233 ( .A(n5512), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7407) );
  AOI22_X1 U7234 ( .A1(n4716), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5716), .B2(
        n7407), .ZN(n5490) );
  NAND2_X1 U7235 ( .A1(n5536), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7236 ( .A1(n5937), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5497) );
  INV_X1 U7237 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7238 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  AND2_X1 U7239 ( .A1(n5505), .A2(n5494), .ZN(n8005) );
  NAND2_X1 U7240 ( .A1(n5812), .A2(n8005), .ZN(n5496) );
  NAND2_X1 U7241 ( .A1(n4389), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5495) );
  NAND4_X1 U7242 ( .A1(n5498), .A2(n5497), .A3(n5496), .A4(n5495), .ZN(n9388)
         );
  NAND2_X1 U7243 ( .A1(n10027), .A2(n9388), .ZN(n8025) );
  NAND2_X1 U7244 ( .A1(n9389), .A2(n10013), .ZN(n5499) );
  NAND2_X1 U7245 ( .A1(n8053), .A2(n5499), .ZN(n7998) );
  NAND2_X1 U7246 ( .A1(n7997), .A2(n7998), .ZN(n5500) );
  NAND2_X1 U7247 ( .A1(n10027), .A2(n8108), .ZN(n5502) );
  NAND2_X1 U7248 ( .A1(n5503), .A2(n5502), .ZN(n8029) );
  NAND2_X1 U7249 ( .A1(n5937), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7250 ( .A1(n5536), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5509) );
  INV_X1 U7251 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7252 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  AND2_X1 U7253 ( .A1(n5538), .A2(n5506), .ZN(n8037) );
  NAND2_X1 U7254 ( .A1(n5812), .A2(n8037), .ZN(n5508) );
  NAND2_X1 U7255 ( .A1(n4389), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5507) );
  INV_X1 U7256 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7257 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  NAND2_X1 U7258 ( .A1(n5513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5515) );
  INV_X1 U7259 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5514) );
  XNOR2_X1 U7260 ( .A(n5515), .B(n5514), .ZN(n7408) );
  NAND2_X1 U7261 ( .A1(n5518), .A2(n5517), .ZN(n5520) );
  NAND2_X1 U7262 ( .A1(n5520), .A2(n5519), .ZN(n7315) );
  OR2_X1 U7263 ( .A1(n7315), .A2(n5563), .ZN(n5522) );
  INV_X1 U7264 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7308) );
  OR2_X1 U7265 ( .A1(n6565), .A2(n7308), .ZN(n5521) );
  OAI211_X1 U7266 ( .C1(n7320), .C2(n7408), .A(n5522), .B(n5521), .ZN(n8113)
         );
  NAND2_X1 U7267 ( .A1(n10040), .A2(n8113), .ZN(n8169) );
  NAND2_X1 U7268 ( .A1(n9387), .A2(n10033), .ZN(n6576) );
  NAND2_X1 U7269 ( .A1(n8169), .A2(n6576), .ZN(n8030) );
  NAND2_X1 U7270 ( .A1(n8029), .A2(n8030), .ZN(n5524) );
  NAND2_X1 U7271 ( .A1(n10040), .A2(n10033), .ZN(n5523) );
  NAND2_X1 U7272 ( .A1(n5524), .A2(n5523), .ZN(n8166) );
  XNOR2_X1 U7273 ( .A(n5526), .B(n5525), .ZN(n7310) );
  NAND2_X1 U7274 ( .A1(n7310), .A2(n5923), .ZN(n5535) );
  INV_X1 U7275 ( .A(n5528), .ZN(n5530) );
  NOR2_X1 U7276 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5529) );
  NAND2_X1 U7277 ( .A1(n5530), .A2(n5529), .ZN(n5532) );
  NAND2_X1 U7278 ( .A1(n5532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5531) );
  MUX2_X1 U7279 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5531), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5533) );
  AOI22_X1 U7280 ( .A1(n5488), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5716), .B2(
        n7680), .ZN(n5534) );
  NAND2_X1 U7281 ( .A1(n5937), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7282 ( .A1(n5536), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7283 ( .A1(n5538), .A2(n5537), .ZN(n5539) );
  AND2_X1 U7284 ( .A1(n5553), .A2(n5539), .ZN(n9199) );
  NAND2_X1 U7285 ( .A1(n5812), .A2(n9199), .ZN(n5541) );
  NAND2_X1 U7286 ( .A1(n4388), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5540) );
  NAND4_X1 U7287 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(n10052)
         );
  NAND2_X1 U7288 ( .A1(n9204), .A2(n10052), .ZN(n8140) );
  INV_X1 U7289 ( .A(n10052), .ZN(n9294) );
  NAND2_X1 U7290 ( .A1(n8140), .A2(n6465), .ZN(n8171) );
  NAND2_X1 U7291 ( .A1(n9204), .A2(n9294), .ZN(n5544) );
  NAND2_X1 U7292 ( .A1(n7345), .A2(n5923), .ZN(n5551) );
  NAND2_X1 U7293 ( .A1(n5548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5547) );
  MUX2_X1 U7294 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5547), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5549) );
  NAND2_X1 U7295 ( .A1(n5549), .A2(n5564), .ZN(n7681) );
  INV_X1 U7296 ( .A(n7681), .ZN(n7848) );
  AOI22_X1 U7297 ( .A1(n4716), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5716), .B2(
        n7848), .ZN(n5550) );
  NAND2_X1 U7298 ( .A1(n5536), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7299 ( .A1(n5937), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5558) );
  INV_X1 U7300 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7301 ( .A1(n5553), .A2(n5552), .ZN(n5554) );
  AND2_X1 U7302 ( .A1(n5568), .A2(n5554), .ZN(n9292) );
  NAND2_X1 U7303 ( .A1(n5812), .A2(n9292), .ZN(n5557) );
  NAND2_X1 U7304 ( .A1(n4388), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7305 ( .A1(n10054), .A2(n10039), .ZN(n6481) );
  NAND2_X1 U7306 ( .A1(n6470), .A2(n6481), .ZN(n8142) );
  INV_X1 U7307 ( .A(n10039), .ZN(n9386) );
  NAND2_X1 U7308 ( .A1(n4463), .A2(n5560), .ZN(n5561) );
  NAND2_X1 U7309 ( .A1(n5562), .A2(n5561), .ZN(n7344) );
  OR2_X1 U7310 ( .A1(n7344), .A2(n5563), .ZN(n5566) );
  NAND2_X1 U7311 ( .A1(n5564), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5579) );
  XNOR2_X1 U7312 ( .A(n5579), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7983) );
  AOI22_X1 U7313 ( .A1(n4716), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5716), .B2(
        n7983), .ZN(n5565) );
  NAND2_X1 U7314 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  AND2_X1 U7315 ( .A1(n5584), .A2(n5569), .ZN(n9158) );
  NAND2_X1 U7316 ( .A1(n5812), .A2(n9158), .ZN(n5573) );
  NAND2_X1 U7317 ( .A1(n5937), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7318 ( .A1(n4388), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5571) );
  NAND2_X1 U7319 ( .A1(n5536), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5570) );
  OR2_X1 U7320 ( .A1(n10062), .A2(n9331), .ZN(n6657) );
  NAND2_X1 U7321 ( .A1(n10062), .A2(n9331), .ZN(n9980) );
  NAND2_X1 U7322 ( .A1(n8227), .A2(n8230), .ZN(n5575) );
  INV_X1 U7323 ( .A(n9331), .ZN(n9987) );
  OR2_X1 U7324 ( .A1(n10062), .A2(n9987), .ZN(n5574) );
  NAND2_X1 U7325 ( .A1(n5575), .A2(n5574), .ZN(n9973) );
  XNOR2_X1 U7326 ( .A(n5577), .B(n5576), .ZN(n7350) );
  NAND2_X1 U7327 ( .A1(n7350), .A2(n5923), .ZN(n5583) );
  NAND2_X1 U7328 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  NAND2_X1 U7329 ( .A1(n5580), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5581) );
  AOI22_X1 U7330 ( .A1(n4716), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5716), .B2(
        n8122), .ZN(n5582) );
  NAND2_X1 U7331 ( .A1(n5583), .A2(n5582), .ZN(n9333) );
  NAND2_X1 U7332 ( .A1(n5937), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7333 ( .A1(n5536), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5588) );
  INV_X1 U7334 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U7335 ( .A1(n5584), .A2(n10278), .ZN(n5585) );
  AND2_X1 U7336 ( .A1(n5603), .A2(n5585), .ZN(n9992) );
  NAND2_X1 U7337 ( .A1(n5812), .A2(n9992), .ZN(n5587) );
  NAND2_X1 U7338 ( .A1(n4389), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5586) );
  OR2_X1 U7339 ( .A1(n9333), .A2(n10083), .ZN(n6473) );
  NAND2_X1 U7340 ( .A1(n9333), .A2(n10083), .ZN(n6476) );
  NAND2_X1 U7341 ( .A1(n6473), .A2(n6476), .ZN(n9981) );
  NAND2_X1 U7342 ( .A1(n9973), .A2(n9981), .ZN(n5591) );
  INV_X1 U7343 ( .A(n10083), .ZN(n9385) );
  OR2_X1 U7344 ( .A1(n9333), .A2(n9385), .ZN(n5590) );
  NAND2_X1 U7345 ( .A1(n5591), .A2(n5590), .ZN(n8276) );
  NAND2_X1 U7346 ( .A1(n5611), .A2(n5592), .ZN(n5593) );
  NAND2_X1 U7347 ( .A1(n5594), .A2(n5593), .ZN(n5595) );
  NAND2_X1 U7348 ( .A1(n7416), .A2(n5923), .ZN(n5601) );
  INV_X1 U7349 ( .A(n5666), .ZN(n5596) );
  NAND2_X1 U7350 ( .A1(n5668), .A2(n5596), .ZN(n5598) );
  NAND2_X1 U7351 ( .A1(n5598), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5597) );
  MUX2_X1 U7352 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5597), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5599) );
  AOI22_X1 U7353 ( .A1(n4716), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5716), .B2(
        n8297), .ZN(n5600) );
  NAND2_X1 U7354 ( .A1(n5937), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7355 ( .A1(n5536), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7356 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  AND2_X1 U7357 ( .A1(n5625), .A2(n5604), .ZN(n9226) );
  NAND2_X1 U7358 ( .A1(n5812), .A2(n9226), .ZN(n5606) );
  NAND2_X1 U7359 ( .A1(n4388), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5605) );
  NAND4_X1 U7360 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .ZN(n9985)
         );
  NAND2_X1 U7361 ( .A1(n8282), .A2(n9985), .ZN(n6474) );
  NAND2_X1 U7362 ( .A1(n10079), .A2(n9757), .ZN(n6666) );
  NAND2_X1 U7363 ( .A1(n6474), .A2(n6666), .ZN(n8277) );
  NAND2_X1 U7364 ( .A1(n8276), .A2(n8277), .ZN(n5610) );
  NAND2_X1 U7365 ( .A1(n8282), .A2(n9757), .ZN(n5609) );
  NAND2_X1 U7366 ( .A1(n5610), .A2(n5609), .ZN(n9750) );
  NAND2_X1 U7367 ( .A1(n5612), .A2(n5611), .ZN(n5616) );
  NAND2_X1 U7368 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  NAND2_X1 U7369 ( .A1(n7512), .A2(n5923), .ZN(n5623) );
  NAND2_X1 U7370 ( .A1(n5618), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5617) );
  MUX2_X1 U7371 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5617), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5621) );
  INV_X1 U7372 ( .A(n5618), .ZN(n5620) );
  NAND2_X1 U7373 ( .A1(n5620), .A2(n5619), .ZN(n5650) );
  NAND2_X1 U7374 ( .A1(n5621), .A2(n5650), .ZN(n7514) );
  AOI22_X1 U7375 ( .A1(n4716), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5716), .B2(
        n9453), .ZN(n5622) );
  NAND2_X1 U7376 ( .A1(n5536), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7377 ( .A1(n5937), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7378 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  AND2_X1 U7379 ( .A1(n5639), .A2(n5626), .ZN(n9760) );
  NAND2_X1 U7380 ( .A1(n5812), .A2(n9760), .ZN(n5628) );
  NAND2_X1 U7381 ( .A1(n4388), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5627) );
  XNOR2_X1 U7382 ( .A(n9902), .B(n9139), .ZN(n9754) );
  INV_X1 U7383 ( .A(n9139), .ZN(n9892) );
  OR2_X1 U7384 ( .A1(n9902), .A2(n9892), .ZN(n5631) );
  XNOR2_X1 U7385 ( .A(n5632), .B(SI_14_), .ZN(n5633) );
  XNOR2_X1 U7386 ( .A(n5634), .B(n5633), .ZN(n7490) );
  NAND2_X1 U7387 ( .A1(n7490), .A2(n5923), .ZN(n5637) );
  NAND2_X1 U7388 ( .A1(n5650), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5635) );
  XNOR2_X1 U7389 ( .A(n5635), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9466) );
  AOI22_X1 U7390 ( .A1(n4716), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5716), .B2(
        n9466), .ZN(n5636) );
  NAND2_X1 U7391 ( .A1(n5937), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7392 ( .A1(n4389), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5643) );
  INV_X1 U7393 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7394 ( .A1(n5639), .A2(n5638), .ZN(n5640) );
  AND2_X1 U7395 ( .A1(n5655), .A2(n5640), .ZN(n9737) );
  NAND2_X1 U7396 ( .A1(n5812), .A2(n9737), .ZN(n5642) );
  NAND2_X1 U7397 ( .A1(n5536), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5641) );
  NAND4_X1 U7398 ( .A1(n5644), .A2(n5643), .A3(n5642), .A4(n5641), .ZN(n9882)
         );
  NAND2_X1 U7399 ( .A1(n9746), .A2(n9882), .ZN(n5645) );
  XNOR2_X1 U7400 ( .A(n5648), .B(SI_15_), .ZN(n5649) );
  XNOR2_X1 U7401 ( .A(n5647), .B(n5649), .ZN(n7704) );
  NAND2_X1 U7402 ( .A1(n7704), .A2(n5923), .ZN(n5653) );
  OAI21_X1 U7403 ( .B1(n5650), .B2(P1_IR_REG_14__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5651) );
  XNOR2_X1 U7404 ( .A(n5651), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U7405 ( .A1(n4716), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5716), .B2(
        n9954), .ZN(n5652) );
  NAND2_X1 U7406 ( .A1(n5937), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5660) );
  INV_X1 U7407 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7408 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  AND2_X1 U7409 ( .A1(n5673), .A2(n5656), .ZN(n9722) );
  NAND2_X1 U7410 ( .A1(n9722), .A2(n5812), .ZN(n5659) );
  NAND2_X1 U7411 ( .A1(n4388), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7412 ( .A1(n5536), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5657) );
  NAND4_X1 U7413 ( .A1(n5660), .A2(n5659), .A3(n5658), .A4(n5657), .ZN(n9891)
         );
  OR2_X1 U7414 ( .A1(n5860), .A2(n9891), .ZN(n5661) );
  XNOR2_X1 U7415 ( .A(n5662), .B(SI_16_), .ZN(n5663) );
  XNOR2_X1 U7416 ( .A(n5664), .B(n5663), .ZN(n7779) );
  NAND2_X1 U7417 ( .A1(n7779), .A2(n5923), .ZN(n5671) );
  NAND2_X1 U7418 ( .A1(n5683), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5669) );
  XNOR2_X1 U7419 ( .A(n5669), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9485) );
  AOI22_X1 U7420 ( .A1(n4716), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5716), .B2(
        n9485), .ZN(n5670) );
  NAND2_X1 U7421 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  AND2_X1 U7422 ( .A1(n9260), .A2(n5674), .ZN(n9708) );
  NAND2_X1 U7423 ( .A1(n9708), .A2(n5812), .ZN(n5679) );
  NAND2_X1 U7424 ( .A1(n5937), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7425 ( .A1(n5536), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5675) );
  AND2_X1 U7426 ( .A1(n5676), .A2(n5675), .ZN(n5678) );
  NAND2_X1 U7427 ( .A1(n4389), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7428 ( .A1(n9877), .A2(n9725), .ZN(n6487) );
  XNOR2_X1 U7429 ( .A(n5695), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9499) );
  AOI22_X1 U7430 ( .A1(n4716), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5716), .B2(
        n9499), .ZN(n5685) );
  XNOR2_X1 U7431 ( .A(n9260), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9686) );
  NAND2_X1 U7432 ( .A1(n9686), .A2(n5812), .ZN(n5691) );
  INV_X1 U7433 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U7434 ( .A1(n5937), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7435 ( .A1(n5536), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5687) );
  OAI211_X1 U7436 ( .C1(n5829), .C2(n9689), .A(n5688), .B(n5687), .ZN(n5689)
         );
  INV_X1 U7437 ( .A(n5689), .ZN(n5690) );
  NOR2_X1 U7438 ( .A1(n9869), .A2(n9675), .ZN(n9665) );
  NAND2_X1 U7439 ( .A1(n7934), .A2(n5923), .ZN(n5700) );
  INV_X1 U7440 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7441 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  NAND2_X1 U7442 ( .A1(n5696), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5697) );
  OR2_X1 U7443 ( .A1(n5697), .A2(n10416), .ZN(n5698) );
  NAND2_X1 U7444 ( .A1(n5697), .A2(n10416), .ZN(n5714) );
  AND2_X1 U7445 ( .A1(n5714), .A2(n5698), .ZN(n9967) );
  AOI22_X1 U7446 ( .A1(n4716), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5716), .B2(
        n9967), .ZN(n5699) );
  INV_X1 U7447 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5705) );
  INV_X1 U7448 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10413) );
  INV_X1 U7449 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5701) );
  OAI21_X1 U7450 ( .B1(n9260), .B2(n10413), .A(n5701), .ZN(n5702) );
  NAND2_X1 U7451 ( .A1(n5719), .A2(n5702), .ZN(n9672) );
  OR2_X1 U7452 ( .A1(n9672), .A2(n5872), .ZN(n5704) );
  AOI22_X1 U7453 ( .A1(n4389), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5937), .B2(
        P1_REG1_REG_18__SCAN_IN), .ZN(n5703) );
  OAI211_X1 U7454 ( .C1(n5875), .C2(n5705), .A(n5704), .B(n5703), .ZN(n9850)
         );
  NAND2_X1 U7455 ( .A1(n9877), .A2(n9883), .ZN(n9664) );
  NAND2_X1 U7456 ( .A1(n9664), .A2(n9874), .ZN(n5706) );
  NAND2_X1 U7457 ( .A1(n9869), .A2(n5706), .ZN(n5707) );
  OAI21_X1 U7458 ( .B1(n9874), .B2(n9664), .A(n5707), .ZN(n5708) );
  AOI21_X1 U7459 ( .B1(n9863), .B2(n9850), .A(n5708), .ZN(n5709) );
  OR2_X1 U7460 ( .A1(n9863), .A2(n9850), .ZN(n5710) );
  NAND2_X1 U7461 ( .A1(n5711), .A2(n5710), .ZN(n9648) );
  XNOR2_X1 U7462 ( .A(n5712), .B(n5713), .ZN(n8116) );
  NAND2_X1 U7463 ( .A1(n8116), .A2(n5923), .ZN(n5718) );
  AOI22_X1 U7464 ( .A1(n5488), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9610), .B2(
        n5716), .ZN(n5717) );
  NAND2_X1 U7465 ( .A1(n5719), .A2(n9171), .ZN(n5720) );
  NAND2_X1 U7466 ( .A1(n5726), .A2(n5720), .ZN(n9652) );
  AOI22_X1 U7467 ( .A1(n4388), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n5937), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U7468 ( .A1(n5536), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5721) );
  OAI211_X1 U7469 ( .C1(n9652), .C2(n5872), .A(n5722), .B(n5721), .ZN(n9638)
         );
  NAND2_X1 U7470 ( .A1(n9657), .A2(n9638), .ZN(n5723) );
  XNOR2_X1 U7471 ( .A(n5735), .B(SI_20_), .ZN(n5724) );
  OR2_X1 U7472 ( .A1(n6565), .A2(n8211), .ZN(n5725) );
  INV_X1 U7473 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U7474 ( .A1(n5726), .A2(n10314), .ZN(n5727) );
  NAND2_X1 U7475 ( .A1(n5746), .A2(n5727), .ZN(n9636) );
  OR2_X1 U7476 ( .A1(n9636), .A2(n5872), .ZN(n5732) );
  INV_X1 U7477 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U7478 ( .A1(n4389), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U7479 ( .A1(n5937), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5728) );
  OAI211_X1 U7480 ( .C1(n5875), .C2(n10254), .A(n5729), .B(n5728), .ZN(n5730)
         );
  INV_X1 U7481 ( .A(n5730), .ZN(n5731) );
  NAND2_X1 U7482 ( .A1(n5732), .A2(n5731), .ZN(n9851) );
  AND2_X1 U7483 ( .A1(n9845), .A2(n9851), .ZN(n5734) );
  OAI21_X1 U7484 ( .B1(n5737), .B2(n5736), .A(n5735), .ZN(n5739) );
  NAND2_X1 U7485 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  NAND2_X1 U7486 ( .A1(n5739), .A2(n5738), .ZN(n5742) );
  XNOR2_X1 U7487 ( .A(n5740), .B(SI_21_), .ZN(n5741) );
  OR2_X1 U7488 ( .A1(n6565), .A2(n8267), .ZN(n5743) );
  NAND2_X1 U7489 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  AND2_X1 U7490 ( .A1(n5759), .A2(n5747), .ZN(n9623) );
  NAND2_X1 U7491 ( .A1(n9623), .A2(n5812), .ZN(n5752) );
  INV_X1 U7492 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U7493 ( .A1(n5937), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7494 ( .A1(n5536), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5748) );
  OAI211_X1 U7495 ( .C1(n10250), .C2(n5829), .A(n5749), .B(n5748), .ZN(n5750)
         );
  INV_X1 U7496 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U7497 ( .A1(n5752), .A2(n5751), .ZN(n9824) );
  NOR2_X1 U7498 ( .A1(n9837), .A2(n9824), .ZN(n5754) );
  NAND2_X1 U7499 ( .A1(n9837), .A2(n9824), .ZN(n5753) );
  XNOR2_X1 U7500 ( .A(n5756), .B(n5755), .ZN(n8270) );
  NAND2_X1 U7501 ( .A1(n8270), .A2(n5923), .ZN(n5758) );
  OR2_X1 U7502 ( .A1(n6565), .A2(n8275), .ZN(n5757) );
  INV_X1 U7503 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U7504 ( .A1(n5759), .A2(n9317), .ZN(n5760) );
  NAND2_X1 U7505 ( .A1(n5771), .A2(n5760), .ZN(n9612) );
  INV_X1 U7506 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U7507 ( .A1(n5937), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7508 ( .A1(n5536), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5761) );
  OAI211_X1 U7509 ( .C1(n5829), .C2(n9611), .A(n5762), .B(n5761), .ZN(n5763)
         );
  INV_X1 U7510 ( .A(n5763), .ZN(n5764) );
  AND2_X1 U7511 ( .A1(n9320), .A2(n9815), .ZN(n5766) );
  NAND2_X1 U7512 ( .A1(n8306), .A2(n5923), .ZN(n5770) );
  OR2_X1 U7513 ( .A1(n6565), .A2(n8309), .ZN(n5769) );
  NAND2_X1 U7514 ( .A1(n5771), .A2(n9147), .ZN(n5772) );
  AND2_X1 U7515 ( .A1(n5786), .A2(n5772), .ZN(n9595) );
  NAND2_X1 U7516 ( .A1(n9595), .A2(n5812), .ZN(n5778) );
  INV_X1 U7517 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10417) );
  NAND2_X1 U7518 ( .A1(n4388), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U7519 ( .A1(n5536), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5773) );
  OAI211_X1 U7520 ( .C1(n5775), .C2(n10417), .A(n5774), .B(n5773), .ZN(n5776)
         );
  INV_X1 U7521 ( .A(n5776), .ZN(n5777) );
  NAND2_X1 U7522 ( .A1(n9600), .A2(n9825), .ZN(n5779) );
  XNOR2_X1 U7523 ( .A(n5781), .B(n5782), .ZN(n8310) );
  NAND2_X1 U7524 ( .A1(n8310), .A2(n5923), .ZN(n5784) );
  OR2_X1 U7525 ( .A1(n6565), .A2(n8313), .ZN(n5783) );
  INV_X1 U7526 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7527 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  NAND2_X1 U7528 ( .A1(n5798), .A2(n5787), .ZN(n9585) );
  INV_X1 U7529 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U7530 ( .A1(n5536), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7531 ( .A1(n5937), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5788) );
  OAI211_X1 U7532 ( .C1(n9584), .C2(n5829), .A(n5789), .B(n5788), .ZN(n5790)
         );
  INV_X1 U7533 ( .A(n5790), .ZN(n5791) );
  AND2_X1 U7534 ( .A1(n9812), .A2(n9816), .ZN(n5793) );
  XNOR2_X1 U7535 ( .A(n5794), .B(n5795), .ZN(n9129) );
  NAND2_X1 U7536 ( .A1(n9129), .A2(n5923), .ZN(n5797) );
  OR2_X1 U7537 ( .A1(n6565), .A2(n9941), .ZN(n5796) );
  NAND2_X1 U7538 ( .A1(n5798), .A2(n10310), .ZN(n5799) );
  NAND2_X1 U7539 ( .A1(n5810), .A2(n5799), .ZN(n9564) );
  INV_X1 U7540 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10202) );
  NAND2_X1 U7541 ( .A1(n4389), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7542 ( .A1(n4391), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5800) );
  OAI211_X1 U7543 ( .C1(n5875), .C2(n10202), .A(n5801), .B(n5800), .ZN(n5802)
         );
  INV_X1 U7544 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U7545 ( .A1(n9808), .A2(n9577), .ZN(n5805) );
  NAND2_X1 U7546 ( .A1(n9126), .A2(n5923), .ZN(n5809) );
  OR2_X1 U7547 ( .A1(n6565), .A2(n9937), .ZN(n5808) );
  NAND2_X1 U7548 ( .A1(n5810), .A2(n9363), .ZN(n5811) );
  NAND2_X1 U7549 ( .A1(n9548), .A2(n5812), .ZN(n5818) );
  INV_X1 U7550 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7551 ( .A1(n5937), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7552 ( .A1(n5536), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5813) );
  OAI211_X1 U7553 ( .C1(n5815), .C2(n5829), .A(n5814), .B(n5813), .ZN(n5816)
         );
  INV_X1 U7554 ( .A(n5816), .ZN(n5817) );
  NAND2_X1 U7555 ( .A1(n9554), .A2(n9553), .ZN(n5820) );
  NAND2_X1 U7556 ( .A1(n9801), .A2(n9788), .ZN(n5819) );
  NAND2_X1 U7557 ( .A1(n9124), .A2(n5923), .ZN(n5824) );
  OR2_X1 U7558 ( .A1(n6565), .A2(n9936), .ZN(n5823) );
  INV_X1 U7559 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10201) );
  NAND2_X1 U7560 ( .A1(n5825), .A2(n10201), .ZN(n5826) );
  NAND2_X1 U7561 ( .A1(n5943), .A2(n5826), .ZN(n9536) );
  INV_X1 U7562 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U7563 ( .A1(n5536), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U7564 ( .A1(n5937), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5827) );
  OAI211_X1 U7565 ( .C1(n9535), .C2(n5829), .A(n5828), .B(n5827), .ZN(n5830)
         );
  INV_X1 U7566 ( .A(n5830), .ZN(n5831) );
  AND2_X2 U7567 ( .A1(n5832), .A2(n5831), .ZN(n9798) );
  NAND2_X1 U7568 ( .A1(n9540), .A2(n9798), .ZN(n6439) );
  AOI21_X1 U7569 ( .B1(n6594), .B2(n5834), .A(n9786), .ZN(n9519) );
  INV_X1 U7570 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7571 ( .A1(n5835), .A2(n5836), .ZN(n5837) );
  OAI21_X1 U7572 ( .B1(n5838), .B2(n5837), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5840) );
  INV_X1 U7573 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7574 ( .A1(n5843), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5845) );
  INV_X1 U7575 ( .A(n8269), .ZN(n6645) );
  INV_X1 U7576 ( .A(n7318), .ZN(n7117) );
  OR2_X1 U7577 ( .A1(n7120), .A2(n7117), .ZN(n8320) );
  INV_X1 U7578 ( .A(n7478), .ZN(n8319) );
  NAND2_X1 U7579 ( .A1(n7120), .A2(n6917), .ZN(n5847) );
  NAND3_X1 U7580 ( .A1(n8320), .A2(n8319), .A3(n5847), .ZN(n9979) );
  INV_X1 U7581 ( .A(n8325), .ZN(n6579) );
  NAND2_X1 U7582 ( .A1(n4648), .A2(n5848), .ZN(n5849) );
  INV_X1 U7583 ( .A(n9389), .ZN(n8049) );
  NAND2_X1 U7584 ( .A1(n9389), .A2(n9281), .ZN(n6448) );
  INV_X1 U7585 ( .A(n6445), .ZN(n8058) );
  INV_X1 U7586 ( .A(n8053), .ZN(n8059) );
  NAND2_X1 U7587 ( .A1(n8058), .A2(n8059), .ZN(n5851) );
  NAND2_X1 U7588 ( .A1(n6470), .A2(n8140), .ZN(n6584) );
  INV_X1 U7589 ( .A(n8026), .ZN(n5852) );
  NAND2_X1 U7590 ( .A1(n8025), .A2(n6576), .ZN(n5853) );
  NOR2_X1 U7591 ( .A1(n6584), .A2(n5853), .ZN(n5854) );
  INV_X1 U7592 ( .A(n9980), .ZN(n5857) );
  NOR2_X1 U7593 ( .A1(n9981), .A2(n5857), .ZN(n5858) );
  INV_X1 U7594 ( .A(n8277), .ZN(n8278) );
  INV_X1 U7595 ( .A(n9891), .ZN(n9873) );
  INV_X1 U7596 ( .A(n9882), .ZN(n9756) );
  NAND2_X1 U7597 ( .A1(n6575), .A2(n9717), .ZN(n5861) );
  INV_X1 U7598 ( .A(n5861), .ZN(n5859) );
  NAND2_X1 U7599 ( .A1(n6671), .A2(n5859), .ZN(n5865) );
  NAND2_X1 U7600 ( .A1(n9746), .A2(n9756), .ZN(n6586) );
  NAND2_X1 U7601 ( .A1(n9902), .A2(n9139), .ZN(n9731) );
  NAND2_X1 U7602 ( .A1(n5860), .A2(n9873), .ZN(n9700) );
  OAI21_X1 U7603 ( .B1(n5861), .B2(n9698), .A(n9700), .ZN(n5862) );
  NAND2_X1 U7604 ( .A1(n5862), .A2(n6671), .ZN(n5863) );
  AND2_X1 U7605 ( .A1(n5863), .A2(n6487), .ZN(n5864) );
  INV_X1 U7606 ( .A(n9692), .ZN(n5867) );
  NAND2_X1 U7607 ( .A1(n9869), .A2(n9874), .ZN(n6501) );
  INV_X1 U7608 ( .A(n9850), .ZN(n9261) );
  NAND2_X1 U7609 ( .A1(n9863), .A2(n9261), .ZN(n6517) );
  INV_X1 U7610 ( .A(n6517), .ZN(n5868) );
  INV_X1 U7611 ( .A(n9638), .ZN(n9860) );
  OR2_X1 U7612 ( .A1(n9657), .A2(n9860), .ZN(n6505) );
  NAND2_X1 U7613 ( .A1(n9657), .A2(n9860), .ZN(n6640) );
  NAND2_X1 U7614 ( .A1(n6505), .A2(n6640), .ZN(n9650) );
  XNOR2_X1 U7615 ( .A(n9845), .B(n9851), .ZN(n9644) );
  INV_X1 U7616 ( .A(n9851), .ZN(n9833) );
  NAND2_X1 U7617 ( .A1(n9643), .A2(n6507), .ZN(n9629) );
  INV_X1 U7618 ( .A(n9824), .ZN(n9842) );
  OR2_X1 U7619 ( .A1(n9320), .A2(n9834), .ZN(n6524) );
  NAND2_X1 U7620 ( .A1(n9320), .A2(n9834), .ZN(n6526) );
  OR2_X1 U7621 ( .A1(n9600), .A2(n9613), .ZN(n6528) );
  NAND2_X1 U7622 ( .A1(n9600), .A2(n9613), .ZN(n9576) );
  NAND2_X1 U7623 ( .A1(n9812), .A2(n9598), .ZN(n6607) );
  NAND2_X1 U7624 ( .A1(n9808), .A2(n9797), .ZN(n6611) );
  INV_X1 U7625 ( .A(n6611), .ZN(n6532) );
  INV_X1 U7626 ( .A(n6612), .ZN(n6536) );
  NAND2_X1 U7627 ( .A1(n9610), .A2(n6914), .ZN(n6569) );
  NAND2_X1 U7628 ( .A1(n4530), .A2(n6645), .ZN(n6635) );
  INV_X1 U7629 ( .A(n5391), .ZN(n9189) );
  NAND2_X1 U7630 ( .A1(n7692), .A2(n6579), .ZN(n7698) );
  NAND2_X1 U7631 ( .A1(n7874), .A2(n9281), .ZN(n8054) );
  NAND2_X1 U7632 ( .A1(n8003), .A2(n10033), .ZN(n8175) );
  INV_X1 U7633 ( .A(n10062), .ZN(n8235) );
  INV_X1 U7634 ( .A(n9333), .ZN(n10072) );
  NAND2_X1 U7635 ( .A1(n8233), .A2(n10072), .ZN(n8281) );
  OR2_X2 U7636 ( .A1(n8281), .A2(n10079), .ZN(n9759) );
  INV_X1 U7637 ( .A(n5860), .ZN(n9886) );
  NOR2_X4 U7638 ( .A1(n9685), .A2(n9863), .ZN(n9670) );
  AND2_X2 U7639 ( .A1(n9608), .A2(n9828), .ZN(n9593) );
  INV_X1 U7640 ( .A(n9801), .ZN(n9547) );
  AND2_X2 U7641 ( .A1(n9563), .A2(n9547), .ZN(n9545) );
  INV_X1 U7642 ( .A(n9975), .ZN(n9768) );
  AOI21_X1 U7643 ( .B1(n9534), .B2(n5391), .A(n9768), .ZN(n5870) );
  OR2_X2 U7644 ( .A1(n9534), .A2(n5391), .ZN(n5947) );
  NAND2_X1 U7645 ( .A1(n5870), .A2(n5947), .ZN(n9528) );
  INV_X1 U7646 ( .A(n8317), .ZN(n9405) );
  INV_X1 U7647 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9186) );
  INV_X1 U7648 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10309) );
  NAND2_X1 U7649 ( .A1(n4388), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7650 ( .A1(n5937), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5873) );
  OAI211_X1 U7651 ( .C1(n5875), .C2(n10309), .A(n5874), .B(n5873), .ZN(n5876)
         );
  INV_X1 U7652 ( .A(n5876), .ZN(n5877) );
  NAND2_X1 U7653 ( .A1(n5878), .A2(n5877), .ZN(n9383) );
  AOI22_X1 U7654 ( .A1(n9384), .A2(n10053), .B1(n9986), .B2(n9383), .ZN(n5879)
         );
  OAI211_X1 U7655 ( .C1(n9189), .C2(n10071), .A(n9528), .B(n5879), .ZN(n5880)
         );
  NAND2_X1 U7656 ( .A1(n5881), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7657 ( .A1(n9944), .A2(P1_B_REG_SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7658 ( .A1(n5884), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5885) );
  MUX2_X1 U7659 ( .A(P1_B_REG_SCAN_IN), .B(n5887), .S(n8315), .Z(n5891) );
  INV_X1 U7660 ( .A(n9939), .ZN(n5890) );
  NAND2_X1 U7661 ( .A1(n9944), .A2(n9939), .ZN(n9925) );
  OAI21_X1 U7662 ( .B1(n9924), .B2(P1_D_REG_1__SCAN_IN), .A(n9925), .ZN(n5928)
         );
  NOR4_X1 U7663 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5899) );
  NOR4_X1 U7664 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5898) );
  INV_X1 U7665 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10199) );
  INV_X1 U7666 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10238) );
  INV_X1 U7667 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10435) );
  INV_X1 U7668 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10463) );
  NAND4_X1 U7669 ( .A1(n10199), .A2(n10238), .A3(n10435), .A4(n10463), .ZN(
        n10354) );
  NOR4_X1 U7670 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5895) );
  NOR4_X1 U7671 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5894) );
  NOR4_X1 U7672 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n5893) );
  NOR4_X1 U7673 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5892) );
  NAND4_X1 U7674 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(n5896)
         );
  NOR4_X1 U7675 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n10354), .A4(n5896), .ZN(n5897) );
  NAND3_X1 U7676 ( .A1(n5899), .A2(n5898), .A3(n5897), .ZN(n5900) );
  NAND2_X1 U7677 ( .A1(n5902), .A2(n5900), .ZN(n5927) );
  NAND2_X1 U7678 ( .A1(n9610), .A2(n9975), .ZN(n5932) );
  INV_X1 U7679 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7680 ( .A1(n5902), .A2(n5901), .ZN(n5903) );
  NAND2_X1 U7681 ( .A1(n9939), .A2(n8315), .ZN(n9926) );
  NAND2_X1 U7682 ( .A1(n5903), .A2(n9926), .ZN(n7115) );
  NAND2_X1 U7683 ( .A1(n7120), .A2(n7318), .ZN(n7132) );
  INV_X1 U7684 ( .A(n9944), .ZN(n5904) );
  NAND2_X1 U7685 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7686 ( .A1(n5907), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5909) );
  XNOR2_X1 U7687 ( .A(n5909), .B(n5908), .ZN(n7317) );
  NAND2_X1 U7688 ( .A1(n7132), .A2(n9923), .ZN(n5911) );
  NOR2_X1 U7689 ( .A1(n7115), .A2(n5911), .ZN(n5910) );
  INV_X1 U7690 ( .A(n5911), .ZN(n5912) );
  NAND2_X1 U7691 ( .A1(n5914), .A2(n10090), .ZN(n5916) );
  NAND2_X1 U7692 ( .A1(n10088), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7693 ( .A1(n5916), .A2(n5915), .ZN(P1_U3518) );
  AND2_X1 U7694 ( .A1(n5391), .A2(n9789), .ZN(n9773) );
  NOR2_X1 U7695 ( .A1(n9786), .A2(n9773), .ZN(n5926) );
  INV_X1 U7696 ( .A(SI_28_), .ZN(n5919) );
  NAND2_X1 U7697 ( .A1(n5920), .A2(n5919), .ZN(n5921) );
  INV_X1 U7698 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5922) );
  INV_X1 U7699 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10469) );
  MUX2_X1 U7700 ( .A(n5922), .B(n10469), .S(n4815), .Z(n6544) );
  OR2_X1 U7701 ( .A1(n6565), .A2(n10469), .ZN(n5924) );
  NAND2_X1 U7702 ( .A1(n9779), .A2(n9521), .ZN(n6620) );
  XNOR2_X1 U7703 ( .A(n5926), .B(n9782), .ZN(n5936) );
  INV_X1 U7704 ( .A(n5927), .ZN(n5929) );
  INV_X1 U7705 ( .A(n7116), .ZN(n5931) );
  NAND2_X1 U7706 ( .A1(n5931), .A2(n5930), .ZN(n5949) );
  INV_X1 U7707 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U7708 ( .A1(n9979), .A2(n8036), .ZN(n5935) );
  NAND2_X1 U7709 ( .A1(n5936), .A2(n9704), .ZN(n5957) );
  AND2_X1 U7710 ( .A1(n4530), .A2(n7478), .ZN(n7128) );
  NAND2_X1 U7711 ( .A1(n9997), .A2(n10053), .ZN(n9522) );
  INV_X2 U7712 ( .A(n9997), .ZN(n9993) );
  NAND2_X1 U7713 ( .A1(n5937), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7714 ( .A1(n4389), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7715 ( .A1(n5536), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5938) );
  NAND3_X1 U7716 ( .A1(n5940), .A2(n5939), .A3(n5938), .ZN(n9382) );
  INV_X1 U7717 ( .A(P1_B_REG_SCAN_IN), .ZN(n5941) );
  OR2_X1 U7718 ( .A1(n9935), .A2(n5941), .ZN(n5942) );
  AND2_X1 U7719 ( .A1(n9986), .A2(n5942), .ZN(n9510) );
  NAND2_X1 U7720 ( .A1(n9382), .A2(n9510), .ZN(n9776) );
  NOR2_X1 U7721 ( .A1(n9993), .A2(n9776), .ZN(n5945) );
  NOR3_X1 U7722 ( .A1(n5943), .A2(n9186), .A3(n9671), .ZN(n5944) );
  AOI211_X1 U7723 ( .C1(n9993), .C2(P1_REG2_REG_29__SCAN_IN), .A(n5945), .B(
        n5944), .ZN(n5946) );
  OAI21_X1 U7724 ( .B1(n9777), .B2(n9522), .A(n5946), .ZN(n5952) );
  AOI21_X1 U7725 ( .B1(n9779), .B2(n5947), .A(n9768), .ZN(n5948) );
  INV_X1 U7726 ( .A(n5949), .ZN(n5950) );
  NOR2_X1 U7727 ( .A1(n9785), .A2(n9743), .ZN(n5951) );
  AOI211_X1 U7728 ( .C1(n9747), .C2(n9779), .A(n5952), .B(n5951), .ZN(n5956)
         );
  INV_X1 U7729 ( .A(n6440), .ZN(n5953) );
  NAND2_X1 U7730 ( .A1(n9997), .A2(n10061), .ZN(n9715) );
  INV_X1 U7731 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7732 ( .A1(n6206), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7733 ( .A1(n6216), .A2(n5970), .ZN(n8853) );
  NOR2_X1 U7734 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5973) );
  NAND4_X1 U7735 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n6354), .ZN(n6362)
         );
  NAND2_X1 U7736 ( .A1(n6008), .A2(n5974), .ZN(n5975) );
  INV_X2 U7737 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10479) );
  NAND4_X1 U7738 ( .A1(n5981), .A2(n10479), .A3(n5980), .A4(n5979), .ZN(n6007)
         );
  INV_X1 U7739 ( .A(n6007), .ZN(n5985) );
  NAND4_X1 U7740 ( .A1(n10243), .A2(n6185), .A3(n6128), .A4(n5982), .ZN(n6006)
         );
  INV_X1 U7741 ( .A(n6006), .ZN(n5984) );
  NOR2_X1 U7742 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5983) );
  NOR2_X1 U7743 ( .A1(n5986), .A2(n9111), .ZN(n5987) );
  NAND2_X1 U7744 ( .A1(n5987), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5992) );
  INV_X1 U7745 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5988) );
  NOR2_X1 U7746 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  NAND2_X1 U7747 ( .A1(n8853), .A2(n6246), .ZN(n5999) );
  INV_X1 U7748 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U7749 ( .A1(n4399), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7750 ( .A1(n6827), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5995) );
  OAI211_X1 U7751 ( .C1(n6830), .C2(n10341), .A(n5996), .B(n5995), .ZN(n5997)
         );
  INV_X1 U7752 ( .A(n5997), .ZN(n5998) );
  NAND2_X1 U7753 ( .A1(n6000), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6002) );
  INV_X1 U7754 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6001) );
  XNOR2_X2 U7755 ( .A(n6002), .B(n6001), .ZN(n6342) );
  NAND2_X1 U7756 ( .A1(n6003), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n6004) );
  INV_X4 U7757 ( .A(n6127), .ZN(n6844) );
  NAND2_X1 U7758 ( .A1(n7864), .A2(n6844), .ZN(n6011) );
  NAND2_X2 U7759 ( .A1(n6034), .A2(n4815), .ZN(n6189) );
  INV_X1 U7760 ( .A(n6189), .ZN(n6014) );
  NAND2_X1 U7761 ( .A1(n6363), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6009) );
  XNOR2_X1 U7762 ( .A(n6009), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8674) );
  AOI22_X1 U7763 ( .A1(n6213), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8674), .B2(
        n6227), .ZN(n6010) );
  INV_X1 U7764 ( .A(n9077), .ZN(n8437) );
  NAND2_X1 U7765 ( .A1(n6013), .A2(n6039), .ZN(n6016) );
  NAND2_X1 U7766 ( .A1(n6014), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7767 ( .A1(n4415), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7768 ( .A1(n4415), .A2(n6018), .ZN(n6022) );
  NAND2_X1 U7769 ( .A1(n6036), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7770 ( .A1(n4399), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7771 ( .A1(n6035), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6019) );
  NAND4_X2 U7772 ( .A1(n6022), .A2(n6021), .A3(n6020), .A4(n6019), .ZN(n8996)
         );
  NAND2_X1 U7773 ( .A1(n10104), .A2(n8996), .ZN(n6029) );
  NOR2_X1 U7774 ( .A1(n7302), .A2(n6127), .ZN(n6027) );
  NAND2_X1 U7775 ( .A1(n7433), .A2(n6023), .ZN(n6057) );
  NAND2_X1 U7776 ( .A1(n6057), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6025) );
  XNOR2_X1 U7777 ( .A(n6025), .B(n6024), .ZN(n7506) );
  OAI22_X1 U7778 ( .A1(n6189), .A2(n4703), .B1(n7506), .B2(n7392), .ZN(n6026)
         );
  INV_X1 U7779 ( .A(n10140), .ZN(n10114) );
  NOR2_X1 U7780 ( .A1(n8996), .A2(n6397), .ZN(n6028) );
  AOI22_X1 U7781 ( .A1(n6029), .A2(n10114), .B1(n6028), .B2(n6398), .ZN(n6051)
         );
  NAND2_X1 U7782 ( .A1(n6035), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7783 ( .A1(n4398), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7784 ( .A1(n6036), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7785 ( .A1(n5243), .A2(SI_0_), .ZN(n6033) );
  XNOR2_X1 U7786 ( .A(n6033), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9134) );
  MUX2_X1 U7787 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9134), .S(n6034), .Z(n10136)
         );
  NAND2_X1 U7788 ( .A1(n6723), .A2(n10136), .ZN(n8916) );
  NAND2_X1 U7789 ( .A1(n6036), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7790 ( .A1(n4398), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7791 ( .A1(n6039), .A2(n7307), .ZN(n6045) );
  NAND2_X1 U7792 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6040) );
  NAND2_X1 U7793 ( .A1(n6043), .A2(n7599), .ZN(n6044) );
  OAI211_X2 U7794 ( .C1(n6189), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n6045), .B(
        n6044), .ZN(n6396) );
  OAI21_X1 U7795 ( .B1(n8916), .B2(n8999), .A(n6396), .ZN(n6047) );
  NAND2_X1 U7796 ( .A1(n8916), .A2(n8999), .ZN(n6046) );
  NAND2_X1 U7797 ( .A1(n6047), .A2(n6046), .ZN(n8994) );
  NAND2_X1 U7798 ( .A1(n8994), .A2(n6049), .ZN(n6050) );
  NAND2_X1 U7799 ( .A1(n6051), .A2(n6050), .ZN(n7743) );
  NAND2_X1 U7800 ( .A1(n6847), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7801 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6052) );
  NAND2_X1 U7802 ( .A1(n6070), .A2(n6052), .ZN(n8459) );
  NAND2_X1 U7803 ( .A1(n4415), .A2(n8459), .ZN(n6055) );
  NAND2_X1 U7804 ( .A1(n6083), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7805 ( .A1(n4399), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6053) );
  NAND4_X1 U7806 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n10109)
         );
  NAND2_X1 U7807 ( .A1(n7300), .A2(n6844), .ZN(n6060) );
  NAND2_X1 U7808 ( .A1(n6064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6058) );
  AOI22_X1 U7809 ( .A1(n6014), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7555), .B2(
        n6043), .ZN(n6059) );
  NAND2_X1 U7810 ( .A1(n10109), .A2(n8458), .ZN(n6061) );
  NAND2_X1 U7811 ( .A1(n7743), .A2(n6061), .ZN(n6063) );
  INV_X1 U7812 ( .A(n10109), .ZN(n7531) );
  NAND2_X1 U7813 ( .A1(n7531), .A2(n10147), .ZN(n6062) );
  OR2_X1 U7814 ( .A1(n8332), .A2(n6127), .ZN(n6069) );
  INV_X1 U7815 ( .A(n6064), .ZN(n6066) );
  INV_X1 U7816 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7817 ( .A1(n6066), .A2(n6065), .ZN(n6077) );
  NAND2_X1 U7818 ( .A1(n6077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7819 ( .A(n6067), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7553) );
  AOI22_X1 U7820 ( .A1(n6213), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7553), .B2(
        n6227), .ZN(n6068) );
  INV_X1 U7821 ( .A(n10152), .ZN(n7761) );
  NAND2_X1 U7822 ( .A1(n6847), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7823 ( .A1(n6070), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7824 ( .A1(n6081), .A2(n6071), .ZN(n7764) );
  NAND2_X1 U7825 ( .A1(n6246), .A2(n7764), .ZN(n6074) );
  NAND2_X1 U7826 ( .A1(n6083), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7827 ( .A1(n4399), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6072) );
  NAND4_X1 U7828 ( .A1(n6075), .A2(n6074), .A3(n6073), .A4(n6072), .ZN(n8552)
         );
  NAND2_X1 U7829 ( .A1(n7761), .A2(n8552), .ZN(n6867) );
  NAND2_X1 U7830 ( .A1(n7754), .A2(n6867), .ZN(n6076) );
  INV_X1 U7831 ( .A(n8552), .ZN(n7838) );
  NAND2_X1 U7832 ( .A1(n10152), .A2(n7838), .ZN(n6868) );
  NAND2_X1 U7833 ( .A1(n7312), .A2(n6844), .ZN(n6080) );
  OAI21_X1 U7834 ( .B1(n6077), .B2(P2_IR_REG_5__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6078) );
  AOI22_X1 U7835 ( .A1(n6213), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7604), .B2(
        n6227), .ZN(n6079) );
  NAND2_X1 U7836 ( .A1(n6847), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7837 ( .A1(n6081), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7838 ( .A1(n6096), .A2(n6082), .ZN(n7857) );
  NAND2_X1 U7839 ( .A1(n4415), .A2(n7857), .ZN(n6087) );
  NAND2_X1 U7840 ( .A1(n6083), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7841 ( .A1(n4399), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6085) );
  NAND4_X1 U7842 ( .A1(n6088), .A2(n6087), .A3(n6086), .A4(n6085), .ZN(n8551)
         );
  NAND2_X1 U7843 ( .A1(n7732), .A2(n8551), .ZN(n6089) );
  OR2_X1 U7844 ( .A1(n7315), .A2(n6127), .ZN(n6095) );
  INV_X1 U7845 ( .A(n6090), .ZN(n6092) );
  NAND2_X1 U7846 ( .A1(n6092), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6091) );
  MUX2_X1 U7847 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6091), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6093) );
  AOI22_X1 U7848 ( .A1(n6213), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7611), .B2(
        n6227), .ZN(n6094) );
  AND2_X2 U7849 ( .A1(n6095), .A2(n6094), .ZN(n7906) );
  NAND2_X1 U7850 ( .A1(n6847), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7851 ( .A1(n6096), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7852 ( .A1(n6106), .A2(n6097), .ZN(n7973) );
  NAND2_X1 U7853 ( .A1(n6246), .A2(n7973), .ZN(n6100) );
  NAND2_X1 U7854 ( .A1(n6083), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7855 ( .A1(n4399), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7856 ( .A1(n7906), .A2(n8550), .ZN(n7881) );
  INV_X1 U7857 ( .A(n7906), .ZN(n7972) );
  NAND2_X1 U7858 ( .A1(n7886), .A2(n7972), .ZN(n6756) );
  NAND2_X1 U7859 ( .A1(n7906), .A2(n7886), .ZN(n6102) );
  NAND2_X1 U7860 ( .A1(n7310), .A2(n6844), .ZN(n6105) );
  NAND2_X1 U7861 ( .A1(n6114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6103) );
  XNOR2_X1 U7862 ( .A(n6103), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7794) );
  AOI22_X1 U7863 ( .A1(n6213), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7794), .B2(
        n6227), .ZN(n6104) );
  NAND2_X1 U7864 ( .A1(n6105), .A2(n6104), .ZN(n8391) );
  NAND2_X1 U7865 ( .A1(n6847), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7866 ( .A1(n6106), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7867 ( .A1(n6119), .A2(n6107), .ZN(n8393) );
  NAND2_X1 U7868 ( .A1(n6246), .A2(n8393), .ZN(n6110) );
  NAND2_X1 U7869 ( .A1(n6083), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7870 ( .A1(n4399), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6108) );
  NAND4_X1 U7871 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n8549)
         );
  NAND2_X1 U7872 ( .A1(n8391), .A2(n8549), .ZN(n6112) );
  OR2_X1 U7873 ( .A1(n8391), .A2(n8549), .ZN(n6113) );
  NAND2_X1 U7874 ( .A1(n7345), .A2(n6844), .ZN(n6118) );
  INV_X1 U7875 ( .A(n6114), .ZN(n6116) );
  INV_X1 U7876 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7877 ( .A1(n6116), .A2(n6115), .ZN(n6142) );
  NAND2_X1 U7878 ( .A1(n6142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U7879 ( .A(n6129), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7911) );
  AOI22_X1 U7880 ( .A1(n6213), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7911), .B2(
        n6227), .ZN(n6117) );
  NAND2_X1 U7881 ( .A1(n6847), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7882 ( .A1(n6119), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7883 ( .A1(n6134), .A2(n6120), .ZN(n8224) );
  NAND2_X1 U7884 ( .A1(n6246), .A2(n8224), .ZN(n6123) );
  NAND2_X1 U7885 ( .A1(n4399), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7886 ( .A1(n6827), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6121) );
  NAND4_X1 U7887 ( .A1(n6124), .A2(n6123), .A3(n6122), .A4(n6121), .ZN(n8548)
         );
  NAND2_X1 U7888 ( .A1(n8044), .A2(n8548), .ZN(n6125) );
  OR2_X1 U7889 ( .A1(n8044), .A2(n8548), .ZN(n6126) );
  OR2_X1 U7890 ( .A1(n7344), .A2(n6127), .ZN(n6133) );
  NAND2_X1 U7891 ( .A1(n6129), .A2(n6128), .ZN(n6130) );
  NAND2_X1 U7892 ( .A1(n6130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6131) );
  XNOR2_X1 U7893 ( .A(n6131), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8185) );
  AOI22_X1 U7894 ( .A1(n6213), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8185), .B2(
        n6227), .ZN(n6132) );
  NAND2_X1 U7895 ( .A1(n6847), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7896 ( .A1(n6134), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7897 ( .A1(n6148), .A2(n6135), .ZN(n8373) );
  NAND2_X1 U7898 ( .A1(n6246), .A2(n8373), .ZN(n6138) );
  NAND2_X1 U7899 ( .A1(n6083), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7900 ( .A1(n4399), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6136) );
  NAND4_X1 U7901 ( .A1(n6139), .A2(n6138), .A3(n6137), .A4(n6136), .ZN(n8547)
         );
  NAND2_X1 U7902 ( .A1(n8983), .A2(n8547), .ZN(n6140) );
  OR2_X1 U7903 ( .A1(n8983), .A2(n8547), .ZN(n6141) );
  NAND2_X1 U7904 ( .A1(n7350), .A2(n6844), .ZN(n6147) );
  INV_X1 U7905 ( .A(n6142), .ZN(n6144) );
  NOR2_X1 U7906 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6143) );
  NAND2_X1 U7907 ( .A1(n6144), .A2(n6143), .ZN(n6156) );
  NAND2_X1 U7908 ( .A1(n6156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6145) );
  XNOR2_X1 U7909 ( .A(n6145), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8243) );
  AOI22_X1 U7910 ( .A1(n6213), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8243), .B2(
        n6227), .ZN(n6146) );
  NAND2_X1 U7911 ( .A1(n6847), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7912 ( .A1(n6148), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7913 ( .A1(n6160), .A2(n6149), .ZN(n8506) );
  NAND2_X1 U7914 ( .A1(n6246), .A2(n8506), .ZN(n6152) );
  NAND2_X1 U7915 ( .A1(n6083), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7916 ( .A1(n4399), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6150) );
  NAND4_X1 U7917 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n8546)
         );
  NOR2_X1 U7918 ( .A1(n8494), .A2(n8546), .ZN(n6155) );
  NAND2_X1 U7919 ( .A1(n8494), .A2(n8546), .ZN(n6154) );
  NAND2_X1 U7920 ( .A1(n7416), .A2(n6844), .ZN(n6159) );
  NAND2_X1 U7921 ( .A1(n6166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6157) );
  XNOR2_X1 U7922 ( .A(n6157), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8258) );
  AOI22_X1 U7923 ( .A1(n6213), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8258), .B2(
        n6227), .ZN(n6158) );
  NAND2_X1 U7924 ( .A1(n6847), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7925 ( .A1(n6160), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7926 ( .A1(n6169), .A2(n6161), .ZN(n8415) );
  NAND2_X1 U7927 ( .A1(n6246), .A2(n8415), .ZN(n6164) );
  NAND2_X1 U7928 ( .A1(n6827), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7929 ( .A1(n4399), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6162) );
  NAND4_X1 U7930 ( .A1(n6165), .A2(n6164), .A3(n6163), .A4(n6162), .ZN(n8904)
         );
  NAND2_X1 U7931 ( .A1(n7512), .A2(n6844), .ZN(n6168) );
  OAI21_X1 U7932 ( .B1(n6166), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6175) );
  XNOR2_X1 U7933 ( .A(n6175), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8572) );
  AOI22_X1 U7934 ( .A1(n6213), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8572), .B2(
        n6227), .ZN(n6167) );
  NAND2_X1 U7935 ( .A1(n6847), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7936 ( .A1(n6169), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7937 ( .A1(n6179), .A2(n6170), .ZN(n8908) );
  NAND2_X1 U7938 ( .A1(n6246), .A2(n8908), .ZN(n6173) );
  NAND2_X1 U7939 ( .A1(n6827), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7940 ( .A1(n4399), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7941 ( .A1(n8900), .A2(n8887), .ZN(n6771) );
  NAND2_X1 U7942 ( .A1(n6772), .A2(n6771), .ZN(n8901) );
  NAND2_X1 U7943 ( .A1(n8900), .A2(n8545), .ZN(n8870) );
  NAND2_X1 U7944 ( .A1(n7490), .A2(n6844), .ZN(n6178) );
  NAND2_X1 U7945 ( .A1(n6175), .A2(n10479), .ZN(n6176) );
  NAND2_X1 U7946 ( .A1(n6176), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6186) );
  XNOR2_X1 U7947 ( .A(n6186), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8587) );
  AOI22_X1 U7948 ( .A1(n8587), .A2(n6227), .B1(n6213), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7949 ( .A1(n6179), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7950 ( .A1(n6193), .A2(n6180), .ZN(n8895) );
  NAND2_X1 U7951 ( .A1(n8895), .A2(n6246), .ZN(n6184) );
  NAND2_X1 U7952 ( .A1(n6847), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7953 ( .A1(n6827), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7954 ( .A1(n4399), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6181) );
  NAND4_X1 U7955 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n8903)
         );
  NAND2_X1 U7956 ( .A1(n9093), .A2(n8903), .ZN(n8872) );
  NAND2_X1 U7957 ( .A1(n8869), .A2(n5236), .ZN(n6200) );
  NAND2_X1 U7958 ( .A1(n7704), .A2(n6844), .ZN(n6192) );
  NAND2_X1 U7959 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  NAND2_X1 U7960 ( .A1(n6187), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6188) );
  XNOR2_X1 U7961 ( .A(n6188), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8618) );
  INV_X1 U7962 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10451) );
  NOR2_X1 U7963 ( .A1(n6189), .A2(n10451), .ZN(n6190) );
  AOI21_X1 U7964 ( .B1(n8618), .B2(n6227), .A(n6190), .ZN(n6191) );
  NAND2_X1 U7965 ( .A1(n6193), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7966 ( .A1(n6204), .A2(n6194), .ZN(n8879) );
  NAND2_X1 U7967 ( .A1(n8879), .A2(n6246), .ZN(n6197) );
  AOI22_X1 U7968 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n6847), .B1(n6083), .B2(
        P2_REG0_REG_15__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7969 ( .A1(n4399), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7970 ( .A1(n8963), .A2(n8889), .ZN(n6408) );
  NAND2_X1 U7971 ( .A1(n6779), .A2(n6408), .ZN(n8871) );
  INV_X1 U7972 ( .A(n8903), .ZN(n8536) );
  NAND2_X1 U7973 ( .A1(n9093), .A2(n8536), .ZN(n6776) );
  NAND2_X1 U7974 ( .A1(n6775), .A2(n6776), .ZN(n8897) );
  NAND2_X1 U7975 ( .A1(n6200), .A2(n5235), .ZN(n8875) );
  INV_X1 U7976 ( .A(n8963), .ZN(n9088) );
  NAND2_X1 U7977 ( .A1(n7779), .A2(n6844), .ZN(n6203) );
  NAND2_X1 U7978 ( .A1(n4502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6201) );
  XNOR2_X1 U7979 ( .A(n6201), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8636) );
  AOI22_X1 U7980 ( .A1(n6213), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8636), .B2(
        n6227), .ZN(n6202) );
  NAND2_X1 U7981 ( .A1(n6204), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7982 ( .A1(n6206), .A2(n6205), .ZN(n8865) );
  NAND2_X1 U7983 ( .A1(n8865), .A2(n6246), .ZN(n6209) );
  AOI22_X1 U7984 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n6847), .B1(n6827), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7985 ( .A1(n4399), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7986 ( .A1(n9083), .A2(n8878), .ZN(n6785) );
  NAND2_X1 U7987 ( .A1(n6784), .A2(n6785), .ZN(n8858) );
  INV_X1 U7988 ( .A(n9083), .ZN(n8429) );
  NAND2_X1 U7989 ( .A1(n7934), .A2(n6844), .ZN(n6215) );
  NAND2_X1 U7990 ( .A1(n6334), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6211) );
  INV_X1 U7991 ( .A(n6211), .ZN(n6210) );
  NAND2_X1 U7992 ( .A1(n6210), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7993 ( .A1(n6211), .A2(n6332), .ZN(n6225) );
  AND2_X1 U7994 ( .A1(n6212), .A2(n6225), .ZN(n8709) );
  AOI22_X1 U7995 ( .A1(n6213), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8709), .B2(
        n6227), .ZN(n6214) );
  NAND2_X1 U7996 ( .A1(n6216), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7997 ( .A1(n6232), .A2(n6217), .ZN(n8836) );
  NAND2_X1 U7998 ( .A1(n8836), .A2(n6246), .ZN(n6222) );
  INV_X1 U7999 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10231) );
  NAND2_X1 U8000 ( .A1(n4399), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U8001 ( .A1(n6827), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6218) );
  OAI211_X1 U8002 ( .C1(n6830), .C2(n10231), .A(n6219), .B(n6218), .ZN(n6220)
         );
  INV_X1 U8003 ( .A(n6220), .ZN(n6221) );
  NAND2_X1 U8004 ( .A1(n7219), .A2(n7222), .ZN(n6224) );
  NAND2_X1 U8005 ( .A1(n8116), .A2(n6844), .ZN(n6229) );
  AOI22_X1 U8006 ( .A1(n6213), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7164), .B2(
        n6227), .ZN(n6228) );
  INV_X1 U8007 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U8008 ( .A1(n6232), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U8009 ( .A1(n6241), .A2(n6233), .ZN(n8827) );
  NAND2_X1 U8010 ( .A1(n8827), .A2(n6246), .ZN(n6238) );
  INV_X1 U8011 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10374) );
  NAND2_X1 U8012 ( .A1(n6083), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U8013 ( .A1(n4399), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6234) );
  OAI211_X1 U8014 ( .C1(n6830), .C2(n10374), .A(n6235), .B(n6234), .ZN(n6236)
         );
  INV_X1 U8015 ( .A(n6236), .ZN(n6237) );
  NAND2_X1 U8016 ( .A1(n9068), .A2(n8835), .ZN(n6796) );
  INV_X1 U8017 ( .A(n9068), .ZN(n8383) );
  NAND2_X1 U8018 ( .A1(n8210), .A2(n6844), .ZN(n6240) );
  NAND2_X1 U8019 ( .A1(n6213), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U8020 ( .A1(n6241), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U8021 ( .A1(n6249), .A2(n6242), .ZN(n8815) );
  INV_X1 U8022 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U8023 ( .A1(n6827), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U8024 ( .A1(n4399), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6243) );
  OAI211_X1 U8025 ( .C1(n6830), .C2(n10320), .A(n6244), .B(n6243), .ZN(n6245)
         );
  NAND2_X1 U8026 ( .A1(n9062), .A2(n8402), .ZN(n6795) );
  NAND2_X1 U8027 ( .A1(n8265), .A2(n6844), .ZN(n6248) );
  NAND2_X1 U8028 ( .A1(n6213), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U8029 ( .A1(n6249), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U8030 ( .A1(n6258), .A2(n6250), .ZN(n8805) );
  NAND2_X1 U8031 ( .A1(n8805), .A2(n6246), .ZN(n6255) );
  INV_X1 U8032 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10267) );
  NAND2_X1 U8033 ( .A1(n6827), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U8034 ( .A1(n4399), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6251) );
  OAI211_X1 U8035 ( .C1(n6830), .C2(n10267), .A(n6252), .B(n6251), .ZN(n6253)
         );
  INV_X1 U8036 ( .A(n6253), .ZN(n6254) );
  NAND2_X1 U8037 ( .A1(n9056), .A2(n8468), .ZN(n6800) );
  NAND2_X1 U8038 ( .A1(n6789), .A2(n6800), .ZN(n8800) );
  NAND2_X1 U8039 ( .A1(n7227), .A2(n8468), .ZN(n8786) );
  NAND2_X1 U8040 ( .A1(n8270), .A2(n6844), .ZN(n6257) );
  NAND2_X1 U8041 ( .A1(n6213), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U8042 ( .A1(n6258), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U8043 ( .A1(n6268), .A2(n6259), .ZN(n8793) );
  NAND2_X1 U8044 ( .A1(n8793), .A2(n6246), .ZN(n6264) );
  INV_X1 U8045 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U8046 ( .A1(n6847), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U8047 ( .A1(n6827), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6260) );
  OAI211_X1 U8048 ( .C1(n8792), .C2(n6327), .A(n6261), .B(n6260), .ZN(n6262)
         );
  INV_X1 U8049 ( .A(n6262), .ZN(n6263) );
  NAND2_X1 U8050 ( .A1(n9050), .A2(n8777), .ZN(n6804) );
  NAND2_X1 U8051 ( .A1(n6805), .A2(n6804), .ZN(n8785) );
  NAND2_X1 U8052 ( .A1(n8306), .A2(n6844), .ZN(n6267) );
  NAND2_X1 U8053 ( .A1(n6213), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U8054 ( .A1(n6268), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U8055 ( .A1(n6282), .A2(n6269), .ZN(n8781) );
  NAND2_X1 U8056 ( .A1(n8781), .A2(n6246), .ZN(n6274) );
  INV_X1 U8057 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U8058 ( .A1(n6847), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U8059 ( .A1(n6827), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6270) );
  OAI211_X1 U8060 ( .C1(n8780), .C2(n6327), .A(n6271), .B(n6270), .ZN(n6272)
         );
  INV_X1 U8061 ( .A(n6272), .ZN(n6273) );
  NAND2_X1 U8062 ( .A1(n6416), .A2(n8790), .ZN(n6277) );
  NAND2_X1 U8063 ( .A1(n9044), .A2(n8761), .ZN(n6275) );
  NAND2_X1 U8064 ( .A1(n8310), .A2(n6844), .ZN(n6279) );
  NAND2_X1 U8065 ( .A1(n6213), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6278) );
  INV_X1 U8066 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U8067 ( .A1(n6282), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U8068 ( .A1(n6291), .A2(n6283), .ZN(n8764) );
  NAND2_X1 U8069 ( .A1(n8764), .A2(n6246), .ZN(n6288) );
  INV_X1 U8070 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U8071 ( .A1(n6827), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U8072 ( .A1(n4399), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6284) );
  OAI211_X1 U8073 ( .C1(n6830), .C2(n10470), .A(n6285), .B(n6284), .ZN(n6286)
         );
  INV_X1 U8074 ( .A(n6286), .ZN(n6287) );
  NAND2_X1 U8075 ( .A1(n9129), .A2(n6844), .ZN(n6290) );
  NAND2_X1 U8076 ( .A1(n6213), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U8077 ( .A1(n6291), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6292) );
  NAND2_X1 U8078 ( .A1(n6300), .A2(n6292), .ZN(n8749) );
  NAND2_X1 U8079 ( .A1(n8749), .A2(n6246), .ZN(n6297) );
  INV_X1 U8080 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U8081 ( .A1(n6847), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U8082 ( .A1(n6827), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6293) );
  OAI211_X1 U8083 ( .C1(n8754), .C2(n6327), .A(n6294), .B(n6293), .ZN(n6295)
         );
  INV_X1 U8084 ( .A(n6295), .ZN(n6296) );
  NAND2_X1 U8085 ( .A1(n9033), .A2(n8739), .ZN(n6810) );
  NOR2_X1 U8086 ( .A1(n9033), .A2(n8739), .ZN(n6812) );
  NAND2_X1 U8087 ( .A1(n9126), .A2(n6844), .ZN(n6299) );
  NAND2_X1 U8088 ( .A1(n6213), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U8089 ( .A1(n6300), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U8090 ( .A1(n6312), .A2(n6301), .ZN(n8742) );
  NAND2_X1 U8091 ( .A1(n8742), .A2(n6246), .ZN(n6306) );
  INV_X1 U8092 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n10441) );
  NAND2_X1 U8093 ( .A1(n6847), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U8094 ( .A1(n6083), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6302) );
  OAI211_X1 U8095 ( .C1(n10441), .C2(n6327), .A(n6303), .B(n6302), .ZN(n6304)
         );
  INV_X1 U8096 ( .A(n6304), .ZN(n6305) );
  NAND2_X1 U8097 ( .A1(n7243), .A2(n8422), .ZN(n6307) );
  NAND2_X1 U8098 ( .A1(n9124), .A2(n6844), .ZN(n6309) );
  NAND2_X1 U8099 ( .A1(n6213), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6308) );
  INV_X1 U8100 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U8101 ( .A1(n6312), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U8102 ( .A1(n6323), .A2(n6313), .ZN(n8732) );
  NAND2_X1 U8103 ( .A1(n8732), .A2(n6246), .ZN(n6318) );
  INV_X1 U8104 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U8105 ( .A1(n6847), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U8106 ( .A1(n6827), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6314) );
  OAI211_X1 U8107 ( .C1(n8731), .C2(n6327), .A(n6315), .B(n6314), .ZN(n6316)
         );
  INV_X1 U8108 ( .A(n6316), .ZN(n6317) );
  NAND2_X1 U8109 ( .A1(n9021), .A2(n8740), .ZN(n6320) );
  INV_X1 U8110 ( .A(n9021), .ZN(n6319) );
  NAND2_X1 U8111 ( .A1(n8316), .A2(n6844), .ZN(n6322) );
  NAND2_X1 U8112 ( .A1(n6213), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U8113 ( .A1(n6323), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U8114 ( .A1(n8334), .A2(n6324), .ZN(n7277) );
  NAND2_X1 U8115 ( .A1(n7277), .A2(n6246), .ZN(n6330) );
  NAND2_X1 U8116 ( .A1(n6847), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U8117 ( .A1(n6827), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6325) );
  OAI211_X1 U8118 ( .C1(n6712), .C2(n6327), .A(n6326), .B(n6325), .ZN(n6328)
         );
  INV_X1 U8119 ( .A(n6328), .ZN(n6329) );
  XNOR2_X1 U8120 ( .A(n7144), .B(n6883), .ZN(n6352) );
  NAND2_X1 U8121 ( .A1(n6332), .A2(n6331), .ZN(n6333) );
  NAND2_X1 U8122 ( .A1(n6353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U8123 ( .A1(n6910), .A2(n7164), .ZN(n6424) );
  INV_X1 U8124 ( .A(n6338), .ZN(n6339) );
  INV_X1 U8125 ( .A(n8215), .ZN(n7162) );
  NAND2_X1 U8126 ( .A1(n6724), .A2(n7162), .ZN(n6896) );
  INV_X1 U8127 ( .A(n6342), .ZN(n7390) );
  XNOR2_X1 U8128 ( .A(n7390), .B(n4387), .ZN(n7262) );
  INV_X1 U8129 ( .A(n7262), .ZN(n7263) );
  INV_X1 U8130 ( .A(n8334), .ZN(n6343) );
  INV_X1 U8131 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U8132 ( .A1(n6827), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U8133 ( .A1(n4399), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6344) );
  OAI211_X1 U8134 ( .C1(n6830), .C2(n6346), .A(n6345), .B(n6344), .ZN(n6347)
         );
  INV_X1 U8135 ( .A(n6347), .ZN(n6348) );
  OAI21_X1 U8136 ( .B1(n6352), .B2(n10132), .A(n6351), .ZN(n6708) );
  OAI21_X1 U8137 ( .B1(n6353), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U8138 ( .A(n6355), .B(n6354), .ZN(n7399) );
  AND2_X1 U8139 ( .A1(n6357), .A2(n6356), .ZN(n6364) );
  INV_X1 U8140 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U8141 ( .A1(n6364), .A2(n6358), .ZN(n6368) );
  NAND2_X1 U8142 ( .A1(n6368), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6359) );
  MUX2_X1 U8143 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6359), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6360) );
  AND2_X1 U8144 ( .A1(n6361), .A2(n6360), .ZN(n6376) );
  INV_X1 U8145 ( .A(n6364), .ZN(n6366) );
  NAND2_X1 U8146 ( .A1(n6366), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6367) );
  MUX2_X1 U8147 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6367), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6369) );
  NAND2_X1 U8148 ( .A1(n6369), .A2(n6368), .ZN(n9133) );
  INV_X1 U8149 ( .A(n9133), .ZN(n6370) );
  NAND3_X1 U8150 ( .A1(n6376), .A2(n6371), .A3(n6370), .ZN(n7292) );
  XNOR2_X1 U8151 ( .A(n8312), .B(P2_B_REG_SCAN_IN), .ZN(n6372) );
  NAND2_X1 U8152 ( .A1(n6372), .A2(n9133), .ZN(n6373) );
  INV_X1 U8153 ( .A(n6376), .ZN(n9128) );
  NAND2_X1 U8154 ( .A1(n9128), .A2(n8312), .ZN(n7334) );
  OR2_X1 U8155 ( .A1(n6377), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U8156 ( .A1(n9128), .A2(n9133), .ZN(n7336) );
  NAND2_X1 U8157 ( .A1(n6702), .A2(n6430), .ZN(n6427) );
  NOR2_X1 U8158 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .ZN(
        n10351) );
  NOR4_X1 U8159 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6381) );
  NOR4_X1 U8160 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6380) );
  NOR4_X1 U8161 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6379) );
  NAND4_X1 U8162 ( .A1(n10351), .A2(n6381), .A3(n6380), .A4(n6379), .ZN(n6387)
         );
  NOR4_X1 U8163 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6385) );
  NOR4_X1 U8164 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6384) );
  NOR4_X1 U8165 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6383) );
  NOR4_X1 U8166 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6382) );
  NAND4_X1 U8167 ( .A1(n6385), .A2(n6384), .A3(n6383), .A4(n6382), .ZN(n6386)
         );
  NOR2_X1 U8168 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  NAND2_X1 U8169 ( .A1(n8704), .A2(n8215), .ZN(n6856) );
  NAND2_X1 U8170 ( .A1(n7293), .A2(n6856), .ZN(n7268) );
  NAND4_X1 U8171 ( .A1(n7333), .A2(n6427), .A3(n6426), .A4(n7268), .ZN(n6705)
         );
  NAND2_X1 U8172 ( .A1(n6910), .A2(n8704), .ZN(n6419) );
  OR2_X1 U8173 ( .A1(n6419), .A2(n8215), .ZN(n6389) );
  NAND2_X1 U8174 ( .A1(n9008), .A2(n8266), .ZN(n6706) );
  NAND2_X1 U8175 ( .A1(n6706), .A2(n6702), .ZN(n6390) );
  NAND2_X1 U8176 ( .A1(n6703), .A2(n6390), .ZN(n6393) );
  INV_X1 U8177 ( .A(n6703), .ZN(n6391) );
  INV_X1 U8178 ( .A(n6430), .ZN(n6700) );
  NAND2_X1 U8179 ( .A1(n6391), .A2(n6700), .ZN(n6392) );
  NAND2_X1 U8180 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  MUX2_X1 U8181 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n6708), .S(n10166), .Z(n6395) );
  INV_X1 U8182 ( .A(n6395), .ZN(n6423) );
  INV_X1 U8183 ( .A(n6730), .ZN(n6400) );
  NAND2_X1 U8184 ( .A1(n7530), .A2(n9004), .ZN(n6731) );
  XNOR2_X1 U8185 ( .A(n8996), .B(n10140), .ZN(n10112) );
  NAND2_X1 U8186 ( .A1(n10113), .A2(n10112), .ZN(n6401) );
  INV_X1 U8187 ( .A(n8996), .ZN(n7468) );
  NAND2_X1 U8188 ( .A1(n7468), .A2(n10140), .ZN(n6739) );
  NAND2_X1 U8189 ( .A1(n6401), .A2(n6739), .ZN(n7741) );
  NAND2_X1 U8190 ( .A1(n10109), .A2(n10147), .ZN(n7748) );
  AND2_X1 U8191 ( .A1(n6742), .A2(n7748), .ZN(n6737) );
  NAND2_X1 U8192 ( .A1(n7761), .A2(n7838), .ZN(n6740) );
  OR2_X1 U8193 ( .A1(n7732), .A2(n7772), .ZN(n6743) );
  NAND2_X1 U8194 ( .A1(n7732), .A2(n7772), .ZN(n6749) );
  OR2_X1 U8195 ( .A1(n8391), .A2(n8221), .ZN(n6865) );
  AND2_X1 U8196 ( .A1(n6865), .A2(n7881), .ZN(n6754) );
  NAND2_X1 U8197 ( .A1(n7820), .A2(n6754), .ZN(n6402) );
  NAND2_X1 U8198 ( .A1(n8391), .A2(n8221), .ZN(n6864) );
  NAND2_X1 U8199 ( .A1(n8983), .A2(n8504), .ZN(n8146) );
  INV_X1 U8200 ( .A(n8548), .ZN(n8369) );
  NAND2_X1 U8201 ( .A1(n8044), .A2(n8369), .ZN(n6859) );
  NAND2_X1 U8202 ( .A1(n8146), .A2(n6859), .ZN(n6757) );
  OR2_X1 U8203 ( .A1(n8494), .A2(n8412), .ZN(n6763) );
  INV_X1 U8204 ( .A(n8044), .ZN(n8218) );
  NAND2_X1 U8205 ( .A1(n8012), .A2(n8504), .ZN(n6403) );
  AOI22_X1 U8206 ( .A1(n8370), .A2(n6403), .B1(n6861), .B2(n8547), .ZN(n6404)
         );
  XNOR2_X1 U8207 ( .A(n8160), .B(n8478), .ZN(n8163) );
  NAND2_X1 U8208 ( .A1(n8978), .A2(n8904), .ZN(n6767) );
  INV_X1 U8209 ( .A(n6775), .ZN(n6407) );
  INV_X1 U8210 ( .A(n6408), .ZN(n6782) );
  NAND2_X1 U8211 ( .A1(n9077), .A2(n8861), .ZN(n6790) );
  NAND2_X1 U8212 ( .A1(n8954), .A2(n7222), .ZN(n6791) );
  NAND2_X1 U8213 ( .A1(n8820), .A2(n6791), .ZN(n8832) );
  AND2_X1 U8214 ( .A1(n6788), .A2(n8820), .ZN(n6793) );
  NAND2_X1 U8215 ( .A1(n6411), .A2(n6796), .ZN(n8808) );
  INV_X1 U8216 ( .A(n6795), .ZN(n6412) );
  NAND2_X1 U8217 ( .A1(n8797), .A2(n6800), .ZN(n6413) );
  NAND2_X1 U8218 ( .A1(n6413), .A2(n6789), .ZN(n8784) );
  NAND2_X1 U8219 ( .A1(n8784), .A2(n6804), .ZN(n6414) );
  NAND2_X1 U8220 ( .A1(n9039), .A2(n8778), .ZN(n8758) );
  NAND2_X1 U8221 ( .A1(n6416), .A2(n8761), .ZN(n8771) );
  NOR2_X1 U8222 ( .A1(n9033), .A2(n8762), .ZN(n6814) );
  NAND2_X1 U8223 ( .A1(n9033), .A2(n8762), .ZN(n6813) );
  NAND2_X1 U8224 ( .A1(n9021), .A2(n7280), .ZN(n6817) );
  XNOR2_X1 U8225 ( .A(n6888), .B(n6883), .ZN(n6710) );
  INV_X1 U8226 ( .A(n6856), .ZN(n6418) );
  NAND2_X1 U8227 ( .A1(n7293), .A2(n6418), .ZN(n6909) );
  AND2_X1 U8228 ( .A1(n6909), .A2(n10151), .ZN(n7736) );
  NAND2_X1 U8229 ( .A1(n6419), .A2(n6856), .ZN(n6420) );
  INV_X1 U8230 ( .A(n9008), .ZN(n10153) );
  OAI22_X1 U8231 ( .A1(n6710), .A2(n8972), .B1(n7147), .B2(n8971), .ZN(n6421)
         );
  INV_X1 U8232 ( .A(n6421), .ZN(n6422) );
  NAND2_X1 U8233 ( .A1(n8266), .A2(n7162), .ZN(n6425) );
  AND2_X1 U8234 ( .A1(n7271), .A2(n6909), .ZN(n6428) );
  INV_X1 U8235 ( .A(n6426), .ZN(n6429) );
  NOR2_X1 U8236 ( .A1(n6427), .A2(n6429), .ZN(n7265) );
  NAND2_X1 U8237 ( .A1(n7265), .A2(n7333), .ZN(n7258) );
  NOR2_X1 U8238 ( .A1(n6430), .A2(n6429), .ZN(n6432) );
  INV_X1 U8239 ( .A(n6702), .ZN(n6431) );
  NAND3_X1 U8240 ( .A1(n7271), .A2(n4402), .A3(n10151), .ZN(n7251) );
  NAND2_X1 U8241 ( .A1(n7251), .A2(n10121), .ZN(n7266) );
  NAND2_X1 U8242 ( .A1(n7261), .A2(n7266), .ZN(n6433) );
  MUX2_X1 U8243 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n6708), .S(n10157), .Z(n6435) );
  INV_X1 U8244 ( .A(n6435), .ZN(n6438) );
  OAI22_X1 U8245 ( .A1(n6710), .A2(n9102), .B1(n7147), .B2(n9100), .ZN(n6436)
         );
  INV_X1 U8246 ( .A(n6436), .ZN(n6437) );
  NAND2_X1 U8247 ( .A1(n6440), .A2(n6439), .ZN(n6539) );
  INV_X1 U8248 ( .A(n6608), .ZN(n6513) );
  AND2_X1 U8249 ( .A1(n6513), .A2(n6630), .ZN(n6520) );
  INV_X1 U8250 ( .A(n6507), .ZN(n6441) );
  AOI21_X1 U8251 ( .B1(n6520), .B2(n6442), .A(n9606), .ZN(n6523) );
  NOR2_X1 U8252 ( .A1(n6443), .A2(n6630), .ZN(n6514) );
  INV_X1 U8253 ( .A(n9700), .ZN(n6444) );
  NAND2_X1 U8254 ( .A1(n6671), .A2(n6444), .ZN(n6491) );
  NAND2_X1 U8255 ( .A1(n6445), .A2(n6630), .ZN(n6451) );
  INV_X1 U8256 ( .A(n7869), .ZN(n6449) );
  NAND2_X1 U8257 ( .A1(n6451), .A2(n6450), .ZN(n6462) );
  NAND2_X1 U8258 ( .A1(n6459), .A2(n6452), .ZN(n6654) );
  OAI211_X1 U8259 ( .C1(n6462), .C2(n6654), .A(n6653), .B(n8025), .ZN(n6453)
         );
  NAND3_X1 U8260 ( .A1(n6453), .A2(n6634), .A3(n8026), .ZN(n6456) );
  NAND2_X1 U8261 ( .A1(n8140), .A2(n6576), .ZN(n6463) );
  NAND2_X1 U8262 ( .A1(n6463), .A2(n6630), .ZN(n6454) );
  NAND2_X1 U8263 ( .A1(n6454), .A2(n8030), .ZN(n6455) );
  NAND2_X1 U8264 ( .A1(n6456), .A2(n6455), .ZN(n6458) );
  OR2_X1 U8265 ( .A1(n8139), .A2(n6630), .ZN(n6457) );
  INV_X1 U8266 ( .A(n6653), .ZN(n6461) );
  AND4_X1 U8267 ( .A1(n6481), .A2(n6630), .A3(n6465), .A4(n6459), .ZN(n6460)
         );
  OAI211_X1 U8268 ( .C1(n6462), .C2(n6461), .A(n6460), .B(n8026), .ZN(n6468)
         );
  INV_X1 U8269 ( .A(n6463), .ZN(n6464) );
  NAND2_X1 U8270 ( .A1(n6464), .A2(n8025), .ZN(n6466) );
  NAND4_X1 U8271 ( .A1(n6466), .A2(n6630), .A3(n6465), .A4(n6481), .ZN(n6467)
         );
  OAI211_X1 U8272 ( .C1(n6630), .C2(n6584), .A(n6468), .B(n6467), .ZN(n6469)
         );
  NAND2_X1 U8273 ( .A1(n6482), .A2(n6470), .ZN(n6472) );
  NAND2_X1 U8274 ( .A1(n6476), .A2(n9980), .ZN(n6663) );
  INV_X1 U8275 ( .A(n6663), .ZN(n6471) );
  NAND2_X1 U8276 ( .A1(n6472), .A2(n6471), .ZN(n6480) );
  NAND2_X1 U8277 ( .A1(n6474), .A2(n6473), .ZN(n6661) );
  INV_X1 U8278 ( .A(n6657), .ZN(n6475) );
  AND2_X1 U8279 ( .A1(n6476), .A2(n6475), .ZN(n6477) );
  NOR2_X1 U8280 ( .A1(n6661), .A2(n6477), .ZN(n6479) );
  INV_X1 U8281 ( .A(n6666), .ZN(n6478) );
  OAI21_X1 U8282 ( .B1(n6483), .B2(n6661), .A(n6666), .ZN(n6484) );
  NAND2_X1 U8283 ( .A1(n6487), .A2(n9700), .ZN(n6641) );
  INV_X1 U8284 ( .A(n9698), .ZN(n6486) );
  NOR2_X1 U8285 ( .A1(n6641), .A2(n6486), .ZN(n6489) );
  INV_X1 U8286 ( .A(n6575), .ZN(n6488) );
  INV_X1 U8287 ( .A(n6492), .ZN(n6494) );
  NAND3_X1 U8288 ( .A1(n9698), .A2(n5073), .A3(n9892), .ZN(n6493) );
  AND2_X1 U8289 ( .A1(n6493), .A2(n9717), .ZN(n6497) );
  NAND2_X1 U8290 ( .A1(n6497), .A2(n6575), .ZN(n6642) );
  AOI21_X1 U8291 ( .B1(n6494), .B2(n9698), .A(n6642), .ZN(n6496) );
  XNOR2_X1 U8292 ( .A(n6671), .B(n6634), .ZN(n6495) );
  OAI21_X1 U8293 ( .B1(n6496), .B2(n5680), .A(n6495), .ZN(n6498) );
  AND2_X1 U8294 ( .A1(n6517), .A2(n6501), .ZN(n6677) );
  NAND2_X1 U8295 ( .A1(n6516), .A2(n6677), .ZN(n6502) );
  AND2_X1 U8296 ( .A1(n6505), .A2(n6515), .ZN(n6674) );
  NAND2_X1 U8297 ( .A1(n6502), .A2(n6674), .ZN(n6511) );
  NAND2_X1 U8298 ( .A1(n6507), .A2(n9854), .ZN(n6503) );
  NAND2_X1 U8299 ( .A1(n6503), .A2(n6634), .ZN(n6504) );
  OR2_X1 U8300 ( .A1(n9845), .A2(n9833), .ZN(n6512) );
  INV_X1 U8301 ( .A(n6505), .ZN(n6506) );
  NAND2_X1 U8302 ( .A1(n6507), .A2(n6634), .ZN(n6508) );
  NAND2_X1 U8303 ( .A1(n6509), .A2(n9860), .ZN(n6510) );
  NAND2_X1 U8304 ( .A1(n6513), .A2(n6512), .ZN(n6615) );
  NAND2_X1 U8305 ( .A1(n6514), .A2(n6615), .ZN(n6522) );
  NAND3_X1 U8306 ( .A1(n6518), .A2(n6517), .A3(n6640), .ZN(n6519) );
  NAND2_X1 U8307 ( .A1(n6528), .A2(n6524), .ZN(n6600) );
  NAND2_X1 U8308 ( .A1(n6600), .A2(n6630), .ZN(n6525) );
  AND2_X1 U8309 ( .A1(n6526), .A2(n9576), .ZN(n6606) );
  INV_X1 U8310 ( .A(n6606), .ZN(n6527) );
  OAI21_X1 U8311 ( .B1(n6630), .B2(n6528), .A(n9575), .ZN(n6529) );
  MUX2_X1 U8312 ( .A(n6602), .B(n6607), .S(n6634), .Z(n6531) );
  AND2_X1 U8313 ( .A1(n6598), .A2(n6605), .ZN(n6533) );
  INV_X1 U8314 ( .A(n6533), .ZN(n6534) );
  AOI21_X1 U8315 ( .B1(n6535), .B2(n6611), .A(n6534), .ZN(n6538) );
  OR3_X1 U8316 ( .A1(n6539), .A2(n6536), .A3(n6634), .ZN(n6537) );
  AND2_X1 U8317 ( .A1(n6539), .A2(n6634), .ZN(n6541) );
  MUX2_X1 U8318 ( .A(n6541), .B(n6630), .S(n6540), .Z(n6543) );
  MUX2_X1 U8319 ( .A(n6620), .B(n6618), .S(n6634), .Z(n6542) );
  INV_X1 U8320 ( .A(SI_29_), .ZN(n6547) );
  INV_X1 U8321 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8341) );
  INV_X1 U8322 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6549) );
  MUX2_X1 U8323 ( .A(n8341), .B(n6549), .S(n4397), .Z(n6550) );
  INV_X1 U8324 ( .A(SI_30_), .ZN(n10359) );
  NAND2_X1 U8325 ( .A1(n6550), .A2(n10359), .ZN(n6558) );
  INV_X1 U8326 ( .A(n6550), .ZN(n6551) );
  NAND2_X1 U8327 ( .A1(n6551), .A2(SI_30_), .ZN(n6552) );
  NAND2_X1 U8328 ( .A1(n6558), .A2(n6552), .ZN(n6559) );
  NAND2_X1 U8329 ( .A1(n8339), .A2(n5923), .ZN(n6554) );
  OR2_X1 U8330 ( .A1(n6565), .A2(n8341), .ZN(n6553) );
  NAND2_X1 U8331 ( .A1(n9772), .A2(n9382), .ZN(n6685) );
  NAND2_X1 U8332 ( .A1(n4391), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U8333 ( .A1(n4388), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8334 ( .A1(n5536), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6555) );
  NAND3_X1 U8335 ( .A1(n6557), .A2(n6556), .A3(n6555), .ZN(n9511) );
  NAND2_X1 U8336 ( .A1(n6685), .A2(n9511), .ZN(n6568) );
  INV_X1 U8337 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6564) );
  MUX2_X1 U8338 ( .A(n6564), .B(n10340), .S(n4397), .Z(n6561) );
  XNOR2_X1 U8339 ( .A(n6561), .B(SI_31_), .ZN(n6562) );
  NAND2_X1 U8340 ( .A1(n9109), .A2(n5923), .ZN(n6567) );
  OR2_X1 U8341 ( .A1(n6565), .A2(n6564), .ZN(n6566) );
  INV_X1 U8342 ( .A(n9511), .ZN(n6574) );
  AOI21_X1 U8343 ( .B1(n9772), .B2(n6574), .A(n9766), .ZN(n6570) );
  XOR2_X1 U8344 ( .A(n9382), .B(n9507), .Z(n6597) );
  INV_X1 U8345 ( .A(n9782), .ZN(n6595) );
  INV_X1 U8346 ( .A(n9575), .ZN(n9571) );
  INV_X1 U8347 ( .A(n7784), .ZN(n7868) );
  NAND3_X1 U8348 ( .A1(n7868), .A2(n6576), .A3(n8269), .ZN(n6582) );
  INV_X1 U8349 ( .A(n6577), .ZN(n7668) );
  NAND2_X1 U8350 ( .A1(n6578), .A2(n6579), .ZN(n6644) );
  NAND2_X1 U8351 ( .A1(n7668), .A2(n6644), .ZN(n8321) );
  INV_X1 U8352 ( .A(n6580), .ZN(n7669) );
  NOR4_X1 U8353 ( .A1(n6582), .A2(n8321), .A3(n7669), .A4(n6581), .ZN(n6583)
         );
  XNOR2_X1 U8354 ( .A(n9389), .B(n10013), .ZN(n7871) );
  NAND2_X1 U8355 ( .A1(n6585), .A2(n8278), .ZN(n6587) );
  NAND2_X1 U8356 ( .A1(n9717), .A2(n6586), .ZN(n9736) );
  NAND4_X1 U8357 ( .A1(n9681), .A2(n9702), .A3(n9719), .A4(n6588), .ZN(n6589)
         );
  NOR4_X1 U8358 ( .A1(n9606), .A2(n9667), .A3(n9650), .A4(n6589), .ZN(n6590)
         );
  NAND4_X1 U8359 ( .A1(n9591), .A2(n6590), .A3(n9628), .A4(n9644), .ZN(n6591)
         );
  NAND4_X1 U8360 ( .A1(n6595), .A2(n6594), .A3(n6593), .A4(n6592), .ZN(n6596)
         );
  NOR2_X1 U8361 ( .A1(n6629), .A2(n7117), .ZN(n6625) );
  AND2_X1 U8362 ( .A1(n6599), .A2(n6598), .ZN(n6679) );
  NAND2_X1 U8363 ( .A1(n6600), .A2(n9576), .ZN(n6601) );
  NAND2_X1 U8364 ( .A1(n6602), .A2(n6601), .ZN(n6603) );
  NAND2_X1 U8365 ( .A1(n6603), .A2(n6607), .ZN(n6604) );
  NAND2_X1 U8366 ( .A1(n6605), .A2(n6604), .ZN(n6616) );
  OAI211_X1 U8367 ( .C1(n6609), .C2(n6608), .A(n6607), .B(n6606), .ZN(n6610)
         );
  INV_X1 U8368 ( .A(n6610), .ZN(n6613) );
  OAI211_X1 U8369 ( .C1(n6616), .C2(n6613), .A(n6612), .B(n6611), .ZN(n6614)
         );
  AOI21_X1 U8370 ( .B1(n6679), .B2(n6614), .A(n6539), .ZN(n6684) );
  NOR2_X1 U8371 ( .A1(n6616), .A2(n6615), .ZN(n6678) );
  NAND3_X1 U8372 ( .A1(n6679), .A2(n6678), .A3(n9645), .ZN(n6619) );
  NAND2_X1 U8373 ( .A1(n6618), .A2(n6617), .ZN(n6682) );
  AOI21_X1 U8374 ( .B1(n6684), .B2(n6619), .A(n6682), .ZN(n6621) );
  OAI21_X1 U8375 ( .B1(n9772), .B2(n9382), .A(n6620), .ZN(n6687) );
  NAND2_X1 U8376 ( .A1(n9511), .A2(n9382), .ZN(n6631) );
  OAI22_X1 U8377 ( .A1(n6621), .A2(n6687), .B1(n9507), .B2(n6631), .ZN(n6622)
         );
  OAI211_X1 U8378 ( .C1(n9772), .C2(n9511), .A(n6622), .B(n6689), .ZN(n6624)
         );
  AOI21_X1 U8379 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(n6626) );
  INV_X2 U8380 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U8381 ( .A1(n7317), .A2(P1_U3086), .ZN(n8307) );
  INV_X1 U8382 ( .A(n8307), .ZN(n7321) );
  OAI21_X1 U8383 ( .B1(n6628), .B2(n6627), .A(n5216), .ZN(n6699) );
  OR3_X1 U8384 ( .A1(n8307), .A2(n6914), .A3(n6635), .ZN(n6636) );
  AOI21_X1 U8385 ( .B1(n6637), .B2(n9610), .A(n6636), .ZN(n6638) );
  NAND2_X1 U8386 ( .A1(n6639), .A2(n6638), .ZN(n6698) );
  INV_X1 U8387 ( .A(n6640), .ZN(n6681) );
  INV_X1 U8388 ( .A(n6641), .ZN(n6670) );
  INV_X1 U8389 ( .A(n6642), .ZN(n6668) );
  OAI211_X1 U8390 ( .C1(n4648), .C2(n5848), .A(n6645), .B(n6644), .ZN(n6647)
         );
  NAND2_X1 U8391 ( .A1(n6647), .A2(n6646), .ZN(n6649) );
  OAI21_X1 U8392 ( .B1(n6643), .B2(n6649), .A(n6648), .ZN(n6652) );
  INV_X1 U8393 ( .A(n6650), .ZN(n6651) );
  AOI21_X1 U8394 ( .B1(n6652), .B2(n7869), .A(n6651), .ZN(n6655) );
  OAI21_X1 U8395 ( .B1(n6655), .B2(n6654), .A(n6653), .ZN(n6660) );
  NAND2_X1 U8396 ( .A1(n6658), .A2(n6657), .ZN(n6659) );
  AOI21_X1 U8397 ( .B1(n6660), .B2(n4670), .A(n6659), .ZN(n6664) );
  INV_X1 U8398 ( .A(n6661), .ZN(n6662) );
  OAI21_X1 U8399 ( .B1(n6664), .B2(n6663), .A(n6662), .ZN(n6665) );
  NAND3_X1 U8400 ( .A1(n9698), .A2(n6666), .A3(n6665), .ZN(n6667) );
  NAND2_X1 U8401 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  NAND2_X1 U8402 ( .A1(n6670), .A2(n6669), .ZN(n6672) );
  NAND3_X1 U8403 ( .A1(n6673), .A2(n6672), .A3(n6671), .ZN(n6676) );
  INV_X1 U8404 ( .A(n6674), .ZN(n6675) );
  AOI21_X1 U8405 ( .B1(n6677), .B2(n6676), .A(n6675), .ZN(n6680) );
  OAI211_X1 U8406 ( .C1(n6681), .C2(n6680), .A(n6679), .B(n6678), .ZN(n6683)
         );
  AOI21_X1 U8407 ( .B1(n6684), .B2(n6683), .A(n6682), .ZN(n6688) );
  OAI211_X1 U8408 ( .C1(n6688), .C2(n6687), .A(n6686), .B(n6685), .ZN(n6690)
         );
  NAND2_X1 U8409 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  XNOR2_X1 U8410 ( .A(n6691), .B(n5846), .ZN(n6692) );
  NAND3_X1 U8411 ( .A1(n6692), .A2(n7321), .A3(n8212), .ZN(n6696) );
  INV_X1 U8412 ( .A(n8320), .ZN(n6693) );
  AND2_X1 U8413 ( .A1(n6693), .A2(n9923), .ZN(n7129) );
  NOR2_X1 U8414 ( .A1(n8317), .A2(n9935), .ZN(n7358) );
  NAND2_X1 U8415 ( .A1(n7129), .A2(n7358), .ZN(n6694) );
  OAI211_X1 U8416 ( .C1(n6914), .C2(n8307), .A(n6694), .B(P1_B_REG_SCAN_IN), 
        .ZN(n6695) );
  NAND2_X1 U8417 ( .A1(n6703), .A2(n6700), .ZN(n6701) );
  OAI21_X1 U8418 ( .B1(n6703), .B2(n6702), .A(n6701), .ZN(n6704) );
  INV_X1 U8419 ( .A(n6706), .ZN(n6707) );
  NAND2_X1 U8420 ( .A1(n6708), .A2(n10128), .ZN(n6716) );
  NAND2_X1 U8421 ( .A1(n6724), .A2(n6857), .ZN(n10120) );
  NAND2_X1 U8422 ( .A1(n7945), .A2(n10120), .ZN(n6709) );
  AOI22_X1 U8423 ( .A1(n7285), .A2(n8925), .B1(n8924), .B2(n7277), .ZN(n6713)
         );
  AND2_X1 U8424 ( .A1(n6713), .A2(n5218), .ZN(n6714) );
  NAND2_X1 U8425 ( .A1(n6716), .A2(n5230), .ZN(P2_U3205) );
  NAND2_X1 U8426 ( .A1(n6213), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6717) );
  INV_X1 U8427 ( .A(n6837), .ZN(n8543) );
  MUX2_X1 U8428 ( .A(n6817), .B(n4449), .S(n4402), .Z(n6719) );
  INV_X1 U8429 ( .A(n6719), .ZN(n6823) );
  NAND3_X1 U8430 ( .A1(n6789), .A2(n7293), .A3(n6720), .ZN(n6722) );
  NAND3_X1 U8431 ( .A1(n6800), .A2(n4402), .A3(n6795), .ZN(n6721) );
  OAI211_X1 U8432 ( .C1(n6789), .C2(n7293), .A(n6722), .B(n6721), .ZN(n6799)
         );
  MUX2_X1 U8433 ( .A(n8987), .B(n6725), .S(n4402), .Z(n6729) );
  XNOR2_X1 U8434 ( .A(n6397), .B(n9004), .ZN(n8992) );
  AND2_X1 U8435 ( .A1(n8987), .A2(n6726), .ZN(n8918) );
  NAND3_X1 U8436 ( .A1(n6727), .A2(n8918), .A3(n6862), .ZN(n6728) );
  NAND2_X1 U8437 ( .A1(n8996), .A2(n10114), .ZN(n6746) );
  NAND2_X1 U8438 ( .A1(n6730), .A2(n6746), .ZN(n6733) );
  NAND2_X1 U8439 ( .A1(n6739), .A2(n6731), .ZN(n6732) );
  MUX2_X1 U8440 ( .A(n6733), .B(n6732), .S(n4402), .Z(n6734) );
  INV_X1 U8441 ( .A(n6734), .ZN(n6736) );
  INV_X1 U8442 ( .A(n7748), .ZN(n6735) );
  INV_X1 U8443 ( .A(n6737), .ZN(n6738) );
  AOI21_X1 U8444 ( .B1(n6747), .B2(n6739), .A(n6738), .ZN(n6741) );
  NAND2_X1 U8445 ( .A1(n6749), .A2(n6740), .ZN(n6744) );
  OAI21_X1 U8446 ( .B1(n6741), .B2(n6744), .A(n6743), .ZN(n6751) );
  NAND2_X1 U8447 ( .A1(n6743), .A2(n6742), .ZN(n6748) );
  NAND2_X1 U8448 ( .A1(n6859), .A2(n6864), .ZN(n6753) );
  NAND2_X1 U8449 ( .A1(n8012), .A2(n6865), .ZN(n6752) );
  NAND2_X1 U8450 ( .A1(n8370), .A2(n8547), .ZN(n6760) );
  OAI211_X1 U8451 ( .C1(n6755), .C2(n6754), .A(n6760), .B(n8012), .ZN(n6759)
         );
  AOI21_X1 U8452 ( .B1(n6864), .B2(n6756), .A(n6755), .ZN(n6758) );
  NAND2_X1 U8453 ( .A1(n6764), .A2(n8146), .ZN(n6762) );
  NAND2_X1 U8454 ( .A1(n6763), .A2(n6760), .ZN(n6761) );
  MUX2_X1 U8455 ( .A(n6762), .B(n6761), .S(n7293), .Z(n6766) );
  MUX2_X1 U8456 ( .A(n6764), .B(n6763), .S(n4402), .Z(n6765) );
  INV_X1 U8457 ( .A(n8901), .ZN(n8909) );
  NAND2_X1 U8458 ( .A1(n8160), .A2(n8478), .ZN(n6768) );
  MUX2_X1 U8459 ( .A(n6768), .B(n6767), .S(n7293), .Z(n6769) );
  NAND3_X1 U8460 ( .A1(n6770), .A2(n8909), .A3(n6769), .ZN(n6774) );
  MUX2_X1 U8461 ( .A(n6772), .B(n6771), .S(n7293), .Z(n6773) );
  NOR2_X1 U8462 ( .A1(n6776), .A2(n7293), .ZN(n6777) );
  AOI211_X1 U8463 ( .C1(n6407), .C2(n7293), .A(n6777), .B(n8871), .ZN(n6778)
         );
  INV_X1 U8464 ( .A(n6785), .ZN(n6781) );
  AOI21_X1 U8465 ( .B1(n6784), .B2(n6779), .A(n7293), .ZN(n6780) );
  AOI211_X1 U8466 ( .C1(n7293), .C2(n6782), .A(n6781), .B(n6780), .ZN(n6783)
         );
  MUX2_X1 U8467 ( .A(n6785), .B(n6784), .S(n7293), .Z(n6787) );
  OAI21_X1 U8468 ( .B1(n8861), .B2(n9077), .A(n8820), .ZN(n6786) );
  NAND3_X1 U8469 ( .A1(n6792), .A2(n6791), .A3(n6790), .ZN(n6794) );
  NAND2_X1 U8470 ( .A1(n6794), .A2(n6793), .ZN(n6797) );
  INV_X1 U8471 ( .A(n8785), .ZN(n8787) );
  NAND2_X1 U8472 ( .A1(n6803), .A2(n6802), .ZN(n6808) );
  AND2_X1 U8473 ( .A1(n8771), .A2(n6804), .ZN(n6806) );
  INV_X1 U8474 ( .A(n6810), .ZN(n6811) );
  MUX2_X1 U8475 ( .A(n6814), .B(n4831), .S(n4402), .Z(n6815) );
  INV_X1 U8476 ( .A(n6820), .ZN(n6816) );
  INV_X1 U8477 ( .A(n6818), .ZN(n6819) );
  MUX2_X1 U8478 ( .A(n6820), .B(n6819), .S(n4402), .Z(n6821) );
  NAND2_X1 U8479 ( .A1(n8339), .A2(n6844), .ZN(n6826) );
  NAND2_X1 U8480 ( .A1(n6213), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6825) );
  INV_X1 U8481 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10400) );
  NAND2_X1 U8482 ( .A1(n6827), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U8483 ( .A1(n4399), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6828) );
  OAI211_X1 U8484 ( .C1(n6830), .C2(n10400), .A(n6829), .B(n6828), .ZN(n6831)
         );
  INV_X1 U8485 ( .A(n6831), .ZN(n6832) );
  NAND2_X1 U8486 ( .A1(n6852), .A2(n6832), .ZN(n8542) );
  INV_X1 U8487 ( .A(n8542), .ZN(n6833) );
  NAND2_X1 U8488 ( .A1(n6890), .A2(n6833), .ZN(n6835) );
  NAND2_X1 U8489 ( .A1(n6838), .A2(n6837), .ZN(n7140) );
  NAND2_X1 U8490 ( .A1(n6835), .A2(n7140), .ZN(n6889) );
  AOI211_X1 U8491 ( .C1(n7148), .C2(n6842), .A(n6889), .B(n6840), .ZN(n6855)
         );
  NAND2_X1 U8492 ( .A1(n6835), .A2(n7293), .ZN(n6836) );
  NAND2_X1 U8493 ( .A1(n6839), .A2(n6836), .ZN(n6854) );
  NAND3_X1 U8494 ( .A1(n6839), .A2(n7293), .A3(n7141), .ZN(n6841) );
  AOI211_X1 U8495 ( .C1(n7147), .C2(n6842), .A(n6841), .B(n6840), .ZN(n6843)
         );
  INV_X1 U8496 ( .A(n6843), .ZN(n6853) );
  NAND2_X1 U8497 ( .A1(n9109), .A2(n6844), .ZN(n6846) );
  NAND2_X1 U8498 ( .A1(n6014), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U8499 ( .A1(n6847), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U8500 ( .A1(n4399), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U8501 ( .A1(n6827), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6848) );
  AND3_X1 U8502 ( .A1(n6850), .A2(n6849), .A3(n6848), .ZN(n6851) );
  OAI211_X1 U8503 ( .C1(n6855), .C2(n6854), .A(n6853), .B(n4450), .ZN(n6858)
         );
  NAND2_X1 U8504 ( .A1(n6894), .A2(n6891), .ZN(n6901) );
  NAND3_X1 U8505 ( .A1(n6858), .A2(n6857), .A3(n6901), .ZN(n6907) );
  INV_X1 U8506 ( .A(n8800), .ZN(n8798) );
  INV_X1 U8507 ( .A(n6859), .ZN(n6860) );
  INV_X1 U8508 ( .A(n6862), .ZN(n6863) );
  NOR2_X1 U8509 ( .A1(n8914), .A2(n6863), .ZN(n10131) );
  AND4_X1 U8510 ( .A1(n10131), .A2(n8918), .A3(n10112), .A4(n8992), .ZN(n6870)
         );
  AND2_X1 U8511 ( .A1(n6865), .A2(n6864), .ZN(n7883) );
  INV_X1 U8512 ( .A(n7742), .ZN(n6866) );
  AND2_X1 U8513 ( .A1(n6866), .A2(n7824), .ZN(n6869) );
  NAND2_X1 U8514 ( .A1(n6868), .A2(n6867), .ZN(n7750) );
  NAND4_X1 U8515 ( .A1(n6870), .A2(n7883), .A3(n6869), .A4(n7750), .ZN(n6871)
         );
  INV_X1 U8516 ( .A(n7729), .ZN(n7724) );
  NOR3_X1 U8517 ( .A1(n7940), .A2(n6871), .A3(n7724), .ZN(n6872) );
  XNOR2_X1 U8518 ( .A(n8983), .B(n8547), .ZN(n8014) );
  NAND3_X1 U8519 ( .A1(n8148), .A2(n6872), .A3(n8014), .ZN(n6873) );
  NOR2_X1 U8520 ( .A1(n8163), .A2(n6873), .ZN(n6874) );
  NAND3_X1 U8521 ( .A1(n6198), .A2(n8909), .A3(n6874), .ZN(n6875) );
  NAND3_X1 U8522 ( .A1(n8810), .A2(n8823), .A3(n6877), .ZN(n6878) );
  NOR2_X1 U8523 ( .A1(n8785), .A2(n6878), .ZN(n6879) );
  AND4_X1 U8524 ( .A1(n4480), .A2(n6880), .A3(n8798), .A4(n6879), .ZN(n6881)
         );
  AND2_X1 U8525 ( .A1(n8738), .A2(n6882), .ZN(n6885) );
  INV_X1 U8526 ( .A(n6883), .ZN(n6884) );
  NAND4_X1 U8527 ( .A1(n6902), .A2(n7162), .A3(n7164), .A4(n6901), .ZN(n6900)
         );
  NOR2_X1 U8528 ( .A1(n7147), .A2(n8730), .ZN(n6887) );
  INV_X1 U8529 ( .A(n7141), .ZN(n6893) );
  INV_X1 U8530 ( .A(n6891), .ZN(n8720) );
  OAI21_X1 U8531 ( .B1(n6890), .B2(n8720), .A(n9015), .ZN(n6892) );
  OAI211_X1 U8532 ( .C1(n7142), .C2(n6893), .A(n6886), .B(n6892), .ZN(n6898)
         );
  NAND2_X1 U8533 ( .A1(n6895), .A2(n6894), .ZN(n6897) );
  AOI21_X1 U8534 ( .B1(n6898), .B2(n6897), .A(n6896), .ZN(n6899) );
  MUX2_X1 U8535 ( .A(n6900), .B(n7164), .S(n6899), .Z(n6906) );
  INV_X1 U8536 ( .A(n6901), .ZN(n6904) );
  OR2_X1 U8537 ( .A1(n7399), .A2(P2_U3151), .ZN(n8291) );
  NOR3_X1 U8538 ( .A1(n6902), .A2(n7164), .A3(n8215), .ZN(n6903) );
  AOI211_X1 U8539 ( .C1(n6904), .C2(n8704), .A(n8291), .B(n6903), .ZN(n6905)
         );
  INV_X1 U8540 ( .A(n6909), .ZN(n7260) );
  NAND2_X1 U8541 ( .A1(n7333), .A2(n7260), .ZN(n7273) );
  INV_X1 U8542 ( .A(n4387), .ZN(n8694) );
  NOR3_X1 U8543 ( .A1(n7273), .A2(n8694), .A3(n6342), .ZN(n6912) );
  OAI21_X1 U8544 ( .B1(n8291), .B2(n6910), .A(P2_B_REG_SCAN_IN), .ZN(n6911) );
  OR2_X1 U8545 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  NAND2_X2 U8546 ( .A1(n7291), .A2(n6915), .ZN(n9176) );
  INV_X1 U8547 ( .A(n6915), .ZN(n6916) );
  OAI22_X1 U8548 ( .A1(n4648), .A2(n9183), .B1(n7692), .B2(n9176), .ZN(n6918)
         );
  INV_X1 U8549 ( .A(n7291), .ZN(n6923) );
  NAND2_X1 U8550 ( .A1(n6923), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U8551 ( .A1(n6578), .A2(n6941), .ZN(n6922) );
  NAND2_X1 U8552 ( .A1(n6578), .A2(n7092), .ZN(n6925) );
  AOI22_X1 U8553 ( .A1(n8325), .A2(n6941), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6923), .ZN(n6924) );
  NAND2_X1 U8554 ( .A1(n6925), .A2(n6924), .ZN(n7507) );
  AND2_X1 U8555 ( .A1(n6926), .A2(n9179), .ZN(n6927) );
  XNOR2_X1 U8556 ( .A(n6928), .B(n7040), .ZN(n6931) );
  OAI22_X1 U8557 ( .A1(n9212), .A2(n4647), .B1(n6929), .B2(n9176), .ZN(n6930)
         );
  NAND2_X1 U8558 ( .A1(n6931), .A2(n6930), .ZN(n6932) );
  OAI22_X1 U8559 ( .A1(n10011), .A2(n9176), .B1(n10006), .B2(n6965), .ZN(n6933) );
  XNOR2_X1 U8560 ( .A(n6933), .B(n7040), .ZN(n6940) );
  OAI22_X1 U8561 ( .A1(n10011), .A2(n4647), .B1(n10006), .B2(n9176), .ZN(n6939) );
  XNOR2_X1 U8562 ( .A(n6940), .B(n6939), .ZN(n7889) );
  OAI22_X1 U8563 ( .A1(n6936), .A2(n9176), .B1(n10021), .B2(n6965), .ZN(n6935)
         );
  XNOR2_X1 U8564 ( .A(n6935), .B(n7040), .ZN(n8073) );
  OR2_X1 U8565 ( .A1(n6936), .A2(n4647), .ZN(n6938) );
  NAND2_X1 U8566 ( .A1(n4394), .A2(n9181), .ZN(n6937) );
  NAND2_X1 U8567 ( .A1(n6938), .A2(n6937), .ZN(n8072) );
  OR2_X1 U8568 ( .A1(n6940), .A2(n6939), .ZN(n8068) );
  NAND2_X1 U8569 ( .A1(n9389), .A2(n9181), .ZN(n6943) );
  NAND2_X1 U8570 ( .A1(n10013), .A2(n9175), .ZN(n6942) );
  NAND2_X1 U8571 ( .A1(n6943), .A2(n6942), .ZN(n6944) );
  NAND2_X1 U8572 ( .A1(n9389), .A2(n7092), .ZN(n6946) );
  NAND2_X1 U8573 ( .A1(n10013), .A2(n9181), .ZN(n6945) );
  AND2_X1 U8574 ( .A1(n6946), .A2(n6945), .ZN(n8069) );
  NAND2_X1 U8575 ( .A1(n8070), .A2(n8069), .ZN(n6947) );
  OAI211_X1 U8576 ( .C1(n8073), .C2(n8072), .A(n8068), .B(n6947), .ZN(n6953)
         );
  NOR2_X1 U8577 ( .A1(n8070), .A2(n8069), .ZN(n8071) );
  OAI21_X1 U8578 ( .B1(n8071), .B2(n8072), .A(n8073), .ZN(n6951) );
  INV_X1 U8579 ( .A(n8070), .ZN(n6949) );
  INV_X1 U8580 ( .A(n8069), .ZN(n6948) );
  NAND3_X1 U8581 ( .A1(n6949), .A2(n8072), .A3(n6948), .ZN(n6950) );
  NAND2_X1 U8582 ( .A1(n9388), .A2(n9181), .ZN(n6954) );
  OAI21_X1 U8583 ( .B1(n10027), .B2(n6965), .A(n6954), .ZN(n6955) );
  XNOR2_X1 U8584 ( .A(n6955), .B(n7040), .ZN(n6960) );
  OR2_X1 U8585 ( .A1(n10027), .A2(n9176), .ZN(n6957) );
  NAND2_X1 U8586 ( .A1(n9388), .A2(n7092), .ZN(n6956) );
  NAND2_X1 U8587 ( .A1(n6957), .A2(n6956), .ZN(n6959) );
  NOR2_X1 U8588 ( .A1(n6960), .A2(n6959), .ZN(n7960) );
  INV_X1 U8589 ( .A(n7960), .ZN(n6958) );
  NAND2_X1 U8590 ( .A1(n6960), .A2(n6959), .ZN(n7959) );
  OAI22_X1 U8591 ( .A1(n10040), .A2(n4647), .B1(n10033), .B2(n9176), .ZN(n6963) );
  AOI22_X1 U8592 ( .A1(n9387), .A2(n9181), .B1(n8113), .B2(n9175), .ZN(n6962)
         );
  XOR2_X1 U8593 ( .A(n7040), .B(n6962), .Z(n8106) );
  NAND2_X1 U8594 ( .A1(n10052), .A2(n9181), .ZN(n6964) );
  OAI21_X1 U8595 ( .B1(n9204), .B2(n6965), .A(n6964), .ZN(n6966) );
  XNOR2_X1 U8596 ( .A(n6966), .B(n7040), .ZN(n9195) );
  OR2_X1 U8597 ( .A1(n9204), .A2(n9176), .ZN(n6968) );
  NAND2_X1 U8598 ( .A1(n10052), .A2(n7092), .ZN(n6967) );
  NAND2_X1 U8599 ( .A1(n6968), .A2(n6967), .ZN(n6974) );
  NAND2_X1 U8600 ( .A1(n10054), .A2(n9175), .ZN(n6970) );
  OR2_X1 U8601 ( .A1(n10039), .A2(n9176), .ZN(n6969) );
  NAND2_X1 U8602 ( .A1(n6970), .A2(n6969), .ZN(n6971) );
  XNOR2_X1 U8603 ( .A(n6971), .B(n9179), .ZN(n6978) );
  NAND2_X1 U8604 ( .A1(n10054), .A2(n9181), .ZN(n6973) );
  OR2_X1 U8605 ( .A1(n10039), .A2(n4647), .ZN(n6972) );
  NAND2_X1 U8606 ( .A1(n6973), .A2(n6972), .ZN(n6979) );
  XNOR2_X1 U8607 ( .A(n6978), .B(n6979), .ZN(n9286) );
  INV_X1 U8608 ( .A(n6974), .ZN(n9198) );
  AND2_X1 U8609 ( .A1(n9286), .A2(n6975), .ZN(n6976) );
  NAND2_X1 U8610 ( .A1(n10062), .A2(n9175), .ZN(n6983) );
  OR2_X1 U8611 ( .A1(n9331), .A2(n9176), .ZN(n6982) );
  NAND2_X1 U8612 ( .A1(n6983), .A2(n6982), .ZN(n6984) );
  XNOR2_X1 U8613 ( .A(n6984), .B(n7040), .ZN(n9153) );
  NAND2_X1 U8614 ( .A1(n10062), .A2(n9181), .ZN(n6986) );
  OR2_X1 U8615 ( .A1(n9331), .A2(n4647), .ZN(n6985) );
  NAND2_X1 U8616 ( .A1(n6986), .A2(n6985), .ZN(n9157) );
  NOR2_X1 U8617 ( .A1(n9153), .A2(n9157), .ZN(n6992) );
  NAND2_X1 U8618 ( .A1(n9333), .A2(n9175), .ZN(n6988) );
  OR2_X1 U8619 ( .A1(n10083), .A2(n9176), .ZN(n6987) );
  NAND2_X1 U8620 ( .A1(n6988), .A2(n6987), .ZN(n6989) );
  XNOR2_X1 U8621 ( .A(n6989), .B(n9179), .ZN(n6994) );
  NOR2_X1 U8622 ( .A1(n10083), .A2(n4647), .ZN(n6990) );
  AOI21_X1 U8623 ( .B1(n9333), .B2(n9181), .A(n6990), .ZN(n6993) );
  NOR2_X1 U8624 ( .A1(n6994), .A2(n6993), .ZN(n9326) );
  AOI21_X1 U8625 ( .B1(n9153), .B2(n9157), .A(n9326), .ZN(n6991) );
  AOI22_X1 U8626 ( .A1(n10079), .A2(n9175), .B1(n9181), .B2(n9985), .ZN(n6995)
         );
  XNOR2_X1 U8627 ( .A(n6995), .B(n7040), .ZN(n6996) );
  OAI22_X1 U8628 ( .A1(n8282), .A2(n9176), .B1(n9757), .B2(n4647), .ZN(n6997)
         );
  XNOR2_X1 U8629 ( .A(n6996), .B(n6997), .ZN(n9224) );
  INV_X1 U8630 ( .A(n6997), .ZN(n6998) );
  NAND2_X1 U8631 ( .A1(n9902), .A2(n9175), .ZN(n7000) );
  OR2_X1 U8632 ( .A1(n9139), .A2(n9176), .ZN(n6999) );
  NAND2_X1 U8633 ( .A1(n7000), .A2(n6999), .ZN(n7001) );
  XNOR2_X1 U8634 ( .A(n7001), .B(n7040), .ZN(n7002) );
  OAI22_X1 U8635 ( .A1(n5073), .A2(n9176), .B1(n9139), .B2(n4647), .ZN(n7003)
         );
  XOR2_X1 U8636 ( .A(n7002), .B(n7003), .Z(n9306) );
  INV_X1 U8637 ( .A(n7002), .ZN(n7005) );
  INV_X1 U8638 ( .A(n7003), .ZN(n7004) );
  NAND2_X1 U8639 ( .A1(n9746), .A2(n9175), .ZN(n7007) );
  NAND2_X1 U8640 ( .A1(n9882), .A2(n9181), .ZN(n7006) );
  NAND2_X1 U8641 ( .A1(n7007), .A2(n7006), .ZN(n7008) );
  XNOR2_X1 U8642 ( .A(n7008), .B(n9179), .ZN(n9135) );
  AOI22_X1 U8643 ( .A1(n9746), .A2(n9181), .B1(n7092), .B2(n9882), .ZN(n9137)
         );
  NAND2_X1 U8644 ( .A1(n9877), .A2(n9175), .ZN(n7010) );
  NAND2_X1 U8645 ( .A1(n9883), .A2(n9181), .ZN(n7009) );
  NAND2_X1 U8646 ( .A1(n7010), .A2(n7009), .ZN(n7011) );
  XNOR2_X1 U8647 ( .A(n7011), .B(n7040), .ZN(n9247) );
  NAND2_X1 U8648 ( .A1(n9877), .A2(n9181), .ZN(n7013) );
  NAND2_X1 U8649 ( .A1(n9883), .A2(n7092), .ZN(n7012) );
  NAND2_X1 U8650 ( .A1(n7013), .A2(n7012), .ZN(n7022) );
  NAND2_X1 U8651 ( .A1(n5860), .A2(n9175), .ZN(n7015) );
  NAND2_X1 U8652 ( .A1(n9891), .A2(n9181), .ZN(n7014) );
  NAND2_X1 U8653 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  XNOR2_X1 U8654 ( .A(n7016), .B(n7040), .ZN(n9243) );
  NAND2_X1 U8655 ( .A1(n5860), .A2(n9181), .ZN(n7018) );
  NAND2_X1 U8656 ( .A1(n9891), .A2(n7092), .ZN(n7017) );
  NAND2_X1 U8657 ( .A1(n7018), .A2(n7017), .ZN(n9370) );
  OAI22_X1 U8658 ( .A1(n9247), .A2(n7022), .B1(n9243), .B2(n9370), .ZN(n7019)
         );
  AOI21_X1 U8659 ( .B1(n9135), .B2(n9137), .A(n7019), .ZN(n7028) );
  INV_X1 U8660 ( .A(n7022), .ZN(n9246) );
  AND2_X1 U8661 ( .A1(n9243), .A2(n9370), .ZN(n7023) );
  INV_X1 U8662 ( .A(n7023), .ZN(n7026) );
  INV_X1 U8663 ( .A(n7019), .ZN(n7021) );
  INV_X1 U8664 ( .A(n9135), .ZN(n9241) );
  INV_X1 U8665 ( .A(n9137), .ZN(n7020) );
  NAND3_X1 U8666 ( .A1(n7021), .A2(n9241), .A3(n7020), .ZN(n7025) );
  OAI21_X1 U8667 ( .B1(n7023), .B2(n7022), .A(n9247), .ZN(n7024) );
  OAI211_X1 U8668 ( .C1(n9246), .C2(n7026), .A(n7025), .B(n7024), .ZN(n7027)
         );
  NAND2_X1 U8669 ( .A1(n9869), .A2(n9175), .ZN(n7030) );
  NAND2_X1 U8670 ( .A1(n9675), .A2(n9181), .ZN(n7029) );
  NAND2_X1 U8671 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  XNOR2_X1 U8672 ( .A(n7031), .B(n9179), .ZN(n7034) );
  INV_X1 U8673 ( .A(n7034), .ZN(n7036) );
  NOR2_X1 U8674 ( .A1(n9874), .A2(n4647), .ZN(n7032) );
  AOI21_X1 U8675 ( .B1(n9869), .B2(n9181), .A(n7032), .ZN(n7033) );
  INV_X1 U8676 ( .A(n7033), .ZN(n7035) );
  AND2_X1 U8677 ( .A1(n7034), .A2(n7033), .ZN(n7037) );
  AOI21_X1 U8678 ( .B1(n7036), .B2(n7035), .A(n7037), .ZN(n9256) );
  NAND2_X1 U8679 ( .A1(n9255), .A2(n9256), .ZN(n9254) );
  INV_X1 U8680 ( .A(n7037), .ZN(n7038) );
  AOI22_X1 U8681 ( .A1(n9863), .A2(n9175), .B1(n9181), .B2(n9850), .ZN(n7039)
         );
  XOR2_X1 U8682 ( .A(n7040), .B(n7039), .Z(n9165) );
  NAND2_X1 U8683 ( .A1(n9863), .A2(n9181), .ZN(n7042) );
  NAND2_X1 U8684 ( .A1(n9850), .A2(n7092), .ZN(n7041) );
  NAND2_X1 U8685 ( .A1(n7042), .A2(n7041), .ZN(n9348) );
  NOR2_X1 U8686 ( .A1(n9165), .A2(n9348), .ZN(n7049) );
  NAND2_X1 U8687 ( .A1(n9657), .A2(n9175), .ZN(n7044) );
  NAND2_X1 U8688 ( .A1(n9638), .A2(n9181), .ZN(n7043) );
  NAND2_X1 U8689 ( .A1(n7044), .A2(n7043), .ZN(n7045) );
  XNOR2_X1 U8690 ( .A(n7045), .B(n7040), .ZN(n7050) );
  AND2_X1 U8691 ( .A1(n9638), .A2(n7092), .ZN(n7046) );
  AOI21_X1 U8692 ( .B1(n9657), .B2(n9181), .A(n7046), .ZN(n7051) );
  XNOR2_X1 U8693 ( .A(n7050), .B(n7051), .ZN(n9169) );
  NAND2_X1 U8694 ( .A1(n9165), .A2(n9348), .ZN(n7047) );
  INV_X1 U8695 ( .A(n7050), .ZN(n7052) );
  NAND2_X1 U8696 ( .A1(n7052), .A2(n7051), .ZN(n7053) );
  NAND2_X1 U8697 ( .A1(n9845), .A2(n9175), .ZN(n7055) );
  NAND2_X1 U8698 ( .A1(n9851), .A2(n9181), .ZN(n7054) );
  NAND2_X1 U8699 ( .A1(n7055), .A2(n7054), .ZN(n7056) );
  XNOR2_X1 U8700 ( .A(n7056), .B(n7040), .ZN(n7062) );
  INV_X1 U8701 ( .A(n7062), .ZN(n7060) );
  NAND2_X1 U8702 ( .A1(n9845), .A2(n9181), .ZN(n7058) );
  NAND2_X1 U8703 ( .A1(n9851), .A2(n7092), .ZN(n7057) );
  NAND2_X1 U8704 ( .A1(n7058), .A2(n7057), .ZN(n7061) );
  INV_X1 U8705 ( .A(n7061), .ZN(n7059) );
  AND2_X1 U8706 ( .A1(n7062), .A2(n7061), .ZN(n9299) );
  NAND2_X1 U8707 ( .A1(n9837), .A2(n9175), .ZN(n7064) );
  NAND2_X1 U8708 ( .A1(n9824), .A2(n9181), .ZN(n7063) );
  NAND2_X1 U8709 ( .A1(n7064), .A2(n7063), .ZN(n7065) );
  XNOR2_X1 U8710 ( .A(n7065), .B(n7040), .ZN(n7066) );
  AOI22_X1 U8711 ( .A1(n9837), .A2(n9181), .B1(n7092), .B2(n9824), .ZN(n7067)
         );
  XNOR2_X1 U8712 ( .A(n7066), .B(n7067), .ZN(n9218) );
  INV_X1 U8713 ( .A(n7066), .ZN(n7068) );
  NAND2_X1 U8714 ( .A1(n7068), .A2(n7067), .ZN(n7069) );
  NAND2_X1 U8715 ( .A1(n9216), .A2(n7069), .ZN(n7074) );
  INV_X1 U8716 ( .A(n7074), .ZN(n7072) );
  AOI22_X1 U8717 ( .A1(n9320), .A2(n9175), .B1(n9181), .B2(n9815), .ZN(n7070)
         );
  XNOR2_X1 U8718 ( .A(n7070), .B(n7040), .ZN(n7073) );
  INV_X1 U8719 ( .A(n7073), .ZN(n7071) );
  NAND2_X1 U8720 ( .A1(n7072), .A2(n7071), .ZN(n9314) );
  AOI22_X1 U8721 ( .A1(n9320), .A2(n9181), .B1(n7092), .B2(n9815), .ZN(n9315)
         );
  NAND2_X1 U8722 ( .A1(n9314), .A2(n9315), .ZN(n7075) );
  NAND2_X1 U8723 ( .A1(n7074), .A2(n7073), .ZN(n9313) );
  AOI22_X1 U8724 ( .A1(n9600), .A2(n9175), .B1(n9181), .B2(n9825), .ZN(n7076)
         );
  XOR2_X1 U8725 ( .A(n7040), .B(n7076), .Z(n7077) );
  OAI22_X1 U8726 ( .A1(n9819), .A2(n9176), .B1(n9613), .B2(n4647), .ZN(n7078)
         );
  NAND2_X1 U8727 ( .A1(n7077), .A2(n7078), .ZN(n9145) );
  INV_X1 U8728 ( .A(n7077), .ZN(n7080) );
  INV_X1 U8729 ( .A(n7078), .ZN(n7079) );
  NAND2_X1 U8730 ( .A1(n7080), .A2(n7079), .ZN(n9144) );
  NAND2_X1 U8731 ( .A1(n9812), .A2(n9175), .ZN(n7082) );
  NAND2_X1 U8732 ( .A1(n9816), .A2(n9181), .ZN(n7081) );
  NAND2_X1 U8733 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  XNOR2_X1 U8734 ( .A(n7083), .B(n7040), .ZN(n7087) );
  NAND2_X1 U8735 ( .A1(n9812), .A2(n9181), .ZN(n7085) );
  NAND2_X1 U8736 ( .A1(n9816), .A2(n7092), .ZN(n7084) );
  NAND2_X1 U8737 ( .A1(n7085), .A2(n7084), .ZN(n7086) );
  NOR2_X1 U8738 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  AOI21_X1 U8739 ( .B1(n7087), .B2(n7086), .A(n7088), .ZN(n9269) );
  NAND2_X1 U8740 ( .A1(n9808), .A2(n9175), .ZN(n7090) );
  NAND2_X1 U8741 ( .A1(n9577), .A2(n9181), .ZN(n7089) );
  NAND2_X1 U8742 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  XNOR2_X1 U8743 ( .A(n7091), .B(n7040), .ZN(n7099) );
  AOI22_X1 U8744 ( .A1(n9808), .A2(n9181), .B1(n7092), .B2(n9577), .ZN(n7097)
         );
  XNOR2_X1 U8745 ( .A(n7099), .B(n7097), .ZN(n9234) );
  NOR2_X1 U8746 ( .A1(n9562), .A2(n4647), .ZN(n7093) );
  AOI21_X1 U8747 ( .B1(n9801), .B2(n9181), .A(n7093), .ZN(n7101) );
  NAND2_X1 U8748 ( .A1(n9801), .A2(n9175), .ZN(n7095) );
  NAND2_X1 U8749 ( .A1(n9788), .A2(n9181), .ZN(n7094) );
  NAND2_X1 U8750 ( .A1(n7095), .A2(n7094), .ZN(n7096) );
  XNOR2_X1 U8751 ( .A(n7096), .B(n7040), .ZN(n7103) );
  XOR2_X1 U8752 ( .A(n7101), .B(n7103), .Z(n9355) );
  INV_X1 U8753 ( .A(n7097), .ZN(n7098) );
  NOR2_X1 U8754 ( .A1(n7099), .A2(n7098), .ZN(n9356) );
  NOR2_X1 U8755 ( .A1(n9355), .A2(n9356), .ZN(n7100) );
  INV_X1 U8756 ( .A(n7101), .ZN(n7102) );
  NAND2_X1 U8757 ( .A1(n9540), .A2(n9175), .ZN(n7105) );
  NAND2_X1 U8758 ( .A1(n9384), .A2(n9181), .ZN(n7104) );
  NAND2_X1 U8759 ( .A1(n7105), .A2(n7104), .ZN(n7106) );
  XNOR2_X1 U8760 ( .A(n7106), .B(n9179), .ZN(n7109) );
  INV_X1 U8761 ( .A(n7109), .ZN(n7111) );
  NOR2_X1 U8762 ( .A1(n9798), .A2(n4647), .ZN(n7107) );
  AOI21_X1 U8763 ( .B1(n9540), .B2(n9181), .A(n7107), .ZN(n7108) );
  INV_X1 U8764 ( .A(n7108), .ZN(n7110) );
  AOI21_X1 U8765 ( .B1(n7111), .B2(n7110), .A(n9192), .ZN(n7112) );
  INV_X1 U8766 ( .A(n7112), .ZN(n7113) );
  NOR2_X1 U8767 ( .A1(n7113), .A2(n4436), .ZN(n7114) );
  NOR2_X1 U8768 ( .A1(n7116), .A2(n7115), .ZN(n7126) );
  AND2_X1 U8769 ( .A1(n10071), .A2(n7117), .ZN(n7127) );
  INV_X1 U8770 ( .A(n7122), .ZN(n7125) );
  INV_X1 U8771 ( .A(n7128), .ZN(n7118) );
  OR2_X1 U8772 ( .A1(n7125), .A2(n7118), .ZN(n7119) );
  INV_X1 U8773 ( .A(n7120), .ZN(n7123) );
  AND2_X1 U8774 ( .A1(n7123), .A2(n9986), .ZN(n7121) );
  NAND2_X1 U8775 ( .A1(n7123), .A2(n10053), .ZN(n7124) );
  NOR2_X1 U8776 ( .A1(n9562), .A2(n9349), .ZN(n7136) );
  INV_X1 U8777 ( .A(n7126), .ZN(n7131) );
  OR3_X1 U8778 ( .A1(n7129), .A2(n7128), .A3(n7127), .ZN(n7130) );
  NAND2_X1 U8779 ( .A1(n7131), .A2(n7130), .ZN(n7134) );
  AND3_X1 U8780 ( .A1(n7132), .A2(n7317), .A3(n7291), .ZN(n7133) );
  NAND2_X1 U8781 ( .A1(n7134), .A2(n7133), .ZN(n7509) );
  NAND2_X1 U8782 ( .A1(n7509), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9350) );
  OAI22_X1 U8783 ( .A1(n9536), .A2(n9350), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10201), .ZN(n7135) );
  AOI211_X1 U8784 ( .C1(n9789), .C2(n9365), .A(n7136), .B(n7135), .ZN(n7137)
         );
  OAI21_X1 U8785 ( .B1(n9792), .B2(n9368), .A(n7137), .ZN(n7138) );
  INV_X1 U8786 ( .A(n7138), .ZN(n7139) );
  NAND2_X1 U8787 ( .A1(n8333), .A2(n8990), .ZN(n7156) );
  NAND2_X1 U8788 ( .A1(n7144), .A2(n7143), .ZN(n7153) );
  INV_X1 U8789 ( .A(n7151), .ZN(n7145) );
  NAND2_X1 U8790 ( .A1(n7285), .A2(n8730), .ZN(n7146) );
  NOR2_X1 U8791 ( .A1(n7148), .A2(n8998), .ZN(n7150) );
  AOI21_X1 U8792 ( .B1(P2_B_REG_SCAN_IN), .B2(n7392), .A(n8888), .ZN(n8719) );
  AND2_X1 U8793 ( .A1(n8542), .A2(n8719), .ZN(n7149) );
  NAND2_X1 U8794 ( .A1(n8333), .A2(n9008), .ZN(n7157) );
  NOR2_X1 U8795 ( .A1(n8336), .A2(n8971), .ZN(n7158) );
  INV_X1 U8796 ( .A(n7158), .ZN(n7159) );
  OR2_X1 U8797 ( .A1(n10157), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7160) );
  NAND2_X1 U8798 ( .A1(n7161), .A2(n5221), .ZN(P2_U3456) );
  NAND4_X1 U8799 ( .A1(n7163), .A2(n7162), .A3(n8266), .A4(n7334), .ZN(n7167)
         );
  NAND2_X1 U8800 ( .A1(n7165), .A2(n8215), .ZN(n7166) );
  INV_X1 U8801 ( .A(n7484), .ZN(n7168) );
  XNOR2_X1 U8802 ( .A(n7171), .B(n7530), .ZN(n7472) );
  INV_X1 U8803 ( .A(n7171), .ZN(n7172) );
  NAND2_X1 U8804 ( .A1(n7172), .A2(n7530), .ZN(n7173) );
  XNOR2_X1 U8805 ( .A(n7175), .B(n7468), .ZN(n7535) );
  NAND2_X1 U8806 ( .A1(n7175), .A2(n8996), .ZN(n7176) );
  NAND2_X1 U8807 ( .A1(n7534), .A2(n7176), .ZN(n8455) );
  INV_X1 U8808 ( .A(n8455), .ZN(n7179) );
  XNOR2_X1 U8809 ( .A(n7249), .B(n8458), .ZN(n7177) );
  NAND2_X1 U8810 ( .A1(n7177), .A2(n7531), .ZN(n7766) );
  OAI21_X1 U8811 ( .B1(n7177), .B2(n7531), .A(n7766), .ZN(n8454) );
  NAND2_X1 U8812 ( .A1(n7179), .A2(n7178), .ZN(n7765) );
  NAND2_X1 U8813 ( .A1(n7181), .A2(n7838), .ZN(n7182) );
  INV_X2 U8814 ( .A(n7174), .ZN(n7242) );
  XNOR2_X1 U8815 ( .A(n7183), .B(n8551), .ZN(n7835) );
  INV_X1 U8816 ( .A(n7183), .ZN(n7184) );
  XNOR2_X1 U8817 ( .A(n7906), .B(n7174), .ZN(n7185) );
  NAND2_X1 U8818 ( .A1(n7185), .A2(n7886), .ZN(n8384) );
  INV_X1 U8819 ( .A(n7185), .ZN(n7186) );
  NAND2_X1 U8820 ( .A1(n7186), .A2(n8550), .ZN(n7187) );
  NAND2_X1 U8821 ( .A1(n8384), .A2(n7187), .ZN(n7969) );
  INV_X1 U8822 ( .A(n7969), .ZN(n7188) );
  XNOR2_X1 U8823 ( .A(n8391), .B(n7242), .ZN(n7190) );
  XNOR2_X1 U8824 ( .A(n7190), .B(n8549), .ZN(n8385) );
  NAND2_X1 U8825 ( .A1(n7190), .A2(n8221), .ZN(n7191) );
  XNOR2_X1 U8826 ( .A(n8044), .B(n7242), .ZN(n7192) );
  XNOR2_X1 U8827 ( .A(n7192), .B(n8548), .ZN(n8217) );
  INV_X1 U8828 ( .A(n7192), .ZN(n7193) );
  XNOR2_X1 U8829 ( .A(n8148), .B(n7174), .ZN(n8496) );
  INV_X1 U8830 ( .A(n8496), .ZN(n7195) );
  XNOR2_X1 U8831 ( .A(n8370), .B(n7242), .ZN(n8366) );
  NAND2_X1 U8832 ( .A1(n7195), .A2(n7194), .ZN(n7202) );
  NOR3_X1 U8833 ( .A1(n8370), .A2(n7174), .A3(n8547), .ZN(n7196) );
  INV_X1 U8834 ( .A(n8148), .ZN(n8150) );
  AOI211_X1 U8835 ( .C1(n8412), .C2(n7174), .A(n7196), .B(n8150), .ZN(n7199)
         );
  NOR3_X1 U8836 ( .A1(n8983), .A2(n8547), .A3(n7242), .ZN(n7197) );
  AOI211_X1 U8837 ( .C1(n8412), .C2(n7242), .A(n7197), .B(n8148), .ZN(n7198)
         );
  XNOR2_X1 U8838 ( .A(n8160), .B(n7242), .ZN(n7203) );
  NAND2_X1 U8839 ( .A1(n7203), .A2(n8478), .ZN(n8406) );
  OAI21_X1 U8840 ( .B1(n7199), .B2(n7198), .A(n8406), .ZN(n7200) );
  INV_X1 U8841 ( .A(n7203), .ZN(n7204) );
  NAND2_X1 U8842 ( .A1(n7204), .A2(n8904), .ZN(n8407) );
  NAND2_X1 U8843 ( .A1(n7205), .A2(n8407), .ZN(n8476) );
  XNOR2_X1 U8844 ( .A(n8900), .B(n7242), .ZN(n8474) );
  NAND2_X1 U8845 ( .A1(n8474), .A2(n8887), .ZN(n7207) );
  INV_X1 U8846 ( .A(n8474), .ZN(n7206) );
  XNOR2_X1 U8847 ( .A(n9093), .B(n7242), .ZN(n7208) );
  XNOR2_X1 U8848 ( .A(n7208), .B(n8903), .ZN(n8352) );
  NAND2_X1 U8849 ( .A1(n8353), .A2(n8352), .ZN(n8351) );
  NAND2_X1 U8850 ( .A1(n7208), .A2(n8536), .ZN(n7209) );
  NAND2_X1 U8851 ( .A1(n8351), .A2(n7209), .ZN(n8530) );
  XNOR2_X1 U8852 ( .A(n8963), .B(n7242), .ZN(n7212) );
  XNOR2_X1 U8853 ( .A(n7212), .B(n8889), .ZN(n8531) );
  INV_X1 U8854 ( .A(n7212), .ZN(n7213) );
  INV_X1 U8855 ( .A(n8889), .ZN(n8544) );
  XNOR2_X1 U8856 ( .A(n8429), .B(n7242), .ZN(n8426) );
  INV_X1 U8857 ( .A(n8878), .ZN(n8848) );
  NAND2_X1 U8858 ( .A1(n8426), .A2(n8848), .ZN(n7216) );
  INV_X1 U8859 ( .A(n8426), .ZN(n7215) );
  XNOR2_X1 U8860 ( .A(n9077), .B(n7242), .ZN(n7217) );
  XNOR2_X1 U8861 ( .A(n7217), .B(n8861), .ZN(n8434) );
  INV_X1 U8862 ( .A(n7217), .ZN(n7218) );
  XNOR2_X1 U8863 ( .A(n7219), .B(n7242), .ZN(n7220) );
  XNOR2_X1 U8864 ( .A(n7220), .B(n7222), .ZN(n8509) );
  INV_X1 U8865 ( .A(n7220), .ZN(n7221) );
  XNOR2_X1 U8866 ( .A(n9068), .B(n7242), .ZN(n7223) );
  XOR2_X1 U8867 ( .A(n8835), .B(n7223), .Z(n8377) );
  XNOR2_X1 U8868 ( .A(n9062), .B(n7242), .ZN(n7225) );
  XNOR2_X1 U8869 ( .A(n7225), .B(n8402), .ZN(n8467) );
  INV_X1 U8870 ( .A(n7225), .ZN(n7226) );
  XNOR2_X1 U8871 ( .A(n7227), .B(n7242), .ZN(n7228) );
  XNOR2_X1 U8872 ( .A(n7228), .B(n8468), .ZN(n8399) );
  INV_X1 U8873 ( .A(n7228), .ZN(n7229) );
  NAND2_X1 U8874 ( .A1(n7229), .A2(n8468), .ZN(n7230) );
  NAND2_X1 U8875 ( .A1(n7231), .A2(n7230), .ZN(n8484) );
  XNOR2_X1 U8876 ( .A(n9050), .B(n7242), .ZN(n7234) );
  XNOR2_X1 U8877 ( .A(n7234), .B(n8777), .ZN(n8483) );
  INV_X1 U8878 ( .A(n8483), .ZN(n7232) );
  INV_X1 U8879 ( .A(n7234), .ZN(n7235) );
  NAND2_X1 U8880 ( .A1(n7235), .A2(n8802), .ZN(n7236) );
  XNOR2_X1 U8881 ( .A(n9039), .B(n7249), .ZN(n8445) );
  INV_X1 U8882 ( .A(n8443), .ZN(n7237) );
  OAI22_X1 U8883 ( .A1(n8445), .A2(n8778), .B1(n8761), .B2(n7237), .ZN(n7241)
         );
  OAI21_X1 U8884 ( .B1(n8443), .B2(n8790), .A(n8746), .ZN(n7239) );
  NOR2_X1 U8885 ( .A1(n8746), .A2(n8790), .ZN(n7238) );
  AOI22_X1 U8886 ( .A1(n8445), .A2(n7239), .B1(n7238), .B2(n7237), .ZN(n7240)
         );
  XNOR2_X1 U8887 ( .A(n9033), .B(n7242), .ZN(n7244) );
  XNOR2_X1 U8888 ( .A(n7244), .B(n8739), .ZN(n8419) );
  XNOR2_X1 U8889 ( .A(n7243), .B(n7242), .ZN(n8518) );
  NAND2_X1 U8890 ( .A1(n7244), .A2(n8762), .ZN(n8516) );
  INV_X1 U8891 ( .A(n7245), .ZN(n7246) );
  NAND2_X1 U8892 ( .A1(n8518), .A2(n8747), .ZN(n7247) );
  NAND2_X1 U8893 ( .A1(n7248), .A2(n7247), .ZN(n8344) );
  XNOR2_X1 U8894 ( .A(n9021), .B(n7242), .ZN(n7281) );
  NOR2_X1 U8895 ( .A1(n7281), .A2(n7280), .ZN(n7256) );
  AOI21_X1 U8896 ( .B1(n7280), .B2(n7281), .A(n7256), .ZN(n8343) );
  NAND2_X1 U8897 ( .A1(n8344), .A2(n8343), .ZN(n8342) );
  XNOR2_X1 U8898 ( .A(n8730), .B(n7242), .ZN(n7250) );
  XNOR2_X1 U8899 ( .A(n7285), .B(n7250), .ZN(n7282) );
  INV_X1 U8900 ( .A(n7282), .ZN(n7255) );
  OR2_X1 U8901 ( .A1(n7258), .A2(n7251), .ZN(n7254) );
  INV_X1 U8902 ( .A(n7271), .ZN(n7252) );
  NAND2_X1 U8903 ( .A1(n7261), .A2(n7252), .ZN(n7253) );
  NAND2_X1 U8904 ( .A1(n7255), .A2(n8500), .ZN(n7288) );
  INV_X1 U8905 ( .A(n7256), .ZN(n7257) );
  NAND2_X1 U8906 ( .A1(n8342), .A2(n5228), .ZN(n7287) );
  OR2_X1 U8907 ( .A1(n7258), .A2(n10151), .ZN(n7259) );
  AND2_X1 U8908 ( .A1(n7261), .A2(n7260), .ZN(n7264) );
  NAND2_X1 U8909 ( .A1(n7264), .A2(n7262), .ZN(n8535) );
  NAND2_X1 U8910 ( .A1(n8543), .A2(n8533), .ZN(n7279) );
  INV_X1 U8911 ( .A(n7265), .ZN(n7267) );
  NAND2_X1 U8912 ( .A1(n7267), .A2(n7266), .ZN(n7270) );
  AND3_X1 U8913 ( .A1(n7268), .A2(n7399), .A3(n7292), .ZN(n7269) );
  OAI211_X1 U8914 ( .C1(n7274), .C2(n7271), .A(n7270), .B(n7269), .ZN(n7272)
         );
  NAND2_X1 U8915 ( .A1(n7272), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7276) );
  OR2_X1 U8916 ( .A1(n7274), .A2(n7273), .ZN(n7275) );
  NAND2_X2 U8917 ( .A1(n7276), .A2(n7275), .ZN(n8538) );
  AOI22_X1 U8918 ( .A1(n7277), .A2(n8538), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7278) );
  OAI211_X1 U8919 ( .C1(n7280), .C2(n8535), .A(n7279), .B(n7278), .ZN(n7284)
         );
  NOR4_X1 U8920 ( .A1(n7282), .A2(n7281), .A3(n7280), .A4(n8529), .ZN(n7283)
         );
  AOI211_X1 U8921 ( .C1(n7285), .C2(n8524), .A(n7284), .B(n7283), .ZN(n7286)
         );
  OAI211_X1 U8922 ( .C1(n8342), .C2(n7288), .A(n7287), .B(n7286), .ZN(P2_U3160) );
  INV_X1 U8923 ( .A(n7289), .ZN(n7290) );
  OR2_X2 U8924 ( .A1(n7291), .A2(n7290), .ZN(n9391) );
  INV_X1 U8925 ( .A(n7292), .ZN(n7398) );
  OAI21_X1 U8926 ( .B1(n7293), .B2(n7398), .A(n7399), .ZN(n7394) );
  NAND2_X1 U8927 ( .A1(n7394), .A2(n7392), .ZN(n7294) );
  NAND2_X1 U8928 ( .A1(n7294), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X2 U8929 ( .A1(n7338), .A2(n7398), .ZN(P2_U3893) );
  INV_X1 U8930 ( .A(n7295), .ZN(n7296) );
  NAND2_X1 U8931 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), .ZN(
        n10353) );
  OAI21_X1 U8932 ( .B1(n7296), .B2(P1_STATE_REG_SCAN_IN), .A(n10353), .ZN(
        P1_U3355) );
  NAND2_X1 U8933 ( .A1(n4397), .A2(P1_U3086), .ZN(n9940) );
  NAND2_X1 U8934 ( .A1(n4725), .A2(P1_U3086), .ZN(n9943) );
  INV_X1 U8935 ( .A(n9943), .ZN(n8305) );
  INV_X1 U8936 ( .A(n8305), .ZN(n9934) );
  OAI222_X1 U8937 ( .A1(n9940), .A2(n7298), .B1(n9934), .B2(n7306), .C1(
        P1_U3086), .C2(n4728), .ZN(P1_U3353) );
  OAI222_X1 U8938 ( .A1(n9943), .A2(n7302), .B1(n9940), .B2(n7299), .C1(
        P1_U3086), .C2(n9422), .ZN(P1_U3352) );
  OAI222_X1 U8939 ( .A1(n9943), .A2(n7307), .B1(n9940), .B2(n10311), .C1(
        P1_U3086), .C2(n7360), .ZN(P1_U3354) );
  INV_X1 U8940 ( .A(n7300), .ZN(n7304) );
  OAI222_X1 U8941 ( .A1(n9940), .A2(n7301), .B1(n9934), .B2(n7304), .C1(
        P1_U3086), .C2(n7366), .ZN(P1_U3351) );
  NOR2_X1 U8942 ( .A1(n4397), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9121) );
  INV_X2 U8943 ( .A(n9121), .ZN(n9130) );
  OAI222_X1 U8944 ( .A1(n7506), .A2(P2_U3151), .B1(n9132), .B2(n7302), .C1(
        n4703), .C2(n9130), .ZN(P2_U3292) );
  INV_X1 U8945 ( .A(n7555), .ZN(n7538) );
  OAI222_X1 U8946 ( .A1(P2_U3151), .A2(n7538), .B1(n9132), .B2(n7304), .C1(
        n7303), .C2(n9130), .ZN(P2_U3291) );
  OAI222_X1 U8947 ( .A1(P2_U3151), .A2(n7599), .B1(n9130), .B2(n5239), .C1(
        n9132), .C2(n7307), .ZN(P2_U3294) );
  OAI222_X1 U8948 ( .A1(n9940), .A2(n7308), .B1(n9934), .B2(n7315), .C1(n7408), 
        .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U8949 ( .A(n7553), .ZN(n7633) );
  OAI222_X1 U8950 ( .A1(n7633), .A2(P2_U3151), .B1(n9132), .B2(n8332), .C1(
        n7309), .C2(n9130), .ZN(P2_U3290) );
  INV_X1 U8951 ( .A(n7310), .ZN(n7316) );
  INV_X1 U8952 ( .A(n9940), .ZN(n9928) );
  AOI22_X1 U8953 ( .A1(n7680), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9928), .ZN(n7311) );
  OAI21_X1 U8954 ( .B1(n7316), .B2(n9943), .A(n7311), .ZN(P1_U3347) );
  INV_X1 U8955 ( .A(n7312), .ZN(n7324) );
  AOI22_X1 U8956 ( .A1(n7407), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9928), .ZN(n7313) );
  OAI21_X1 U8957 ( .B1(n7324), .B2(n9934), .A(n7313), .ZN(P1_U3349) );
  INV_X1 U8958 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7314) );
  OAI222_X1 U8959 ( .A1(n7640), .A2(P2_U3151), .B1(n9132), .B2(n7315), .C1(
        n7314), .C2(n9130), .ZN(P2_U3288) );
  INV_X1 U8960 ( .A(n7794), .ZN(n7797) );
  OAI222_X1 U8961 ( .A1(P2_U3151), .A2(n7797), .B1(n9132), .B2(n7316), .C1(
        n4635), .C2(n9130), .ZN(P2_U3287) );
  NAND2_X1 U8962 ( .A1(n7318), .A2(n7317), .ZN(n7319) );
  AND2_X1 U8963 ( .A1(n7320), .A2(n7319), .ZN(n7329) );
  INV_X1 U8964 ( .A(n7329), .ZN(n7322) );
  OR2_X1 U8965 ( .A1(n9923), .A2(n7321), .ZN(n7330) );
  NAND2_X1 U8966 ( .A1(n7322), .A2(n7330), .ZN(n9972) );
  INV_X1 U8967 ( .A(n9972), .ZN(n9506) );
  NOR2_X1 U8968 ( .A1(n9506), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8969 ( .A(n7604), .ZN(n7600) );
  OAI222_X1 U8970 ( .A1(P2_U3151), .A2(n7600), .B1(n9132), .B2(n7324), .C1(
        n7323), .C2(n9130), .ZN(P2_U3289) );
  NAND2_X1 U8971 ( .A1(P2_U3893), .A2(n6723), .ZN(n7325) );
  OAI21_X1 U8972 ( .B1(P2_U3893), .B2(n5413), .A(n7325), .ZN(P2_U3491) );
  INV_X1 U8973 ( .A(n9935), .ZN(n7327) );
  INV_X1 U8974 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7326) );
  AOI21_X1 U8975 ( .B1(n7327), .B2(n7326), .A(n8317), .ZN(n9408) );
  OAI21_X1 U8976 ( .B1(n7327), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9408), .ZN(
        n7328) );
  XOR2_X1 U8977 ( .A(P1_IR_REG_0__SCAN_IN), .B(n7328), .Z(n7332) );
  NAND2_X1 U8978 ( .A1(n7330), .A2(n7329), .ZN(n7371) );
  AOI22_X1 U8979 ( .A1(n9506), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n7331) );
  OAI21_X1 U8980 ( .B1(n7332), .B2(n7371), .A(n7331), .ZN(P1_U3243) );
  AND2_X1 U8981 ( .A1(n7341), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8982 ( .A1(n7341), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8983 ( .A1(n7341), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8984 ( .A1(n7341), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8985 ( .A1(n7341), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8986 ( .A1(n7341), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8987 ( .A1(n7341), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8988 ( .A1(n7341), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8989 ( .A1(n7341), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8990 ( .A1(n7341), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8991 ( .A1(n7341), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8992 ( .A1(n7341), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8993 ( .A1(n7341), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8994 ( .A1(n7341), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8995 ( .A1(n7341), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8996 ( .A1(n7341), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8997 ( .A1(n7341), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8998 ( .A1(n7341), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8999 ( .A1(n7341), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U9000 ( .A1(n7341), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U9001 ( .A1(n7341), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U9002 ( .A1(n7341), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U9003 ( .A1(n7341), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U9004 ( .A1(n7341), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U9005 ( .A1(n7341), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U9006 ( .A(n7334), .ZN(n7335) );
  AOI22_X1 U9007 ( .A1(n7341), .A2(n6374), .B1(n7338), .B2(n7335), .ZN(
        P2_U3376) );
  INV_X1 U9008 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7339) );
  INV_X1 U9009 ( .A(n7336), .ZN(n7337) );
  AOI22_X1 U9010 ( .A1(n7341), .A2(n7339), .B1(n7338), .B2(n7337), .ZN(
        P2_U3377) );
  AOI22_X1 U9011 ( .A1(n7983), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9928), .ZN(n7340) );
  OAI21_X1 U9012 ( .B1(n7344), .B2(n9934), .A(n7340), .ZN(P1_U3345) );
  INV_X1 U9013 ( .A(n7341), .ZN(n7342) );
  INV_X1 U9014 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10406) );
  NOR2_X1 U9015 ( .A1(n7342), .A2(n10406), .ZN(P2_U3239) );
  INV_X1 U9016 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10292) );
  NOR2_X1 U9017 ( .A1(n7342), .A2(n10292), .ZN(P2_U3250) );
  INV_X1 U9018 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10391) );
  NOR2_X1 U9019 ( .A1(n7342), .A2(n10391), .ZN(P2_U3260) );
  INV_X1 U9020 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10290) );
  NOR2_X1 U9021 ( .A1(n7342), .A2(n10290), .ZN(P2_U3262) );
  INV_X1 U9022 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10252) );
  NOR2_X1 U9023 ( .A1(n7342), .A2(n10252), .ZN(P2_U3245) );
  INV_X1 U9024 ( .A(n8185), .ZN(n8181) );
  INV_X1 U9025 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7343) );
  OAI222_X1 U9026 ( .A1(n8181), .A2(P2_U3151), .B1(n9132), .B2(n7344), .C1(
        n7343), .C2(n9130), .ZN(P2_U3285) );
  INV_X1 U9027 ( .A(n7911), .ZN(n7806) );
  INV_X1 U9028 ( .A(n7345), .ZN(n7346) );
  OAI222_X1 U9029 ( .A1(n7806), .A2(P2_U3151), .B1(n9132), .B2(n7346), .C1(
        n10440), .C2(n9130), .ZN(P2_U3286) );
  OAI222_X1 U9030 ( .A1(n9940), .A2(n7347), .B1(n9934), .B2(n7346), .C1(n7681), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U9031 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U9032 ( .A1(n9511), .A2(P1_U3973), .ZN(n7348) );
  OAI21_X1 U9033 ( .B1(P1_U3973), .B2(n10340), .A(n7348), .ZN(P1_U3585) );
  NAND2_X1 U9034 ( .A1(n6578), .A2(P1_U3973), .ZN(n7349) );
  OAI21_X1 U9035 ( .B1(P1_U3973), .B2(n5240), .A(n7349), .ZN(P1_U3554) );
  INV_X1 U9036 ( .A(n7350), .ZN(n7389) );
  AOI22_X1 U9037 ( .A1(n8122), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9928), .ZN(n7351) );
  OAI21_X1 U9038 ( .B1(n7389), .B2(n9934), .A(n7351), .ZN(P1_U3344) );
  AND2_X1 U9039 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9404) );
  NAND2_X1 U9040 ( .A1(n4632), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7352) );
  INV_X1 U9041 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7353) );
  OR2_X1 U9042 ( .A1(n4728), .A2(n7353), .ZN(n7354) );
  XNOR2_X1 U9043 ( .A(n9422), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9428) );
  INV_X1 U9044 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7786) );
  OR2_X1 U9045 ( .A1(n9422), .A2(n7786), .ZN(n7355) );
  XNOR2_X1 U9046 ( .A(n7366), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9442) );
  INV_X1 U9047 ( .A(n7366), .ZN(n9445) );
  NAND2_X1 U9048 ( .A1(n9445), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7356) );
  INV_X1 U9049 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7357) );
  INV_X1 U9050 ( .A(n7371), .ZN(n7368) );
  NAND2_X1 U9051 ( .A1(n7368), .A2(n7358), .ZN(n9963) );
  AOI211_X1 U9052 ( .C1(n5237), .C2(n7359), .A(n7379), .B(n9963), .ZN(n7375)
         );
  INV_X1 U9053 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10375) );
  AND2_X1 U9054 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9396) );
  NAND2_X1 U9055 ( .A1(n4632), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7361) );
  NAND2_X1 U9056 ( .A1(n9395), .A2(n7361), .ZN(n9417) );
  INV_X1 U9057 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7703) );
  OR2_X1 U9058 ( .A1(n4728), .A2(n7703), .ZN(n7363) );
  XNOR2_X1 U9059 ( .A(n9422), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9431) );
  INV_X1 U9060 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7364) );
  OR2_X1 U9061 ( .A1(n9422), .A2(n7364), .ZN(n7365) );
  XNOR2_X1 U9062 ( .A(n7366), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9439) );
  INV_X1 U9063 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7367) );
  MUX2_X1 U9064 ( .A(n7367), .B(P1_REG1_REG_5__SCAN_IN), .S(n8330), .Z(n7369)
         );
  NAND2_X1 U9065 ( .A1(n7368), .A2(n9935), .ZN(n9959) );
  AOI211_X1 U9066 ( .C1(n7370), .C2(n7369), .A(n4518), .B(n9959), .ZN(n7374)
         );
  INV_X1 U9067 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10204) );
  NOR2_X2 U9068 ( .A1(n7371), .A2(n9405), .ZN(n9968) );
  NAND2_X1 U9069 ( .A1(n9968), .A2(n8330), .ZN(n7372) );
  NAND2_X1 U9070 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n8077) );
  OAI211_X1 U9071 ( .C1(n10204), .C2(n9972), .A(n7372), .B(n8077), .ZN(n7373)
         );
  OR3_X1 U9072 ( .A1(n7375), .A2(n7374), .A3(n7373), .ZN(P1_U3248) );
  INV_X1 U9073 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7376) );
  MUX2_X1 U9074 ( .A(n7376), .B(P1_REG1_REG_6__SCAN_IN), .S(n7407), .Z(n7377)
         );
  AOI211_X1 U9075 ( .C1(n7378), .C2(n7377), .A(n9959), .B(n7403), .ZN(n7387)
         );
  INV_X1 U9076 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7380) );
  MUX2_X1 U9077 ( .A(n7380), .B(P1_REG2_REG_6__SCAN_IN), .S(n7407), .Z(n7381)
         );
  NOR2_X1 U9078 ( .A1(n7382), .A2(n7381), .ZN(n7406) );
  AOI211_X1 U9079 ( .C1(n7382), .C2(n7381), .A(n9963), .B(n7406), .ZN(n7386)
         );
  INV_X1 U9080 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7384) );
  NAND2_X1 U9081 ( .A1(n9968), .A2(n7407), .ZN(n7383) );
  NAND2_X1 U9082 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7962) );
  OAI211_X1 U9083 ( .C1(n7384), .C2(n9972), .A(n7383), .B(n7962), .ZN(n7385)
         );
  OR3_X1 U9084 ( .A1(n7387), .A2(n7386), .A3(n7385), .ZN(P1_U3249) );
  INV_X1 U9085 ( .A(n8243), .ZN(n8202) );
  INV_X1 U9086 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7388) );
  OAI222_X1 U9087 ( .A1(P2_U3151), .A2(n8202), .B1(n9132), .B2(n7389), .C1(
        n7388), .C2(n9130), .ZN(P2_U3284) );
  AND2_X1 U9088 ( .A1(n7394), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7391) );
  MUX2_X1 U9089 ( .A(n7391), .B(P2_U3893), .S(n7390), .Z(n7393) );
  NAND2_X1 U9090 ( .A1(n7393), .A2(n7392), .ZN(n8705) );
  INV_X1 U9091 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7432) );
  AND2_X1 U9092 ( .A1(P2_U3893), .A2(n6342), .ZN(n8707) );
  NOR2_X1 U9093 ( .A1(n6342), .A2(P2_U3151), .ZN(n9120) );
  AND2_X1 U9094 ( .A1(n7394), .A2(n9120), .ZN(n7418) );
  INV_X1 U9095 ( .A(n7418), .ZN(n7447) );
  MUX2_X1 U9096 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n9125), .Z(n7395) );
  NOR2_X1 U9097 ( .A1(n7395), .A2(n7432), .ZN(n7587) );
  AOI21_X1 U9098 ( .B1(n7432), .B2(n7395), .A(n7587), .ZN(n7396) );
  AOI21_X1 U9099 ( .B1(n8683), .B2(n7447), .A(n7396), .ZN(n7397) );
  AOI21_X1 U9100 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n7397), .ZN(
        n7402) );
  AND2_X1 U9101 ( .A1(n7399), .A2(n7398), .ZN(n7400) );
  INV_X1 U9102 ( .A(n8622), .ZN(n8701) );
  NAND2_X1 U9103 ( .A1(n8701), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n7401) );
  OAI211_X1 U9104 ( .C1(n8705), .C2(n7432), .A(n7402), .B(n7401), .ZN(P2_U3182) );
  XOR2_X1 U9105 ( .A(n7408), .B(P1_REG1_REG_7__SCAN_IN), .Z(n7404) );
  AOI211_X1 U9106 ( .C1(n7405), .C2(n7404), .A(n9959), .B(n7518), .ZN(n7415)
         );
  INV_X1 U9107 ( .A(n7408), .ZN(n7522) );
  XNOR2_X1 U9108 ( .A(n7522), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7409) );
  NOR2_X1 U9109 ( .A1(n7410), .A2(n7409), .ZN(n7521) );
  AOI211_X1 U9110 ( .C1(n7410), .C2(n7409), .A(n9963), .B(n7521), .ZN(n7414)
         );
  INV_X1 U9111 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7412) );
  NAND2_X1 U9112 ( .A1(n9968), .A2(n7522), .ZN(n7411) );
  NAND2_X1 U9113 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n8110) );
  OAI211_X1 U9114 ( .C1(n7412), .C2(n9972), .A(n7411), .B(n8110), .ZN(n7413)
         );
  OR3_X1 U9115 ( .A1(n7415), .A2(n7414), .A3(n7413), .ZN(P1_U3250) );
  INV_X1 U9116 ( .A(n7416), .ZN(n7467) );
  AOI22_X1 U9117 ( .A1(n8297), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9928), .ZN(n7417) );
  OAI21_X1 U9118 ( .B1(n7467), .B2(n9934), .A(n7417), .ZN(P1_U3343) );
  INV_X1 U9119 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7431) );
  INV_X1 U9120 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7419) );
  MUX2_X1 U9121 ( .A(n7419), .B(P2_REG1_REG_4__SCAN_IN), .S(n7555), .Z(n7428)
         );
  INV_X1 U9122 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7420) );
  NAND2_X1 U9123 ( .A1(n7432), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7422) );
  INV_X1 U9124 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U9125 ( .A1(n7433), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U9126 ( .A1(n7599), .A2(n7423), .ZN(n7421) );
  OAI21_X1 U9127 ( .B1(n7433), .B2(n7422), .A(n7421), .ZN(n7592) );
  NAND2_X1 U9128 ( .A1(n7592), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7424) );
  INV_X1 U9129 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U9130 ( .A1(n7427), .A2(n7428), .ZN(n7551) );
  OAI21_X1 U9131 ( .B1(n7428), .B2(n7427), .A(n7551), .ZN(n7429) );
  NAND2_X1 U9132 ( .A1(n8714), .A2(n7429), .ZN(n7430) );
  OAI21_X1 U9133 ( .B1(n8622), .B2(n7431), .A(n7430), .ZN(n7450) );
  INV_X1 U9134 ( .A(n7599), .ZN(n7435) );
  NAND2_X1 U9135 ( .A1(n7432), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7434) );
  AND2_X1 U9136 ( .A1(n7433), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7436) );
  AOI21_X1 U9137 ( .B1(n7435), .B2(n7434), .A(n7436), .ZN(n7590) );
  NAND2_X1 U9138 ( .A1(n7590), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7589) );
  INV_X1 U9139 ( .A(n7436), .ZN(n7437) );
  NAND2_X1 U9140 ( .A1(n7589), .A2(n7437), .ZN(n7574) );
  INV_X1 U9141 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7438) );
  NAND2_X1 U9142 ( .A1(n7574), .A2(n7575), .ZN(n7573) );
  INV_X1 U9143 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10119) );
  XNOR2_X1 U9144 ( .A(n7555), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7444) );
  INV_X1 U9145 ( .A(n7444), .ZN(n7446) );
  NAND3_X1 U9146 ( .A1(n7443), .A2(n7446), .A3(n7445), .ZN(n7448) );
  OR2_X1 U9147 ( .A1(n7447), .A2(n4387), .ZN(n8717) );
  AOI21_X1 U9148 ( .B1(n7557), .B2(n7448), .A(n8717), .ZN(n7449) );
  AND2_X1 U9149 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8457) );
  NOR3_X1 U9150 ( .A1(n7450), .A2(n7449), .A3(n8457), .ZN(n7463) );
  XNOR2_X1 U9151 ( .A(n7451), .B(n7599), .ZN(n7588) );
  NAND2_X1 U9152 ( .A1(n7451), .A2(n7599), .ZN(n7452) );
  MUX2_X1 U9153 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9125), .Z(n7453) );
  XNOR2_X1 U9154 ( .A(n7453), .B(n4395), .ZN(n7571) );
  INV_X1 U9155 ( .A(n7453), .ZN(n7454) );
  NOR2_X1 U9156 ( .A1(n7454), .A2(n4395), .ZN(n7455) );
  AOI21_X1 U9157 ( .B1(n7572), .B2(n7571), .A(n7455), .ZN(n7502) );
  MUX2_X1 U9158 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n4705), .Z(n7456) );
  XNOR2_X1 U9159 ( .A(n7456), .B(n4644), .ZN(n7501) );
  NAND2_X1 U9160 ( .A1(n7502), .A2(n7501), .ZN(n7500) );
  INV_X1 U9161 ( .A(n7500), .ZN(n7457) );
  NOR2_X1 U9162 ( .A1(n7456), .A2(n7506), .ZN(n7458) );
  MUX2_X1 U9163 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4705), .Z(n7539) );
  XNOR2_X1 U9164 ( .A(n7539), .B(n7538), .ZN(n7459) );
  OAI21_X1 U9165 ( .B1(n7457), .B2(n7458), .A(n7459), .ZN(n7461) );
  NOR2_X1 U9166 ( .A1(n7459), .A2(n7458), .ZN(n7460) );
  NAND2_X1 U9167 ( .A1(n7500), .A2(n7460), .ZN(n7541) );
  NAND3_X1 U9168 ( .A1(n7461), .A2(n8707), .A3(n7541), .ZN(n7462) );
  OAI211_X1 U9169 ( .C1(n8705), .C2(n7538), .A(n7463), .B(n7462), .ZN(P2_U3186) );
  INV_X1 U9170 ( .A(n8538), .ZN(n7777) );
  NAND2_X1 U9171 ( .A1(n7777), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7487) );
  NAND2_X1 U9172 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n7487), .ZN(n7465) );
  INV_X1 U9173 ( .A(n10131), .ZN(n7737) );
  AOI22_X1 U9174 ( .A1(n7737), .A2(n8500), .B1(n8524), .B2(n10136), .ZN(n7464)
         );
  OAI211_X1 U9175 ( .C1(n8489), .C2(n8999), .A(n7465), .B(n7464), .ZN(P2_U3172) );
  INV_X1 U9176 ( .A(n8258), .ZN(n8554) );
  INV_X1 U9177 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7466) );
  OAI222_X1 U9178 ( .A1(n8554), .A2(P2_U3151), .B1(n9132), .B2(n7467), .C1(
        n7466), .C2(n9130), .ZN(P2_U3283) );
  INV_X1 U9179 ( .A(n7487), .ZN(n7477) );
  INV_X1 U9180 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7476) );
  OAI22_X1 U9181 ( .A1(n8489), .A2(n7468), .B1(n8999), .B2(n8535), .ZN(n7469)
         );
  AOI21_X1 U9182 ( .B1(n9004), .B2(n8524), .A(n7469), .ZN(n7475) );
  OAI21_X1 U9183 ( .B1(n7472), .B2(n7470), .A(n7471), .ZN(n7473) );
  NAND2_X1 U9184 ( .A1(n7473), .A2(n8500), .ZN(n7474) );
  OAI211_X1 U9185 ( .C1(n7477), .C2(n7476), .A(n7475), .B(n7474), .ZN(P2_U3177) );
  NAND2_X1 U9186 ( .A1(n10057), .A2(n9881), .ZN(n7479) );
  AOI222_X1 U9187 ( .A1(n7479), .A2(n8321), .B1(n8325), .B2(n7478), .C1(n4646), 
        .C2(n9986), .ZN(n10004) );
  NAND2_X1 U9188 ( .A1(n10101), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7480) );
  OAI21_X1 U9189 ( .B1(n10004), .B2(n10101), .A(n7480), .ZN(P1_U3522) );
  INV_X1 U9190 ( .A(n7481), .ZN(n7482) );
  AOI21_X1 U9191 ( .B1(n7484), .B2(n7483), .A(n7482), .ZN(n7489) );
  AOI22_X1 U9192 ( .A1(n8487), .A2(n6723), .B1(n8533), .B2(n6397), .ZN(n7485)
         );
  OAI21_X1 U9193 ( .B1(n8541), .B2(n6396), .A(n7485), .ZN(n7486) );
  AOI21_X1 U9194 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7487), .A(n7486), .ZN(
        n7488) );
  OAI21_X1 U9195 ( .B1(n8529), .B2(n7489), .A(n7488), .ZN(P2_U3162) );
  INV_X1 U9196 ( .A(n7490), .ZN(n7517) );
  AOI22_X1 U9197 ( .A1(n9466), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9928), .ZN(n7491) );
  OAI21_X1 U9198 ( .B1(n7517), .B2(n9934), .A(n7491), .ZN(P1_U3341) );
  INV_X1 U9199 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7495) );
  INV_X1 U9200 ( .A(n7443), .ZN(n7492) );
  AOI21_X1 U9201 ( .B1(n10119), .B2(n7493), .A(n7492), .ZN(n7494) );
  OAI22_X1 U9202 ( .A1(n8622), .A2(n7495), .B1(n8717), .B2(n7494), .ZN(n7499)
         );
  XNOR2_X1 U9203 ( .A(n7496), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n7497) );
  NOR2_X1 U9204 ( .A1(n8690), .A2(n7497), .ZN(n7498) );
  AOI211_X1 U9205 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3151), .A(n7499), .B(
        n7498), .ZN(n7505) );
  OAI21_X1 U9206 ( .B1(n7502), .B2(n7501), .A(n7500), .ZN(n7503) );
  NAND2_X1 U9207 ( .A1(n7503), .A2(n8707), .ZN(n7504) );
  OAI211_X1 U9208 ( .C1(n8705), .C2(n7506), .A(n7505), .B(n7504), .ZN(P2_U3185) );
  XNOR2_X1 U9209 ( .A(n7508), .B(n7507), .ZN(n9403) );
  INV_X1 U9210 ( .A(n7509), .ZN(n9259) );
  NAND2_X1 U9211 ( .A1(n9259), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9341) );
  AOI22_X1 U9212 ( .A1(n9378), .A2(n8325), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9341), .ZN(n7511) );
  NAND2_X1 U9213 ( .A1(n9365), .A2(n4646), .ZN(n7510) );
  OAI211_X1 U9214 ( .C1(n9403), .C2(n9380), .A(n7511), .B(n7510), .ZN(P1_U3232) );
  INV_X1 U9215 ( .A(n7512), .ZN(n7515) );
  OAI222_X1 U9216 ( .A1(P2_U3151), .A2(n4984), .B1(n9132), .B2(n7515), .C1(
        n7513), .C2(n9130), .ZN(P2_U3282) );
  OAI222_X1 U9217 ( .A1(n9940), .A2(n7516), .B1(n9934), .B2(n7515), .C1(
        P1_U3086), .C2(n7514), .ZN(P1_U3342) );
  INV_X1 U9218 ( .A(n8587), .ZN(n8597) );
  INV_X1 U9219 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10277) );
  OAI222_X1 U9220 ( .A1(P2_U3151), .A2(n8597), .B1(n9132), .B2(n7517), .C1(
        n10277), .C2(n9130), .ZN(P2_U3281) );
  AOI21_X1 U9221 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n7522), .A(n7518), .ZN(
        n7520) );
  XNOR2_X1 U9222 ( .A(n7680), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7519) );
  AOI211_X1 U9223 ( .C1(n7520), .C2(n7519), .A(n9959), .B(n7679), .ZN(n7529)
         );
  XNOR2_X1 U9224 ( .A(n7680), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7523) );
  AOI211_X1 U9225 ( .C1(n7524), .C2(n7523), .A(n9963), .B(n7674), .ZN(n7528)
         );
  INV_X1 U9226 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7526) );
  NAND2_X1 U9227 ( .A1(n9968), .A2(n7680), .ZN(n7525) );
  NAND2_X1 U9228 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9200) );
  OAI211_X1 U9229 ( .C1(n7526), .C2(n9972), .A(n7525), .B(n9200), .ZN(n7527)
         );
  OR3_X1 U9230 ( .A1(n7529), .A2(n7528), .A3(n7527), .ZN(P1_U3251) );
  MUX2_X1 U9231 ( .A(n8538), .B(P2_U3151), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n7533) );
  OAI22_X1 U9232 ( .A1(n8489), .A2(n7531), .B1(n7530), .B2(n8535), .ZN(n7532)
         );
  AOI211_X1 U9233 ( .C1(n10140), .C2(n8524), .A(n7533), .B(n7532), .ZN(n7537)
         );
  NAND2_X1 U9234 ( .A1(n7537), .A2(n7536), .ZN(P2_U3158) );
  NAND2_X1 U9235 ( .A1(n7539), .A2(n7538), .ZN(n7540) );
  NAND2_X1 U9236 ( .A1(n7541), .A2(n7540), .ZN(n7627) );
  MUX2_X1 U9237 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4387), .Z(n7542) );
  XNOR2_X1 U9238 ( .A(n7542), .B(n7553), .ZN(n7626) );
  NAND2_X1 U9239 ( .A1(n7627), .A2(n7626), .ZN(n7544) );
  NAND2_X1 U9240 ( .A1(n7542), .A2(n7633), .ZN(n7543) );
  NAND2_X1 U9241 ( .A1(n7544), .A2(n7543), .ZN(n7550) );
  INV_X1 U9242 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7603) );
  INV_X1 U9243 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7727) );
  MUX2_X1 U9244 ( .A(n7603), .B(n7727), .S(n4387), .Z(n7545) );
  NAND2_X1 U9245 ( .A1(n7545), .A2(n7604), .ZN(n7618) );
  INV_X1 U9246 ( .A(n7545), .ZN(n7546) );
  NAND2_X1 U9247 ( .A1(n7546), .A2(n7600), .ZN(n7547) );
  NAND2_X1 U9248 ( .A1(n7618), .A2(n7547), .ZN(n7549) );
  INV_X1 U9249 ( .A(n7619), .ZN(n7548) );
  AOI21_X1 U9250 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n7570) );
  INV_X1 U9251 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7554) );
  XNOR2_X1 U9252 ( .A(n7604), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7601) );
  XNOR2_X1 U9253 ( .A(n7602), .B(n7601), .ZN(n7568) );
  INV_X1 U9254 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7745) );
  OR2_X1 U9255 ( .A1(n7555), .A2(n7745), .ZN(n7556) );
  NAND2_X1 U9256 ( .A1(n7629), .A2(n7561), .ZN(n7559) );
  XNOR2_X1 U9257 ( .A(n7604), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7560) );
  INV_X1 U9258 ( .A(n7560), .ZN(n7562) );
  NAND3_X1 U9259 ( .A1(n7629), .A2(n7562), .A3(n7561), .ZN(n7563) );
  AOI21_X1 U9260 ( .B1(n7606), .B2(n7563), .A(n8717), .ZN(n7567) );
  INV_X1 U9261 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U9262 ( .A1(n8634), .A2(n7604), .ZN(n7564) );
  NAND2_X1 U9263 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7836) );
  OAI211_X1 U9264 ( .C1(n7565), .C2(n8622), .A(n7564), .B(n7836), .ZN(n7566)
         );
  AOI211_X1 U9265 ( .C1(n8714), .C2(n7568), .A(n7567), .B(n7566), .ZN(n7569)
         );
  OAI21_X1 U9266 ( .B1(n7570), .B2(n8683), .A(n7569), .ZN(P2_U3188) );
  XNOR2_X1 U9267 ( .A(n7572), .B(n7571), .ZN(n7586) );
  INV_X1 U9268 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7582) );
  OAI21_X1 U9269 ( .B1(n7575), .B2(n7574), .A(n7573), .ZN(n7576) );
  AOI22_X1 U9270 ( .A1(n8670), .A2(n7576), .B1(P2_U3151), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7581) );
  XNOR2_X1 U9271 ( .A(n7578), .B(n7577), .ZN(n7579) );
  NAND2_X1 U9272 ( .A1(n8714), .A2(n7579), .ZN(n7580) );
  OAI211_X1 U9273 ( .C1(n7582), .C2(n8622), .A(n7581), .B(n7580), .ZN(n7583)
         );
  AOI21_X1 U9274 ( .B1(n4395), .B2(n8634), .A(n7583), .ZN(n7585) );
  OAI21_X1 U9275 ( .B1(n8683), .B2(n7586), .A(n7585), .ZN(P2_U3184) );
  XOR2_X1 U9276 ( .A(n7588), .B(n7587), .Z(n7597) );
  INV_X1 U9277 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10171) );
  OAI21_X1 U9278 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n7590), .A(n7589), .ZN(
        n7591) );
  AOI22_X1 U9279 ( .A1(n8670), .A2(n7591), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n7595) );
  XNOR2_X1 U9280 ( .A(n7592), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9281 ( .A1(n8714), .A2(n7593), .ZN(n7594) );
  OAI211_X1 U9282 ( .C1(n10171), .C2(n8622), .A(n7595), .B(n7594), .ZN(n7596)
         );
  AOI21_X1 U9283 ( .B1(n8707), .B2(n7597), .A(n7596), .ZN(n7598) );
  OAI21_X1 U9284 ( .B1(n7599), .B2(n8705), .A(n7598), .ZN(P2_U3183) );
  INV_X1 U9285 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7904) );
  XNOR2_X1 U9286 ( .A(n7641), .B(n7904), .ZN(n7625) );
  OR2_X1 U9287 ( .A1(n7604), .A2(n7603), .ZN(n7605) );
  INV_X1 U9288 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7610) );
  OAI21_X1 U9289 ( .B1(n4508), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7655), .ZN(
        n7623) );
  INV_X1 U9290 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9291 ( .A1(n8634), .A2(n7611), .ZN(n7608) );
  AND2_X1 U9292 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7971) );
  INV_X1 U9293 ( .A(n7971), .ZN(n7607) );
  OAI211_X1 U9294 ( .C1(n7609), .C2(n8622), .A(n7608), .B(n7607), .ZN(n7622)
         );
  NAND2_X1 U9295 ( .A1(n7619), .A2(n7618), .ZN(n7616) );
  MUX2_X1 U9296 ( .A(n7610), .B(n7904), .S(n4387), .Z(n7612) );
  NAND2_X1 U9297 ( .A1(n7612), .A2(n7611), .ZN(n7648) );
  INV_X1 U9298 ( .A(n7612), .ZN(n7613) );
  NAND2_X1 U9299 ( .A1(n7613), .A2(n7640), .ZN(n7614) );
  NAND2_X1 U9300 ( .A1(n7648), .A2(n7614), .ZN(n7617) );
  INV_X1 U9301 ( .A(n7617), .ZN(n7615) );
  NAND3_X1 U9302 ( .A1(n7619), .A2(n7618), .A3(n7617), .ZN(n7620) );
  AOI21_X1 U9303 ( .B1(n7649), .B2(n7620), .A(n8683), .ZN(n7621) );
  AOI211_X1 U9304 ( .C1(n8670), .C2(n7623), .A(n7622), .B(n7621), .ZN(n7624)
         );
  OAI21_X1 U9305 ( .B1(n7625), .B2(n8690), .A(n7624), .ZN(P2_U3189) );
  XNOR2_X1 U9306 ( .A(n7627), .B(n7626), .ZN(n7637) );
  XOR2_X1 U9307 ( .A(n7628), .B(P2_REG1_REG_5__SCAN_IN), .Z(n7635) );
  OAI21_X1 U9308 ( .B1(n5233), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7629), .ZN(
        n7631) );
  AND2_X1 U9309 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7774) );
  INV_X1 U9310 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10454) );
  NOR2_X1 U9311 ( .A1(n8622), .A2(n10454), .ZN(n7630) );
  AOI211_X1 U9312 ( .C1(n8670), .C2(n7631), .A(n7774), .B(n7630), .ZN(n7632)
         );
  OAI21_X1 U9313 ( .B1(n7633), .B2(n8705), .A(n7632), .ZN(n7634) );
  AOI21_X1 U9314 ( .B1(n8714), .B2(n7635), .A(n7634), .ZN(n7636) );
  OAI21_X1 U9315 ( .B1(n8683), .B2(n7637), .A(n7636), .ZN(P2_U3187) );
  XOR2_X1 U9316 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7794), .Z(n7795) );
  INV_X1 U9317 ( .A(n7638), .ZN(n7639) );
  XOR2_X1 U9318 ( .A(n7795), .B(n7796), .Z(n7662) );
  NAND2_X1 U9319 ( .A1(n7649), .A2(n7648), .ZN(n7646) );
  INV_X1 U9320 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7952) );
  INV_X1 U9321 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10293) );
  MUX2_X1 U9322 ( .A(n7952), .B(n10293), .S(n4387), .Z(n7642) );
  NAND2_X1 U9323 ( .A1(n7642), .A2(n7794), .ZN(n7812) );
  INV_X1 U9324 ( .A(n7642), .ZN(n7643) );
  NAND2_X1 U9325 ( .A1(n7643), .A2(n7797), .ZN(n7644) );
  NAND2_X1 U9326 ( .A1(n7812), .A2(n7644), .ZN(n7647) );
  INV_X1 U9327 ( .A(n7647), .ZN(n7645) );
  NAND3_X1 U9328 ( .A1(n7649), .A2(n7648), .A3(n7647), .ZN(n7650) );
  AOI21_X1 U9329 ( .B1(n7813), .B2(n7650), .A(n8683), .ZN(n7660) );
  XNOR2_X1 U9330 ( .A(n7794), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7652) );
  INV_X1 U9331 ( .A(n7652), .ZN(n7654) );
  NAND3_X1 U9332 ( .A1(n7655), .A2(n7654), .A3(n7653), .ZN(n7656) );
  AOI21_X1 U9333 ( .B1(n7799), .B2(n7656), .A(n8717), .ZN(n7659) );
  AND2_X1 U9334 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8392) );
  AOI21_X1 U9335 ( .B1(n8701), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8392), .ZN(
        n7657) );
  OAI21_X1 U9336 ( .B1(n7797), .B2(n8705), .A(n7657), .ZN(n7658) );
  NOR3_X1 U9337 ( .A1(n7660), .A2(n7659), .A3(n7658), .ZN(n7661) );
  OAI21_X1 U9338 ( .B1(n7662), .B2(n8690), .A(n7661), .ZN(P2_U3190) );
  NOR2_X1 U9339 ( .A1(n6580), .A2(n7663), .ZN(n7691) );
  INV_X1 U9340 ( .A(n7691), .ZN(n7664) );
  OAI21_X1 U9341 ( .B1(n7669), .B2(n7665), .A(n7664), .ZN(n7714) );
  AOI22_X1 U9342 ( .A1(n6578), .A2(n10053), .B1(n10078), .B2(n5848), .ZN(n7667) );
  NAND2_X1 U9343 ( .A1(n5848), .A2(n8325), .ZN(n7666) );
  NAND3_X1 U9344 ( .A1(n7698), .A2(n9975), .A3(n7666), .ZN(n7718) );
  OAI211_X1 U9345 ( .C1(n9212), .C2(n10065), .A(n7667), .B(n7718), .ZN(n7672)
         );
  NAND2_X1 U9346 ( .A1(n7669), .A2(n7668), .ZN(n7671) );
  AOI21_X1 U9347 ( .B1(n7671), .B2(n7670), .A(n9881), .ZN(n7720) );
  AOI211_X1 U9348 ( .C1(n10087), .C2(n7714), .A(n7672), .B(n7720), .ZN(n7688)
         );
  NAND2_X1 U9349 ( .A1(n10101), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7673) );
  OAI21_X1 U9350 ( .B1(n7688), .B2(n10101), .A(n7673), .ZN(P1_U3523) );
  XNOR2_X1 U9351 ( .A(n7681), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7675) );
  OAI21_X1 U9352 ( .B1(n7675), .B2(n4514), .A(n7843), .ZN(n7678) );
  INV_X1 U9353 ( .A(n9963), .ZN(n9496) );
  NAND2_X1 U9354 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U9355 ( .A1(n9506), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n7676) );
  OAI211_X1 U9356 ( .C1(n4733), .C2(n7681), .A(n9293), .B(n7676), .ZN(n7677)
         );
  AOI21_X1 U9357 ( .B1(n7678), .B2(n9496), .A(n7677), .ZN(n7687) );
  INV_X1 U9358 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7682) );
  MUX2_X1 U9359 ( .A(n7682), .B(P1_REG1_REG_9__SCAN_IN), .S(n7681), .Z(n7683)
         );
  OAI21_X1 U9360 ( .B1(n7684), .B2(n7683), .A(n7847), .ZN(n7685) );
  INV_X1 U9361 ( .A(n9959), .ZN(n9502) );
  NAND2_X1 U9362 ( .A1(n7685), .A2(n9502), .ZN(n7686) );
  NAND2_X1 U9363 ( .A1(n7687), .A2(n7686), .ZN(P1_U3252) );
  INV_X1 U9364 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7690) );
  OR2_X1 U9365 ( .A1(n7688), .A2(n10088), .ZN(n7689) );
  OAI21_X1 U9366 ( .B1(n10090), .B2(n7690), .A(n7689), .ZN(P1_U3456) );
  INV_X1 U9367 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10467) );
  AOI21_X1 U9368 ( .B1(n4648), .B2(n7692), .A(n7691), .ZN(n7693) );
  XNOR2_X1 U9369 ( .A(n6581), .B(n7693), .ZN(n7713) );
  INV_X1 U9370 ( .A(n6581), .ZN(n7694) );
  XNOR2_X1 U9371 ( .A(n6643), .B(n7694), .ZN(n7696) );
  OAI22_X1 U9372 ( .A1(n10011), .A2(n10065), .B1(n4648), .B2(n10082), .ZN(
        n7695) );
  AOI21_X1 U9373 ( .B1(n7696), .B2(n10061), .A(n7695), .ZN(n7710) );
  INV_X1 U9374 ( .A(n7697), .ZN(n7788) );
  AOI21_X1 U9375 ( .B1(n10078), .B2(n9342), .A(n7707), .ZN(n7699) );
  OAI211_X1 U9376 ( .C1(n7713), .C2(n10057), .A(n7710), .B(n7699), .ZN(n7701)
         );
  NAND2_X1 U9377 ( .A1(n7701), .A2(n10090), .ZN(n7700) );
  OAI21_X1 U9378 ( .B1(n10090), .B2(n10467), .A(n7700), .ZN(P1_U3459) );
  NAND2_X1 U9379 ( .A1(n7701), .A2(n10103), .ZN(n7702) );
  OAI21_X1 U9380 ( .B1(n10103), .B2(n7703), .A(n7702), .ZN(P1_U3524) );
  INV_X1 U9381 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7705) );
  INV_X1 U9382 ( .A(n7704), .ZN(n7706) );
  INV_X1 U9383 ( .A(n9954), .ZN(n9467) );
  OAI222_X1 U9384 ( .A1(n9940), .A2(n7705), .B1(n9934), .B2(n7706), .C1(
        P1_U3086), .C2(n9467), .ZN(P1_U3340) );
  OAI222_X1 U9385 ( .A1(P2_U3151), .A2(n4897), .B1(n9132), .B2(n7706), .C1(
        n10451), .C2(n9130), .ZN(P2_U3280) );
  INV_X1 U9386 ( .A(n7707), .ZN(n7708) );
  INV_X1 U9387 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9409) );
  OAI22_X1 U9388 ( .A1(n7708), .A2(n9743), .B1(n9409), .B2(n9671), .ZN(n7709)
         );
  AOI21_X1 U9389 ( .B1(n9747), .B2(n9342), .A(n7709), .ZN(n7712) );
  MUX2_X1 U9390 ( .A(n7353), .B(n7710), .S(n9997), .Z(n7711) );
  OAI211_X1 U9391 ( .C1(n9765), .C2(n7713), .A(n7712), .B(n7711), .ZN(P1_U3291) );
  INV_X1 U9392 ( .A(n7714), .ZN(n7723) );
  INV_X1 U9393 ( .A(n9522), .ZN(n9738) );
  AOI22_X1 U9394 ( .A1(n9738), .A2(n6578), .B1(n9747), .B2(n5848), .ZN(n7722)
         );
  INV_X1 U9395 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9392) );
  OAI22_X1 U9396 ( .A1(n9997), .A2(n10344), .B1(n9392), .B2(n9671), .ZN(n7715)
         );
  INV_X1 U9397 ( .A(n7715), .ZN(n7717) );
  NAND2_X1 U9398 ( .A1(n9997), .A2(n9986), .ZN(n9741) );
  OR2_X1 U9399 ( .A1(n9741), .A2(n9212), .ZN(n7716) );
  OAI211_X1 U9400 ( .C1(n7718), .C2(n9743), .A(n7717), .B(n7716), .ZN(n7719)
         );
  AOI21_X1 U9401 ( .B1(n7720), .B2(n9997), .A(n7719), .ZN(n7721) );
  OAI211_X1 U9402 ( .C1(n9765), .C2(n7723), .A(n7722), .B(n7721), .ZN(P1_U3292) );
  XNOR2_X1 U9403 ( .A(n7725), .B(n7724), .ZN(n7726) );
  AOI222_X1 U9404 ( .A1(n10111), .A2(n7726), .B1(n8550), .B2(n10108), .C1(
        n8552), .C2(n10107), .ZN(n7863) );
  MUX2_X1 U9405 ( .A(n7727), .B(n7863), .S(n10166), .Z(n7731) );
  XNOR2_X1 U9406 ( .A(n7728), .B(n7729), .ZN(n7861) );
  INV_X1 U9407 ( .A(n8972), .ZN(n8968) );
  AOI22_X1 U9408 ( .A1(n7861), .A2(n8968), .B1(n8967), .B2(n7732), .ZN(n7730)
         );
  NAND2_X1 U9409 ( .A1(n7731), .A2(n7730), .ZN(P2_U3465) );
  INV_X1 U9410 ( .A(n9102), .ZN(n9095) );
  INV_X1 U9411 ( .A(n7732), .ZN(n7856) );
  INV_X1 U9412 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7733) );
  OAI22_X1 U9413 ( .A1(n9100), .A2(n7856), .B1(n10157), .B2(n7733), .ZN(n7734)
         );
  AOI21_X1 U9414 ( .B1(n7861), .B2(n9095), .A(n7734), .ZN(n7735) );
  OAI21_X1 U9415 ( .B1(n7863), .B2(n10159), .A(n7735), .ZN(P2_U3408) );
  NOR2_X1 U9416 ( .A1(n8999), .A2(n8888), .ZN(n10135) );
  AOI21_X1 U9417 ( .B1(n7737), .B2(n7736), .A(n10135), .ZN(n7740) );
  AOI22_X1 U9418 ( .A1(n8925), .A2(n10136), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8924), .ZN(n7739) );
  INV_X1 U9419 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U9420 ( .A1(n10130), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7738) );
  OAI211_X1 U9421 ( .C1(n10130), .C2(n7740), .A(n7739), .B(n7738), .ZN(
        P2_U3233) );
  XNOR2_X1 U9422 ( .A(n7741), .B(n7742), .ZN(n10145) );
  XNOR2_X1 U9423 ( .A(n7743), .B(n7742), .ZN(n7744) );
  AOI222_X1 U9424 ( .A1(n10111), .A2(n7744), .B1(n8552), .B2(n10108), .C1(
        n8996), .C2(n10107), .ZN(n10146) );
  MUX2_X1 U9425 ( .A(n7745), .B(n10146), .S(n10128), .Z(n7747) );
  AOI22_X1 U9426 ( .A1(n8925), .A2(n8458), .B1(n8924), .B2(n8459), .ZN(n7746)
         );
  OAI211_X1 U9427 ( .C1(n8883), .C2(n10145), .A(n7747), .B(n7746), .ZN(
        P2_U3229) );
  NAND2_X1 U9428 ( .A1(n7749), .A2(n7748), .ZN(n7751) );
  INV_X1 U9429 ( .A(n7750), .ZN(n7753) );
  XNOR2_X1 U9430 ( .A(n7751), .B(n7753), .ZN(n7752) );
  INV_X1 U9431 ( .A(n7752), .ZN(n10154) );
  NOR2_X1 U9432 ( .A1(n10130), .A2(n10120), .ZN(n8926) );
  INV_X1 U9433 ( .A(n8926), .ZN(n8047) );
  NAND2_X1 U9434 ( .A1(n7752), .A2(n8990), .ZN(n7759) );
  XNOR2_X1 U9435 ( .A(n7754), .B(n7753), .ZN(n7757) );
  NAND2_X1 U9436 ( .A1(n10107), .A2(n10109), .ZN(n7755) );
  OAI21_X1 U9437 ( .B1(n7772), .B2(n8888), .A(n7755), .ZN(n7756) );
  AOI21_X1 U9438 ( .B1(n7757), .B2(n10111), .A(n7756), .ZN(n7758) );
  NAND2_X1 U9439 ( .A1(n7759), .A2(n7758), .ZN(n10155) );
  MUX2_X1 U9440 ( .A(n10155), .B(P2_REG2_REG_5__SCAN_IN), .S(n10130), .Z(n7760) );
  INV_X1 U9441 ( .A(n7760), .ZN(n7763) );
  AOI22_X1 U9442 ( .A1(n8925), .A2(n7761), .B1(n8924), .B2(n7764), .ZN(n7762)
         );
  OAI211_X1 U9443 ( .C1(n10154), .C2(n8047), .A(n7763), .B(n7762), .ZN(
        P2_U3228) );
  INV_X1 U9444 ( .A(n7764), .ZN(n7778) );
  INV_X1 U9445 ( .A(n7765), .ZN(n8453) );
  INV_X1 U9446 ( .A(n7766), .ZN(n7768) );
  NOR3_X1 U9447 ( .A1(n8453), .A2(n7768), .A3(n7767), .ZN(n7771) );
  INV_X1 U9448 ( .A(n7769), .ZN(n7770) );
  OAI21_X1 U9449 ( .B1(n7771), .B2(n7770), .A(n8500), .ZN(n7776) );
  OAI22_X1 U9450 ( .A1(n8489), .A2(n7772), .B1(n10152), .B2(n8541), .ZN(n7773)
         );
  AOI211_X1 U9451 ( .C1(n8487), .C2(n10109), .A(n7774), .B(n7773), .ZN(n7775)
         );
  OAI211_X1 U9452 ( .C1(n7778), .C2(n7777), .A(n7776), .B(n7775), .ZN(P2_U3167) );
  INV_X1 U9453 ( .A(n7779), .ZN(n7781) );
  INV_X1 U9454 ( .A(n9485), .ZN(n9477) );
  OAI222_X1 U9455 ( .A1(n9940), .A2(n10386), .B1(n9934), .B2(n7781), .C1(n9477), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U9456 ( .A(n8636), .ZN(n8647) );
  OAI222_X1 U9457 ( .A1(n8647), .A2(P2_U3151), .B1(n9132), .B2(n7781), .C1(
        n7780), .C2(n9130), .ZN(P2_U3279) );
  OAI21_X1 U9458 ( .B1(n7782), .B2(n7784), .A(n7783), .ZN(n10009) );
  INV_X1 U9459 ( .A(n10009), .ZN(n7793) );
  XNOR2_X1 U9460 ( .A(n6446), .B(n7784), .ZN(n7785) );
  OAI222_X1 U9461 ( .A1(n10065), .A2(n8049), .B1(n10082), .B2(n9212), .C1(
        n7785), .C2(n9881), .ZN(n10007) );
  NAND2_X1 U9462 ( .A1(n10007), .A2(n9997), .ZN(n7792) );
  OAI22_X1 U9463 ( .A1(n9997), .A2(n7786), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9671), .ZN(n7790) );
  INV_X1 U9464 ( .A(n7874), .ZN(n7787) );
  OAI211_X1 U9465 ( .C1(n10006), .C2(n7788), .A(n7787), .B(n9975), .ZN(n10005)
         );
  NOR2_X1 U9466 ( .A1(n10005), .A2(n9743), .ZN(n7789) );
  AOI211_X1 U9467 ( .C1(n9747), .C2(n7894), .A(n7790), .B(n7789), .ZN(n7791)
         );
  OAI211_X1 U9468 ( .C1(n7793), .C2(n9765), .A(n7792), .B(n7791), .ZN(P1_U3290) );
  XNOR2_X1 U9469 ( .A(n7912), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U9470 ( .A1(n7797), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7798) );
  NAND2_X1 U9471 ( .A1(n7800), .A2(n7806), .ZN(n7914) );
  INV_X1 U9472 ( .A(n7800), .ZN(n7801) );
  INV_X1 U9473 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7804) );
  OAI21_X1 U9474 ( .B1(n5232), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7916), .ZN(
        n7817) );
  INV_X1 U9475 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U9476 ( .A1(n8634), .A2(n7911), .ZN(n7803) );
  NAND2_X1 U9477 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8219) );
  OAI211_X1 U9478 ( .C1(n10275), .C2(n8622), .A(n7803), .B(n8219), .ZN(n7816)
         );
  NAND2_X1 U9479 ( .A1(n7813), .A2(n7812), .ZN(n7810) );
  INV_X1 U9480 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10264) );
  MUX2_X1 U9481 ( .A(n7804), .B(n10264), .S(n4387), .Z(n7805) );
  NAND2_X1 U9482 ( .A1(n7805), .A2(n7911), .ZN(n7927) );
  INV_X1 U9483 ( .A(n7805), .ZN(n7807) );
  NAND2_X1 U9484 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U9485 ( .A1(n7927), .A2(n7808), .ZN(n7811) );
  INV_X1 U9486 ( .A(n7811), .ZN(n7809) );
  NAND2_X1 U9487 ( .A1(n7810), .A2(n7809), .ZN(n7928) );
  NAND3_X1 U9488 ( .A1(n7813), .A2(n7812), .A3(n7811), .ZN(n7814) );
  AOI21_X1 U9489 ( .B1(n7928), .B2(n7814), .A(n8683), .ZN(n7815) );
  AOI211_X1 U9490 ( .C1(n8670), .C2(n7817), .A(n7816), .B(n7815), .ZN(n7818)
         );
  OAI21_X1 U9491 ( .B1(n7819), .B2(n8690), .A(n7818), .ZN(P2_U3191) );
  NAND2_X1 U9492 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  NAND2_X1 U9493 ( .A1(n7820), .A2(n7823), .ZN(n7902) );
  INV_X1 U9494 ( .A(n7902), .ZN(n7831) );
  AOI22_X1 U9495 ( .A1(n10107), .A2(n8551), .B1(n10108), .B2(n8549), .ZN(n7830) );
  NAND2_X1 U9496 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  NAND2_X1 U9497 ( .A1(n7827), .A2(n7826), .ZN(n7828) );
  NAND2_X1 U9498 ( .A1(n7828), .A2(n10111), .ZN(n7829) );
  OAI211_X1 U9499 ( .C1(n7902), .C2(n7945), .A(n7830), .B(n7829), .ZN(n7898)
         );
  AOI21_X1 U9500 ( .B1(n9008), .B2(n7831), .A(n7898), .ZN(n7903) );
  INV_X1 U9501 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10453) );
  OAI22_X1 U9502 ( .A1(n9100), .A2(n7906), .B1(n10157), .B2(n10453), .ZN(n7832) );
  INV_X1 U9503 ( .A(n7832), .ZN(n7833) );
  OAI21_X1 U9504 ( .B1(n7903), .B2(n10159), .A(n7833), .ZN(P2_U3411) );
  OAI211_X1 U9505 ( .C1(n4515), .C2(n7835), .A(n7834), .B(n8500), .ZN(n7842)
         );
  NOR2_X1 U9506 ( .A1(n8541), .A2(n7856), .ZN(n7840) );
  NAND2_X1 U9507 ( .A1(n8533), .A2(n8550), .ZN(n7837) );
  OAI211_X1 U9508 ( .C1(n7838), .C2(n8535), .A(n7837), .B(n7836), .ZN(n7839)
         );
  AOI211_X1 U9509 ( .C1(n7857), .C2(n8538), .A(n7840), .B(n7839), .ZN(n7841)
         );
  NAND2_X1 U9510 ( .A1(n7842), .A2(n7841), .ZN(P2_U3179) );
  XNOR2_X1 U9511 ( .A(n7983), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7845) );
  AOI211_X1 U9512 ( .C1(n7845), .C2(n7844), .A(n9963), .B(n7979), .ZN(n7855)
         );
  INV_X1 U9513 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7846) );
  MUX2_X1 U9514 ( .A(n7846), .B(P1_REG1_REG_10__SCAN_IN), .S(n7983), .Z(n7850)
         );
  AOI211_X1 U9515 ( .C1(n7850), .C2(n7849), .A(n9959), .B(n7982), .ZN(n7854)
         );
  INV_X1 U9516 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7852) );
  NAND2_X1 U9517 ( .A1(n9968), .A2(n7983), .ZN(n7851) );
  NAND2_X1 U9518 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9159) );
  OAI211_X1 U9519 ( .C1(n7852), .C2(n9972), .A(n7851), .B(n9159), .ZN(n7853)
         );
  OR3_X1 U9520 ( .A1(n7855), .A2(n7854), .A3(n7853), .ZN(P1_U3253) );
  INV_X1 U9521 ( .A(n8883), .ZN(n10117) );
  INV_X1 U9522 ( .A(n8880), .ZN(n10115) );
  NOR2_X1 U9523 ( .A1(n10115), .A2(n7856), .ZN(n7860) );
  INV_X1 U9524 ( .A(n7857), .ZN(n7858) );
  OAI22_X1 U9525 ( .A1(n10128), .A2(n7603), .B1(n7858), .B2(n10122), .ZN(n7859) );
  AOI211_X1 U9526 ( .C1(n7861), .C2(n10117), .A(n7860), .B(n7859), .ZN(n7862)
         );
  OAI21_X1 U9527 ( .B1(n7863), .B2(n10130), .A(n7862), .ZN(P2_U3227) );
  INV_X1 U9528 ( .A(n7864), .ZN(n7908) );
  AOI22_X1 U9529 ( .A1(n9499), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9928), .ZN(n7865) );
  OAI21_X1 U9530 ( .B1(n7908), .B2(n9934), .A(n7865), .ZN(P1_U3338) );
  XNOR2_X1 U9531 ( .A(n7867), .B(n7871), .ZN(n10016) );
  NAND2_X1 U9532 ( .A1(n6446), .A2(n7868), .ZN(n7870) );
  NAND2_X1 U9533 ( .A1(n7870), .A2(n7869), .ZN(n7872) );
  XNOR2_X1 U9534 ( .A(n7872), .B(n7871), .ZN(n10018) );
  NAND2_X1 U9535 ( .A1(n10018), .A2(n9729), .ZN(n7880) );
  INV_X1 U9536 ( .A(n9741), .ZN(n7878) );
  OAI22_X1 U9537 ( .A1(n9995), .A2(n9281), .B1(n10011), .B2(n9522), .ZN(n7877)
         );
  OAI211_X1 U9538 ( .C1(n7874), .C2(n9281), .A(n8054), .B(n9975), .ZN(n10014)
         );
  INV_X1 U9539 ( .A(n9671), .ZN(n9991) );
  AOI22_X1 U9540 ( .A1(n9993), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9280), .B2(
        n9991), .ZN(n7875) );
  OAI21_X1 U9541 ( .B1(n10014), .B2(n9743), .A(n7875), .ZN(n7876) );
  AOI211_X1 U9542 ( .C1(n7878), .C2(n7873), .A(n7877), .B(n7876), .ZN(n7879)
         );
  OAI211_X1 U9543 ( .C1(n10016), .C2(n9765), .A(n7880), .B(n7879), .ZN(
        P1_U3289) );
  NAND2_X1 U9544 ( .A1(n7820), .A2(n7881), .ZN(n7882) );
  XOR2_X1 U9545 ( .A(n7882), .B(n7883), .Z(n7949) );
  XNOR2_X1 U9546 ( .A(n7884), .B(n7883), .ZN(n7885) );
  OAI222_X1 U9547 ( .A1(n8998), .A2(n7886), .B1(n8888), .B2(n8369), .C1(n10132), .C2(n7885), .ZN(n7950) );
  AOI21_X1 U9548 ( .B1(n10149), .B2(n7949), .A(n7950), .ZN(n7992) );
  AOI22_X1 U9549 ( .A1(n9094), .A2(n8391), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n10159), .ZN(n7887) );
  OAI21_X1 U9550 ( .B1(n7992), .B2(n10159), .A(n7887), .ZN(P2_U3414) );
  AOI21_X1 U9551 ( .B1(n7890), .B2(n7889), .A(n7888), .ZN(n7897) );
  AOI22_X1 U9552 ( .A1(n9373), .A2(n7891), .B1(n9365), .B2(n9389), .ZN(n7896)
         );
  NAND2_X1 U9553 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9423) );
  INV_X1 U9554 ( .A(n9423), .ZN(n7893) );
  NOR2_X1 U9555 ( .A1(n9349), .A2(n9212), .ZN(n7892) );
  AOI211_X1 U9556 ( .C1(n7894), .C2(n9378), .A(n7893), .B(n7892), .ZN(n7895)
         );
  OAI211_X1 U9557 ( .C1(n7897), .C2(n9380), .A(n7896), .B(n7895), .ZN(P1_U3218) );
  MUX2_X1 U9558 ( .A(n7898), .B(P2_REG2_REG_7__SCAN_IN), .S(n10130), .Z(n7899)
         );
  INV_X1 U9559 ( .A(n7899), .ZN(n7901) );
  AOI22_X1 U9560 ( .A1(n8925), .A2(n7972), .B1(n8924), .B2(n7973), .ZN(n7900)
         );
  OAI211_X1 U9561 ( .C1(n7902), .C2(n8047), .A(n7901), .B(n7900), .ZN(P2_U3226) );
  MUX2_X1 U9562 ( .A(n7904), .B(n7903), .S(n10166), .Z(n7905) );
  OAI21_X1 U9563 ( .B1(n7906), .B2(n8971), .A(n7905), .ZN(P2_U3466) );
  OAI222_X1 U9564 ( .A1(P2_U3151), .A2(n4895), .B1(n9132), .B2(n7908), .C1(
        n7907), .C2(n9130), .ZN(P2_U3278) );
  XNOR2_X1 U9565 ( .A(n8185), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n8182) );
  INV_X1 U9566 ( .A(n7909), .ZN(n7910) );
  XOR2_X1 U9567 ( .A(n8183), .B(n8182), .Z(n7933) );
  INV_X1 U9568 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U9569 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8367) );
  OAI21_X1 U9570 ( .B1(n8622), .B2(n10403), .A(n8367), .ZN(n7919) );
  XNOR2_X1 U9571 ( .A(n8185), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7913) );
  INV_X1 U9572 ( .A(n7913), .ZN(n7915) );
  NAND3_X1 U9573 ( .A1(n7916), .A2(n7915), .A3(n7914), .ZN(n7917) );
  AOI21_X1 U9574 ( .B1(n8187), .B2(n7917), .A(n8717), .ZN(n7918) );
  AOI211_X1 U9575 ( .C1(n8634), .C2(n8185), .A(n7919), .B(n7918), .ZN(n7932)
         );
  NAND2_X1 U9576 ( .A1(n7928), .A2(n7927), .ZN(n7925) );
  INV_X1 U9577 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8184) );
  INV_X1 U9578 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7920) );
  MUX2_X1 U9579 ( .A(n8184), .B(n7920), .S(n4387), .Z(n7921) );
  NAND2_X1 U9580 ( .A1(n7921), .A2(n8185), .ZN(n8198) );
  INV_X1 U9581 ( .A(n7921), .ZN(n7922) );
  NAND2_X1 U9582 ( .A1(n7922), .A2(n8181), .ZN(n7923) );
  NAND2_X1 U9583 ( .A1(n8198), .A2(n7923), .ZN(n7926) );
  INV_X1 U9584 ( .A(n7926), .ZN(n7924) );
  INV_X1 U9585 ( .A(n8199), .ZN(n7930) );
  AND3_X1 U9586 ( .A1(n7928), .A2(n7927), .A3(n7926), .ZN(n7929) );
  OAI21_X1 U9587 ( .B1(n7930), .B2(n7929), .A(n8707), .ZN(n7931) );
  OAI211_X1 U9588 ( .C1(n7933), .C2(n8690), .A(n7932), .B(n7931), .ZN(P2_U3192) );
  INV_X1 U9589 ( .A(n7934), .ZN(n7957) );
  AOI22_X1 U9590 ( .A1(n9967), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9928), .ZN(n7935) );
  OAI21_X1 U9591 ( .B1(n7957), .B2(n9934), .A(n7935), .ZN(P1_U3337) );
  INV_X1 U9592 ( .A(n7936), .ZN(n7938) );
  INV_X1 U9593 ( .A(n7940), .ZN(n7937) );
  NAND2_X1 U9594 ( .A1(n7938), .A2(n7937), .ZN(n8013) );
  NAND2_X1 U9595 ( .A1(n7936), .A2(n7940), .ZN(n7939) );
  NAND2_X1 U9596 ( .A1(n8013), .A2(n7939), .ZN(n8048) );
  INV_X1 U9597 ( .A(n8048), .ZN(n7946) );
  AOI22_X1 U9598 ( .A1(n10108), .A2(n8547), .B1(n10107), .B2(n8549), .ZN(n7944) );
  XNOR2_X1 U9599 ( .A(n7941), .B(n7940), .ZN(n7942) );
  NAND2_X1 U9600 ( .A1(n7942), .A2(n10111), .ZN(n7943) );
  OAI211_X1 U9601 ( .C1(n8048), .C2(n7945), .A(n7944), .B(n7943), .ZN(n8042)
         );
  AOI21_X1 U9602 ( .B1(n9008), .B2(n7946), .A(n8042), .ZN(n8066) );
  OR2_X1 U9603 ( .A1(n9100), .A2(n8218), .ZN(n7948) );
  NAND2_X1 U9604 ( .A1(n10159), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7947) );
  OAI211_X1 U9605 ( .C1(n8066), .C2(n10159), .A(n7948), .B(n7947), .ZN(
        P2_U3417) );
  INV_X1 U9606 ( .A(n7949), .ZN(n7955) );
  INV_X1 U9607 ( .A(n7950), .ZN(n7951) );
  MUX2_X1 U9608 ( .A(n7952), .B(n7951), .S(n10128), .Z(n7954) );
  AOI22_X1 U9609 ( .A1(n8925), .A2(n8391), .B1(n8924), .B2(n8393), .ZN(n7953)
         );
  OAI211_X1 U9610 ( .C1(n7955), .C2(n8883), .A(n7954), .B(n7953), .ZN(P2_U3225) );
  INV_X1 U9611 ( .A(n8709), .ZN(n8698) );
  OAI222_X1 U9612 ( .A1(n8698), .A2(P2_U3151), .B1(n9132), .B2(n7957), .C1(
        n7956), .C2(n9130), .ZN(P2_U3277) );
  NOR2_X1 U9613 ( .A1(n7960), .A2(n5120), .ZN(n7961) );
  XNOR2_X1 U9614 ( .A(n7958), .B(n7961), .ZN(n7967) );
  AOI22_X1 U9615 ( .A1(n9373), .A2(n8005), .B1(n9365), .B2(n9387), .ZN(n7966)
         );
  INV_X1 U9616 ( .A(n7962), .ZN(n7964) );
  NOR2_X1 U9617 ( .A1(n9349), .A2(n6936), .ZN(n7963) );
  AOI211_X1 U9618 ( .C1(n8006), .C2(n9378), .A(n7964), .B(n7963), .ZN(n7965)
         );
  OAI211_X1 U9619 ( .C1(n7967), .C2(n9380), .A(n7966), .B(n7965), .ZN(P1_U3239) );
  INV_X1 U9620 ( .A(n7968), .ZN(n8387) );
  AOI21_X1 U9621 ( .B1(n7970), .B2(n7969), .A(n8387), .ZN(n7978) );
  AOI21_X1 U9622 ( .B1(n8487), .B2(n8551), .A(n7971), .ZN(n7976) );
  AOI22_X1 U9623 ( .A1(n8533), .A2(n8549), .B1(n7972), .B2(n8524), .ZN(n7975)
         );
  NAND2_X1 U9624 ( .A1(n8538), .A2(n7973), .ZN(n7974) );
  AND3_X1 U9625 ( .A1(n7976), .A2(n7975), .A3(n7974), .ZN(n7977) );
  OAI21_X1 U9626 ( .B1(n7978), .B2(n8529), .A(n7977), .ZN(P2_U3153) );
  XNOR2_X1 U9627 ( .A(n8122), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n7980) );
  AOI211_X1 U9628 ( .C1(n7981), .C2(n7980), .A(n9963), .B(n8124), .ZN(n7991)
         );
  INV_X1 U9629 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7984) );
  MUX2_X1 U9630 ( .A(n7984), .B(P1_REG1_REG_11__SCAN_IN), .S(n8122), .Z(n7985)
         );
  AOI211_X1 U9631 ( .C1(n7986), .C2(n7985), .A(n9959), .B(n8117), .ZN(n7990)
         );
  INV_X1 U9632 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U9633 ( .A1(n9968), .A2(n8122), .ZN(n7987) );
  NAND2_X1 U9634 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9329) );
  OAI211_X1 U9635 ( .C1(n7988), .C2(n9972), .A(n7987), .B(n9329), .ZN(n7989)
         );
  OR3_X1 U9636 ( .A1(n7991), .A2(n7990), .A3(n7989), .ZN(P1_U3254) );
  INV_X1 U9637 ( .A(n8391), .ZN(n7994) );
  MUX2_X1 U9638 ( .A(n10293), .B(n7992), .S(n10166), .Z(n7993) );
  OAI21_X1 U9639 ( .B1(n7994), .B2(n8971), .A(n7993), .ZN(P2_U3467) );
  XNOR2_X1 U9640 ( .A(n7995), .B(n8000), .ZN(n7996) );
  OAI222_X1 U9641 ( .A1(n10082), .A2(n6936), .B1(n10065), .B2(n10040), .C1(
        n7996), .C2(n9881), .ZN(n10028) );
  INV_X1 U9642 ( .A(n10028), .ZN(n8011) );
  INV_X1 U9643 ( .A(n7867), .ZN(n7999) );
  OAI21_X1 U9644 ( .B1(n7999), .B2(n7998), .A(n7997), .ZN(n8001) );
  XNOR2_X1 U9645 ( .A(n8000), .B(n8001), .ZN(n10030) );
  INV_X1 U9646 ( .A(n8002), .ZN(n8055) );
  INV_X1 U9647 ( .A(n8003), .ZN(n8004) );
  OAI211_X1 U9648 ( .C1(n10027), .C2(n8002), .A(n8004), .B(n9975), .ZN(n10026)
         );
  AOI22_X1 U9649 ( .A1(n9993), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n8005), .B2(
        n9991), .ZN(n8008) );
  NAND2_X1 U9650 ( .A1(n9747), .A2(n8006), .ZN(n8007) );
  OAI211_X1 U9651 ( .C1(n10026), .C2(n9743), .A(n8008), .B(n8007), .ZN(n8009)
         );
  AOI21_X1 U9652 ( .B1(n10030), .B2(n9704), .A(n8009), .ZN(n8010) );
  OAI21_X1 U9653 ( .B1(n8011), .B2(n9993), .A(n8010), .ZN(P1_U3287) );
  NAND2_X1 U9654 ( .A1(n8013), .A2(n8012), .ZN(n8015) );
  OR2_X1 U9655 ( .A1(n8015), .A2(n8018), .ZN(n8147) );
  NAND2_X1 U9656 ( .A1(n8015), .A2(n8018), .ZN(n8016) );
  NAND2_X1 U9657 ( .A1(n8147), .A2(n8016), .ZN(n8984) );
  INV_X1 U9658 ( .A(n8984), .ZN(n8024) );
  XNOR2_X1 U9659 ( .A(n8017), .B(n8018), .ZN(n8021) );
  NAND2_X1 U9660 ( .A1(n10107), .A2(n8548), .ZN(n8019) );
  OAI21_X1 U9661 ( .B1(n8412), .B2(n8888), .A(n8019), .ZN(n8020) );
  AOI21_X1 U9662 ( .B1(n8021), .B2(n10111), .A(n8020), .ZN(n8985) );
  MUX2_X1 U9663 ( .A(n8184), .B(n8985), .S(n10128), .Z(n8023) );
  AOI22_X1 U9664 ( .A1(n8983), .A2(n8880), .B1(n8924), .B2(n8373), .ZN(n8022)
         );
  OAI211_X1 U9665 ( .C1(n8024), .C2(n8883), .A(n8023), .B(n8022), .ZN(P2_U3223) );
  NAND2_X1 U9666 ( .A1(n7995), .A2(n8025), .ZN(n8027) );
  AOI21_X1 U9667 ( .B1(n8027), .B2(n8026), .A(n8030), .ZN(n8168) );
  AND3_X1 U9668 ( .A1(n8027), .A2(n8026), .A3(n8030), .ZN(n8028) );
  OR2_X1 U9669 ( .A1(n8168), .A2(n8028), .ZN(n8034) );
  INV_X1 U9670 ( .A(n8030), .ZN(n8031) );
  XNOR2_X1 U9671 ( .A(n8029), .B(n8031), .ZN(n8035) );
  AOI22_X1 U9672 ( .A1(n9986), .A2(n10052), .B1(n9388), .B2(n10053), .ZN(n8032) );
  OAI21_X1 U9673 ( .B1(n8035), .B2(n9979), .A(n8032), .ZN(n8033) );
  AOI21_X1 U9674 ( .B1(n8034), .B2(n10061), .A(n8033), .ZN(n10037) );
  INV_X1 U9675 ( .A(n8035), .ZN(n10035) );
  NOR2_X1 U9676 ( .A1(n9993), .A2(n8036), .ZN(n9978) );
  OAI211_X1 U9677 ( .C1(n8003), .C2(n10033), .A(n9975), .B(n8175), .ZN(n10032)
         );
  INV_X1 U9678 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10372) );
  INV_X1 U9679 ( .A(n8037), .ZN(n8109) );
  OAI22_X1 U9680 ( .A1(n9997), .A2(n10372), .B1(n8109), .B2(n9671), .ZN(n8038)
         );
  AOI21_X1 U9681 ( .B1(n9747), .B2(n8113), .A(n8038), .ZN(n8039) );
  OAI21_X1 U9682 ( .B1(n10032), .B2(n9743), .A(n8039), .ZN(n8040) );
  AOI21_X1 U9683 ( .B1(n10035), .B2(n9978), .A(n8040), .ZN(n8041) );
  OAI21_X1 U9684 ( .B1(n10037), .B2(n9993), .A(n8041), .ZN(P1_U3286) );
  MUX2_X1 U9685 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8042), .S(n10128), .Z(n8043)
         );
  INV_X1 U9686 ( .A(n8043), .ZN(n8046) );
  AOI22_X1 U9687 ( .A1(n8880), .A2(n8044), .B1(n8924), .B2(n8224), .ZN(n8045)
         );
  OAI211_X1 U9688 ( .C1(n8048), .C2(n8047), .A(n8046), .B(n8045), .ZN(P2_U3224) );
  OAI21_X1 U9689 ( .B1(n7867), .B2(n9281), .A(n8049), .ZN(n8051) );
  NAND2_X1 U9690 ( .A1(n7867), .A2(n9281), .ZN(n8050) );
  NAND2_X1 U9691 ( .A1(n8051), .A2(n8050), .ZN(n8052) );
  XNOR2_X1 U9692 ( .A(n8053), .B(n8052), .ZN(n10019) );
  AOI21_X1 U9693 ( .B1(n8054), .B2(n4394), .A(n9768), .ZN(n8056) );
  NAND2_X1 U9694 ( .A1(n8056), .A2(n8055), .ZN(n10020) );
  AOI22_X1 U9695 ( .A1(n9747), .A2(n4394), .B1(n9991), .B2(n8076), .ZN(n8057)
         );
  OAI21_X1 U9696 ( .B1(n10020), .B2(n9743), .A(n8057), .ZN(n8064) );
  XNOR2_X1 U9697 ( .A(n8058), .B(n8059), .ZN(n8060) );
  NAND2_X1 U9698 ( .A1(n8060), .A2(n10061), .ZN(n8062) );
  AOI22_X1 U9699 ( .A1(n9986), .A2(n9388), .B1(n9389), .B2(n10053), .ZN(n8061)
         );
  NAND2_X1 U9700 ( .A1(n8062), .A2(n8061), .ZN(n10024) );
  MUX2_X1 U9701 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10024), .S(n9997), .Z(n8063)
         );
  AOI211_X1 U9702 ( .C1(n9704), .C2(n10019), .A(n8064), .B(n8063), .ZN(n8065)
         );
  INV_X1 U9703 ( .A(n8065), .ZN(P1_U3288) );
  MUX2_X1 U9704 ( .A(n10264), .B(n8066), .S(n10166), .Z(n8067) );
  OAI21_X1 U9705 ( .B1(n8218), .B2(n8971), .A(n8067), .ZN(P2_U3468) );
  INV_X1 U9706 ( .A(n8068), .ZN(n9277) );
  XNOR2_X1 U9707 ( .A(n8070), .B(n8069), .ZN(n9276) );
  NOR3_X1 U9708 ( .A1(n7888), .A2(n9277), .A3(n9276), .ZN(n9275) );
  NOR2_X1 U9709 ( .A1(n9275), .A2(n8071), .ZN(n8075) );
  XNOR2_X1 U9710 ( .A(n8073), .B(n8072), .ZN(n8074) );
  XNOR2_X1 U9711 ( .A(n8075), .B(n8074), .ZN(n8081) );
  AOI22_X1 U9712 ( .A1(n8076), .A2(n9373), .B1(n9372), .B2(n9389), .ZN(n8080)
         );
  OAI21_X1 U9713 ( .B1(n9376), .B2(n8108), .A(n8077), .ZN(n8078) );
  AOI21_X1 U9714 ( .B1(n4394), .B2(n9378), .A(n8078), .ZN(n8079) );
  OAI211_X1 U9715 ( .C1(n8081), .C2(n9380), .A(n8080), .B(n8079), .ZN(P1_U3227) );
  NOR2_X1 U9716 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8100) );
  NOR2_X1 U9717 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8098) );
  NOR2_X1 U9718 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8096) );
  NOR2_X1 U9719 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10196) );
  NOR2_X1 U9720 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8082) );
  AOI21_X1 U9721 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8082), .ZN(n10185) );
  NOR2_X1 U9722 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8083) );
  AOI21_X1 U9723 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8083), .ZN(n10188) );
  NOR2_X1 U9724 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8084) );
  AOI21_X1 U9725 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8084), .ZN(n10191) );
  NOR2_X1 U9726 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8085) );
  AOI21_X1 U9727 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8085), .ZN(n10194) );
  NOR2_X1 U9728 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8086) );
  AOI21_X1 U9729 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n8086), .ZN(n10518) );
  NOR2_X1 U9730 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8087) );
  AOI21_X1 U9731 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n8087), .ZN(n10521) );
  NOR2_X1 U9732 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n8088) );
  AOI21_X1 U9733 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n8088), .ZN(n10524) );
  NOR2_X1 U9734 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n8089) );
  AOI21_X1 U9735 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n8089), .ZN(n10509) );
  NOR2_X1 U9736 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8090) );
  AOI21_X1 U9737 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n8090), .ZN(n10512) );
  INV_X1 U9738 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10173) );
  NOR2_X1 U9739 ( .A1(n10212), .A2(n10173), .ZN(n10172) );
  NOR2_X1 U9740 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10172), .ZN(n10168) );
  INV_X1 U9741 ( .A(n10168), .ZN(n10169) );
  NAND3_X1 U9742 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10170) );
  NAND2_X1 U9743 ( .A1(n10171), .A2(n10170), .ZN(n10167) );
  NAND2_X1 U9744 ( .A1(n10169), .A2(n10167), .ZN(n10515) );
  NAND2_X1 U9745 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n8091) );
  OAI21_X1 U9746 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n8091), .ZN(n10514) );
  NOR2_X1 U9747 ( .A1(n10515), .A2(n10514), .ZN(n10513) );
  AOI21_X1 U9748 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10513), .ZN(n10527) );
  NAND2_X1 U9749 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8092) );
  OAI21_X1 U9750 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n8092), .ZN(n10526) );
  NOR2_X1 U9751 ( .A1(n10527), .A2(n10526), .ZN(n10525) );
  AOI21_X1 U9752 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10525), .ZN(n10530) );
  NOR2_X1 U9753 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8093) );
  AOI21_X1 U9754 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n8093), .ZN(n10529) );
  NAND2_X1 U9755 ( .A1(n10530), .A2(n10529), .ZN(n10528) );
  OAI21_X1 U9756 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10528), .ZN(n10511) );
  NAND2_X1 U9757 ( .A1(n10512), .A2(n10511), .ZN(n10510) );
  OAI21_X1 U9758 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10510), .ZN(n10508) );
  NAND2_X1 U9759 ( .A1(n10509), .A2(n10508), .ZN(n10507) );
  OAI21_X1 U9760 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10507), .ZN(n10523) );
  NAND2_X1 U9761 ( .A1(n10524), .A2(n10523), .ZN(n10522) );
  OAI21_X1 U9762 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10522), .ZN(n10520) );
  NAND2_X1 U9763 ( .A1(n10521), .A2(n10520), .ZN(n10519) );
  OAI21_X1 U9764 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10519), .ZN(n10517) );
  NAND2_X1 U9765 ( .A1(n10518), .A2(n10517), .ZN(n10516) );
  OAI21_X1 U9766 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10516), .ZN(n10193) );
  NAND2_X1 U9767 ( .A1(n10194), .A2(n10193), .ZN(n10192) );
  OAI21_X1 U9768 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10192), .ZN(n10190) );
  NAND2_X1 U9769 ( .A1(n10191), .A2(n10190), .ZN(n10189) );
  OAI21_X1 U9770 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10189), .ZN(n10187) );
  NAND2_X1 U9771 ( .A1(n10188), .A2(n10187), .ZN(n10186) );
  OAI21_X1 U9772 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10186), .ZN(n10184) );
  NAND2_X1 U9773 ( .A1(n10185), .A2(n10184), .ZN(n10183) );
  OAI21_X1 U9774 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10183), .ZN(n10505) );
  INV_X1 U9775 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10237) );
  INV_X1 U9776 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9458) );
  NOR2_X1 U9777 ( .A1(n10237), .A2(n9458), .ZN(n10195) );
  INV_X1 U9778 ( .A(n10195), .ZN(n8094) );
  OAI21_X1 U9779 ( .B1(n10196), .B2(n10505), .A(n8094), .ZN(n10182) );
  INV_X1 U9780 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9957) );
  INV_X1 U9781 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U9782 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9957), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10464), .ZN(n10181) );
  NOR2_X1 U9783 ( .A1(n10182), .A2(n10181), .ZN(n8095) );
  NOR2_X1 U9784 ( .A1(n8096), .A2(n8095), .ZN(n10180) );
  XNOR2_X1 U9785 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10179) );
  NOR2_X1 U9786 ( .A1(n10180), .A2(n10179), .ZN(n8097) );
  NOR2_X1 U9787 ( .A1(n8098), .A2(n8097), .ZN(n10178) );
  INV_X1 U9788 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10487) );
  XOR2_X1 U9789 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n10487), .Z(n10177) );
  NOR2_X1 U9790 ( .A1(n10178), .A2(n10177), .ZN(n8099) );
  NOR2_X1 U9791 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  AND2_X1 U9792 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8101), .ZN(n10174) );
  NOR2_X1 U9793 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10174), .ZN(n8102) );
  NOR2_X1 U9794 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8101), .ZN(n10175) );
  NOR2_X1 U9795 ( .A1(n8102), .A2(n10175), .ZN(n8104) );
  XNOR2_X1 U9796 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8103) );
  XNOR2_X1 U9797 ( .A(n8104), .B(n8103), .ZN(ADD_1068_U4) );
  XNOR2_X1 U9798 ( .A(n8106), .B(n5122), .ZN(n8107) );
  XNOR2_X1 U9799 ( .A(n8105), .B(n8107), .ZN(n8115) );
  OAI22_X1 U9800 ( .A1(n9350), .A2(n8109), .B1(n9349), .B2(n8108), .ZN(n8112)
         );
  OAI21_X1 U9801 ( .B1(n9376), .B2(n9294), .A(n8110), .ZN(n8111) );
  AOI211_X1 U9802 ( .C1(n8113), .C2(n9378), .A(n8112), .B(n8111), .ZN(n8114)
         );
  OAI21_X1 U9803 ( .B1(n8115), .B2(n9380), .A(n8114), .ZN(P1_U3213) );
  INV_X1 U9804 ( .A(n8116), .ZN(n8209) );
  OAI222_X1 U9805 ( .A1(n9940), .A2(n10371), .B1(n9943), .B2(n8209), .C1(n5846), .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U9806 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8118) );
  MUX2_X1 U9807 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n8118), .S(n8297), .Z(n8119)
         );
  OAI21_X1 U9808 ( .B1(n8120), .B2(n8119), .A(n8296), .ZN(n8121) );
  INV_X1 U9809 ( .A(n8121), .ZN(n8132) );
  XOR2_X1 U9810 ( .A(n8297), .B(P1_REG2_REG_12__SCAN_IN), .Z(n8126) );
  OAI21_X1 U9811 ( .B1(n8126), .B2(n8125), .A(n8293), .ZN(n8130) );
  INV_X1 U9812 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U9813 ( .A1(n9968), .A2(n8297), .ZN(n8127) );
  NAND2_X1 U9814 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9227) );
  OAI211_X1 U9815 ( .C1(n8128), .C2(n9972), .A(n8127), .B(n9227), .ZN(n8129)
         );
  AOI21_X1 U9816 ( .B1(n8130), .B2(n9496), .A(n8129), .ZN(n8131) );
  OAI21_X1 U9817 ( .B1(n8132), .B2(n9959), .A(n8131), .ZN(P1_U3255) );
  XOR2_X1 U9818 ( .A(n8133), .B(n8142), .Z(n10058) );
  AOI22_X1 U9819 ( .A1(n9993), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9292), .B2(
        n9991), .ZN(n8134) );
  OAI21_X1 U9820 ( .B1(n9294), .B2(n9522), .A(n8134), .ZN(n8138) );
  AOI211_X1 U9821 ( .C1(n10054), .C2(n8135), .A(n9768), .B(n4495), .ZN(n8136)
         );
  AOI21_X1 U9822 ( .B1(n9986), .B2(n9987), .A(n8136), .ZN(n10056) );
  NOR2_X1 U9823 ( .A1(n10056), .A2(n9743), .ZN(n8137) );
  AOI211_X1 U9824 ( .C1(n9747), .C2(n10054), .A(n8138), .B(n8137), .ZN(n8145)
         );
  INV_X1 U9825 ( .A(n8139), .ZN(n8141) );
  OAI21_X1 U9826 ( .B1(n8168), .B2(n8141), .A(n8140), .ZN(n8143) );
  XNOR2_X1 U9827 ( .A(n8143), .B(n8142), .ZN(n10060) );
  NAND2_X1 U9828 ( .A1(n10060), .A2(n9729), .ZN(n8144) );
  OAI211_X1 U9829 ( .C1(n10058), .C2(n9765), .A(n8145), .B(n8144), .ZN(
        P1_U3284) );
  NAND2_X1 U9830 ( .A1(n8147), .A2(n8146), .ZN(n8149) );
  XNOR2_X1 U9831 ( .A(n8149), .B(n8148), .ZN(n8979) );
  INV_X1 U9832 ( .A(n8979), .ZN(n8155) );
  INV_X1 U9833 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8191) );
  XNOR2_X1 U9834 ( .A(n8151), .B(n8150), .ZN(n8152) );
  AOI222_X1 U9835 ( .A1(n10111), .A2(n8152), .B1(n8904), .B2(n10108), .C1(
        n8547), .C2(n10107), .ZN(n8981) );
  MUX2_X1 U9836 ( .A(n8191), .B(n8981), .S(n10128), .Z(n8154) );
  AOI22_X1 U9837 ( .A1(n8494), .A2(n8925), .B1(n8924), .B2(n8506), .ZN(n8153)
         );
  OAI211_X1 U9838 ( .C1(n8155), .C2(n8883), .A(n8154), .B(n8153), .ZN(P2_U3222) );
  XNOR2_X1 U9839 ( .A(n8156), .B(n6406), .ZN(n8157) );
  AOI222_X1 U9840 ( .A1(n10111), .A2(n8157), .B1(n8545), .B2(n10108), .C1(
        n8546), .C2(n10107), .ZN(n8977) );
  INV_X1 U9841 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8257) );
  INV_X1 U9842 ( .A(n8415), .ZN(n8158) );
  OAI22_X1 U9843 ( .A1(n10128), .A2(n8257), .B1(n8158), .B2(n10122), .ZN(n8159) );
  AOI21_X1 U9844 ( .B1(n8160), .B2(n8880), .A(n8159), .ZN(n8165) );
  NAND2_X1 U9845 ( .A1(n8162), .A2(n8163), .ZN(n8975) );
  NAND3_X1 U9846 ( .A1(n8161), .A2(n8975), .A3(n10117), .ZN(n8164) );
  OAI211_X1 U9847 ( .C1(n8977), .C2(n10130), .A(n8165), .B(n8164), .ZN(
        P2_U3221) );
  XOR2_X1 U9848 ( .A(n8167), .B(n8171), .Z(n10046) );
  INV_X1 U9849 ( .A(n8168), .ZN(n8170) );
  NAND2_X1 U9850 ( .A1(n8170), .A2(n8169), .ZN(n8172) );
  XNOR2_X1 U9851 ( .A(n8172), .B(n8171), .ZN(n8173) );
  NOR2_X1 U9852 ( .A1(n8173), .A2(n9881), .ZN(n10048) );
  NAND2_X1 U9853 ( .A1(n10048), .A2(n9997), .ZN(n8180) );
  INV_X1 U9854 ( .A(n8135), .ZN(n8174) );
  AOI211_X1 U9855 ( .C1(n10043), .C2(n8175), .A(n9768), .B(n8174), .ZN(n10041)
         );
  AOI22_X1 U9856 ( .A1(n9993), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9199), .B2(
        n9991), .ZN(n8176) );
  OAI21_X1 U9857 ( .B1(n9995), .B2(n9204), .A(n8176), .ZN(n8178) );
  OAI22_X1 U9858 ( .A1(n10040), .A2(n9522), .B1(n9741), .B2(n10039), .ZN(n8177) );
  AOI211_X1 U9859 ( .C1(n10041), .C2(n9977), .A(n8178), .B(n8177), .ZN(n8179)
         );
  OAI211_X1 U9860 ( .C1(n10046), .C2(n9765), .A(n8180), .B(n8179), .ZN(
        P1_U3285) );
  XNOR2_X1 U9861 ( .A(n8244), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n8207) );
  OR2_X1 U9862 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  OAI21_X1 U9863 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n8190), .A(n8260), .ZN(
        n8205) );
  NAND2_X1 U9864 ( .A1(n8199), .A2(n8198), .ZN(n8196) );
  INV_X1 U9865 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10343) );
  MUX2_X1 U9866 ( .A(n8191), .B(n10343), .S(n4387), .Z(n8192) );
  NAND2_X1 U9867 ( .A1(n8192), .A2(n8243), .ZN(n8252) );
  INV_X1 U9868 ( .A(n8192), .ZN(n8193) );
  NAND2_X1 U9869 ( .A1(n8193), .A2(n8202), .ZN(n8194) );
  NAND2_X1 U9870 ( .A1(n8252), .A2(n8194), .ZN(n8197) );
  INV_X1 U9871 ( .A(n8197), .ZN(n8195) );
  NAND3_X1 U9872 ( .A1(n8199), .A2(n8198), .A3(n8197), .ZN(n8200) );
  AOI21_X1 U9873 ( .B1(n8253), .B2(n8200), .A(n8683), .ZN(n8204) );
  NAND2_X1 U9874 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U9875 ( .A1(n8701), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n8201) );
  OAI211_X1 U9876 ( .C1(n8705), .C2(n8202), .A(n8502), .B(n8201), .ZN(n8203)
         );
  AOI211_X1 U9877 ( .C1(n8205), .C2(n8670), .A(n8204), .B(n8203), .ZN(n8206)
         );
  OAI21_X1 U9878 ( .B1(n8207), .B2(n8690), .A(n8206), .ZN(P2_U3193) );
  OAI222_X1 U9879 ( .A1(P2_U3151), .A2(n8704), .B1(n9132), .B2(n8209), .C1(
        n8208), .C2(n9130), .ZN(P2_U3276) );
  INV_X1 U9880 ( .A(n8210), .ZN(n8214) );
  OAI222_X1 U9881 ( .A1(n8212), .A2(P1_U3086), .B1(n9934), .B2(n8214), .C1(
        n8211), .C2(n9940), .ZN(P1_U3335) );
  OAI222_X1 U9882 ( .A1(P2_U3151), .A2(n8215), .B1(n9132), .B2(n8214), .C1(
        n8213), .C2(n9130), .ZN(P2_U3275) );
  OAI211_X1 U9883 ( .C1(n4504), .C2(n8217), .A(n8216), .B(n8500), .ZN(n8226)
         );
  NOR2_X1 U9884 ( .A1(n8541), .A2(n8218), .ZN(n8223) );
  NAND2_X1 U9885 ( .A1(n8533), .A2(n8547), .ZN(n8220) );
  OAI211_X1 U9886 ( .C1(n8221), .C2(n8535), .A(n8220), .B(n8219), .ZN(n8222)
         );
  AOI211_X1 U9887 ( .C1(n8224), .C2(n8538), .A(n8223), .B(n8222), .ZN(n8225)
         );
  NAND2_X1 U9888 ( .A1(n8226), .A2(n8225), .ZN(P2_U3171) );
  XNOR2_X1 U9889 ( .A(n8227), .B(n8230), .ZN(n10068) );
  INV_X1 U9890 ( .A(n10068), .ZN(n8241) );
  INV_X1 U9891 ( .A(n8228), .ZN(n8229) );
  AOI21_X1 U9892 ( .B1(n8231), .B2(n8230), .A(n8229), .ZN(n8232) );
  OAI22_X1 U9893 ( .A1(n8232), .A2(n9881), .B1(n10039), .B2(n10082), .ZN(
        n10066) );
  INV_X1 U9894 ( .A(n8233), .ZN(n8234) );
  OAI211_X1 U9895 ( .C1(n8235), .C2(n4495), .A(n8234), .B(n9975), .ZN(n10064)
         );
  AOI22_X1 U9896 ( .A1(n9993), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9158), .B2(
        n9991), .ZN(n8236) );
  OAI21_X1 U9897 ( .B1(n10083), .B2(n9741), .A(n8236), .ZN(n8237) );
  AOI21_X1 U9898 ( .B1(n9747), .B2(n10062), .A(n8237), .ZN(n8238) );
  OAI21_X1 U9899 ( .B1(n10064), .B2(n9743), .A(n8238), .ZN(n8239) );
  AOI21_X1 U9900 ( .B1(n10066), .B2(n9997), .A(n8239), .ZN(n8240) );
  OAI21_X1 U9901 ( .B1(n8241), .B2(n9765), .A(n8240), .ZN(P1_U3283) );
  XNOR2_X1 U9902 ( .A(n8258), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8553) );
  XOR2_X1 U9903 ( .A(n8553), .B(n4503), .Z(n8264) );
  INV_X1 U9904 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U9905 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8410) );
  OAI21_X1 U9906 ( .B1(n8622), .B2(n8245), .A(n8410), .ZN(n8256) );
  NAND2_X1 U9907 ( .A1(n8253), .A2(n8252), .ZN(n8250) );
  INV_X1 U9908 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10448) );
  MUX2_X1 U9909 ( .A(n8257), .B(n10448), .S(n4387), .Z(n8246) );
  NAND2_X1 U9910 ( .A1(n8246), .A2(n8258), .ZN(n8561) );
  INV_X1 U9911 ( .A(n8246), .ZN(n8247) );
  NAND2_X1 U9912 ( .A1(n8247), .A2(n8554), .ZN(n8248) );
  NAND2_X1 U9913 ( .A1(n8561), .A2(n8248), .ZN(n8251) );
  INV_X1 U9914 ( .A(n8251), .ZN(n8249) );
  NAND3_X1 U9915 ( .A1(n8253), .A2(n8252), .A3(n8251), .ZN(n8254) );
  AOI21_X1 U9916 ( .B1(n8562), .B2(n8254), .A(n8683), .ZN(n8255) );
  AOI211_X1 U9917 ( .C1(n8634), .C2(n8258), .A(n8256), .B(n8255), .ZN(n8263)
         );
  XNOR2_X1 U9918 ( .A(n8258), .B(n8257), .ZN(n8259) );
  AND3_X1 U9919 ( .A1(n8260), .A2(n8259), .A3(n5231), .ZN(n8261) );
  OAI21_X1 U9920 ( .B1(n4506), .B2(n8261), .A(n8670), .ZN(n8262) );
  OAI211_X1 U9921 ( .C1(n8264), .C2(n8690), .A(n8263), .B(n8262), .ZN(P2_U3194) );
  INV_X1 U9922 ( .A(n8265), .ZN(n8268) );
  OAI222_X1 U9923 ( .A1(n8266), .A2(P2_U3151), .B1(n9132), .B2(n8268), .C1(
        n10438), .C2(n9130), .ZN(P2_U3274) );
  OAI222_X1 U9924 ( .A1(n8269), .A2(P1_U3086), .B1(n9934), .B2(n8268), .C1(
        n8267), .C2(n9940), .ZN(P1_U3334) );
  INV_X1 U9925 ( .A(n8270), .ZN(n8274) );
  OAI222_X1 U9926 ( .A1(P2_U3151), .A2(n8272), .B1(n9132), .B2(n8274), .C1(
        n8271), .C2(n9130), .ZN(P2_U3273) );
  OAI222_X1 U9927 ( .A1(n9940), .A2(n8275), .B1(n9934), .B2(n8274), .C1(n8273), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  XNOR2_X1 U9928 ( .A(n8276), .B(n8277), .ZN(n10086) );
  INV_X1 U9929 ( .A(n10086), .ZN(n8289) );
  XNOR2_X1 U9930 ( .A(n8279), .B(n8278), .ZN(n8280) );
  OAI22_X1 U9931 ( .A1(n8280), .A2(n9881), .B1(n9139), .B2(n10065), .ZN(n10084) );
  INV_X1 U9932 ( .A(n9974), .ZN(n8283) );
  OAI211_X1 U9933 ( .C1(n8283), .C2(n8282), .A(n9975), .B(n9759), .ZN(n10081)
         );
  AOI22_X1 U9934 ( .A1(n9993), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9226), .B2(
        n9991), .ZN(n8284) );
  OAI21_X1 U9935 ( .B1(n10083), .B2(n9522), .A(n8284), .ZN(n8285) );
  AOI21_X1 U9936 ( .B1(n10079), .B2(n9747), .A(n8285), .ZN(n8286) );
  OAI21_X1 U9937 ( .B1(n10081), .B2(n9743), .A(n8286), .ZN(n8287) );
  AOI21_X1 U9938 ( .B1(n10084), .B2(n9997), .A(n8287), .ZN(n8288) );
  OAI21_X1 U9939 ( .B1(n8289), .B2(n9765), .A(n8288), .ZN(P1_U3281) );
  INV_X1 U9940 ( .A(n8306), .ZN(n8292) );
  NAND2_X1 U9941 ( .A1(n9121), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8290) );
  OAI211_X1 U9942 ( .C1(n8292), .C2(n9132), .A(n8291), .B(n8290), .ZN(P2_U3272) );
  XNOR2_X1 U9943 ( .A(n9453), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n8295) );
  AOI211_X1 U9944 ( .C1(n8295), .C2(n8294), .A(n9963), .B(n4416), .ZN(n8304)
         );
  XNOR2_X1 U9945 ( .A(n9453), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n8299) );
  AOI211_X1 U9946 ( .C1(n8299), .C2(n8298), .A(n9959), .B(n9452), .ZN(n8303)
         );
  INV_X1 U9947 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U9948 ( .A1(n9968), .A2(n9453), .ZN(n8300) );
  NAND2_X1 U9949 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9308) );
  OAI211_X1 U9950 ( .C1(n8301), .C2(n9972), .A(n8300), .B(n9308), .ZN(n8302)
         );
  OR3_X1 U9951 ( .A1(n8304), .A2(n8303), .A3(n8302), .ZN(P1_U3256) );
  NAND2_X1 U9952 ( .A1(n8306), .A2(n8305), .ZN(n8308) );
  OAI211_X1 U9953 ( .C1(n8309), .C2(n9940), .A(n8308), .B(n8307), .ZN(P1_U3332) );
  INV_X1 U9954 ( .A(n8310), .ZN(n8314) );
  OAI222_X1 U9955 ( .A1(n8312), .A2(P2_U3151), .B1(n9132), .B2(n8314), .C1(
        n8311), .C2(n9130), .ZN(P2_U3271) );
  OAI222_X1 U9956 ( .A1(n8315), .A2(P1_U3086), .B1(n9934), .B2(n8314), .C1(
        n8313), .C2(n9940), .ZN(P1_U3331) );
  INV_X1 U9957 ( .A(n8316), .ZN(n9123) );
  OAI222_X1 U9958 ( .A1(n9940), .A2(n8318), .B1(P1_U3086), .B2(n8317), .C1(
        n9934), .C2(n9123), .ZN(P1_U3327) );
  INV_X1 U9959 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8323) );
  NAND4_X1 U9960 ( .A1(n9997), .A2(n8321), .A3(n8320), .A4(n8319), .ZN(n8322)
         );
  OAI21_X1 U9961 ( .B1(n9671), .B2(n8323), .A(n8322), .ZN(n8324) );
  AOI21_X1 U9962 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n9993), .A(n8324), .ZN(
        n8328) );
  NAND2_X1 U9963 ( .A1(n9977), .A2(n9975), .ZN(n9514) );
  INV_X1 U9964 ( .A(n9514), .ZN(n8326) );
  OAI21_X1 U9965 ( .B1(n8326), .B2(n9747), .A(n8325), .ZN(n8327) );
  OAI211_X1 U9966 ( .C1(n4648), .C2(n9741), .A(n8328), .B(n8327), .ZN(P1_U3293) );
  AOI22_X1 U9967 ( .A1(n8330), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9928), .ZN(n8331) );
  OAI21_X1 U9968 ( .B1(n8332), .B2(n9934), .A(n8331), .ZN(P1_U3350) );
  NOR2_X1 U9969 ( .A1(n8334), .A2(n10122), .ZN(n8721) );
  AOI21_X1 U9970 ( .B1(n10130), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8721), .ZN(
        n8335) );
  OAI21_X1 U9971 ( .B1(n8336), .B2(n10115), .A(n8335), .ZN(n8337) );
  AOI21_X1 U9972 ( .B1(n8333), .B2(n8926), .A(n8337), .ZN(n8338) );
  INV_X1 U9973 ( .A(n8339), .ZN(n9116) );
  OAI222_X1 U9974 ( .A1(n9940), .A2(n8341), .B1(n9934), .B2(n9116), .C1(n8340), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  INV_X1 U9975 ( .A(n8342), .ZN(n8350) );
  OAI21_X1 U9976 ( .B1(n8344), .B2(n8343), .A(n8500), .ZN(n8349) );
  NAND2_X1 U9977 ( .A1(n8730), .A2(n8533), .ZN(n8346) );
  AOI22_X1 U9978 ( .A1(n8732), .A2(n8538), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8345) );
  OAI211_X1 U9979 ( .C1(n8422), .C2(n8535), .A(n8346), .B(n8345), .ZN(n8347)
         );
  AOI21_X1 U9980 ( .B1(n9021), .B2(n8524), .A(n8347), .ZN(n8348) );
  OAI21_X1 U9981 ( .B1(n8350), .B2(n8349), .A(n8348), .ZN(P2_U3154) );
  INV_X1 U9982 ( .A(n9093), .ZN(n8884) );
  OAI21_X1 U9983 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8354) );
  NAND2_X1 U9984 ( .A1(n8354), .A2(n8500), .ZN(n8358) );
  NAND2_X1 U9985 ( .A1(n8533), .A2(n8544), .ZN(n8355) );
  NAND2_X1 U9986 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8575) );
  OAI211_X1 U9987 ( .C1(n8887), .C2(n8535), .A(n8355), .B(n8575), .ZN(n8356)
         );
  AOI21_X1 U9988 ( .B1(n8895), .B2(n8538), .A(n8356), .ZN(n8357) );
  OAI211_X1 U9989 ( .C1(n8884), .C2(n8541), .A(n8358), .B(n8357), .ZN(P2_U3155) );
  XNOR2_X1 U9990 ( .A(n8444), .B(n8761), .ZN(n8363) );
  AOI22_X1 U9991 ( .A1(n8802), .A2(n8487), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8360) );
  NAND2_X1 U9992 ( .A1(n8781), .A2(n8538), .ZN(n8359) );
  OAI211_X1 U9993 ( .C1(n8778), .C2(n8489), .A(n8360), .B(n8359), .ZN(n8361)
         );
  AOI21_X1 U9994 ( .B1(n6416), .B2(n8524), .A(n8361), .ZN(n8362) );
  OAI21_X1 U9995 ( .B1(n8363), .B2(n8529), .A(n8362), .ZN(P2_U3156) );
  XNOR2_X1 U9996 ( .A(n8364), .B(n8547), .ZN(n8365) );
  NOR2_X1 U9997 ( .A1(n8365), .A2(n8366), .ZN(n8498) );
  AOI21_X1 U9998 ( .B1(n8366), .B2(n8365), .A(n8498), .ZN(n8375) );
  NAND2_X1 U9999 ( .A1(n8533), .A2(n8546), .ZN(n8368) );
  OAI211_X1 U10000 ( .C1(n8369), .C2(n8535), .A(n8368), .B(n8367), .ZN(n8372)
         );
  NOR2_X1 U10001 ( .A1(n8370), .A2(n8541), .ZN(n8371) );
  AOI211_X1 U10002 ( .C1(n8373), .C2(n8538), .A(n8372), .B(n8371), .ZN(n8374)
         );
  OAI21_X1 U10003 ( .B1(n8375), .B2(n8529), .A(n8374), .ZN(P2_U3157) );
  OAI211_X1 U10004 ( .C1(n8378), .C2(n8377), .A(n8376), .B(n8500), .ZN(n8382)
         );
  NAND2_X1 U10005 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U10006 ( .A1(n8849), .A2(n8487), .ZN(n8379) );
  OAI211_X1 U10007 ( .C1(n8402), .C2(n8489), .A(n8703), .B(n8379), .ZN(n8380)
         );
  AOI21_X1 U10008 ( .B1(n8827), .B2(n8538), .A(n8380), .ZN(n8381) );
  OAI211_X1 U10009 ( .C1(n8383), .C2(n8541), .A(n8382), .B(n8381), .ZN(
        P2_U3159) );
  INV_X1 U10010 ( .A(n8384), .ZN(n8386) );
  NOR3_X1 U10011 ( .A1(n8387), .A2(n8386), .A3(n8385), .ZN(n8390) );
  INV_X1 U10012 ( .A(n8388), .ZN(n8389) );
  OAI21_X1 U10013 ( .B1(n8390), .B2(n8389), .A(n8500), .ZN(n8397) );
  AOI22_X1 U10014 ( .A1(n8533), .A2(n8548), .B1(n8391), .B2(n8524), .ZN(n8396)
         );
  AOI21_X1 U10015 ( .B1(n8487), .B2(n8550), .A(n8392), .ZN(n8395) );
  NAND2_X1 U10016 ( .A1(n8538), .A2(n8393), .ZN(n8394) );
  NAND4_X1 U10017 ( .A1(n8397), .A2(n8396), .A3(n8395), .A4(n8394), .ZN(
        P2_U3161) );
  XOR2_X1 U10018 ( .A(n8399), .B(n8398), .Z(n8405) );
  AOI22_X1 U10019 ( .A1(n8802), .A2(n8533), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8401) );
  NAND2_X1 U10020 ( .A1(n8805), .A2(n8538), .ZN(n8400) );
  OAI211_X1 U10021 ( .C1(n8402), .C2(n8535), .A(n8401), .B(n8400), .ZN(n8403)
         );
  AOI21_X1 U10022 ( .B1(n9056), .B2(n8524), .A(n8403), .ZN(n8404) );
  OAI21_X1 U10023 ( .B1(n8405), .B2(n8529), .A(n8404), .ZN(P2_U3163) );
  NOR2_X1 U10024 ( .A1(n8364), .A2(n8547), .ZN(n8497) );
  NOR3_X1 U10025 ( .A1(n8498), .A2(n8497), .A3(n8496), .ZN(n8495) );
  AOI21_X1 U10026 ( .B1(n8546), .B2(n8496), .A(n8495), .ZN(n8409) );
  NAND2_X1 U10027 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  XNOR2_X1 U10028 ( .A(n8409), .B(n8408), .ZN(n8417) );
  NAND2_X1 U10029 ( .A1(n8533), .A2(n8545), .ZN(n8411) );
  OAI211_X1 U10030 ( .C1(n8412), .C2(n8535), .A(n8411), .B(n8410), .ZN(n8414)
         );
  NOR2_X1 U10031 ( .A1(n8978), .A2(n8541), .ZN(n8413) );
  AOI211_X1 U10032 ( .C1(n8415), .C2(n8538), .A(n8414), .B(n8413), .ZN(n8416)
         );
  OAI21_X1 U10033 ( .B1(n8417), .B2(n8529), .A(n8416), .ZN(P2_U3164) );
  XOR2_X1 U10034 ( .A(n8419), .B(n8418), .Z(n8425) );
  AOI22_X1 U10035 ( .A1(n8749), .A2(n8538), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8421) );
  NAND2_X1 U10036 ( .A1(n8746), .A2(n8487), .ZN(n8420) );
  OAI211_X1 U10037 ( .C1(n8422), .C2(n8489), .A(n8421), .B(n8420), .ZN(n8423)
         );
  AOI21_X1 U10038 ( .B1(n9033), .B2(n8524), .A(n8423), .ZN(n8424) );
  OAI21_X1 U10039 ( .B1(n8425), .B2(n8529), .A(n8424), .ZN(P2_U3165) );
  XNOR2_X1 U10040 ( .A(n8426), .B(n8848), .ZN(n8427) );
  XNOR2_X1 U10041 ( .A(n4477), .B(n8427), .ZN(n8433) );
  NAND2_X1 U10042 ( .A1(n8533), .A2(n5041), .ZN(n8428) );
  NAND2_X1 U10043 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8620) );
  OAI211_X1 U10044 ( .C1(n8889), .C2(n8535), .A(n8428), .B(n8620), .ZN(n8431)
         );
  NOR2_X1 U10045 ( .A1(n8429), .A2(n8541), .ZN(n8430) );
  AOI211_X1 U10046 ( .C1(n8865), .C2(n8538), .A(n8431), .B(n8430), .ZN(n8432)
         );
  OAI21_X1 U10047 ( .B1(n8433), .B2(n8529), .A(n8432), .ZN(P2_U3166) );
  XOR2_X1 U10048 ( .A(n8435), .B(n8434), .Z(n8441) );
  NAND2_X1 U10049 ( .A1(n8849), .A2(n8533), .ZN(n8436) );
  NAND2_X1 U10050 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8657) );
  OAI211_X1 U10051 ( .C1(n8878), .C2(n8535), .A(n8436), .B(n8657), .ZN(n8439)
         );
  NOR2_X1 U10052 ( .A1(n8437), .A2(n8541), .ZN(n8438) );
  AOI211_X1 U10053 ( .C1(n8853), .C2(n8538), .A(n8439), .B(n8438), .ZN(n8440)
         );
  OAI21_X1 U10054 ( .B1(n8441), .B2(n8529), .A(n8440), .ZN(P2_U3168) );
  XNOR2_X1 U10055 ( .A(n8445), .B(n8778), .ZN(n8446) );
  XNOR2_X1 U10056 ( .A(n8447), .B(n8446), .ZN(n8452) );
  AOI22_X1 U10057 ( .A1(n8790), .A2(n8487), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8449) );
  NAND2_X1 U10058 ( .A1(n8764), .A2(n8538), .ZN(n8448) );
  OAI211_X1 U10059 ( .C1(n8762), .C2(n8489), .A(n8449), .B(n8448), .ZN(n8450)
         );
  AOI21_X1 U10060 ( .B1(n9039), .B2(n8524), .A(n8450), .ZN(n8451) );
  OAI21_X1 U10061 ( .B1(n8452), .B2(n8529), .A(n8451), .ZN(P2_U3169) );
  AOI21_X1 U10062 ( .B1(n8455), .B2(n8454), .A(n8453), .ZN(n8456) );
  OR2_X1 U10063 ( .A1(n8456), .A2(n8529), .ZN(n8463) );
  AOI21_X1 U10064 ( .B1(n8533), .B2(n8552), .A(n8457), .ZN(n8462) );
  AOI22_X1 U10065 ( .A1(n8487), .A2(n8996), .B1(n8458), .B2(n8524), .ZN(n8461)
         );
  NAND2_X1 U10066 ( .A1(n8538), .A2(n8459), .ZN(n8460) );
  NAND4_X1 U10067 ( .A1(n8463), .A2(n8462), .A3(n8461), .A4(n8460), .ZN(
        P2_U3170) );
  INV_X1 U10068 ( .A(n8464), .ZN(n8465) );
  AOI21_X1 U10069 ( .B1(n8467), .B2(n8466), .A(n8465), .ZN(n8473) );
  AOI22_X1 U10070 ( .A1(n8812), .A2(n8533), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8470) );
  NAND2_X1 U10071 ( .A1(n8815), .A2(n8538), .ZN(n8469) );
  OAI211_X1 U10072 ( .C1(n8835), .C2(n8535), .A(n8470), .B(n8469), .ZN(n8471)
         );
  AOI21_X1 U10073 ( .B1(n9062), .B2(n8524), .A(n8471), .ZN(n8472) );
  OAI21_X1 U10074 ( .B1(n8473), .B2(n8529), .A(n8472), .ZN(P2_U3173) );
  XNOR2_X1 U10075 ( .A(n8474), .B(n8545), .ZN(n8475) );
  XNOR2_X1 U10076 ( .A(n8476), .B(n8475), .ZN(n8482) );
  NAND2_X1 U10077 ( .A1(n8533), .A2(n8903), .ZN(n8477) );
  NAND2_X1 U10078 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8565) );
  OAI211_X1 U10079 ( .C1(n8478), .C2(n8535), .A(n8477), .B(n8565), .ZN(n8479)
         );
  AOI21_X1 U10080 ( .B1(n8908), .B2(n8538), .A(n8479), .ZN(n8481) );
  NAND2_X1 U10081 ( .A1(n8900), .A2(n8524), .ZN(n8480) );
  OAI211_X1 U10082 ( .C1(n8482), .C2(n8529), .A(n8481), .B(n8480), .ZN(
        P2_U3174) );
  INV_X1 U10083 ( .A(n9050), .ZN(n8493) );
  AOI21_X1 U10084 ( .B1(n8484), .B2(n8483), .A(n8529), .ZN(n8486) );
  NAND2_X1 U10085 ( .A1(n8486), .A2(n8485), .ZN(n8492) );
  AOI22_X1 U10086 ( .A1(n8812), .A2(n8487), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8488) );
  OAI21_X1 U10087 ( .B1(n8761), .B2(n8489), .A(n8488), .ZN(n8490) );
  AOI21_X1 U10088 ( .B1(n8793), .B2(n8538), .A(n8490), .ZN(n8491) );
  OAI211_X1 U10089 ( .C1(n8493), .C2(n8541), .A(n8492), .B(n8491), .ZN(
        P2_U3175) );
  INV_X1 U10090 ( .A(n8494), .ZN(n8982) );
  INV_X1 U10091 ( .A(n8495), .ZN(n8501) );
  OAI21_X1 U10092 ( .B1(n8498), .B2(n8497), .A(n8496), .ZN(n8499) );
  NAND3_X1 U10093 ( .A1(n8501), .A2(n8500), .A3(n8499), .ZN(n8508) );
  NAND2_X1 U10094 ( .A1(n8533), .A2(n8904), .ZN(n8503) );
  OAI211_X1 U10095 ( .C1(n8504), .C2(n8535), .A(n8503), .B(n8502), .ZN(n8505)
         );
  AOI21_X1 U10096 ( .B1(n8506), .B2(n8538), .A(n8505), .ZN(n8507) );
  OAI211_X1 U10097 ( .C1(n8982), .C2(n8541), .A(n8508), .B(n8507), .ZN(
        P2_U3176) );
  XOR2_X1 U10098 ( .A(n8510), .B(n8509), .Z(n8515) );
  INV_X1 U10099 ( .A(n8835), .ZN(n8811) );
  AND2_X1 U10100 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8688) );
  AOI21_X1 U10101 ( .B1(n8811), .B2(n8533), .A(n8688), .ZN(n8512) );
  NAND2_X1 U10102 ( .A1(n8538), .A2(n8836), .ZN(n8511) );
  OAI211_X1 U10103 ( .C1(n8861), .C2(n8535), .A(n8512), .B(n8511), .ZN(n8513)
         );
  AOI21_X1 U10104 ( .B1(n8954), .B2(n8524), .A(n8513), .ZN(n8514) );
  OAI21_X1 U10105 ( .B1(n8515), .B2(n8529), .A(n8514), .ZN(P2_U3178) );
  NAND2_X1 U10106 ( .A1(n8517), .A2(n8516), .ZN(n8520) );
  XNOR2_X1 U10107 ( .A(n8518), .B(n8747), .ZN(n8519) );
  XNOR2_X1 U10108 ( .A(n8520), .B(n8519), .ZN(n8526) );
  NAND2_X1 U10109 ( .A1(n8740), .A2(n8533), .ZN(n8522) );
  AOI22_X1 U10110 ( .A1(n8742), .A2(n8538), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8521) );
  OAI211_X1 U10111 ( .C1(n8762), .C2(n8535), .A(n8522), .B(n8521), .ZN(n8523)
         );
  AOI21_X1 U10112 ( .B1(n9027), .B2(n8524), .A(n8523), .ZN(n8525) );
  OAI21_X1 U10113 ( .B1(n8526), .B2(n8529), .A(n8525), .ZN(P2_U3180) );
  AOI211_X1 U10114 ( .C1(n8531), .C2(n8530), .A(n8529), .B(n8528), .ZN(n8532)
         );
  INV_X1 U10115 ( .A(n8532), .ZN(n8540) );
  NAND2_X1 U10116 ( .A1(n8533), .A2(n8848), .ZN(n8534) );
  NAND2_X1 U10117 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8610) );
  OAI211_X1 U10118 ( .C1(n8536), .C2(n8535), .A(n8534), .B(n8610), .ZN(n8537)
         );
  AOI21_X1 U10119 ( .B1(n8879), .B2(n8538), .A(n8537), .ZN(n8539) );
  OAI211_X1 U10120 ( .C1(n9088), .C2(n8541), .A(n8540), .B(n8539), .ZN(
        P2_U3181) );
  MUX2_X1 U10121 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8720), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8542), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10123 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8543), .S(P2_U3893), .Z(
        P2_U3520) );
  INV_X1 U10124 ( .A(P2_U3893), .ZN(n8681) );
  MUX2_X1 U10125 ( .A(n8730), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8681), .Z(
        P2_U3519) );
  MUX2_X1 U10126 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8740), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10127 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8747), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10128 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8739), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10129 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8746), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10130 ( .A(n8790), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8681), .Z(
        P2_U3514) );
  MUX2_X1 U10131 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8802), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10132 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8812), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10133 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8824), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10134 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8811), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10135 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8849), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10136 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n5041), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10137 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8848), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10138 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8544), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10139 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8903), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10140 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8545), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10141 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8904), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10142 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8546), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10143 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8547), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10144 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8548), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10145 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8549), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10146 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8550), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10147 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8551), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10148 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8552), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10149 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n10109), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10150 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8996), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6397), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10152 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n4392), .S(P2_U3893), .Z(
        P2_U3492) );
  XNOR2_X1 U10153 ( .A(n8574), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U10154 ( .A1(n8555), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8590) );
  OAI21_X1 U10155 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8555), .A(n8590), .ZN(
        n8568) );
  NAND2_X1 U10156 ( .A1(n8562), .A2(n8561), .ZN(n8559) );
  INV_X1 U10157 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8556) );
  INV_X1 U10158 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8573) );
  MUX2_X1 U10159 ( .A(n8556), .B(n8573), .S(n4387), .Z(n8557) );
  NAND2_X1 U10160 ( .A1(n8557), .A2(n8572), .ZN(n8580) );
  OAI21_X1 U10161 ( .B1(n8572), .B2(n8557), .A(n8580), .ZN(n8560) );
  INV_X1 U10162 ( .A(n8560), .ZN(n8558) );
  NAND2_X1 U10163 ( .A1(n8559), .A2(n8558), .ZN(n8581) );
  NAND3_X1 U10164 ( .A1(n8562), .A2(n8561), .A3(n8560), .ZN(n8563) );
  AOI21_X1 U10165 ( .B1(n8581), .B2(n8563), .A(n8683), .ZN(n8567) );
  NAND2_X1 U10166 ( .A1(n8701), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8564) );
  OAI211_X1 U10167 ( .C1(n8705), .C2(n4984), .A(n8565), .B(n8564), .ZN(n8566)
         );
  AOI211_X1 U10168 ( .C1(n8568), .C2(n8670), .A(n8567), .B(n8566), .ZN(n8569)
         );
  OAI21_X1 U10169 ( .B1(n8570), .B2(n8690), .A(n8569), .ZN(P2_U3195) );
  XNOR2_X1 U10170 ( .A(n8587), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8595) );
  XOR2_X1 U10171 ( .A(n8595), .B(n8596), .Z(n8594) );
  OAI21_X1 U10172 ( .B1(n8622), .B2(n10237), .A(n8575), .ZN(n8584) );
  NAND2_X1 U10173 ( .A1(n8581), .A2(n8580), .ZN(n8578) );
  INV_X1 U10174 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8586) );
  INV_X1 U10175 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8966) );
  MUX2_X1 U10176 ( .A(n8586), .B(n8966), .S(n4387), .Z(n8576) );
  NAND2_X1 U10177 ( .A1(n8587), .A2(n8576), .ZN(n8607) );
  OAI21_X1 U10178 ( .B1(n8587), .B2(n8576), .A(n8607), .ZN(n8579) );
  INV_X1 U10179 ( .A(n8579), .ZN(n8577) );
  NAND3_X1 U10180 ( .A1(n8581), .A2(n8580), .A3(n8579), .ZN(n8582) );
  AOI21_X1 U10181 ( .B1(n8608), .B2(n8582), .A(n8683), .ZN(n8583) );
  AOI211_X1 U10182 ( .C1(n8634), .C2(n8587), .A(n8584), .B(n8583), .ZN(n8593)
         );
  INV_X1 U10183 ( .A(n8585), .ZN(n8588) );
  XNOR2_X1 U10184 ( .A(n8587), .B(n8586), .ZN(n8589) );
  AND3_X1 U10185 ( .A1(n8590), .A2(n8589), .A3(n8588), .ZN(n8591) );
  OAI21_X1 U10186 ( .B1(n8599), .B2(n8591), .A(n8670), .ZN(n8592) );
  OAI211_X1 U10187 ( .C1(n8594), .C2(n8690), .A(n8593), .B(n8592), .ZN(
        P2_U3196) );
  XNOR2_X1 U10188 ( .A(n8619), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n8616) );
  NOR2_X1 U10189 ( .A1(n8599), .A2(n8598), .ZN(n8600) );
  OAI21_X1 U10190 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8601), .A(n8639), .ZN(
        n8614) );
  NAND2_X1 U10191 ( .A1(n8608), .A2(n8607), .ZN(n8604) );
  INV_X1 U10192 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10378) );
  INV_X1 U10193 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8961) );
  MUX2_X1 U10194 ( .A(n10378), .B(n8961), .S(n4387), .Z(n8602) );
  OR2_X1 U10195 ( .A1(n8602), .A2(n8618), .ZN(n8603) );
  NAND2_X1 U10196 ( .A1(n8618), .A2(n8602), .ZN(n8629) );
  AND2_X1 U10197 ( .A1(n8603), .A2(n8629), .ZN(n8605) );
  INV_X1 U10198 ( .A(n8605), .ZN(n8606) );
  NAND3_X1 U10199 ( .A1(n8608), .A2(n8607), .A3(n8606), .ZN(n8609) );
  AOI21_X1 U10200 ( .B1(n8630), .B2(n8609), .A(n8683), .ZN(n8613) );
  NAND2_X1 U10201 ( .A1(n8634), .A2(n8618), .ZN(n8611) );
  OAI211_X1 U10202 ( .C1(n8622), .C2(n10464), .A(n8611), .B(n8610), .ZN(n8612)
         );
  AOI211_X1 U10203 ( .C1(n8614), .C2(n8670), .A(n8613), .B(n8612), .ZN(n8615)
         );
  OAI21_X1 U10204 ( .B1(n8616), .B2(n8690), .A(n8615), .ZN(P2_U3197) );
  XNOR2_X1 U10205 ( .A(n8636), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8644) );
  XOR2_X1 U10206 ( .A(n8644), .B(n8645), .Z(n8643) );
  INV_X1 U10207 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8621) );
  OAI21_X1 U10208 ( .B1(n8622), .B2(n8621), .A(n8620), .ZN(n8633) );
  NAND2_X1 U10209 ( .A1(n8630), .A2(n8629), .ZN(n8627) );
  INV_X1 U10210 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10210) );
  INV_X1 U10211 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8958) );
  MUX2_X1 U10212 ( .A(n10210), .B(n8958), .S(n4387), .Z(n8623) );
  NAND2_X1 U10213 ( .A1(n8623), .A2(n8636), .ZN(n8652) );
  INV_X1 U10214 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U10215 ( .A1(n8624), .A2(n8647), .ZN(n8625) );
  NAND2_X1 U10216 ( .A1(n8652), .A2(n8625), .ZN(n8628) );
  INV_X1 U10217 ( .A(n8628), .ZN(n8626) );
  NAND3_X1 U10218 ( .A1(n8630), .A2(n8629), .A3(n8628), .ZN(n8631) );
  AOI21_X1 U10219 ( .B1(n8654), .B2(n8631), .A(n8683), .ZN(n8632) );
  AOI211_X1 U10220 ( .C1(n8634), .C2(n8636), .A(n8633), .B(n8632), .ZN(n8642)
         );
  INV_X1 U10221 ( .A(n8635), .ZN(n8637) );
  XNOR2_X1 U10222 ( .A(n8636), .B(n10210), .ZN(n8638) );
  AND3_X1 U10223 ( .A1(n8639), .A2(n8638), .A3(n8637), .ZN(n8640) );
  OAI21_X1 U10224 ( .B1(n8646), .B2(n8640), .A(n8670), .ZN(n8641) );
  OAI211_X1 U10225 ( .C1(n8643), .C2(n8690), .A(n8642), .B(n8641), .ZN(
        P2_U3198) );
  XOR2_X1 U10226 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8665), .Z(n8662) );
  OAI21_X1 U10227 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8649), .A(n4994), .ZN(
        n8660) );
  NAND2_X1 U10228 ( .A1(n8654), .A2(n8652), .ZN(n8650) );
  MUX2_X1 U10229 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n4387), .Z(n8673) );
  XNOR2_X1 U10230 ( .A(n8673), .B(n8674), .ZN(n8651) );
  NAND2_X1 U10231 ( .A1(n8650), .A2(n8651), .ZN(n8677) );
  INV_X1 U10232 ( .A(n8651), .ZN(n8653) );
  NAND3_X1 U10233 ( .A1(n8654), .A2(n8653), .A3(n8652), .ZN(n8655) );
  AOI21_X1 U10234 ( .B1(n8677), .B2(n8655), .A(n8683), .ZN(n8659) );
  NAND2_X1 U10235 ( .A1(n8701), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8656) );
  OAI211_X1 U10236 ( .C1(n8705), .C2(n4895), .A(n8657), .B(n8656), .ZN(n8658)
         );
  OAI21_X1 U10237 ( .B1(n8662), .B2(n8690), .A(n8661), .ZN(P2_U3199) );
  XOR2_X1 U10238 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8709), .Z(n8710) );
  INV_X1 U10239 ( .A(n8663), .ZN(n8664) );
  NAND2_X1 U10240 ( .A1(n8698), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8691) );
  INV_X1 U10241 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U10242 ( .A1(n8709), .A2(n8838), .ZN(n8666) );
  AND2_X1 U10243 ( .A1(n8691), .A2(n8666), .ZN(n8668) );
  INV_X1 U10244 ( .A(n8692), .ZN(n8672) );
  INV_X1 U10245 ( .A(n8673), .ZN(n8675) );
  NAND2_X1 U10246 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  NAND2_X1 U10247 ( .A1(n8677), .A2(n8676), .ZN(n8679) );
  MUX2_X1 U10248 ( .A(n8838), .B(n10231), .S(n4387), .Z(n8678) );
  NOR2_X1 U10249 ( .A1(n8679), .A2(n8678), .ZN(n8696) );
  NAND2_X1 U10250 ( .A1(n8679), .A2(n8678), .ZN(n8697) );
  INV_X1 U10251 ( .A(n8697), .ZN(n8680) );
  NOR2_X1 U10252 ( .A1(n8696), .A2(n8680), .ZN(n8684) );
  INV_X1 U10253 ( .A(n8684), .ZN(n8682) );
  OAI21_X1 U10254 ( .B1(n8682), .B2(n8681), .A(n8705), .ZN(n8686) );
  NOR2_X1 U10255 ( .A1(n8684), .A2(n8683), .ZN(n8685) );
  MUX2_X1 U10256 ( .A(n8686), .B(n8685), .S(n8698), .Z(n8687) );
  XNOR2_X1 U10257 ( .A(n8704), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8695) );
  XNOR2_X1 U10258 ( .A(n8693), .B(n8695), .ZN(n8718) );
  XNOR2_X1 U10259 ( .A(n8704), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8713) );
  MUX2_X1 U10260 ( .A(n8713), .B(n8695), .S(n8694), .Z(n8700) );
  AOI21_X1 U10261 ( .B1(n8698), .B2(n8697), .A(n8696), .ZN(n8699) );
  XOR2_X1 U10262 ( .A(n8700), .B(n8699), .Z(n8708) );
  NAND2_X1 U10263 ( .A1(n8701), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8702) );
  OAI211_X1 U10264 ( .C1(n8705), .C2(n8704), .A(n8703), .B(n8702), .ZN(n8706)
         );
  AOI21_X1 U10265 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8716) );
  OAI211_X1 U10266 ( .C1(n8718), .C2(n8717), .A(n8716), .B(n8715), .ZN(
        P2_U3201) );
  NAND2_X1 U10267 ( .A1(n10130), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U10268 ( .A1(n8720), .A2(n8719), .ZN(n9013) );
  INV_X1 U10269 ( .A(n9013), .ZN(n8722) );
  OAI21_X1 U10270 ( .B1(n8722), .B2(n8721), .A(n10128), .ZN(n8724) );
  OAI211_X1 U10271 ( .C1(n9015), .C2(n10115), .A(n8723), .B(n8724), .ZN(
        P2_U3202) );
  NAND2_X1 U10272 ( .A1(n10130), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8725) );
  OAI211_X1 U10273 ( .C1(n9018), .C2(n10115), .A(n8725), .B(n8724), .ZN(
        P2_U3203) );
  XNOR2_X1 U10274 ( .A(n8727), .B(n8726), .ZN(n9024) );
  MUX2_X1 U10275 ( .A(n8731), .B(n9019), .S(n10128), .Z(n8734) );
  AOI22_X1 U10276 ( .A1(n9021), .A2(n8925), .B1(n8924), .B2(n8732), .ZN(n8733)
         );
  OAI211_X1 U10277 ( .C1(n9024), .C2(n8883), .A(n8734), .B(n8733), .ZN(
        P2_U3206) );
  XNOR2_X1 U10278 ( .A(n8736), .B(n8735), .ZN(n9030) );
  XNOR2_X1 U10279 ( .A(n8737), .B(n8738), .ZN(n8741) );
  AOI222_X1 U10280 ( .A1(n10111), .A2(n8741), .B1(n8740), .B2(n10108), .C1(
        n8739), .C2(n10107), .ZN(n9025) );
  MUX2_X1 U10281 ( .A(n10441), .B(n9025), .S(n10128), .Z(n8744) );
  AOI22_X1 U10282 ( .A1(n9027), .A2(n8925), .B1(n8924), .B2(n8742), .ZN(n8743)
         );
  OAI211_X1 U10283 ( .C1(n9030), .C2(n8883), .A(n8744), .B(n8743), .ZN(
        P2_U3207) );
  XOR2_X1 U10284 ( .A(n8753), .B(n8745), .Z(n8748) );
  AOI222_X1 U10285 ( .A1(n10111), .A2(n8748), .B1(n8747), .B2(n10108), .C1(
        n8746), .C2(n10107), .ZN(n9031) );
  INV_X1 U10286 ( .A(n10121), .ZN(n8750) );
  AOI22_X1 U10287 ( .A1(n9033), .A2(n8750), .B1(n8924), .B2(n8749), .ZN(n8751)
         );
  AOI21_X1 U10288 ( .B1(n9031), .B2(n8751), .A(n10130), .ZN(n8756) );
  XNOR2_X1 U10289 ( .A(n8752), .B(n8753), .ZN(n9036) );
  OAI22_X1 U10290 ( .A1(n9036), .A2(n8883), .B1(n8754), .B2(n10128), .ZN(n8755) );
  OR2_X1 U10291 ( .A1(n8756), .A2(n8755), .ZN(P2_U3208) );
  NOR2_X1 U10292 ( .A1(n8757), .A2(n10121), .ZN(n8763) );
  NAND2_X1 U10293 ( .A1(n8759), .A2(n8758), .ZN(n8767) );
  AOI211_X1 U10294 ( .C1(n8924), .C2(n8764), .A(n8763), .B(n8939), .ZN(n8769)
         );
  NAND2_X1 U10295 ( .A1(n8765), .A2(n8771), .ZN(n8766) );
  XOR2_X1 U10296 ( .A(n8767), .B(n8766), .Z(n9040) );
  AOI22_X1 U10297 ( .A1(n9040), .A2(n10117), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10130), .ZN(n8768) );
  OAI21_X1 U10298 ( .B1(n8769), .B2(n10130), .A(n8768), .ZN(P2_U3209) );
  INV_X1 U10299 ( .A(n8771), .ZN(n8772) );
  NOR2_X1 U10300 ( .A1(n8773), .A2(n8772), .ZN(n8775) );
  XNOR2_X1 U10301 ( .A(n8770), .B(n8775), .ZN(n9045) );
  XNOR2_X1 U10302 ( .A(n8774), .B(n8775), .ZN(n8776) );
  OAI222_X1 U10303 ( .A1(n8888), .A2(n8778), .B1(n8998), .B2(n8777), .C1(
        n10132), .C2(n8776), .ZN(n9043) );
  INV_X1 U10304 ( .A(n9043), .ZN(n8779) );
  MUX2_X1 U10305 ( .A(n8780), .B(n8779), .S(n10128), .Z(n8783) );
  AOI22_X1 U10306 ( .A1(n6416), .A2(n8880), .B1(n8924), .B2(n8781), .ZN(n8782)
         );
  OAI211_X1 U10307 ( .C1(n9045), .C2(n8883), .A(n8783), .B(n8782), .ZN(
        P2_U3210) );
  XNOR2_X1 U10308 ( .A(n8784), .B(n8785), .ZN(n9051) );
  INV_X1 U10309 ( .A(n9051), .ZN(n8796) );
  NAND3_X1 U10310 ( .A1(n8799), .A2(n8787), .A3(n8786), .ZN(n8788) );
  NAND2_X1 U10311 ( .A1(n8789), .A2(n8788), .ZN(n8791) );
  AOI222_X1 U10312 ( .A1(n10111), .A2(n8791), .B1(n8790), .B2(n10108), .C1(
        n8812), .C2(n10107), .ZN(n9048) );
  MUX2_X1 U10313 ( .A(n8792), .B(n9048), .S(n10128), .Z(n8795) );
  AOI22_X1 U10314 ( .A1(n9050), .A2(n8880), .B1(n8924), .B2(n8793), .ZN(n8794)
         );
  OAI211_X1 U10315 ( .C1(n8796), .C2(n8883), .A(n8795), .B(n8794), .ZN(
        P2_U3211) );
  XNOR2_X1 U10316 ( .A(n8797), .B(n8798), .ZN(n9059) );
  INV_X1 U10317 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8804) );
  OAI21_X1 U10318 ( .B1(n8801), .B2(n8800), .A(n8799), .ZN(n8803) );
  AOI222_X1 U10319 ( .A1(n10111), .A2(n8803), .B1(n8802), .B2(n10108), .C1(
        n8824), .C2(n10107), .ZN(n9054) );
  MUX2_X1 U10320 ( .A(n8804), .B(n9054), .S(n10128), .Z(n8807) );
  AOI22_X1 U10321 ( .A1(n9056), .A2(n8880), .B1(n8924), .B2(n8805), .ZN(n8806)
         );
  OAI211_X1 U10322 ( .C1(n9059), .C2(n8883), .A(n8807), .B(n8806), .ZN(
        P2_U3212) );
  XNOR2_X1 U10323 ( .A(n8808), .B(n8810), .ZN(n9063) );
  INV_X1 U10324 ( .A(n9063), .ZN(n8818) );
  INV_X1 U10325 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8814) );
  XNOR2_X1 U10326 ( .A(n8809), .B(n8810), .ZN(n8813) );
  AOI222_X1 U10327 ( .A1(n10111), .A2(n8813), .B1(n8812), .B2(n10108), .C1(
        n8811), .C2(n10107), .ZN(n9060) );
  MUX2_X1 U10328 ( .A(n8814), .B(n9060), .S(n10128), .Z(n8817) );
  AOI22_X1 U10329 ( .A1(n9062), .A2(n8880), .B1(n8924), .B2(n8815), .ZN(n8816)
         );
  OAI211_X1 U10330 ( .C1(n8818), .C2(n8883), .A(n8817), .B(n8816), .ZN(
        P2_U3213) );
  NAND2_X1 U10331 ( .A1(n8819), .A2(n8820), .ZN(n8821) );
  XNOR2_X1 U10332 ( .A(n8823), .B(n8821), .ZN(n9071) );
  INV_X1 U10333 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8826) );
  XOR2_X1 U10334 ( .A(n8823), .B(n8822), .Z(n8825) );
  AOI222_X1 U10335 ( .A1(n10111), .A2(n8825), .B1(n8824), .B2(n10108), .C1(
        n8849), .C2(n10107), .ZN(n9066) );
  MUX2_X1 U10336 ( .A(n8826), .B(n9066), .S(n10128), .Z(n8829) );
  AOI22_X1 U10337 ( .A1(n9068), .A2(n8880), .B1(n8924), .B2(n8827), .ZN(n8828)
         );
  OAI211_X1 U10338 ( .C1(n9071), .C2(n8883), .A(n8829), .B(n8828), .ZN(
        P2_U3214) );
  NAND2_X1 U10339 ( .A1(n8830), .A2(n8832), .ZN(n8831) );
  NAND2_X1 U10340 ( .A1(n8819), .A2(n8831), .ZN(n9075) );
  XNOR2_X1 U10341 ( .A(n8833), .B(n8832), .ZN(n8834) );
  OAI222_X1 U10342 ( .A1(n8888), .A2(n8835), .B1(n8998), .B2(n8861), .C1(n8834), .C2(n10132), .ZN(n8953) );
  NAND2_X1 U10343 ( .A1(n8953), .A2(n10128), .ZN(n8841) );
  INV_X1 U10344 ( .A(n8836), .ZN(n8837) );
  OAI22_X1 U10345 ( .A1(n10128), .A2(n8838), .B1(n8837), .B2(n10122), .ZN(
        n8839) );
  AOI21_X1 U10346 ( .B1(n8954), .B2(n8880), .A(n8839), .ZN(n8840) );
  OAI211_X1 U10347 ( .C1(n9075), .C2(n8883), .A(n8841), .B(n8840), .ZN(
        P2_U3215) );
  INV_X1 U10348 ( .A(n8843), .ZN(n8844) );
  AOI21_X1 U10349 ( .B1(n8846), .B2(n8842), .A(n8844), .ZN(n9080) );
  OAI211_X1 U10350 ( .C1(n8847), .C2(n8846), .A(n8845), .B(n10111), .ZN(n8851)
         );
  AOI22_X1 U10351 ( .A1(n8849), .A2(n10108), .B1(n10107), .B2(n8848), .ZN(
        n8850) );
  AND2_X1 U10352 ( .A1(n8851), .A2(n8850), .ZN(n9076) );
  INV_X1 U10353 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8852) );
  MUX2_X1 U10354 ( .A(n9076), .B(n8852), .S(n10130), .Z(n8855) );
  AOI22_X1 U10355 ( .A1(n9077), .A2(n8925), .B1(n8924), .B2(n8853), .ZN(n8854)
         );
  OAI211_X1 U10356 ( .C1(n9080), .C2(n8883), .A(n8855), .B(n8854), .ZN(
        P2_U3216) );
  XOR2_X1 U10357 ( .A(n8856), .B(n8858), .Z(n9086) );
  INV_X1 U10358 ( .A(n8857), .ZN(n8860) );
  INV_X1 U10359 ( .A(n8858), .ZN(n8859) );
  AOI21_X1 U10360 ( .B1(n8860), .B2(n8859), .A(n10132), .ZN(n8864) );
  OAI22_X1 U10361 ( .A1(n8861), .A2(n8888), .B1(n8889), .B2(n8998), .ZN(n8862)
         );
  AOI21_X1 U10362 ( .B1(n8864), .B2(n8863), .A(n8862), .ZN(n9081) );
  MUX2_X1 U10363 ( .A(n10210), .B(n9081), .S(n10128), .Z(n8867) );
  AOI22_X1 U10364 ( .A1(n9083), .A2(n8925), .B1(n8924), .B2(n8865), .ZN(n8866)
         );
  OAI211_X1 U10365 ( .C1(n9086), .C2(n8883), .A(n8867), .B(n8866), .ZN(
        P2_U3217) );
  XNOR2_X1 U10366 ( .A(n8868), .B(n8871), .ZN(n9089) );
  NAND2_X1 U10367 ( .A1(n8869), .A2(n8870), .ZN(n8885) );
  NAND2_X1 U10368 ( .A1(n8885), .A2(n8897), .ZN(n8891) );
  INV_X1 U10369 ( .A(n8871), .ZN(n8873) );
  NAND3_X1 U10370 ( .A1(n8891), .A2(n8873), .A3(n8872), .ZN(n8874) );
  NAND3_X1 U10371 ( .A1(n8875), .A2(n10111), .A3(n8874), .ZN(n8877) );
  NAND2_X1 U10372 ( .A1(n10107), .A2(n8903), .ZN(n8876) );
  OAI211_X1 U10373 ( .C1(n8878), .C2(n8888), .A(n8877), .B(n8876), .ZN(n9087)
         );
  INV_X1 U10374 ( .A(n9087), .ZN(n8962) );
  MUX2_X1 U10375 ( .A(n8962), .B(n10378), .S(n10130), .Z(n8882) );
  AOI22_X1 U10376 ( .A1(n8963), .A2(n8880), .B1(n8924), .B2(n8879), .ZN(n8881)
         );
  OAI211_X1 U10377 ( .C1(n9089), .C2(n8883), .A(n8882), .B(n8881), .ZN(
        P2_U3218) );
  NOR2_X1 U10378 ( .A1(n8884), .A2(n10121), .ZN(n8894) );
  INV_X1 U10379 ( .A(n8885), .ZN(n8886) );
  AOI21_X1 U10380 ( .B1(n8886), .B2(n6198), .A(n10132), .ZN(n8892) );
  OAI22_X1 U10381 ( .A1(n8889), .A2(n8888), .B1(n8887), .B2(n8998), .ZN(n8890)
         );
  AOI21_X1 U10382 ( .B1(n8892), .B2(n8891), .A(n8890), .ZN(n9092) );
  INV_X1 U10383 ( .A(n9092), .ZN(n8893) );
  AOI211_X1 U10384 ( .C1(n8924), .C2(n8895), .A(n8894), .B(n8893), .ZN(n8899)
         );
  XNOR2_X1 U10385 ( .A(n8896), .B(n8897), .ZN(n9096) );
  AOI22_X1 U10386 ( .A1(n9096), .A2(n10117), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n10130), .ZN(n8898) );
  OAI21_X1 U10387 ( .B1(n8899), .B2(n10130), .A(n8898), .ZN(P2_U3219) );
  INV_X1 U10388 ( .A(n8900), .ZN(n9101) );
  NOR2_X1 U10389 ( .A1(n9101), .A2(n10121), .ZN(n8907) );
  OAI211_X1 U10390 ( .C1(n8902), .C2(n8901), .A(n8869), .B(n10111), .ZN(n8906)
         );
  AOI22_X1 U10391 ( .A1(n10107), .A2(n8904), .B1(n10108), .B2(n8903), .ZN(
        n8905) );
  NAND2_X1 U10392 ( .A1(n8906), .A2(n8905), .ZN(n9099) );
  AOI211_X1 U10393 ( .C1(n8924), .C2(n8908), .A(n8907), .B(n9099), .ZN(n8913)
         );
  XNOR2_X1 U10394 ( .A(n8910), .B(n8909), .ZN(n9103) );
  INV_X1 U10395 ( .A(n9103), .ZN(n8911) );
  AOI22_X1 U10396 ( .A1(n8911), .A2(n10117), .B1(P2_REG2_REG_13__SCAN_IN), 
        .B2(n10130), .ZN(n8912) );
  OAI21_X1 U10397 ( .B1(n8913), .B2(n10130), .A(n8912), .ZN(P2_U3220) );
  NAND2_X1 U10398 ( .A1(n8918), .A2(n8914), .ZN(n8988) );
  OR2_X1 U10399 ( .A1(n8918), .A2(n8914), .ZN(n8915) );
  NAND2_X1 U10400 ( .A1(n8988), .A2(n8915), .ZN(n9009) );
  NAND2_X1 U10401 ( .A1(n9009), .A2(n8990), .ZN(n8923) );
  AOI22_X1 U10402 ( .A1(n10107), .A2(n6723), .B1(n10108), .B2(n6397), .ZN(
        n8922) );
  INV_X1 U10403 ( .A(n8916), .ZN(n8917) );
  OR2_X1 U10404 ( .A1(n8918), .A2(n8917), .ZN(n8991) );
  NAND2_X1 U10405 ( .A1(n8918), .A2(n8917), .ZN(n8919) );
  NAND2_X1 U10406 ( .A1(n8991), .A2(n8919), .ZN(n8920) );
  NAND2_X1 U10407 ( .A1(n8920), .A2(n10111), .ZN(n8921) );
  AND3_X1 U10408 ( .A1(n8923), .A2(n8922), .A3(n8921), .ZN(n9011) );
  MUX2_X1 U10409 ( .A(n9011), .B(n4712), .S(n10130), .Z(n8929) );
  AOI22_X1 U10410 ( .A1(n8925), .A2(n9007), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8924), .ZN(n8928) );
  NAND2_X1 U10411 ( .A1(n8926), .A2(n9009), .ZN(n8927) );
  NAND3_X1 U10412 ( .A1(n8929), .A2(n8928), .A3(n8927), .ZN(P2_U3232) );
  NOR2_X1 U10413 ( .A1(n9013), .A2(n10164), .ZN(n8931) );
  AOI21_X1 U10414 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10164), .A(n8931), .ZN(
        n8930) );
  OAI21_X1 U10415 ( .B1(n9015), .B2(n8971), .A(n8930), .ZN(P2_U3490) );
  AOI21_X1 U10416 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10164), .A(n8931), .ZN(
        n8932) );
  OAI21_X1 U10417 ( .B1(n9018), .B2(n8971), .A(n8932), .ZN(P2_U3489) );
  INV_X1 U10418 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8933) );
  INV_X1 U10419 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10466) );
  MUX2_X1 U10420 ( .A(n10466), .B(n9025), .S(n10166), .Z(n8935) );
  NAND2_X1 U10421 ( .A1(n9027), .A2(n8967), .ZN(n8934) );
  OAI211_X1 U10422 ( .C1(n8972), .C2(n9030), .A(n8935), .B(n8934), .ZN(
        P2_U3485) );
  INV_X1 U10423 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8936) );
  MUX2_X1 U10424 ( .A(n8936), .B(n9031), .S(n10166), .Z(n8938) );
  NAND2_X1 U10425 ( .A1(n9033), .A2(n8967), .ZN(n8937) );
  OAI211_X1 U10426 ( .C1(n8972), .C2(n9036), .A(n8938), .B(n8937), .ZN(
        P2_U3484) );
  INV_X1 U10427 ( .A(n8939), .ZN(n9037) );
  MUX2_X1 U10428 ( .A(n10470), .B(n9037), .S(n10166), .Z(n8941) );
  AOI22_X1 U10429 ( .A1(n9040), .A2(n8968), .B1(n8967), .B2(n9039), .ZN(n8940)
         );
  NAND2_X1 U10430 ( .A1(n8941), .A2(n8940), .ZN(P2_U3483) );
  MUX2_X1 U10431 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9043), .S(n10166), .Z(
        n8943) );
  OAI22_X1 U10432 ( .A1(n9045), .A2(n8972), .B1(n9044), .B2(n8971), .ZN(n8942)
         );
  OR2_X1 U10433 ( .A1(n8943), .A2(n8942), .ZN(P2_U3482) );
  INV_X1 U10434 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8944) );
  MUX2_X1 U10435 ( .A(n8944), .B(n9048), .S(n10166), .Z(n8946) );
  AOI22_X1 U10436 ( .A1(n9051), .A2(n8968), .B1(n8967), .B2(n9050), .ZN(n8945)
         );
  NAND2_X1 U10437 ( .A1(n8946), .A2(n8945), .ZN(P2_U3481) );
  MUX2_X1 U10438 ( .A(n10267), .B(n9054), .S(n10166), .Z(n8948) );
  NAND2_X1 U10439 ( .A1(n9056), .A2(n8967), .ZN(n8947) );
  OAI211_X1 U10440 ( .C1(n8972), .C2(n9059), .A(n8948), .B(n8947), .ZN(
        P2_U3480) );
  MUX2_X1 U10441 ( .A(n10320), .B(n9060), .S(n10166), .Z(n8950) );
  AOI22_X1 U10442 ( .A1(n9063), .A2(n8968), .B1(n8967), .B2(n9062), .ZN(n8949)
         );
  NAND2_X1 U10443 ( .A1(n8950), .A2(n8949), .ZN(P2_U3479) );
  MUX2_X1 U10444 ( .A(n10374), .B(n9066), .S(n10166), .Z(n8952) );
  NAND2_X1 U10445 ( .A1(n9068), .A2(n8967), .ZN(n8951) );
  OAI211_X1 U10446 ( .C1(n9071), .C2(n8972), .A(n8952), .B(n8951), .ZN(
        P2_U3478) );
  AOI21_X1 U10447 ( .B1(n10141), .B2(n8954), .A(n8953), .ZN(n9072) );
  MUX2_X1 U10448 ( .A(n10231), .B(n9072), .S(n10166), .Z(n8955) );
  OAI21_X1 U10449 ( .B1(n8972), .B2(n9075), .A(n8955), .ZN(P2_U3477) );
  MUX2_X1 U10450 ( .A(n9076), .B(n10341), .S(n10164), .Z(n8957) );
  NAND2_X1 U10451 ( .A1(n9077), .A2(n8967), .ZN(n8956) );
  OAI211_X1 U10452 ( .C1(n9080), .C2(n8972), .A(n8957), .B(n8956), .ZN(
        P2_U3476) );
  MUX2_X1 U10453 ( .A(n8958), .B(n9081), .S(n10166), .Z(n8960) );
  NAND2_X1 U10454 ( .A1(n9083), .A2(n8967), .ZN(n8959) );
  OAI211_X1 U10455 ( .C1(n9086), .C2(n8972), .A(n8960), .B(n8959), .ZN(
        P2_U3475) );
  MUX2_X1 U10456 ( .A(n8962), .B(n8961), .S(n10164), .Z(n8965) );
  NAND2_X1 U10457 ( .A1(n8963), .A2(n8967), .ZN(n8964) );
  OAI211_X1 U10458 ( .C1(n8972), .C2(n9089), .A(n8965), .B(n8964), .ZN(
        P2_U3474) );
  MUX2_X1 U10459 ( .A(n8966), .B(n9092), .S(n10166), .Z(n8970) );
  AOI22_X1 U10460 ( .A1(n9096), .A2(n8968), .B1(n8967), .B2(n9093), .ZN(n8969)
         );
  NAND2_X1 U10461 ( .A1(n8970), .A2(n8969), .ZN(P2_U3473) );
  MUX2_X1 U10462 ( .A(n9099), .B(P2_REG1_REG_13__SCAN_IN), .S(n10164), .Z(
        n8974) );
  OAI22_X1 U10463 ( .A1(n9103), .A2(n8972), .B1(n9101), .B2(n8971), .ZN(n8973)
         );
  OR2_X1 U10464 ( .A1(n8974), .A2(n8973), .ZN(P2_U3472) );
  NAND3_X1 U10465 ( .A1(n8161), .A2(n10149), .A3(n8975), .ZN(n8976) );
  OAI211_X1 U10466 ( .C1(n8978), .C2(n10151), .A(n8977), .B(n8976), .ZN(n9106)
         );
  MUX2_X1 U10467 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9106), .S(n10166), .Z(
        P2_U3471) );
  NAND2_X1 U10468 ( .A1(n8979), .A2(n10149), .ZN(n8980) );
  OAI211_X1 U10469 ( .C1(n8982), .C2(n10151), .A(n8981), .B(n8980), .ZN(n9107)
         );
  MUX2_X1 U10470 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9107), .S(n10166), .Z(
        P2_U3470) );
  AOI22_X1 U10471 ( .A1(n8984), .A2(n10149), .B1(n10141), .B2(n8983), .ZN(
        n8986) );
  NAND2_X1 U10472 ( .A1(n8986), .A2(n8985), .ZN(n9108) );
  MUX2_X1 U10473 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9108), .S(n10166), .Z(
        P2_U3469) );
  NAND2_X1 U10474 ( .A1(n8988), .A2(n8987), .ZN(n8989) );
  XNOR2_X1 U10475 ( .A(n8989), .B(n8992), .ZN(n10126) );
  NAND2_X1 U10476 ( .A1(n10126), .A2(n8990), .ZN(n9003) );
  OAI211_X1 U10477 ( .C1(n9007), .C2(n4392), .A(n8991), .B(n8992), .ZN(n8995)
         );
  INV_X1 U10478 ( .A(n8992), .ZN(n8993) );
  NAND2_X1 U10479 ( .A1(n8994), .A2(n8993), .ZN(n10105) );
  NAND2_X1 U10480 ( .A1(n8995), .A2(n10105), .ZN(n9001) );
  NAND2_X1 U10481 ( .A1(n10108), .A2(n8996), .ZN(n8997) );
  OAI21_X1 U10482 ( .B1(n8999), .B2(n8998), .A(n8997), .ZN(n9000) );
  AOI21_X1 U10483 ( .B1(n9001), .B2(n10111), .A(n9000), .ZN(n9002) );
  AND2_X1 U10484 ( .A1(n9003), .A2(n9002), .ZN(n10123) );
  AOI22_X1 U10485 ( .A1(n10126), .A2(n9008), .B1(n10141), .B2(n9004), .ZN(
        n9005) );
  AND2_X1 U10486 ( .A1(n10123), .A2(n9005), .ZN(n10138) );
  INV_X1 U10487 ( .A(n10138), .ZN(n9006) );
  MUX2_X1 U10488 ( .A(n9006), .B(P2_REG1_REG_2__SCAN_IN), .S(n10164), .Z(
        P2_U3461) );
  AOI22_X1 U10489 ( .A1(n9009), .A2(n9008), .B1(n9007), .B2(n10141), .ZN(n9010) );
  AND2_X1 U10490 ( .A1(n9011), .A2(n9010), .ZN(n10137) );
  INV_X1 U10491 ( .A(n10137), .ZN(n9012) );
  MUX2_X1 U10492 ( .A(n9012), .B(P2_REG1_REG_1__SCAN_IN), .S(n10164), .Z(
        P2_U3460) );
  NOR2_X1 U10493 ( .A1(n9013), .A2(n10159), .ZN(n9016) );
  AOI21_X1 U10494 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n10159), .A(n9016), .ZN(
        n9014) );
  OAI21_X1 U10495 ( .B1(n9015), .B2(n9100), .A(n9014), .ZN(P2_U3458) );
  AOI21_X1 U10496 ( .B1(n10159), .B2(P2_REG0_REG_30__SCAN_IN), .A(n9016), .ZN(
        n9017) );
  OAI21_X1 U10497 ( .B1(n9018), .B2(n9100), .A(n9017), .ZN(P2_U3457) );
  INV_X1 U10498 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9020) );
  MUX2_X1 U10499 ( .A(n9020), .B(n9019), .S(n10157), .Z(n9023) );
  NAND2_X1 U10500 ( .A1(n9021), .A2(n9094), .ZN(n9022) );
  OAI211_X1 U10501 ( .C1(n9024), .C2(n9102), .A(n9023), .B(n9022), .ZN(
        P2_U3454) );
  INV_X1 U10502 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9026) );
  MUX2_X1 U10503 ( .A(n9026), .B(n9025), .S(n10157), .Z(n9029) );
  NAND2_X1 U10504 ( .A1(n9027), .A2(n9094), .ZN(n9028) );
  OAI211_X1 U10505 ( .C1(n9030), .C2(n9102), .A(n9029), .B(n9028), .ZN(
        P2_U3453) );
  INV_X1 U10506 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9032) );
  MUX2_X1 U10507 ( .A(n9032), .B(n9031), .S(n10157), .Z(n9035) );
  NAND2_X1 U10508 ( .A1(n9033), .A2(n9094), .ZN(n9034) );
  OAI211_X1 U10509 ( .C1(n9036), .C2(n9102), .A(n9035), .B(n9034), .ZN(
        P2_U3452) );
  INV_X1 U10510 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9038) );
  MUX2_X1 U10511 ( .A(n9038), .B(n9037), .S(n10157), .Z(n9042) );
  AOI22_X1 U10512 ( .A1(n9040), .A2(n9095), .B1(n9094), .B2(n9039), .ZN(n9041)
         );
  NAND2_X1 U10513 ( .A1(n9042), .A2(n9041), .ZN(P2_U3451) );
  MUX2_X1 U10514 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9043), .S(n10157), .Z(
        n9047) );
  OAI22_X1 U10515 ( .A1(n9045), .A2(n9102), .B1(n9044), .B2(n9100), .ZN(n9046)
         );
  OR2_X1 U10516 ( .A1(n9047), .A2(n9046), .ZN(P2_U3450) );
  INV_X1 U10517 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9049) );
  MUX2_X1 U10518 ( .A(n9049), .B(n9048), .S(n10157), .Z(n9053) );
  AOI22_X1 U10519 ( .A1(n9051), .A2(n9095), .B1(n9094), .B2(n9050), .ZN(n9052)
         );
  NAND2_X1 U10520 ( .A1(n9053), .A2(n9052), .ZN(P2_U3449) );
  INV_X1 U10521 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9055) );
  MUX2_X1 U10522 ( .A(n9055), .B(n9054), .S(n10157), .Z(n9058) );
  NAND2_X1 U10523 ( .A1(n9056), .A2(n9094), .ZN(n9057) );
  OAI211_X1 U10524 ( .C1(n9059), .C2(n9102), .A(n9058), .B(n9057), .ZN(
        P2_U3448) );
  INV_X1 U10525 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9061) );
  MUX2_X1 U10526 ( .A(n9061), .B(n9060), .S(n10157), .Z(n9065) );
  AOI22_X1 U10527 ( .A1(n9063), .A2(n9095), .B1(n9094), .B2(n9062), .ZN(n9064)
         );
  NAND2_X1 U10528 ( .A1(n9065), .A2(n9064), .ZN(P2_U3447) );
  INV_X1 U10529 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9067) );
  MUX2_X1 U10530 ( .A(n9067), .B(n9066), .S(n10157), .Z(n9070) );
  NAND2_X1 U10531 ( .A1(n9068), .A2(n9094), .ZN(n9069) );
  OAI211_X1 U10532 ( .C1(n9071), .C2(n9102), .A(n9070), .B(n9069), .ZN(
        P2_U3446) );
  INV_X1 U10533 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9073) );
  MUX2_X1 U10534 ( .A(n9073), .B(n9072), .S(n10157), .Z(n9074) );
  OAI21_X1 U10535 ( .B1(n9075), .B2(n9102), .A(n9074), .ZN(P2_U3444) );
  INV_X1 U10536 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10404) );
  MUX2_X1 U10537 ( .A(n9076), .B(n10404), .S(n10159), .Z(n9079) );
  NAND2_X1 U10538 ( .A1(n9077), .A2(n9094), .ZN(n9078) );
  OAI211_X1 U10539 ( .C1(n9080), .C2(n9102), .A(n9079), .B(n9078), .ZN(
        P2_U3441) );
  INV_X1 U10540 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9082) );
  MUX2_X1 U10541 ( .A(n9082), .B(n9081), .S(n10157), .Z(n9085) );
  NAND2_X1 U10542 ( .A1(n9083), .A2(n9094), .ZN(n9084) );
  OAI211_X1 U10543 ( .C1(n9086), .C2(n9102), .A(n9085), .B(n9084), .ZN(
        P2_U3438) );
  MUX2_X1 U10544 ( .A(n9087), .B(P2_REG0_REG_15__SCAN_IN), .S(n10159), .Z(
        n9091) );
  OAI22_X1 U10545 ( .A1(n9089), .A2(n9102), .B1(n9088), .B2(n9100), .ZN(n9090)
         );
  OR2_X1 U10546 ( .A1(n9091), .A2(n9090), .ZN(P2_U3435) );
  INV_X1 U10547 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U10548 ( .A(n10226), .B(n9092), .S(n10157), .Z(n9098) );
  AOI22_X1 U10549 ( .A1(n9096), .A2(n9095), .B1(n9094), .B2(n9093), .ZN(n9097)
         );
  NAND2_X1 U10550 ( .A1(n9098), .A2(n9097), .ZN(P2_U3432) );
  MUX2_X1 U10551 ( .A(n9099), .B(P2_REG0_REG_13__SCAN_IN), .S(n10159), .Z(
        n9105) );
  OAI22_X1 U10552 ( .A1(n9103), .A2(n9102), .B1(n9101), .B2(n9100), .ZN(n9104)
         );
  OR2_X1 U10553 ( .A1(n9105), .A2(n9104), .ZN(P2_U3429) );
  MUX2_X1 U10554 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9106), .S(n10157), .Z(
        P2_U3426) );
  MUX2_X1 U10555 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9107), .S(n10157), .Z(
        P2_U3423) );
  MUX2_X1 U10556 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n9108), .S(n10157), .Z(
        P2_U3420) );
  INV_X1 U10557 ( .A(n9109), .ZN(n9930) );
  NOR4_X1 U10558 ( .A1(n9110), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9111), .ZN(n9112) );
  AOI21_X1 U10559 ( .B1(n9121), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9112), .ZN(
        n9113) );
  OAI21_X1 U10560 ( .B1(n9930), .B2(n9132), .A(n9113), .ZN(P2_U3264) );
  AOI22_X1 U10561 ( .A1(n4393), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9121), .ZN(n9115) );
  OAI21_X1 U10562 ( .B1(n9116), .B2(n9132), .A(n9115), .ZN(P2_U3265) );
  INV_X1 U10563 ( .A(n9117), .ZN(n9931) );
  AOI22_X1 U10564 ( .A1(n9118), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9121), .ZN(n9119) );
  OAI21_X1 U10565 ( .B1(n9931), .B2(n9132), .A(n9119), .ZN(P2_U3266) );
  AOI21_X1 U10566 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9121), .A(n9120), .ZN(
        n9122) );
  OAI21_X1 U10567 ( .B1(n9123), .B2(n9132), .A(n9122), .ZN(P2_U3267) );
  INV_X1 U10568 ( .A(n9124), .ZN(n9933) );
  OAI222_X1 U10569 ( .A1(n4387), .A2(P2_U3151), .B1(n9132), .B2(n9933), .C1(
        n10431), .C2(n9130), .ZN(P2_U3268) );
  INV_X1 U10570 ( .A(n9126), .ZN(n9938) );
  OAI222_X1 U10571 ( .A1(n9128), .A2(P2_U3151), .B1(n9132), .B2(n9938), .C1(
        n9127), .C2(n9130), .ZN(P2_U3269) );
  INV_X1 U10572 ( .A(n9129), .ZN(n9942) );
  OAI222_X1 U10573 ( .A1(n9133), .A2(P2_U3151), .B1(n9132), .B2(n9942), .C1(
        n9131), .C2(n9130), .ZN(P2_U3270) );
  MUX2_X1 U10574 ( .A(n9134), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  XNOR2_X1 U10575 ( .A(n9242), .B(n9135), .ZN(n9136) );
  NAND2_X1 U10576 ( .A1(n9136), .A2(n9137), .ZN(n9240) );
  OAI21_X1 U10577 ( .B1(n9137), .B2(n9136), .A(n9240), .ZN(n9138) );
  NAND2_X1 U10578 ( .A1(n9138), .A2(n9359), .ZN(n9143) );
  AND2_X1 U10579 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9455) );
  INV_X1 U10580 ( .A(n9737), .ZN(n9140) );
  OAI22_X1 U10581 ( .A1(n9140), .A2(n9350), .B1(n9349), .B2(n9139), .ZN(n9141)
         );
  AOI211_X1 U10582 ( .C1(n9365), .C2(n9891), .A(n9455), .B(n9141), .ZN(n9142)
         );
  OAI211_X1 U10583 ( .C1(n9895), .C2(n9368), .A(n9143), .B(n9142), .ZN(
        P1_U3215) );
  NAND2_X1 U10584 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  OAI22_X1 U10585 ( .A1(n9598), .A2(n9376), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9147), .ZN(n9150) );
  INV_X1 U10586 ( .A(n9595), .ZN(n9148) );
  OAI22_X1 U10587 ( .A1(n9834), .A2(n9349), .B1(n9148), .B2(n9350), .ZN(n9149)
         );
  AOI211_X1 U10588 ( .C1(n9600), .C2(n9378), .A(n9150), .B(n9149), .ZN(n9151)
         );
  OAI21_X1 U10589 ( .B1(n9152), .B2(n9380), .A(n9151), .ZN(P1_U3216) );
  INV_X1 U10590 ( .A(n9153), .ZN(n9154) );
  NAND2_X1 U10591 ( .A1(n9155), .A2(n9154), .ZN(n9323) );
  OAI21_X1 U10592 ( .B1(n9155), .B2(n9154), .A(n9323), .ZN(n9156) );
  NOR2_X1 U10593 ( .A1(n9156), .A2(n9157), .ZN(n9325) );
  AOI21_X1 U10594 ( .B1(n9157), .B2(n9156), .A(n9325), .ZN(n9163) );
  AOI22_X1 U10595 ( .A1(n9373), .A2(n9158), .B1(n9365), .B2(n9385), .ZN(n9162)
         );
  OAI21_X1 U10596 ( .B1(n9349), .B2(n10039), .A(n9159), .ZN(n9160) );
  AOI21_X1 U10597 ( .B1(n9378), .B2(n10062), .A(n9160), .ZN(n9161) );
  OAI211_X1 U10598 ( .C1(n9163), .C2(n9380), .A(n9162), .B(n9161), .ZN(
        P1_U3217) );
  INV_X1 U10599 ( .A(n9165), .ZN(n9166) );
  NAND2_X1 U10600 ( .A1(n4720), .A2(n9166), .ZN(n9167) );
  OAI21_X1 U10601 ( .B1(n4720), .B2(n9166), .A(n9167), .ZN(n9347) );
  NOR2_X1 U10602 ( .A1(n9347), .A2(n9348), .ZN(n9346) );
  INV_X1 U10603 ( .A(n9167), .ZN(n9168) );
  NOR3_X1 U10604 ( .A1(n9346), .A2(n9169), .A3(n9168), .ZN(n9170) );
  OAI21_X1 U10605 ( .B1(n9170), .B2(n4469), .A(n9359), .ZN(n9174) );
  NOR2_X1 U10606 ( .A1(n9171), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9505) );
  OAI22_X1 U10607 ( .A1(n9833), .A2(n9376), .B1(n9652), .B2(n9350), .ZN(n9172)
         );
  AOI211_X1 U10608 ( .C1(n9372), .C2(n9850), .A(n9505), .B(n9172), .ZN(n9173)
         );
  OAI211_X1 U10609 ( .C1(n9854), .C2(n9368), .A(n9174), .B(n9173), .ZN(
        P1_U3219) );
  NAND2_X1 U10610 ( .A1(n5391), .A2(n9175), .ZN(n9178) );
  OR2_X1 U10611 ( .A1(n9777), .A2(n9176), .ZN(n9177) );
  NAND2_X1 U10612 ( .A1(n9178), .A2(n9177), .ZN(n9180) );
  XNOR2_X1 U10613 ( .A(n9180), .B(n9179), .ZN(n9185) );
  NAND2_X1 U10614 ( .A1(n5391), .A2(n9181), .ZN(n9182) );
  OAI21_X1 U10615 ( .B1(n9777), .B2(n4647), .A(n9182), .ZN(n9184) );
  XNOR2_X1 U10616 ( .A(n9185), .B(n9184), .ZN(n9193) );
  NOR2_X1 U10617 ( .A1(n9186), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9187) );
  AOI21_X1 U10618 ( .B1(n9383), .B2(n9365), .A(n9187), .ZN(n9188) );
  OAI21_X1 U10619 ( .B1(n9798), .B2(n9349), .A(n9188), .ZN(n9191) );
  NOR2_X1 U10620 ( .A1(n9189), .A2(n9368), .ZN(n9190) );
  AOI211_X1 U10621 ( .C1(n9373), .C2(n9525), .A(n9191), .B(n9190), .ZN(n9194)
         );
  NOR2_X1 U10622 ( .A1(n9196), .A2(n9195), .ZN(n9287) );
  AOI21_X1 U10623 ( .B1(n9196), .B2(n9195), .A(n9287), .ZN(n9197) );
  NAND2_X1 U10624 ( .A1(n9197), .A2(n9198), .ZN(n9291) );
  OAI21_X1 U10625 ( .B1(n9198), .B2(n9197), .A(n9291), .ZN(n9206) );
  AOI22_X1 U10626 ( .A1(n9373), .A2(n9199), .B1(n9365), .B2(n9386), .ZN(n9203)
         );
  INV_X1 U10627 ( .A(n9200), .ZN(n9201) );
  AOI21_X1 U10628 ( .B1(n9372), .B2(n9387), .A(n9201), .ZN(n9202) );
  OAI211_X1 U10629 ( .C1(n9204), .C2(n9368), .A(n9203), .B(n9202), .ZN(n9205)
         );
  AOI21_X1 U10630 ( .B1(n9206), .B2(n9359), .A(n9205), .ZN(n9207) );
  INV_X1 U10631 ( .A(n9207), .ZN(P1_U3221) );
  NOR2_X1 U10632 ( .A1(n9209), .A2(n9208), .ZN(n9211) );
  OAI21_X1 U10633 ( .B1(n9211), .B2(n9210), .A(n9359), .ZN(n9215) );
  AOI22_X1 U10634 ( .A1(n9372), .A2(n6578), .B1(n9365), .B2(n5407), .ZN(n9214)
         );
  AOI22_X1 U10635 ( .A1(n9378), .A2(n5848), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9341), .ZN(n9213) );
  NAND3_X1 U10636 ( .A1(n9215), .A2(n9214), .A3(n9213), .ZN(P1_U3222) );
  OAI21_X1 U10637 ( .B1(n9218), .B2(n9217), .A(n9216), .ZN(n9219) );
  NAND2_X1 U10638 ( .A1(n9219), .A2(n9359), .ZN(n9223) );
  AOI22_X1 U10639 ( .A1(n9815), .A2(n9365), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9222) );
  AOI22_X1 U10640 ( .A1(n9373), .A2(n9623), .B1(n9372), .B2(n9851), .ZN(n9221)
         );
  NAND2_X1 U10641 ( .A1(n9837), .A2(n9378), .ZN(n9220) );
  NAND4_X1 U10642 ( .A1(n9223), .A2(n9222), .A3(n9221), .A4(n9220), .ZN(
        P1_U3223) );
  XOR2_X1 U10643 ( .A(n9225), .B(n9224), .Z(n9231) );
  AOI22_X1 U10644 ( .A1(n9373), .A2(n9226), .B1(n9365), .B2(n9892), .ZN(n9228)
         );
  OAI211_X1 U10645 ( .C1(n10083), .C2(n9349), .A(n9228), .B(n9227), .ZN(n9229)
         );
  AOI21_X1 U10646 ( .B1(n10079), .B2(n9378), .A(n9229), .ZN(n9230) );
  OAI21_X1 U10647 ( .B1(n9231), .B2(n9380), .A(n9230), .ZN(P1_U3224) );
  INV_X1 U10648 ( .A(n9808), .ZN(n9568) );
  OAI21_X1 U10649 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9235) );
  NAND2_X1 U10650 ( .A1(n9235), .A2(n9359), .ZN(n9239) );
  AOI22_X1 U10651 ( .A1(n9816), .A2(n9372), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9236) );
  OAI21_X1 U10652 ( .B1(n9564), .B2(n9350), .A(n9236), .ZN(n9237) );
  AOI21_X1 U10653 ( .B1(n9788), .B2(n9365), .A(n9237), .ZN(n9238) );
  OAI211_X1 U10654 ( .C1(n9568), .C2(n9368), .A(n9239), .B(n9238), .ZN(
        P1_U3225) );
  INV_X1 U10655 ( .A(n9243), .ZN(n9245) );
  OAI21_X1 U10656 ( .B1(n9242), .B2(n9241), .A(n9240), .ZN(n9244) );
  XOR2_X1 U10657 ( .A(n9243), .B(n9244), .Z(n9371) );
  NOR2_X1 U10658 ( .A1(n9371), .A2(n9370), .ZN(n9369) );
  AOI21_X1 U10659 ( .B1(n9245), .B2(n9244), .A(n9369), .ZN(n9249) );
  XNOR2_X1 U10660 ( .A(n9247), .B(n9246), .ZN(n9248) );
  XNOR2_X1 U10661 ( .A(n9249), .B(n9248), .ZN(n9253) );
  AOI22_X1 U10662 ( .A1(n9708), .A2(n9373), .B1(n9372), .B2(n9891), .ZN(n9250)
         );
  NAND2_X1 U10663 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9472) );
  OAI211_X1 U10664 ( .C1(n9874), .C2(n9376), .A(n9250), .B(n9472), .ZN(n9251)
         );
  AOI21_X1 U10665 ( .B1(n9877), .B2(n9378), .A(n9251), .ZN(n9252) );
  OAI21_X1 U10666 ( .B1(n9253), .B2(n9380), .A(n9252), .ZN(P1_U3226) );
  OAI21_X1 U10667 ( .B1(n9256), .B2(n9255), .A(n9254), .ZN(n9257) );
  NAND2_X1 U10668 ( .A1(n9257), .A2(n9359), .ZN(n9266) );
  OAI21_X1 U10669 ( .B1(n9259), .B2(n9258), .A(P1_STATE_REG_SCAN_IN), .ZN(
        n9264) );
  NOR3_X1 U10670 ( .A1(n9350), .A2(P1_REG3_REG_17__SCAN_IN), .A3(n9260), .ZN(
        n9263) );
  OAI22_X1 U10671 ( .A1(n9376), .A2(n9261), .B1(n9349), .B2(n9725), .ZN(n9262)
         );
  AOI211_X1 U10672 ( .C1(P1_REG3_REG_17__SCAN_IN), .C2(n9264), .A(n9263), .B(
        n9262), .ZN(n9265) );
  OAI211_X1 U10673 ( .C1(n5866), .C2(n9368), .A(n9266), .B(n9265), .ZN(
        P1_U3228) );
  INV_X1 U10674 ( .A(n9812), .ZN(n9583) );
  OAI21_X1 U10675 ( .B1(n9269), .B2(n9268), .A(n9267), .ZN(n9270) );
  NAND2_X1 U10676 ( .A1(n9270), .A2(n9359), .ZN(n9274) );
  NOR2_X1 U10677 ( .A1(n9613), .A2(n9349), .ZN(n9272) );
  OAI22_X1 U10678 ( .A1(n9797), .A2(n9376), .B1(n9350), .B2(n9585), .ZN(n9271)
         );
  AOI211_X1 U10679 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n9272), 
        .B(n9271), .ZN(n9273) );
  OAI211_X1 U10680 ( .C1(n9583), .C2(n9368), .A(n9274), .B(n9273), .ZN(
        P1_U3229) );
  INV_X1 U10681 ( .A(n9275), .ZN(n9279) );
  OAI21_X1 U10682 ( .B1(n7888), .B2(n9277), .A(n9276), .ZN(n9278) );
  NAND3_X1 U10683 ( .A1(n9279), .A2(n9359), .A3(n9278), .ZN(n9285) );
  AOI22_X1 U10684 ( .A1(n9280), .A2(n9373), .B1(n9372), .B2(n9390), .ZN(n9284)
         );
  AND2_X1 U10685 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9435) );
  NOR2_X1 U10686 ( .A1(n9368), .A2(n9281), .ZN(n9282) );
  AOI211_X1 U10687 ( .C1(n9365), .C2(n7873), .A(n9435), .B(n9282), .ZN(n9283)
         );
  NAND3_X1 U10688 ( .A1(n9285), .A2(n9284), .A3(n9283), .ZN(P1_U3230) );
  NOR2_X1 U10689 ( .A1(n9287), .A2(n9286), .ZN(n9290) );
  INV_X1 U10690 ( .A(n9288), .ZN(n9289) );
  AOI21_X1 U10691 ( .B1(n9291), .B2(n9290), .A(n9289), .ZN(n9298) );
  AOI22_X1 U10692 ( .A1(n9373), .A2(n9292), .B1(n9365), .B2(n9987), .ZN(n9297)
         );
  OAI21_X1 U10693 ( .B1(n9349), .B2(n9294), .A(n9293), .ZN(n9295) );
  AOI21_X1 U10694 ( .B1(n9378), .B2(n10054), .A(n9295), .ZN(n9296) );
  OAI211_X1 U10695 ( .C1(n9298), .C2(n9380), .A(n9297), .B(n9296), .ZN(
        P1_U3231) );
  NOR2_X1 U10696 ( .A1(n4497), .A2(n9299), .ZN(n9300) );
  XNOR2_X1 U10697 ( .A(n9301), .B(n9300), .ZN(n9305) );
  OAI22_X1 U10698 ( .A1(n9860), .A2(n9349), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10314), .ZN(n9303) );
  OAI22_X1 U10699 ( .A1(n9842), .A2(n9376), .B1(n9636), .B2(n9350), .ZN(n9302)
         );
  AOI211_X1 U10700 ( .C1(n9845), .C2(n9378), .A(n9303), .B(n9302), .ZN(n9304)
         );
  OAI21_X1 U10701 ( .B1(n9305), .B2(n9380), .A(n9304), .ZN(P1_U3233) );
  XOR2_X1 U10702 ( .A(n9307), .B(n9306), .Z(n9312) );
  AOI22_X1 U10703 ( .A1(n9373), .A2(n9760), .B1(n9365), .B2(n9882), .ZN(n9309)
         );
  OAI211_X1 U10704 ( .C1(n9757), .C2(n9349), .A(n9309), .B(n9308), .ZN(n9310)
         );
  AOI21_X1 U10705 ( .B1(n9902), .B2(n9378), .A(n9310), .ZN(n9311) );
  OAI21_X1 U10706 ( .B1(n9312), .B2(n9380), .A(n9311), .ZN(P1_U3234) );
  NAND2_X1 U10707 ( .A1(n9314), .A2(n9313), .ZN(n9316) );
  XNOR2_X1 U10708 ( .A(n9316), .B(n9315), .ZN(n9322) );
  OAI22_X1 U10709 ( .A1(n9613), .A2(n9376), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9317), .ZN(n9319) );
  OAI22_X1 U10710 ( .A1(n9842), .A2(n9349), .B1(n9612), .B2(n9350), .ZN(n9318)
         );
  AOI211_X1 U10711 ( .C1(n9320), .C2(n9378), .A(n9319), .B(n9318), .ZN(n9321)
         );
  OAI21_X1 U10712 ( .B1(n9322), .B2(n9380), .A(n9321), .ZN(P1_U3235) );
  INV_X1 U10713 ( .A(n9323), .ZN(n9324) );
  NOR2_X1 U10714 ( .A1(n9325), .A2(n9324), .ZN(n9328) );
  NOR2_X1 U10715 ( .A1(n9326), .A2(n4507), .ZN(n9327) );
  XNOR2_X1 U10716 ( .A(n9328), .B(n9327), .ZN(n9335) );
  AOI22_X1 U10717 ( .A1(n9373), .A2(n9992), .B1(n9365), .B2(n9985), .ZN(n9330)
         );
  OAI211_X1 U10718 ( .C1(n9331), .C2(n9349), .A(n9330), .B(n9329), .ZN(n9332)
         );
  AOI21_X1 U10719 ( .B1(n9333), .B2(n9378), .A(n9332), .ZN(n9334) );
  OAI21_X1 U10720 ( .B1(n9335), .B2(n9380), .A(n9334), .ZN(P1_U3236) );
  INV_X1 U10721 ( .A(n9336), .ZN(n9340) );
  NOR3_X1 U10722 ( .A1(n9210), .A2(n9338), .A3(n9337), .ZN(n9339) );
  OAI21_X1 U10723 ( .B1(n9340), .B2(n9339), .A(n9359), .ZN(n9345) );
  AOI22_X1 U10724 ( .A1(n9372), .A2(n4646), .B1(n9365), .B2(n9390), .ZN(n9344)
         );
  AOI22_X1 U10725 ( .A1(n9378), .A2(n9342), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9341), .ZN(n9343) );
  NAND3_X1 U10726 ( .A1(n9345), .A2(n9344), .A3(n9343), .ZN(P1_U3237) );
  AOI21_X1 U10727 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9354) );
  NAND2_X1 U10728 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9969) );
  OAI21_X1 U10729 ( .B1(n9349), .B2(n9874), .A(n9969), .ZN(n9352) );
  OAI22_X1 U10730 ( .A1(n9376), .A2(n9860), .B1(n9672), .B2(n9350), .ZN(n9351)
         );
  AOI211_X1 U10731 ( .C1(n9863), .C2(n9378), .A(n9352), .B(n9351), .ZN(n9353)
         );
  OAI21_X1 U10732 ( .B1(n9354), .B2(n9380), .A(n9353), .ZN(P1_U3238) );
  INV_X1 U10733 ( .A(n9232), .ZN(n9357) );
  OAI21_X1 U10734 ( .B1(n9357), .B2(n9356), .A(n9355), .ZN(n9360) );
  NAND3_X1 U10735 ( .A1(n9360), .A2(n9359), .A3(n9358), .ZN(n9367) );
  NAND2_X1 U10736 ( .A1(n9577), .A2(n9372), .ZN(n9362) );
  NAND2_X1 U10737 ( .A1(n9548), .A2(n9373), .ZN(n9361) );
  OAI211_X1 U10738 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9363), .A(n9362), .B(
        n9361), .ZN(n9364) );
  AOI21_X1 U10739 ( .B1(n9384), .B2(n9365), .A(n9364), .ZN(n9366) );
  OAI211_X1 U10740 ( .C1(n9547), .C2(n9368), .A(n9367), .B(n9366), .ZN(
        P1_U3240) );
  AOI21_X1 U10741 ( .B1(n9371), .B2(n9370), .A(n9369), .ZN(n9381) );
  AOI22_X1 U10742 ( .A1(n9722), .A2(n9373), .B1(n9372), .B2(n9882), .ZN(n9375)
         );
  NAND2_X1 U10743 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9955) );
  OAI211_X1 U10744 ( .C1(n9725), .C2(n9376), .A(n9375), .B(n9955), .ZN(n9377)
         );
  AOI21_X1 U10745 ( .B1(n5860), .B2(n9378), .A(n9377), .ZN(n9379) );
  OAI21_X1 U10746 ( .B1(n9381), .B2(n9380), .A(n9379), .ZN(P1_U3241) );
  MUX2_X1 U10747 ( .A(n9382), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9391), .Z(
        P1_U3584) );
  MUX2_X1 U10748 ( .A(n9383), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9391), .Z(
        P1_U3583) );
  MUX2_X1 U10749 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9789), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10750 ( .A(n9384), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9391), .Z(
        P1_U3581) );
  MUX2_X1 U10751 ( .A(n9788), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9391), .Z(
        P1_U3580) );
  MUX2_X1 U10752 ( .A(n9577), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9391), .Z(
        P1_U3579) );
  MUX2_X1 U10753 ( .A(n9816), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9391), .Z(
        P1_U3578) );
  MUX2_X1 U10754 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9825), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10755 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9815), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10756 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9824), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10757 ( .A(n9851), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9391), .Z(
        P1_U3574) );
  MUX2_X1 U10758 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9638), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10759 ( .A(n9850), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9391), .Z(
        P1_U3572) );
  MUX2_X1 U10760 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9675), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10761 ( .A(n9883), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9391), .Z(
        P1_U3570) );
  MUX2_X1 U10762 ( .A(n9891), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9391), .Z(
        P1_U3569) );
  MUX2_X1 U10763 ( .A(n9882), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9391), .Z(
        P1_U3568) );
  MUX2_X1 U10764 ( .A(n9892), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9391), .Z(
        P1_U3567) );
  MUX2_X1 U10765 ( .A(n9985), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9391), .Z(
        P1_U3566) );
  MUX2_X1 U10766 ( .A(n9385), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9391), .Z(
        P1_U3565) );
  MUX2_X1 U10767 ( .A(n9987), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9391), .Z(
        P1_U3564) );
  MUX2_X1 U10768 ( .A(n9386), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9391), .Z(
        P1_U3563) );
  MUX2_X1 U10769 ( .A(n10052), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9391), .Z(
        P1_U3562) );
  MUX2_X1 U10770 ( .A(n9387), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9391), .Z(
        P1_U3561) );
  MUX2_X1 U10771 ( .A(n9388), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9391), .Z(
        P1_U3560) );
  MUX2_X1 U10772 ( .A(n7873), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9391), .Z(
        P1_U3559) );
  MUX2_X1 U10773 ( .A(n9389), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9391), .Z(
        P1_U3558) );
  MUX2_X1 U10774 ( .A(n9390), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9391), .Z(
        P1_U3557) );
  MUX2_X1 U10775 ( .A(n5407), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9391), .Z(
        P1_U3556) );
  MUX2_X1 U10776 ( .A(n4646), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9391), .Z(
        P1_U3555) );
  INV_X1 U10777 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9393) );
  OAI22_X1 U10778 ( .A1(n9972), .A2(n9393), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9392), .ZN(n9394) );
  AOI21_X1 U10779 ( .B1(n4632), .B2(n9968), .A(n9394), .ZN(n9402) );
  OAI211_X1 U10780 ( .C1(n9397), .C2(n9396), .A(n9502), .B(n9395), .ZN(n9401)
         );
  OAI211_X1 U10781 ( .C1(n9399), .C2(n9404), .A(n9496), .B(n9398), .ZN(n9400)
         );
  NAND3_X1 U10782 ( .A1(n9402), .A2(n9401), .A3(n9400), .ZN(P1_U3244) );
  MUX2_X1 U10783 ( .A(n9404), .B(n9403), .S(n9935), .Z(n9406) );
  NAND2_X1 U10784 ( .A1(n9406), .A2(n9405), .ZN(n9407) );
  OAI211_X1 U10785 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9408), .A(n9407), .B(
        P1_U3973), .ZN(n9449) );
  INV_X1 U10786 ( .A(n4728), .ZN(n9412) );
  INV_X1 U10787 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9410) );
  OAI22_X1 U10788 ( .A1(n9972), .A2(n9410), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9409), .ZN(n9411) );
  AOI21_X1 U10789 ( .B1(n9412), .B2(n9968), .A(n9411), .ZN(n9421) );
  OAI211_X1 U10790 ( .C1(n9415), .C2(n9414), .A(n9496), .B(n9413), .ZN(n9420)
         );
  OAI211_X1 U10791 ( .C1(n9418), .C2(n9417), .A(n9502), .B(n9416), .ZN(n9419)
         );
  NAND4_X1 U10792 ( .A1(n9449), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(
        P1_U3245) );
  INV_X1 U10793 ( .A(n9422), .ZN(n9425) );
  INV_X1 U10794 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10289) );
  OAI21_X1 U10795 ( .B1(n9972), .B2(n10289), .A(n9423), .ZN(n9424) );
  AOI21_X1 U10796 ( .B1(n9425), .B2(n9968), .A(n9424), .ZN(n9434) );
  OAI211_X1 U10797 ( .C1(n9428), .C2(n9427), .A(n9496), .B(n9426), .ZN(n9433)
         );
  OAI211_X1 U10798 ( .C1(n9431), .C2(n9430), .A(n9502), .B(n9429), .ZN(n9432)
         );
  NAND3_X1 U10799 ( .A1(n9434), .A2(n9433), .A3(n9432), .ZN(P1_U3246) );
  AOI21_X1 U10800 ( .B1(n9506), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9435), .ZN(
        n9448) );
  INV_X1 U10801 ( .A(n9436), .ZN(n9437) );
  OAI211_X1 U10802 ( .C1(n9439), .C2(n9438), .A(n9502), .B(n9437), .ZN(n9444)
         );
  OAI211_X1 U10803 ( .C1(n9442), .C2(n9441), .A(n9496), .B(n9440), .ZN(n9443)
         );
  AND2_X1 U10804 ( .A1(n9444), .A2(n9443), .ZN(n9447) );
  NAND2_X1 U10805 ( .A1(n9968), .A2(n9445), .ZN(n9446) );
  NAND4_X1 U10806 ( .A1(n9449), .A2(n9448), .A3(n9447), .A4(n9446), .ZN(
        P1_U3247) );
  XNOR2_X1 U10807 ( .A(n9466), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n9450) );
  AOI211_X1 U10808 ( .C1(n9451), .C2(n9450), .A(n9963), .B(n9465), .ZN(n9461)
         );
  XNOR2_X1 U10809 ( .A(n9466), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9454) );
  AOI211_X1 U10810 ( .C1(n4540), .C2(n9454), .A(n9959), .B(n9463), .ZN(n9460)
         );
  NAND2_X1 U10811 ( .A1(n9968), .A2(n9466), .ZN(n9457) );
  INV_X1 U10812 ( .A(n9455), .ZN(n9456) );
  OAI211_X1 U10813 ( .C1(n9458), .C2(n9972), .A(n9457), .B(n9456), .ZN(n9459)
         );
  OR3_X1 U10814 ( .A1(n9461), .A2(n9460), .A3(n9459), .ZN(P1_U3257) );
  INV_X1 U10815 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9462) );
  XNOR2_X1 U10816 ( .A(n9485), .B(n9462), .ZN(n9484) );
  XNOR2_X1 U10817 ( .A(n9484), .B(n9483), .ZN(n9475) );
  INV_X1 U10818 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9473) );
  INV_X1 U10819 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9946) );
  XNOR2_X1 U10820 ( .A(n9485), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9468) );
  AOI211_X1 U10821 ( .C1(n9469), .C2(n9468), .A(n4485), .B(n9963), .ZN(n9470)
         );
  INV_X1 U10822 ( .A(n9470), .ZN(n9471) );
  OAI211_X1 U10823 ( .C1(n9972), .C2(n9473), .A(n9472), .B(n9471), .ZN(n9474)
         );
  AOI21_X1 U10824 ( .B1(n9502), .B2(n9475), .A(n9474), .ZN(n9476) );
  OAI21_X1 U10825 ( .B1(n9477), .B2(n4733), .A(n9476), .ZN(P1_U3259) );
  OAI22_X1 U10826 ( .A1(n9972), .A2(n10487), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10413), .ZN(n9491) );
  XNOR2_X1 U10827 ( .A(n9499), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9481) );
  AND2_X1 U10828 ( .A1(n9485), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9478) );
  INV_X1 U10829 ( .A(n9494), .ZN(n9479) );
  AOI21_X1 U10830 ( .B1(n9481), .B2(n9480), .A(n9479), .ZN(n9489) );
  INV_X1 U10831 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9482) );
  XNOR2_X1 U10832 ( .A(n9499), .B(n9482), .ZN(n9497) );
  OR2_X1 U10833 ( .A1(n9485), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9486) );
  XOR2_X1 U10834 ( .A(n9497), .B(n9498), .Z(n9488) );
  OAI22_X1 U10835 ( .A1(n9489), .A2(n9963), .B1(n9959), .B2(n9488), .ZN(n9490)
         );
  AOI211_X1 U10836 ( .C1(n9499), .C2(n9968), .A(n9491), .B(n9490), .ZN(n9492)
         );
  INV_X1 U10837 ( .A(n9492), .ZN(P1_U3260) );
  OR2_X1 U10838 ( .A1(n9499), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U10839 ( .A1(n9967), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9495) );
  OAI21_X1 U10840 ( .B1(n9967), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9495), .ZN(
        n9966) );
  NAND2_X1 U10841 ( .A1(n9967), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9500) );
  OAI21_X1 U10842 ( .B1(n9967), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9500), .ZN(
        n9961) );
  NAND2_X1 U10843 ( .A1(n9958), .A2(n9500), .ZN(n9501) );
  NOR2_X1 U10844 ( .A1(n4418), .A2(n9507), .ZN(n9508) );
  XNOR2_X1 U10845 ( .A(n9509), .B(n9508), .ZN(n9769) );
  NAND2_X1 U10846 ( .A1(n9511), .A2(n9510), .ZN(n9770) );
  NOR2_X1 U10847 ( .A1(n9993), .A2(n9770), .ZN(n9517) );
  AOI21_X1 U10848 ( .B1(n9993), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9517), .ZN(
        n9513) );
  NAND2_X1 U10849 ( .A1(n9766), .A2(n9747), .ZN(n9512) );
  OAI211_X1 U10850 ( .C1(n9769), .C2(n9514), .A(n9513), .B(n9512), .ZN(
        P1_U3263) );
  XNOR2_X1 U10851 ( .A(n4418), .B(n9772), .ZN(n9515) );
  NAND2_X1 U10852 ( .A1(n9515), .A2(n9975), .ZN(n9771) );
  NOR2_X1 U10853 ( .A1(n9772), .A2(n9995), .ZN(n9516) );
  AOI211_X1 U10854 ( .C1(n9993), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9517), .B(
        n9516), .ZN(n9518) );
  OAI21_X1 U10855 ( .B1(n9771), .B2(n9743), .A(n9518), .ZN(P1_U3264) );
  OAI22_X1 U10856 ( .A1(n9521), .A2(n9741), .B1(n9997), .B2(n9520), .ZN(n9524)
         );
  NOR2_X1 U10857 ( .A1(n9798), .A2(n9522), .ZN(n9523) );
  AOI211_X1 U10858 ( .C1(n9991), .C2(n9525), .A(n9524), .B(n9523), .ZN(n9527)
         );
  NAND2_X1 U10859 ( .A1(n5391), .A2(n9747), .ZN(n9526) );
  OAI211_X1 U10860 ( .C1(n9528), .C2(n9743), .A(n9527), .B(n9526), .ZN(n9529)
         );
  AOI21_X1 U10861 ( .B1(n9519), .B2(n9704), .A(n9529), .ZN(n9530) );
  OAI21_X1 U10862 ( .B1(n9531), .B2(n9715), .A(n9530), .ZN(P1_U3265) );
  XNOR2_X1 U10863 ( .A(n9532), .B(n5833), .ZN(n9796) );
  XNOR2_X1 U10864 ( .A(n9533), .B(n5833), .ZN(n9794) );
  OAI211_X1 U10865 ( .C1(n9545), .C2(n9792), .A(n9975), .B(n9534), .ZN(n9791)
         );
  OAI22_X1 U10866 ( .A1(n9536), .A2(n9671), .B1(n9535), .B2(n9997), .ZN(n9537)
         );
  AOI21_X1 U10867 ( .B1(n9738), .B2(n9788), .A(n9537), .ZN(n9538) );
  OAI21_X1 U10868 ( .B1(n9777), .B2(n9741), .A(n9538), .ZN(n9539) );
  AOI21_X1 U10869 ( .B1(n9540), .B2(n9747), .A(n9539), .ZN(n9541) );
  OAI21_X1 U10870 ( .B1(n9791), .B2(n9743), .A(n9541), .ZN(n9542) );
  AOI21_X1 U10871 ( .B1(n9794), .B2(n9729), .A(n9542), .ZN(n9543) );
  OAI21_X1 U10872 ( .B1(n9796), .B2(n9765), .A(n9543), .ZN(P1_U3266) );
  AOI21_X1 U10873 ( .B1(n9544), .B2(n9553), .A(n4484), .ZN(n9805) );
  INV_X1 U10874 ( .A(n9563), .ZN(n9546) );
  AOI211_X1 U10875 ( .C1(n9801), .C2(n9546), .A(n9768), .B(n9545), .ZN(n9799)
         );
  NOR2_X1 U10876 ( .A1(n9547), .A2(n9995), .ZN(n9552) );
  AOI22_X1 U10877 ( .A1(n9548), .A2(n9991), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9993), .ZN(n9550) );
  NAND2_X1 U10878 ( .A1(n9577), .A2(n9738), .ZN(n9549) );
  OAI211_X1 U10879 ( .C1(n9798), .C2(n9741), .A(n9550), .B(n9549), .ZN(n9551)
         );
  AOI211_X1 U10880 ( .C1(n9799), .C2(n9977), .A(n9552), .B(n9551), .ZN(n9556)
         );
  XOR2_X1 U10881 ( .A(n9554), .B(n9553), .Z(n9802) );
  NAND2_X1 U10882 ( .A1(n9802), .A2(n9704), .ZN(n9555) );
  OAI211_X1 U10883 ( .C1(n9805), .C2(n9715), .A(n9556), .B(n9555), .ZN(
        P1_U3267) );
  XOR2_X1 U10884 ( .A(n9557), .B(n9560), .Z(n9809) );
  AOI21_X1 U10885 ( .B1(n9560), .B2(n9559), .A(n9558), .ZN(n9561) );
  OAI222_X1 U10886 ( .A1(n10065), .A2(n9562), .B1(n10082), .B2(n9598), .C1(
        n9881), .C2(n9561), .ZN(n9806) );
  AOI211_X1 U10887 ( .C1(n9808), .C2(n9581), .A(n9768), .B(n9563), .ZN(n9807)
         );
  NAND2_X1 U10888 ( .A1(n9807), .A2(n9977), .ZN(n9567) );
  INV_X1 U10889 ( .A(n9564), .ZN(n9565) );
  AOI22_X1 U10890 ( .A1(n9565), .A2(n9991), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9993), .ZN(n9566) );
  OAI211_X1 U10891 ( .C1(n9568), .C2(n9995), .A(n9567), .B(n9566), .ZN(n9569)
         );
  AOI21_X1 U10892 ( .B1(n9806), .B2(n9997), .A(n9569), .ZN(n9570) );
  OAI21_X1 U10893 ( .B1(n9809), .B2(n9765), .A(n9570), .ZN(P1_U3268) );
  XNOR2_X1 U10894 ( .A(n9572), .B(n9571), .ZN(n9814) );
  NAND2_X1 U10895 ( .A1(n9573), .A2(n10061), .ZN(n9580) );
  AOI21_X1 U10896 ( .B1(n9574), .B2(n9576), .A(n9575), .ZN(n9579) );
  AOI22_X1 U10897 ( .A1(n9577), .A2(n9986), .B1(n10053), .B2(n9825), .ZN(n9578) );
  OAI21_X1 U10898 ( .B1(n9580), .B2(n9579), .A(n9578), .ZN(n9810) );
  NAND2_X1 U10899 ( .A1(n9810), .A2(n9997), .ZN(n9589) );
  INV_X1 U10900 ( .A(n9581), .ZN(n9582) );
  AOI211_X1 U10901 ( .C1(n9812), .C2(n9594), .A(n9768), .B(n9582), .ZN(n9811)
         );
  NOR2_X1 U10902 ( .A1(n9583), .A2(n9995), .ZN(n9587) );
  OAI22_X1 U10903 ( .A1(n9585), .A2(n9671), .B1(n9584), .B2(n9997), .ZN(n9586)
         );
  AOI211_X1 U10904 ( .C1(n9811), .C2(n9977), .A(n9587), .B(n9586), .ZN(n9588)
         );
  OAI211_X1 U10905 ( .C1(n9814), .C2(n9765), .A(n9589), .B(n9588), .ZN(
        P1_U3269) );
  XNOR2_X1 U10906 ( .A(n9590), .B(n9591), .ZN(n9823) );
  OAI21_X1 U10907 ( .B1(n9592), .B2(n9591), .A(n9574), .ZN(n9821) );
  OAI211_X1 U10908 ( .C1(n9593), .C2(n9819), .A(n9975), .B(n9594), .ZN(n9818)
         );
  AOI22_X1 U10909 ( .A1(n9595), .A2(n9991), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9993), .ZN(n9597) );
  NAND2_X1 U10910 ( .A1(n9815), .A2(n9738), .ZN(n9596) );
  OAI211_X1 U10911 ( .C1(n9598), .C2(n9741), .A(n9597), .B(n9596), .ZN(n9599)
         );
  AOI21_X1 U10912 ( .B1(n9600), .B2(n9747), .A(n9599), .ZN(n9601) );
  OAI21_X1 U10913 ( .B1(n9818), .B2(n9743), .A(n9601), .ZN(n9602) );
  AOI21_X1 U10914 ( .B1(n9821), .B2(n9729), .A(n9602), .ZN(n9603) );
  OAI21_X1 U10915 ( .B1(n9823), .B2(n9765), .A(n9603), .ZN(P1_U3270) );
  XNOR2_X1 U10916 ( .A(n9606), .B(n9605), .ZN(n9832) );
  XNOR2_X1 U10917 ( .A(n9606), .B(n9607), .ZN(n9830) );
  INV_X1 U10918 ( .A(n9593), .ZN(n9609) );
  OAI211_X1 U10919 ( .C1(n9828), .C2(n9608), .A(n9609), .B(n9975), .ZN(n9827)
         );
  NOR3_X1 U10920 ( .A1(n9827), .A2(n9610), .A3(n9993), .ZN(n9618) );
  OAI22_X1 U10921 ( .A1(n9612), .A2(n9671), .B1(n9611), .B2(n9997), .ZN(n9615)
         );
  NOR2_X1 U10922 ( .A1(n9613), .A2(n9741), .ZN(n9614) );
  AOI211_X1 U10923 ( .C1(n9738), .C2(n9824), .A(n9615), .B(n9614), .ZN(n9616)
         );
  OAI21_X1 U10924 ( .B1(n9828), .B2(n9995), .A(n9616), .ZN(n9617) );
  AOI211_X1 U10925 ( .C1(n9830), .C2(n9729), .A(n9618), .B(n9617), .ZN(n9619)
         );
  OAI21_X1 U10926 ( .B1(n9765), .B2(n9832), .A(n9619), .ZN(P1_U3271) );
  XNOR2_X1 U10927 ( .A(n9620), .B(n9628), .ZN(n9841) );
  AOI211_X1 U10928 ( .C1(n9837), .C2(n9621), .A(n9768), .B(n9608), .ZN(n9835)
         );
  INV_X1 U10929 ( .A(n9837), .ZN(n9622) );
  NOR2_X1 U10930 ( .A1(n9622), .A2(n9995), .ZN(n9627) );
  AOI22_X1 U10931 ( .A1(n9623), .A2(n9991), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9993), .ZN(n9625) );
  NAND2_X1 U10932 ( .A1(n9851), .A2(n9738), .ZN(n9624) );
  OAI211_X1 U10933 ( .C1(n9834), .C2(n9741), .A(n9625), .B(n9624), .ZN(n9626)
         );
  AOI211_X1 U10934 ( .C1(n9835), .C2(n9977), .A(n9627), .B(n9626), .ZN(n9631)
         );
  XNOR2_X1 U10935 ( .A(n9629), .B(n9628), .ZN(n9838) );
  NAND2_X1 U10936 ( .A1(n9838), .A2(n9729), .ZN(n9630) );
  OAI211_X1 U10937 ( .C1(n9841), .C2(n9765), .A(n9631), .B(n9630), .ZN(
        P1_U3272) );
  XOR2_X1 U10938 ( .A(n9644), .B(n9632), .Z(n9849) );
  INV_X1 U10939 ( .A(n9621), .ZN(n9634) );
  AOI211_X1 U10940 ( .C1(n9845), .C2(n9633), .A(n9768), .B(n9634), .ZN(n9843)
         );
  INV_X1 U10941 ( .A(n9845), .ZN(n9635) );
  NOR2_X1 U10942 ( .A1(n9635), .A2(n9995), .ZN(n9642) );
  INV_X1 U10943 ( .A(n9636), .ZN(n9637) );
  AOI22_X1 U10944 ( .A1(n9637), .A2(n9991), .B1(n9993), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U10945 ( .A1(n9738), .A2(n9638), .ZN(n9639) );
  OAI211_X1 U10946 ( .C1(n9842), .C2(n9741), .A(n9640), .B(n9639), .ZN(n9641)
         );
  AOI211_X1 U10947 ( .C1(n9843), .C2(n9977), .A(n9642), .B(n9641), .ZN(n9647)
         );
  OAI21_X1 U10948 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9846) );
  NAND2_X1 U10949 ( .A1(n9846), .A2(n9729), .ZN(n9646) );
  OAI211_X1 U10950 ( .C1(n9849), .C2(n9765), .A(n9647), .B(n9646), .ZN(
        P1_U3273) );
  XOR2_X1 U10951 ( .A(n9649), .B(n9650), .Z(n9858) );
  XNOR2_X1 U10952 ( .A(n9651), .B(n9650), .ZN(n9856) );
  OAI211_X1 U10953 ( .C1(n9670), .C2(n9854), .A(n9975), .B(n9633), .ZN(n9853)
         );
  INV_X1 U10954 ( .A(n9652), .ZN(n9653) );
  AOI22_X1 U10955 ( .A1(n9993), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9653), .B2(
        n9991), .ZN(n9655) );
  NAND2_X1 U10956 ( .A1(n9738), .A2(n9850), .ZN(n9654) );
  OAI211_X1 U10957 ( .C1(n9833), .C2(n9741), .A(n9655), .B(n9654), .ZN(n9656)
         );
  AOI21_X1 U10958 ( .B1(n9657), .B2(n9747), .A(n9656), .ZN(n9658) );
  OAI21_X1 U10959 ( .B1(n9853), .B2(n9743), .A(n9658), .ZN(n9659) );
  AOI21_X1 U10960 ( .B1(n9856), .B2(n9729), .A(n9659), .ZN(n9660) );
  OAI21_X1 U10961 ( .B1(n9858), .B2(n9765), .A(n9660), .ZN(P1_U3274) );
  AOI21_X1 U10962 ( .B1(n9667), .B2(n9662), .A(n9661), .ZN(n9866) );
  OAI22_X1 U10963 ( .A1(n9682), .A2(n9665), .B1(n5866), .B2(n9874), .ZN(n9666)
         );
  XOR2_X1 U10964 ( .A(n9667), .B(n9666), .Z(n9859) );
  NAND2_X1 U10965 ( .A1(n9859), .A2(n9704), .ZN(n9680) );
  NAND2_X1 U10966 ( .A1(n9685), .A2(n9863), .ZN(n9668) );
  NAND2_X1 U10967 ( .A1(n9668), .A2(n9975), .ZN(n9669) );
  NOR2_X1 U10968 ( .A1(n9670), .A2(n9669), .ZN(n9861) );
  NAND2_X1 U10969 ( .A1(n9863), .A2(n9747), .ZN(n9677) );
  INV_X1 U10970 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9673) );
  OAI22_X1 U10971 ( .A1(n9997), .A2(n9673), .B1(n9672), .B2(n9671), .ZN(n9674)
         );
  AOI21_X1 U10972 ( .B1(n9738), .B2(n9675), .A(n9674), .ZN(n9676) );
  OAI211_X1 U10973 ( .C1(n9860), .C2(n9741), .A(n9677), .B(n9676), .ZN(n9678)
         );
  AOI21_X1 U10974 ( .B1(n9861), .B2(n9977), .A(n9678), .ZN(n9679) );
  OAI211_X1 U10975 ( .C1(n9866), .C2(n9715), .A(n9680), .B(n9679), .ZN(
        P1_U3275) );
  XNOR2_X1 U10976 ( .A(n9682), .B(n9681), .ZN(n9871) );
  AOI21_X1 U10977 ( .B1(n9706), .B2(n9869), .A(n9768), .ZN(n9684) );
  AND2_X1 U10978 ( .A1(n9685), .A2(n9684), .ZN(n9868) );
  NAND2_X1 U10979 ( .A1(n9869), .A2(n9747), .ZN(n9688) );
  NAND2_X1 U10980 ( .A1(n9686), .A2(n9991), .ZN(n9687) );
  OAI211_X1 U10981 ( .C1(n9997), .C2(n9689), .A(n9688), .B(n9687), .ZN(n9690)
         );
  AOI21_X1 U10982 ( .B1(n9868), .B2(n9977), .A(n9690), .ZN(n9697) );
  NAND2_X1 U10983 ( .A1(n9692), .A2(n6499), .ZN(n9693) );
  NAND3_X1 U10984 ( .A1(n9691), .A2(n10061), .A3(n9693), .ZN(n9695) );
  AOI22_X1 U10985 ( .A1(n10053), .A2(n9883), .B1(n9850), .B2(n9986), .ZN(n9694) );
  NAND2_X1 U10986 ( .A1(n9695), .A2(n9694), .ZN(n9867) );
  NAND2_X1 U10987 ( .A1(n9867), .A2(n9997), .ZN(n9696) );
  OAI211_X1 U10988 ( .C1(n9871), .C2(n9765), .A(n9697), .B(n9696), .ZN(
        P1_U3276) );
  AND2_X1 U10989 ( .A1(n9698), .A2(n9717), .ZN(n9699) );
  NAND2_X1 U10990 ( .A1(n9751), .A2(n9699), .ZN(n9733) );
  NAND3_X1 U10991 ( .A1(n9733), .A2(n9719), .A3(n9717), .ZN(n9718) );
  NAND2_X1 U10992 ( .A1(n9718), .A2(n9700), .ZN(n9701) );
  XNOR2_X1 U10993 ( .A(n9701), .B(n5680), .ZN(n9880) );
  NAND2_X1 U10994 ( .A1(n9703), .A2(n9702), .ZN(n9872) );
  NAND3_X1 U10995 ( .A1(n9663), .A2(n9704), .A3(n9872), .ZN(n9714) );
  AOI21_X1 U10996 ( .B1(n9705), .B2(n9877), .A(n9768), .ZN(n9707) );
  AND2_X1 U10997 ( .A1(n9707), .A2(n9706), .ZN(n9875) );
  AOI22_X1 U10998 ( .A1(n9993), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9708), .B2(
        n9991), .ZN(n9709) );
  OAI21_X1 U10999 ( .B1(n9874), .B2(n9741), .A(n9709), .ZN(n9710) );
  AOI21_X1 U11000 ( .B1(n9738), .B2(n9891), .A(n9710), .ZN(n9711) );
  OAI21_X1 U11001 ( .B1(n5070), .B2(n9995), .A(n9711), .ZN(n9712) );
  AOI21_X1 U11002 ( .B1(n9875), .B2(n9977), .A(n9712), .ZN(n9713) );
  OAI211_X1 U11003 ( .C1(n9880), .C2(n9715), .A(n9714), .B(n9713), .ZN(
        P1_U3277) );
  XOR2_X1 U11004 ( .A(n9716), .B(n9719), .Z(n9890) );
  AND2_X1 U11005 ( .A1(n9733), .A2(n9717), .ZN(n9720) );
  OAI21_X1 U11006 ( .B1(n9720), .B2(n9719), .A(n9718), .ZN(n9888) );
  OAI211_X1 U11007 ( .C1(n9721), .C2(n9886), .A(n9975), .B(n9705), .ZN(n9885)
         );
  AOI22_X1 U11008 ( .A1(n9993), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9722), .B2(
        n9991), .ZN(n9724) );
  NAND2_X1 U11009 ( .A1(n9738), .A2(n9882), .ZN(n9723) );
  OAI211_X1 U11010 ( .C1(n9725), .C2(n9741), .A(n9724), .B(n9723), .ZN(n9726)
         );
  AOI21_X1 U11011 ( .B1(n5860), .B2(n9747), .A(n9726), .ZN(n9727) );
  OAI21_X1 U11012 ( .B1(n9885), .B2(n9743), .A(n9727), .ZN(n9728) );
  AOI21_X1 U11013 ( .B1(n9888), .B2(n9729), .A(n9728), .ZN(n9730) );
  OAI21_X1 U11014 ( .B1(n9890), .B2(n9765), .A(n9730), .ZN(P1_U3278) );
  NAND2_X1 U11015 ( .A1(n9751), .A2(n9731), .ZN(n9732) );
  NAND2_X1 U11016 ( .A1(n9732), .A2(n9736), .ZN(n9734) );
  NAND3_X1 U11017 ( .A1(n9734), .A2(n10061), .A3(n9733), .ZN(n9897) );
  XOR2_X1 U11018 ( .A(n9735), .B(n9736), .Z(n9899) );
  OR2_X1 U11019 ( .A1(n9899), .A2(n9765), .ZN(n9749) );
  AOI22_X1 U11020 ( .A1(n9993), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9737), .B2(
        n9991), .ZN(n9740) );
  NAND2_X1 U11021 ( .A1(n9738), .A2(n9892), .ZN(n9739) );
  OAI211_X1 U11022 ( .C1(n9873), .C2(n9741), .A(n9740), .B(n9739), .ZN(n9745)
         );
  OAI21_X1 U11023 ( .B1(n9758), .B2(n9895), .A(n9975), .ZN(n9742) );
  OR2_X1 U11024 ( .A1(n9742), .A2(n9721), .ZN(n9894) );
  NOR2_X1 U11025 ( .A1(n9894), .A2(n9743), .ZN(n9744) );
  AOI211_X1 U11026 ( .C1(n9747), .C2(n9746), .A(n9745), .B(n9744), .ZN(n9748)
         );
  OAI211_X1 U11027 ( .C1(n9993), .C2(n9897), .A(n9749), .B(n9748), .ZN(
        P1_U3279) );
  XOR2_X1 U11028 ( .A(n9750), .B(n9754), .Z(n9904) );
  INV_X1 U11029 ( .A(n9751), .ZN(n9752) );
  AOI21_X1 U11030 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9755) );
  OAI222_X1 U11031 ( .A1(n10082), .A2(n9757), .B1(n10065), .B2(n9756), .C1(
        n9881), .C2(n9755), .ZN(n9900) );
  AOI211_X1 U11032 ( .C1(n9902), .C2(n9759), .A(n9768), .B(n9758), .ZN(n9901)
         );
  NAND2_X1 U11033 ( .A1(n9901), .A2(n9977), .ZN(n9762) );
  AOI22_X1 U11034 ( .A1(n9993), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9760), .B2(
        n9991), .ZN(n9761) );
  OAI211_X1 U11035 ( .C1(n5073), .C2(n9995), .A(n9762), .B(n9761), .ZN(n9763)
         );
  AOI21_X1 U11036 ( .B1(n9900), .B2(n9997), .A(n9763), .ZN(n9764) );
  OAI21_X1 U11037 ( .B1(n9765), .B2(n9904), .A(n9764), .ZN(P1_U3280) );
  NAND2_X1 U11038 ( .A1(n9766), .A2(n10078), .ZN(n9767) );
  OAI211_X1 U11039 ( .C1(n9769), .C2(n9768), .A(n9767), .B(n9770), .ZN(n9905)
         );
  MUX2_X1 U11040 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9905), .S(n10103), .Z(
        P1_U3553) );
  OAI211_X1 U11041 ( .C1(n9772), .C2(n10071), .A(n9771), .B(n9770), .ZN(n9906)
         );
  MUX2_X1 U11042 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9906), .S(n10103), .Z(
        P1_U3552) );
  NOR2_X1 U11043 ( .A1(n9782), .A2(n10057), .ZN(n9775) );
  NAND3_X1 U11044 ( .A1(n5391), .A2(n9789), .A3(n10087), .ZN(n9781) );
  OAI21_X1 U11045 ( .B1(n9777), .B2(n10082), .A(n9776), .ZN(n9778) );
  AOI21_X1 U11046 ( .B1(n9779), .B2(n10078), .A(n9778), .ZN(n9780) );
  MUX2_X1 U11047 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9907), .S(n10103), .Z(
        P1_U3551) );
  AOI22_X1 U11048 ( .A1(n9789), .A2(n9986), .B1(n10053), .B2(n9788), .ZN(n9790) );
  OAI211_X1 U11049 ( .C1(n9792), .C2(n10071), .A(n9791), .B(n9790), .ZN(n9793)
         );
  AOI21_X1 U11050 ( .B1(n9794), .B2(n10061), .A(n9793), .ZN(n9795) );
  OAI21_X1 U11051 ( .B1(n10057), .B2(n9796), .A(n9795), .ZN(n9908) );
  MUX2_X1 U11052 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9908), .S(n10103), .Z(
        P1_U3549) );
  OAI22_X1 U11053 ( .A1(n9798), .A2(n10065), .B1(n9797), .B2(n10082), .ZN(
        n9800) );
  AOI211_X1 U11054 ( .C1(n10078), .C2(n9801), .A(n9800), .B(n9799), .ZN(n9804)
         );
  NAND2_X1 U11055 ( .A1(n9802), .A2(n10087), .ZN(n9803) );
  OAI211_X1 U11056 ( .C1(n9805), .C2(n9881), .A(n9804), .B(n9803), .ZN(n9909)
         );
  MUX2_X1 U11057 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9909), .S(n10103), .Z(
        P1_U3548) );
  MUX2_X1 U11058 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9910), .S(n10103), .Z(
        P1_U3547) );
  AOI211_X1 U11059 ( .C1(n10078), .C2(n9812), .A(n9811), .B(n9810), .ZN(n9813)
         );
  OAI21_X1 U11060 ( .B1(n10057), .B2(n9814), .A(n9813), .ZN(n9911) );
  MUX2_X1 U11061 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9911), .S(n10103), .Z(
        P1_U3546) );
  AOI22_X1 U11062 ( .A1(n9816), .A2(n9986), .B1(n10053), .B2(n9815), .ZN(n9817) );
  OAI211_X1 U11063 ( .C1(n9819), .C2(n10071), .A(n9818), .B(n9817), .ZN(n9820)
         );
  AOI21_X1 U11064 ( .B1(n9821), .B2(n10061), .A(n9820), .ZN(n9822) );
  OAI21_X1 U11065 ( .B1(n9823), .B2(n10057), .A(n9822), .ZN(n9912) );
  MUX2_X1 U11066 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9912), .S(n10103), .Z(
        P1_U3545) );
  AOI22_X1 U11067 ( .A1(n9825), .A2(n9986), .B1(n10053), .B2(n9824), .ZN(n9826) );
  OAI211_X1 U11068 ( .C1(n9828), .C2(n10071), .A(n9827), .B(n9826), .ZN(n9829)
         );
  AOI21_X1 U11069 ( .B1(n9830), .B2(n10061), .A(n9829), .ZN(n9831) );
  OAI21_X1 U11070 ( .B1(n9832), .B2(n10057), .A(n9831), .ZN(n9913) );
  MUX2_X1 U11071 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9913), .S(n10103), .Z(
        P1_U3544) );
  OAI22_X1 U11072 ( .A1(n9834), .A2(n10065), .B1(n9833), .B2(n10082), .ZN(
        n9836) );
  AOI211_X1 U11073 ( .C1(n10078), .C2(n9837), .A(n9836), .B(n9835), .ZN(n9840)
         );
  NAND2_X1 U11074 ( .A1(n9838), .A2(n10061), .ZN(n9839) );
  OAI211_X1 U11075 ( .C1(n10057), .C2(n9841), .A(n9840), .B(n9839), .ZN(n9914)
         );
  MUX2_X1 U11076 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9914), .S(n10103), .Z(
        P1_U3543) );
  OAI22_X1 U11077 ( .A1(n9842), .A2(n10065), .B1(n9860), .B2(n10082), .ZN(
        n9844) );
  AOI211_X1 U11078 ( .C1(n10078), .C2(n9845), .A(n9844), .B(n9843), .ZN(n9848)
         );
  NAND2_X1 U11079 ( .A1(n9846), .A2(n10061), .ZN(n9847) );
  OAI211_X1 U11080 ( .C1(n9849), .C2(n10057), .A(n9848), .B(n9847), .ZN(n9915)
         );
  MUX2_X1 U11081 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9915), .S(n10103), .Z(
        P1_U3542) );
  AOI22_X1 U11082 ( .A1(n9851), .A2(n9986), .B1(n10053), .B2(n9850), .ZN(n9852) );
  OAI211_X1 U11083 ( .C1(n9854), .C2(n10071), .A(n9853), .B(n9852), .ZN(n9855)
         );
  AOI21_X1 U11084 ( .B1(n9856), .B2(n10061), .A(n9855), .ZN(n9857) );
  OAI21_X1 U11085 ( .B1(n9858), .B2(n10057), .A(n9857), .ZN(n9916) );
  MUX2_X1 U11086 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9916), .S(n10103), .Z(
        P1_U3541) );
  NAND2_X1 U11087 ( .A1(n9859), .A2(n10087), .ZN(n9865) );
  OAI22_X1 U11088 ( .A1(n9860), .A2(n10065), .B1(n9874), .B2(n10082), .ZN(
        n9862) );
  AOI211_X1 U11089 ( .C1(n10078), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9864)
         );
  OAI211_X1 U11090 ( .C1(n9881), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9917)
         );
  MUX2_X1 U11091 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9917), .S(n10103), .Z(
        P1_U3540) );
  AOI211_X1 U11092 ( .C1(n10078), .C2(n9869), .A(n9868), .B(n9867), .ZN(n9870)
         );
  OAI21_X1 U11093 ( .B1(n9871), .B2(n10057), .A(n9870), .ZN(n9918) );
  MUX2_X1 U11094 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9918), .S(n10103), .Z(
        P1_U3539) );
  NAND3_X1 U11095 ( .A1(n9663), .A2(n10087), .A3(n9872), .ZN(n9879) );
  OAI22_X1 U11096 ( .A1(n9874), .A2(n10065), .B1(n9873), .B2(n10082), .ZN(
        n9876) );
  AOI211_X1 U11097 ( .C1(n10078), .C2(n9877), .A(n9876), .B(n9875), .ZN(n9878)
         );
  OAI211_X1 U11098 ( .C1(n9881), .C2(n9880), .A(n9879), .B(n9878), .ZN(n9919)
         );
  MUX2_X1 U11099 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9919), .S(n10103), .Z(
        P1_U3538) );
  AOI22_X1 U11100 ( .A1(n9883), .A2(n9986), .B1(n10053), .B2(n9882), .ZN(n9884) );
  OAI211_X1 U11101 ( .C1(n9886), .C2(n10071), .A(n9885), .B(n9884), .ZN(n9887)
         );
  AOI21_X1 U11102 ( .B1(n9888), .B2(n10061), .A(n9887), .ZN(n9889) );
  OAI21_X1 U11103 ( .B1(n9890), .B2(n10057), .A(n9889), .ZN(n9920) );
  MUX2_X1 U11104 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9920), .S(n10103), .Z(
        P1_U3537) );
  AOI22_X1 U11105 ( .A1(n9892), .A2(n10053), .B1(n9986), .B2(n9891), .ZN(n9893) );
  OAI211_X1 U11106 ( .C1(n9895), .C2(n10071), .A(n9894), .B(n9893), .ZN(n9896)
         );
  INV_X1 U11107 ( .A(n9896), .ZN(n9898) );
  OAI211_X1 U11108 ( .C1(n9899), .C2(n10057), .A(n9898), .B(n9897), .ZN(n9921)
         );
  MUX2_X1 U11109 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9921), .S(n10103), .Z(
        P1_U3536) );
  AOI211_X1 U11110 ( .C1(n10078), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9903)
         );
  OAI21_X1 U11111 ( .B1(n10057), .B2(n9904), .A(n9903), .ZN(n9922) );
  MUX2_X1 U11112 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9922), .S(n10103), .Z(
        P1_U3535) );
  MUX2_X1 U11113 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9905), .S(n10090), .Z(
        P1_U3521) );
  MUX2_X1 U11114 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9906), .S(n10090), .Z(
        P1_U3520) );
  MUX2_X1 U11115 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9907), .S(n10090), .Z(
        P1_U3519) );
  MUX2_X1 U11116 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9908), .S(n10090), .Z(
        P1_U3517) );
  MUX2_X1 U11117 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9909), .S(n10090), .Z(
        P1_U3516) );
  MUX2_X1 U11118 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9910), .S(n10090), .Z(
        P1_U3515) );
  MUX2_X1 U11119 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9911), .S(n10090), .Z(
        P1_U3514) );
  MUX2_X1 U11120 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9912), .S(n10090), .Z(
        P1_U3513) );
  MUX2_X1 U11121 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9913), .S(n10090), .Z(
        P1_U3512) );
  MUX2_X1 U11122 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9914), .S(n10090), .Z(
        P1_U3511) );
  MUX2_X1 U11123 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9915), .S(n10090), .Z(
        P1_U3510) );
  MUX2_X1 U11124 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9916), .S(n10090), .Z(
        P1_U3509) );
  MUX2_X1 U11125 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9917), .S(n10090), .Z(
        P1_U3507) );
  MUX2_X1 U11126 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9918), .S(n10090), .Z(
        P1_U3504) );
  MUX2_X1 U11127 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9919), .S(n10090), .Z(
        P1_U3501) );
  MUX2_X1 U11128 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9920), .S(n10090), .Z(
        P1_U3498) );
  MUX2_X1 U11129 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9921), .S(n10090), .Z(
        P1_U3495) );
  MUX2_X1 U11130 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9922), .S(n10090), .Z(
        P1_U3492) );
  MUX2_X1 U11131 ( .A(P1_D_REG_1__SCAN_IN), .B(n9925), .S(n10001), .Z(P1_U3440) );
  MUX2_X1 U11132 ( .A(P1_D_REG_0__SCAN_IN), .B(n9926), .S(n10001), .Z(P1_U3439) );
  NOR4_X1 U11133 ( .A1(n4594), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5369), .A4(
        P1_U3086), .ZN(n9927) );
  AOI21_X1 U11134 ( .B1(n9928), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9927), .ZN(
        n9929) );
  OAI21_X1 U11135 ( .B1(n9930), .B2(n9934), .A(n9929), .ZN(P1_U3324) );
  OAI222_X1 U11136 ( .A1(P1_U3086), .A2(n9932), .B1(n9943), .B2(n9931), .C1(
        n10469), .C2(n9940), .ZN(P1_U3326) );
  OAI222_X1 U11137 ( .A1(n9940), .A2(n9936), .B1(P1_U3086), .B2(n9935), .C1(
        n9934), .C2(n9933), .ZN(P1_U3328) );
  OAI222_X1 U11138 ( .A1(n9939), .A2(P1_U3086), .B1(n9943), .B2(n9938), .C1(
        n9937), .C2(n9940), .ZN(P1_U3329) );
  OAI222_X1 U11139 ( .A1(n9944), .A2(P1_U3086), .B1(n9943), .B2(n9942), .C1(
        n9941), .C2(n9940), .ZN(P1_U3330) );
  XNOR2_X1 U11140 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11141 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI211_X1 U11142 ( .C1(n9947), .C2(n9946), .A(n9945), .B(n9963), .ZN(n9953)
         );
  INV_X1 U11143 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9951) );
  INV_X1 U11144 ( .A(n9948), .ZN(n9950) );
  AOI211_X1 U11145 ( .C1(n9951), .C2(n9950), .A(n9959), .B(n9949), .ZN(n9952)
         );
  AOI211_X1 U11146 ( .C1(n9954), .C2(n9968), .A(n9953), .B(n9952), .ZN(n9956)
         );
  OAI211_X1 U11147 ( .C1(n9972), .C2(n9957), .A(n9956), .B(n9955), .ZN(
        P1_U3258) );
  INV_X1 U11148 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9971) );
  INV_X1 U11149 ( .A(n9962), .ZN(n9964) );
  OAI211_X1 U11150 ( .C1(n9972), .C2(n9971), .A(n9970), .B(n9969), .ZN(
        P1_U3261) );
  XNOR2_X1 U11151 ( .A(n9973), .B(n9981), .ZN(n10075) );
  OAI211_X1 U11152 ( .C1(n8233), .C2(n10072), .A(n9975), .B(n9974), .ZN(n10070) );
  INV_X1 U11153 ( .A(n10070), .ZN(n9976) );
  AOI22_X1 U11154 ( .A1(n10075), .A2(n9978), .B1(n9977), .B2(n9976), .ZN(
        n10000) );
  INV_X1 U11155 ( .A(n9979), .ZN(n10050) );
  NAND2_X1 U11156 ( .A1(n8228), .A2(n9980), .ZN(n9982) );
  NAND2_X1 U11157 ( .A1(n9982), .A2(n9981), .ZN(n9984) );
  NAND3_X1 U11158 ( .A1(n9984), .A2(n9983), .A3(n10061), .ZN(n9989) );
  AOI22_X1 U11159 ( .A1(n9987), .A2(n10053), .B1(n9986), .B2(n9985), .ZN(n9988) );
  NAND2_X1 U11160 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  AOI21_X1 U11161 ( .B1(n10075), .B2(n10050), .A(n9990), .ZN(n10077) );
  INV_X1 U11162 ( .A(n10077), .ZN(n9998) );
  AOI22_X1 U11163 ( .A1(n9993), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9992), .B2(
        n9991), .ZN(n9994) );
  OAI21_X1 U11164 ( .B1(n10072), .B2(n9995), .A(n9994), .ZN(n9996) );
  AOI21_X1 U11165 ( .B1(n9998), .B2(n9997), .A(n9996), .ZN(n9999) );
  NAND2_X1 U11166 ( .A1(n10000), .A2(n9999), .ZN(P1_U3282) );
  AND2_X1 U11167 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10002), .ZN(P1_U3294) );
  AND2_X1 U11168 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10002), .ZN(P1_U3295) );
  NOR2_X1 U11169 ( .A1(n10001), .A2(n10199), .ZN(P1_U3296) );
  AND2_X1 U11170 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10002), .ZN(P1_U3297) );
  NOR2_X1 U11171 ( .A1(n10001), .A2(n10435), .ZN(P1_U3298) );
  AND2_X1 U11172 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10002), .ZN(P1_U3299) );
  AND2_X1 U11173 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10002), .ZN(P1_U3300) );
  INV_X1 U11174 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10450) );
  NOR2_X1 U11175 ( .A1(n10001), .A2(n10450), .ZN(P1_U3301) );
  AND2_X1 U11176 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10002), .ZN(P1_U3302) );
  AND2_X1 U11177 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10002), .ZN(P1_U3303) );
  AND2_X1 U11178 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10002), .ZN(P1_U3304) );
  AND2_X1 U11179 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10002), .ZN(P1_U3305) );
  AND2_X1 U11180 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10002), .ZN(P1_U3306) );
  AND2_X1 U11181 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10002), .ZN(P1_U3307) );
  AND2_X1 U11182 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10002), .ZN(P1_U3308) );
  AND2_X1 U11183 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10002), .ZN(P1_U3309) );
  AND2_X1 U11184 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10002), .ZN(P1_U3310) );
  AND2_X1 U11185 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10002), .ZN(P1_U3311) );
  AND2_X1 U11186 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10002), .ZN(P1_U3312) );
  AND2_X1 U11187 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10002), .ZN(P1_U3313) );
  AND2_X1 U11188 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10002), .ZN(P1_U3314) );
  AND2_X1 U11189 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10002), .ZN(P1_U3315) );
  AND2_X1 U11190 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10002), .ZN(P1_U3316) );
  AND2_X1 U11191 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10002), .ZN(P1_U3317) );
  NOR2_X1 U11192 ( .A1(n10001), .A2(n10238), .ZN(P1_U3318) );
  AND2_X1 U11193 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10002), .ZN(P1_U3319) );
  AND2_X1 U11194 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10002), .ZN(P1_U3320) );
  AND2_X1 U11195 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10002), .ZN(P1_U3321) );
  NOR2_X1 U11196 ( .A1(n10001), .A2(n10463), .ZN(P1_U3322) );
  AND2_X1 U11197 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10002), .ZN(P1_U3323) );
  INV_X1 U11198 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U11199 ( .A1(n10090), .A2(n10004), .B1(n10003), .B2(n10088), .ZN(
        P1_U3453) );
  OAI21_X1 U11200 ( .B1(n10006), .B2(n10071), .A(n10005), .ZN(n10008) );
  AOI211_X1 U11201 ( .C1(n10087), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10091) );
  INV_X1 U11202 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10010) );
  AOI22_X1 U11203 ( .A1(n10090), .A2(n10091), .B1(n10010), .B2(n10088), .ZN(
        P1_U3462) );
  OAI22_X1 U11204 ( .A1(n10011), .A2(n10082), .B1(n6936), .B2(n10065), .ZN(
        n10012) );
  AOI21_X1 U11205 ( .B1(n10078), .B2(n10013), .A(n10012), .ZN(n10015) );
  OAI211_X1 U11206 ( .C1(n10016), .C2(n10057), .A(n10015), .B(n10014), .ZN(
        n10017) );
  AOI21_X1 U11207 ( .B1(n10061), .B2(n10018), .A(n10017), .ZN(n10092) );
  INV_X1 U11208 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U11209 ( .A1(n10090), .A2(n10092), .B1(n10481), .B2(n10088), .ZN(
        P1_U3465) );
  AND2_X1 U11210 ( .A1(n10019), .A2(n10087), .ZN(n10023) );
  OAI21_X1 U11211 ( .B1(n10021), .B2(n10071), .A(n10020), .ZN(n10022) );
  NOR3_X1 U11212 ( .A1(n10024), .A2(n10023), .A3(n10022), .ZN(n10093) );
  INV_X1 U11213 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10025) );
  AOI22_X1 U11214 ( .A1(n10090), .A2(n10093), .B1(n10025), .B2(n10088), .ZN(
        P1_U3468) );
  OAI21_X1 U11215 ( .B1(n10027), .B2(n10071), .A(n10026), .ZN(n10029) );
  AOI211_X1 U11216 ( .C1(n10087), .C2(n10030), .A(n10029), .B(n10028), .ZN(
        n10094) );
  INV_X1 U11217 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10031) );
  AOI22_X1 U11218 ( .A1(n10090), .A2(n10094), .B1(n10031), .B2(n10088), .ZN(
        P1_U3471) );
  INV_X1 U11219 ( .A(n10045), .ZN(n10074) );
  OAI21_X1 U11220 ( .B1(n10033), .B2(n10071), .A(n10032), .ZN(n10034) );
  AOI21_X1 U11221 ( .B1(n10035), .B2(n10074), .A(n10034), .ZN(n10036) );
  AND2_X1 U11222 ( .A1(n10037), .A2(n10036), .ZN(n10096) );
  INV_X1 U11223 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U11224 ( .A1(n10090), .A2(n10096), .B1(n10038), .B2(n10088), .ZN(
        P1_U3474) );
  INV_X1 U11225 ( .A(n10046), .ZN(n10049) );
  OAI22_X1 U11226 ( .A1(n10040), .A2(n10082), .B1(n10039), .B2(n10065), .ZN(
        n10042) );
  AOI211_X1 U11227 ( .C1(n10078), .C2(n10043), .A(n10042), .B(n10041), .ZN(
        n10044) );
  OAI21_X1 U11228 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(n10047) );
  AOI211_X1 U11229 ( .C1(n10050), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n10097) );
  INV_X1 U11230 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10051) );
  AOI22_X1 U11231 ( .A1(n10090), .A2(n10097), .B1(n10051), .B2(n10088), .ZN(
        P1_U3477) );
  AOI22_X1 U11232 ( .A1(n10054), .A2(n10078), .B1(n10053), .B2(n10052), .ZN(
        n10055) );
  OAI211_X1 U11233 ( .C1(n10058), .C2(n10057), .A(n10056), .B(n10055), .ZN(
        n10059) );
  AOI21_X1 U11234 ( .B1(n10061), .B2(n10060), .A(n10059), .ZN(n10098) );
  INV_X1 U11235 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U11236 ( .A1(n10090), .A2(n10098), .B1(n10255), .B2(n10088), .ZN(
        P1_U3480) );
  NAND2_X1 U11237 ( .A1(n10062), .A2(n10078), .ZN(n10063) );
  OAI211_X1 U11238 ( .C1(n10083), .C2(n10065), .A(n10064), .B(n10063), .ZN(
        n10067) );
  AOI211_X1 U11239 ( .C1(n10087), .C2(n10068), .A(n10067), .B(n10066), .ZN(
        n10099) );
  INV_X1 U11240 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10069) );
  AOI22_X1 U11241 ( .A1(n10090), .A2(n10099), .B1(n10069), .B2(n10088), .ZN(
        P1_U3483) );
  OAI21_X1 U11242 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(n10073) );
  AOI21_X1 U11243 ( .B1(n10075), .B2(n10074), .A(n10073), .ZN(n10076) );
  AND2_X1 U11244 ( .A1(n10077), .A2(n10076), .ZN(n10100) );
  INV_X1 U11245 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U11246 ( .A1(n10090), .A2(n10100), .B1(n10334), .B2(n10088), .ZN(
        P1_U3486) );
  NAND2_X1 U11247 ( .A1(n10079), .A2(n10078), .ZN(n10080) );
  OAI211_X1 U11248 ( .C1(n10083), .C2(n10082), .A(n10081), .B(n10080), .ZN(
        n10085) );
  AOI211_X1 U11249 ( .C1(n10087), .C2(n10086), .A(n10085), .B(n10084), .ZN(
        n10102) );
  INV_X1 U11250 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U11251 ( .A1(n10090), .A2(n10102), .B1(n10089), .B2(n10088), .ZN(
        P1_U3489) );
  AOI22_X1 U11252 ( .A1(n10103), .A2(n10091), .B1(n7364), .B2(n10101), .ZN(
        P1_U3525) );
  AOI22_X1 U11253 ( .A1(n10103), .A2(n10092), .B1(n4884), .B2(n10101), .ZN(
        P1_U3526) );
  AOI22_X1 U11254 ( .A1(n10103), .A2(n10093), .B1(n7367), .B2(n10101), .ZN(
        P1_U3527) );
  AOI22_X1 U11255 ( .A1(n10103), .A2(n10094), .B1(n7376), .B2(n10101), .ZN(
        P1_U3528) );
  INV_X1 U11256 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U11257 ( .A1(n10103), .A2(n10096), .B1(n10095), .B2(n10101), .ZN(
        P1_U3529) );
  INV_X1 U11258 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U11259 ( .A1(n10103), .A2(n10097), .B1(n10484), .B2(n10101), .ZN(
        P1_U3530) );
  AOI22_X1 U11260 ( .A1(n10103), .A2(n10098), .B1(n7682), .B2(n10101), .ZN(
        P1_U3531) );
  AOI22_X1 U11261 ( .A1(n10103), .A2(n10099), .B1(n7846), .B2(n10101), .ZN(
        P1_U3532) );
  AOI22_X1 U11262 ( .A1(n10103), .A2(n10100), .B1(n7984), .B2(n10101), .ZN(
        P1_U3533) );
  AOI22_X1 U11263 ( .A1(n10103), .A2(n10102), .B1(n8118), .B2(n10101), .ZN(
        P1_U3534) );
  NAND2_X1 U11264 ( .A1(n10105), .A2(n10104), .ZN(n10106) );
  XOR2_X1 U11265 ( .A(n10112), .B(n10106), .Z(n10110) );
  AOI222_X1 U11266 ( .A1(n10111), .A2(n10110), .B1(n10109), .B2(n10108), .C1(
        n6397), .C2(n10107), .ZN(n10144) );
  XNOR2_X1 U11267 ( .A(n10113), .B(n10112), .ZN(n10142) );
  OAI22_X1 U11268 ( .A1(n10115), .A2(n10114), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n10122), .ZN(n10116) );
  AOI21_X1 U11269 ( .B1(n10117), .B2(n10142), .A(n10116), .ZN(n10118) );
  OAI221_X1 U11270 ( .B1(n10130), .B2(n10144), .C1(n10128), .C2(n10119), .A(
        n10118), .ZN(P2_U3230) );
  INV_X1 U11271 ( .A(n10120), .ZN(n10127) );
  OAI22_X1 U11272 ( .A1(n10122), .A2(n7476), .B1(n6398), .B2(n10121), .ZN(
        n10125) );
  INV_X1 U11273 ( .A(n10123), .ZN(n10124) );
  AOI211_X1 U11274 ( .C1(n10127), .C2(n10126), .A(n10125), .B(n10124), .ZN(
        n10129) );
  AOI22_X1 U11275 ( .A1(n10130), .A2(n7438), .B1(n10129), .B2(n10128), .ZN(
        P2_U3231) );
  INV_X1 U11276 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10455) );
  INV_X1 U11277 ( .A(n10149), .ZN(n10133) );
  AOI21_X1 U11278 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(n10134) );
  AOI211_X1 U11279 ( .C1(n10141), .C2(n10136), .A(n10135), .B(n10134), .ZN(
        n10161) );
  AOI22_X1 U11280 ( .A1(n10159), .A2(n10455), .B1(n10161), .B2(n10157), .ZN(
        P2_U3390) );
  INV_X1 U11281 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U11282 ( .A1(n10159), .A2(n10418), .B1(n10137), .B2(n10157), .ZN(
        P2_U3393) );
  INV_X1 U11283 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U11284 ( .A1(n10159), .A2(n10139), .B1(n10138), .B2(n10157), .ZN(
        P2_U3396) );
  INV_X1 U11285 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U11286 ( .A1(n10142), .A2(n10149), .B1(n10141), .B2(n10140), .ZN(
        n10143) );
  AND2_X1 U11287 ( .A1(n10144), .A2(n10143), .ZN(n10162) );
  AOI22_X1 U11288 ( .A1(n10159), .A2(n10447), .B1(n10162), .B2(n10157), .ZN(
        P2_U3399) );
  INV_X1 U11289 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10434) );
  INV_X1 U11290 ( .A(n10145), .ZN(n10150) );
  OAI21_X1 U11291 ( .B1(n10147), .B2(n10151), .A(n10146), .ZN(n10148) );
  AOI21_X1 U11292 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(n10163) );
  AOI22_X1 U11293 ( .A1(n10159), .A2(n10434), .B1(n10163), .B2(n10157), .ZN(
        P2_U3402) );
  INV_X1 U11294 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10158) );
  OAI22_X1 U11295 ( .A1(n10154), .A2(n10153), .B1(n10152), .B2(n10151), .ZN(
        n10156) );
  NOR2_X1 U11296 ( .A1(n10156), .A2(n10155), .ZN(n10165) );
  AOI22_X1 U11297 ( .A1(n10159), .A2(n10158), .B1(n10165), .B2(n10157), .ZN(
        P2_U3405) );
  AOI22_X1 U11298 ( .A1(n10166), .A2(n10161), .B1(n10160), .B2(n10164), .ZN(
        P2_U3459) );
  AOI22_X1 U11299 ( .A1(n10166), .A2(n10162), .B1(n7426), .B2(n10164), .ZN(
        P2_U3462) );
  AOI22_X1 U11300 ( .A1(n10166), .A2(n10163), .B1(n7419), .B2(n10164), .ZN(
        P2_U3463) );
  AOI22_X1 U11301 ( .A1(n10166), .A2(n10165), .B1(n7554), .B2(n10164), .ZN(
        P2_U3464) );
  OAI222_X1 U11302 ( .A1(n10171), .A2(n10170), .B1(n10171), .B2(n10169), .C1(
        n10168), .C2(n10167), .ZN(ADD_1068_U5) );
  AOI21_X1 U11303 ( .B1(n10212), .B2(n10173), .A(n10172), .ZN(ADD_1068_U46) );
  NOR2_X1 U11304 ( .A1(n10175), .A2(n10174), .ZN(n10176) );
  XOR2_X1 U11305 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10176), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11306 ( .A(n10178), .B(n10177), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11307 ( .A(n10180), .B(n10179), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11308 ( .A(n10182), .B(n10181), .ZN(ADD_1068_U58) );
  OAI21_X1 U11309 ( .B1(n10185), .B2(n10184), .A(n10183), .ZN(ADD_1068_U60) );
  OAI21_X1 U11310 ( .B1(n10188), .B2(n10187), .A(n10186), .ZN(ADD_1068_U61) );
  OAI21_X1 U11311 ( .B1(n10191), .B2(n10190), .A(n10189), .ZN(ADD_1068_U62) );
  OAI21_X1 U11312 ( .B1(n10194), .B2(n10193), .A(n10192), .ZN(ADD_1068_U63) );
  NOR2_X1 U11313 ( .A1(n10196), .A2(n10195), .ZN(n10504) );
  INV_X1 U11314 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U11315 ( .A1(n10344), .A2(keyinput29), .B1(n10339), .B2(keyinput21), 
        .ZN(n10197) );
  OAI221_X1 U11316 ( .B1(n10344), .B2(keyinput29), .C1(n10339), .C2(keyinput21), .A(n10197), .ZN(n10208) );
  AOI22_X1 U11317 ( .A1(n10343), .A2(keyinput87), .B1(n10199), .B2(keyinput86), 
        .ZN(n10198) );
  OAI221_X1 U11318 ( .B1(n10343), .B2(keyinput87), .C1(n10199), .C2(keyinput86), .A(n10198), .ZN(n10207) );
  AOI22_X1 U11319 ( .A1(n10202), .A2(keyinput63), .B1(n10201), .B2(keyinput45), 
        .ZN(n10200) );
  OAI221_X1 U11320 ( .B1(n10202), .B2(keyinput63), .C1(n10201), .C2(keyinput45), .A(n10200), .ZN(n10206) );
  AOI22_X1 U11321 ( .A1(n10204), .A2(keyinput96), .B1(n6310), .B2(keyinput33), 
        .ZN(n10203) );
  OAI221_X1 U11322 ( .B1(n10204), .B2(keyinput96), .C1(n6310), .C2(keyinput33), 
        .A(n10203), .ZN(n10205) );
  NOR4_X1 U11323 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(
        n10502) );
  AOI22_X1 U11324 ( .A1(n10210), .A2(keyinput34), .B1(n4877), .B2(keyinput44), 
        .ZN(n10209) );
  OAI221_X1 U11325 ( .B1(n10210), .B2(keyinput34), .C1(n4877), .C2(keyinput44), 
        .A(n10209), .ZN(n10223) );
  XOR2_X1 U11326 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput84), .Z(n10222) );
  XNOR2_X1 U11327 ( .A(n10211), .B(keyinput28), .ZN(n10218) );
  XNOR2_X1 U11328 ( .A(keyinput43), .B(n10212), .ZN(n10217) );
  INV_X1 U11329 ( .A(SI_0_), .ZN(n10345) );
  NOR2_X1 U11330 ( .A1(keyinput76), .A2(n10345), .ZN(n10216) );
  NAND2_X1 U11331 ( .A1(n10345), .A2(keyinput76), .ZN(n10213) );
  OAI21_X1 U11332 ( .B1(n10214), .B2(keyinput108), .A(n10213), .ZN(n10215) );
  OR4_X1 U11333 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10221) );
  INV_X1 U11334 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n10219) );
  XNOR2_X1 U11335 ( .A(keyinput74), .B(n10219), .ZN(n10220) );
  NOR4_X1 U11336 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10501) );
  INV_X1 U11337 ( .A(SI_16_), .ZN(n10308) );
  OAI22_X1 U11338 ( .A1(n10308), .A2(keyinput58), .B1(n5413), .B2(keyinput101), 
        .ZN(n10224) );
  AOI221_X1 U11339 ( .B1(n10308), .B2(keyinput58), .C1(keyinput101), .C2(n5413), .A(n10224), .ZN(n10235) );
  OAI22_X1 U11340 ( .A1(n10314), .A2(keyinput69), .B1(n10226), .B2(keyinput80), 
        .ZN(n10225) );
  AOI221_X1 U11341 ( .B1(n10314), .B2(keyinput69), .C1(keyinput80), .C2(n10226), .A(n10225), .ZN(n10234) );
  XOR2_X1 U11342 ( .A(P1_REG0_REG_29__SCAN_IN), .B(keyinput99), .Z(n10229) );
  XNOR2_X1 U11343 ( .A(n10227), .B(keyinput47), .ZN(n10228) );
  NOR2_X1 U11344 ( .A1(n10229), .A2(n10228), .ZN(n10233) );
  OAI22_X1 U11345 ( .A1(n5537), .A2(keyinput32), .B1(n10231), .B2(keyinput115), 
        .ZN(n10230) );
  AOI221_X1 U11346 ( .B1(n5537), .B2(keyinput32), .C1(keyinput115), .C2(n10231), .A(n10230), .ZN(n10232) );
  NAND4_X1 U11347 ( .A1(n10235), .A2(n10234), .A3(n10233), .A4(n10232), .ZN(
        n10307) );
  OAI22_X1 U11348 ( .A1(n10238), .A2(keyinput105), .B1(n10237), .B2(keyinput14), .ZN(n10236) );
  AOI221_X1 U11349 ( .B1(n10238), .B2(keyinput105), .C1(keyinput14), .C2(
        n10237), .A(n10236), .ZN(n10248) );
  XNOR2_X1 U11350 ( .A(SI_7_), .B(keyinput16), .ZN(n10242) );
  XNOR2_X1 U11351 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput111), .ZN(n10241) );
  XNOR2_X1 U11352 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput122), .ZN(n10240)
         );
  XNOR2_X1 U11353 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput46), .ZN(n10239) );
  NAND4_X1 U11354 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n10246) );
  XNOR2_X1 U11355 ( .A(n10243), .B(keyinput50), .ZN(n10245) );
  XNOR2_X1 U11356 ( .A(keyinput93), .B(n5815), .ZN(n10244) );
  NOR3_X1 U11357 ( .A1(n10246), .A2(n10245), .A3(n10244), .ZN(n10247) );
  NAND2_X1 U11358 ( .A1(n10248), .A2(n10247), .ZN(n10306) );
  AOI22_X1 U11359 ( .A1(n10250), .A2(keyinput20), .B1(keyinput90), .B2(n10334), 
        .ZN(n10249) );
  OAI221_X1 U11360 ( .B1(n10250), .B2(keyinput20), .C1(n10334), .C2(keyinput90), .A(n10249), .ZN(n10262) );
  AOI22_X1 U11361 ( .A1(n10252), .A2(keyinput56), .B1(keyinput36), .B2(n10319), 
        .ZN(n10251) );
  OAI221_X1 U11362 ( .B1(n10252), .B2(keyinput56), .C1(n10319), .C2(keyinput36), .A(n10251), .ZN(n10261) );
  AOI22_X1 U11363 ( .A1(n10255), .A2(keyinput117), .B1(n10254), .B2(keyinput81), .ZN(n10253) );
  OAI221_X1 U11364 ( .B1(n10255), .B2(keyinput117), .C1(n10254), .C2(
        keyinput81), .A(n10253), .ZN(n10260) );
  INV_X1 U11365 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10256) );
  XOR2_X1 U11366 ( .A(n10256), .B(keyinput123), .Z(n10258) );
  XNOR2_X1 U11367 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput92), .ZN(n10257)
         );
  NAND2_X1 U11368 ( .A1(n10258), .A2(n10257), .ZN(n10259) );
  NOR4_X1 U11369 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10304) );
  AOI22_X1 U11370 ( .A1(n7786), .A2(keyinput82), .B1(keyinput125), .B2(n10264), 
        .ZN(n10263) );
  OAI221_X1 U11371 ( .B1(n7786), .B2(keyinput82), .C1(n10264), .C2(keyinput125), .A(n10263), .ZN(n10273) );
  AOI22_X1 U11372 ( .A1(n10342), .A2(keyinput61), .B1(keyinput11), .B2(n10341), 
        .ZN(n10265) );
  OAI221_X1 U11373 ( .B1(n10342), .B2(keyinput61), .C1(n10341), .C2(keyinput11), .A(n10265), .ZN(n10272) );
  AOI22_X1 U11374 ( .A1(P1_U3086), .A2(keyinput31), .B1(keyinput104), .B2(
        n10267), .ZN(n10266) );
  OAI221_X1 U11375 ( .B1(P1_U3086), .B2(keyinput31), .C1(n10267), .C2(
        keyinput104), .A(n10266), .ZN(n10271) );
  XOR2_X1 U11376 ( .A(n10340), .B(keyinput113), .Z(n10269) );
  XNOR2_X1 U11377 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput110), .ZN(n10268) );
  NAND2_X1 U11378 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  NOR4_X1 U11379 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10303) );
  AOI22_X1 U11380 ( .A1(n10320), .A2(keyinput83), .B1(keyinput118), .B2(n10275), .ZN(n10274) );
  OAI221_X1 U11381 ( .B1(n10320), .B2(keyinput83), .C1(n10275), .C2(
        keyinput118), .A(n10274), .ZN(n10287) );
  AOI22_X1 U11382 ( .A1(n10278), .A2(keyinput66), .B1(n10277), .B2(keyinput98), 
        .ZN(n10276) );
  OAI221_X1 U11383 ( .B1(n10278), .B2(keyinput66), .C1(n10277), .C2(keyinput98), .A(n10276), .ZN(n10286) );
  INV_X1 U11384 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10281) );
  INV_X1 U11385 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U11386 ( .A1(n10281), .A2(keyinput42), .B1(n10280), .B2(keyinput77), 
        .ZN(n10279) );
  OAI221_X1 U11387 ( .B1(n10281), .B2(keyinput42), .C1(n10280), .C2(keyinput77), .A(n10279), .ZN(n10285) );
  XNOR2_X1 U11388 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput22), .ZN(n10283)
         );
  XNOR2_X1 U11389 ( .A(P2_REG0_REG_12__SCAN_IN), .B(keyinput26), .ZN(n10282)
         );
  NAND2_X1 U11390 ( .A1(n10283), .A2(n10282), .ZN(n10284) );
  NOR4_X1 U11391 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n10302) );
  AOI22_X1 U11392 ( .A1(n10290), .A2(keyinput30), .B1(keyinput100), .B2(n10289), .ZN(n10288) );
  OAI221_X1 U11393 ( .B1(n10290), .B2(keyinput30), .C1(n10289), .C2(
        keyinput100), .A(n10288), .ZN(n10300) );
  AOI22_X1 U11394 ( .A1(n10293), .A2(keyinput38), .B1(n10292), .B2(keyinput40), 
        .ZN(n10291) );
  OAI221_X1 U11395 ( .B1(n10293), .B2(keyinput38), .C1(n10292), .C2(keyinput40), .A(n10291), .ZN(n10299) );
  XNOR2_X1 U11396 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput24), .ZN(n10297) );
  XNOR2_X1 U11397 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput72), .ZN(n10296)
         );
  XNOR2_X1 U11398 ( .A(P1_REG3_REG_25__SCAN_IN), .B(keyinput49), .ZN(n10295)
         );
  XNOR2_X1 U11399 ( .A(keyinput79), .B(P2_REG1_REG_0__SCAN_IN), .ZN(n10294) );
  NAND4_X1 U11400 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  NOR3_X1 U11401 ( .A1(n10300), .A2(n10299), .A3(n10298), .ZN(n10301) );
  NAND4_X1 U11402 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10305) );
  NOR3_X1 U11403 ( .A1(n10307), .A2(n10306), .A3(n10305), .ZN(n10500) );
  NAND4_X1 U11404 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .A3(P2_ADDR_REG_14__SCAN_IN), .A4(n10308), .ZN(n10332) );
  NAND4_X1 U11405 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n5413), .A3(n5537), .A4(
        n10309), .ZN(n10331) );
  NOR4_X1 U11406 ( .A1(n10311), .A2(n10310), .A3(P1_REG1_REG_1__SCAN_IN), .A4(
        P1_REG1_REG_14__SCAN_IN), .ZN(n10313) );
  NOR2_X1 U11407 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n10312) );
  NAND4_X1 U11408 ( .A1(n10313), .A2(P1_IR_REG_11__SCAN_IN), .A3(
        P2_REG1_REG_1__SCAN_IN), .A4(n10312), .ZN(n10330) );
  AND4_X1 U11409 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P2_REG0_REG_14__SCAN_IN), 
        .A3(P2_REG1_REG_0__SCAN_IN), .A4(n10314), .ZN(n10318) );
  NOR4_X1 U11410 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(P1_REG2_REG_3__SCAN_IN), 
        .A3(P2_REG1_REG_21__SCAN_IN), .A4(P2_REG1_REG_9__SCAN_IN), .ZN(n10317)
         );
  NOR4_X1 U11411 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(P1_REG0_REG_9__SCAN_IN), .A4(P1_REG2_REG_4__SCAN_IN), .ZN(n10316)
         );
  NOR4_X1 U11412 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P2_DATAO_REG_19__SCAN_IN), 
        .A3(P1_REG1_REG_19__SCAN_IN), .A4(P2_REG2_REG_15__SCAN_IN), .ZN(n10315) );
  NAND4_X1 U11413 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10326) );
  INV_X1 U11414 ( .A(P2_B_REG_SCAN_IN), .ZN(n10392) );
  NOR2_X1 U11415 ( .A1(n10319), .A2(n10392), .ZN(n10324) );
  NOR4_X1 U11416 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .A3(P2_REG1_REG_31__SCAN_IN), .A4(n10320), .ZN(n10323) );
  INV_X1 U11417 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10401) );
  INV_X1 U11418 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10387) );
  NOR4_X1 U11419 ( .A1(P2_REG1_REG_30__SCAN_IN), .A2(n10401), .A3(n10386), 
        .A4(n10387), .ZN(n10322) );
  NOR4_X1 U11420 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_REG2_REG_7__SCAN_IN), 
        .A3(n5908), .A4(n10374), .ZN(n10321) );
  NAND4_X1 U11421 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  NOR4_X1 U11422 ( .A1(n10292), .A2(P2_REG3_REG_20__SCAN_IN), .A3(n10326), 
        .A4(n10325), .ZN(n10328) );
  NOR2_X1 U11423 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(SI_5_), .ZN(n10327) );
  NAND4_X1 U11424 ( .A1(n10328), .A2(P2_REG1_REG_8__SCAN_IN), .A3(
        P2_REG0_REG_12__SCAN_IN), .A4(n10327), .ZN(n10329) );
  OR4_X1 U11425 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10338) );
  NOR4_X1 U11426 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .A3(n10417), .A4(n10406), .ZN(n10333) );
  NAND3_X1 U11427 ( .A1(P1_REG2_REG_28__SCAN_IN), .A2(P2_REG0_REG_17__SCAN_IN), 
        .A3(n10333), .ZN(n10337) );
  NOR4_X1 U11428 ( .A1(SI_7_), .A2(P1_REG2_REG_26__SCAN_IN), .A3(
        P2_IR_REG_17__SCAN_IN), .A4(P2_IR_REG_7__SCAN_IN), .ZN(n10335) );
  NAND3_X1 U11429 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10335), .A3(n10334), .ZN(
        n10336) );
  OR3_X1 U11430 ( .A1(n10338), .A2(n10337), .A3(n10336), .ZN(n10369) );
  NAND4_X1 U11431 ( .A1(P1_REG0_REG_25__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .A3(n10339), .A4(n6310), .ZN(n10349) );
  NAND4_X1 U11432 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n10342), .A3(n10341), .A4(
        n10340), .ZN(n10347) );
  NAND4_X1 U11433 ( .A1(n10344), .A2(P2_REG2_REG_16__SCAN_IN), .A3(
        P2_REG3_REG_11__SCAN_IN), .A4(n10343), .ZN(n10346) );
  OR4_X1 U11434 ( .A1(SI_4_), .A2(n10347), .A3(n10346), .A4(SI_0_), .ZN(n10348) );
  NOR4_X1 U11435 ( .A1(n10349), .A2(n4703), .A3(n10219), .A4(n10348), .ZN(
        n10367) );
  NOR4_X1 U11436 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .A3(P1_ADDR_REG_3__SCAN_IN), .A4(P1_ADDR_REG_0__SCAN_IN), .ZN(n10350)
         );
  NAND4_X1 U11437 ( .A1(n10351), .A2(P1_ADDR_REG_5__SCAN_IN), .A3(n10350), 
        .A4(n10454), .ZN(n10352) );
  NOR4_X1 U11438 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n10354), .A3(n10353), 
        .A4(n10352), .ZN(n10366) );
  NAND4_X1 U11439 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(P1_REG0_REG_4__SCAN_IN), 
        .A3(n10484), .A4(n10487), .ZN(n10358) );
  NAND4_X1 U11440 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_REG2_REG_11__SCAN_IN), 
        .A3(P2_IR_REG_13__SCAN_IN), .A4(P2_REG1_REG_26__SCAN_IN), .ZN(n10356)
         );
  NAND4_X1 U11441 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P2_REG1_REG_24__SCAN_IN), 
        .A3(n10467), .A4(n10469), .ZN(n10355) );
  OR4_X1 U11442 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n10356), .A3(n10355), .A4(
        P2_REG0_REG_3__SCAN_IN), .ZN(n10357) );
  NOR4_X1 U11443 ( .A1(n10358), .A2(P2_ADDR_REG_15__SCAN_IN), .A3(n10448), 
        .A4(n10357), .ZN(n10365) );
  NAND4_X1 U11444 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), .A3(P2_REG3_REG_3__SCAN_IN), .A4(P2_REG0_REG_4__SCAN_IN), .ZN(n10363) );
  NAND4_X1 U11445 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(n10414), .A3(n10413), 
        .A4(n10359), .ZN(n10362) );
  NAND4_X1 U11446 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), 
        .A3(P2_REG0_REG_7__SCAN_IN), .A4(n10455), .ZN(n10361) );
  NAND4_X1 U11447 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n10438), .A3(n10440), 
        .A4(n10441), .ZN(n10360) );
  NOR4_X1 U11448 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10364) );
  NAND4_X1 U11449 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(
        n10368) );
  OAI21_X1 U11450 ( .B1(n10369), .B2(n10368), .A(P2_IR_REG_27__SCAN_IN), .ZN(
        n10498) );
  AOI22_X1 U11451 ( .A1(n10372), .A2(keyinput73), .B1(n10371), .B2(keyinput4), 
        .ZN(n10370) );
  OAI221_X1 U11452 ( .B1(n10372), .B2(keyinput73), .C1(n10371), .C2(keyinput4), 
        .A(n10370), .ZN(n10384) );
  AOI22_X1 U11453 ( .A1(n10375), .A2(keyinput126), .B1(keyinput13), .B2(n10374), .ZN(n10373) );
  OAI221_X1 U11454 ( .B1(n10375), .B2(keyinput126), .C1(n10374), .C2(
        keyinput13), .A(n10373), .ZN(n10383) );
  INV_X1 U11455 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U11456 ( .A1(n10378), .A2(keyinput1), .B1(n10377), .B2(keyinput106), 
        .ZN(n10376) );
  OAI221_X1 U11457 ( .B1(n10378), .B2(keyinput1), .C1(n10377), .C2(keyinput106), .A(n10376), .ZN(n10382) );
  XOR2_X1 U11458 ( .A(n5908), .B(keyinput94), .Z(n10380) );
  XNOR2_X1 U11459 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput18), .ZN(n10379) );
  NAND2_X1 U11460 ( .A1(n10380), .A2(n10379), .ZN(n10381) );
  NOR4_X1 U11461 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10429) );
  AOI22_X1 U11462 ( .A1(n10387), .A2(keyinput60), .B1(n10386), .B2(keyinput97), 
        .ZN(n10385) );
  OAI221_X1 U11463 ( .B1(n10387), .B2(keyinput60), .C1(n10386), .C2(keyinput97), .A(n10385), .ZN(n10390) );
  XOR2_X1 U11464 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput91), .Z(n10389) );
  XOR2_X1 U11465 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput124), .Z(n10388) );
  OR3_X1 U11466 ( .A1(n10390), .A2(n10389), .A3(n10388), .ZN(n10398) );
  XNOR2_X1 U11467 ( .A(n10391), .B(keyinput12), .ZN(n10397) );
  XNOR2_X1 U11468 ( .A(keyinput9), .B(n10392), .ZN(n10396) );
  XNOR2_X1 U11469 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput89), .ZN(n10394)
         );
  XNOR2_X1 U11470 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput62), .ZN(n10393) );
  NAND2_X1 U11471 ( .A1(n10394), .A2(n10393), .ZN(n10395) );
  NOR4_X1 U11472 ( .A1(n10398), .A2(n10397), .A3(n10396), .A4(n10395), .ZN(
        n10428) );
  AOI22_X1 U11473 ( .A1(n10401), .A2(keyinput114), .B1(keyinput15), .B2(n10400), .ZN(n10399) );
  OAI221_X1 U11474 ( .B1(n10401), .B2(keyinput114), .C1(n10400), .C2(
        keyinput15), .A(n10399), .ZN(n10411) );
  AOI22_X1 U11475 ( .A1(n10404), .A2(keyinput6), .B1(keyinput102), .B2(n10403), 
        .ZN(n10402) );
  OAI221_X1 U11476 ( .B1(n10404), .B2(keyinput6), .C1(n10403), .C2(keyinput102), .A(n10402), .ZN(n10410) );
  AOI22_X1 U11477 ( .A1(n9520), .A2(keyinput35), .B1(keyinput51), .B2(n10406), 
        .ZN(n10405) );
  OAI221_X1 U11478 ( .B1(n9520), .B2(keyinput35), .C1(n10406), .C2(keyinput51), 
        .A(n10405), .ZN(n10409) );
  AOI22_X1 U11479 ( .A1(n5701), .A2(keyinput68), .B1(keyinput78), .B2(n4868), 
        .ZN(n10407) );
  OAI221_X1 U11480 ( .B1(n5701), .B2(keyinput68), .C1(n4868), .C2(keyinput78), 
        .A(n10407), .ZN(n10408) );
  NOR4_X1 U11481 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10427) );
  AOI22_X1 U11482 ( .A1(n10414), .A2(keyinput7), .B1(keyinput57), .B2(n10413), 
        .ZN(n10412) );
  OAI221_X1 U11483 ( .B1(n10414), .B2(keyinput7), .C1(n10413), .C2(keyinput57), 
        .A(n10412), .ZN(n10425) );
  AOI22_X1 U11484 ( .A1(n10417), .A2(keyinput10), .B1(n10416), .B2(keyinput127), .ZN(n10415) );
  OAI221_X1 U11485 ( .B1(n10417), .B2(keyinput10), .C1(n10416), .C2(
        keyinput127), .A(n10415), .ZN(n10424) );
  XOR2_X1 U11486 ( .A(n10418), .B(keyinput112), .Z(n10422) );
  XNOR2_X1 U11487 ( .A(SI_30_), .B(keyinput3), .ZN(n10421) );
  XNOR2_X1 U11488 ( .A(SI_5_), .B(keyinput65), .ZN(n10420) );
  XNOR2_X1 U11489 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput41), .ZN(n10419) );
  NAND4_X1 U11490 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10423) );
  NOR3_X1 U11491 ( .A1(n10425), .A2(n10424), .A3(n10423), .ZN(n10426) );
  NAND4_X1 U11492 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10497) );
  INV_X1 U11493 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U11494 ( .A1(n10432), .A2(keyinput25), .B1(n10431), .B2(keyinput23), 
        .ZN(n10430) );
  OAI221_X1 U11495 ( .B1(n10432), .B2(keyinput25), .C1(n10431), .C2(keyinput23), .A(n10430), .ZN(n10445) );
  AOI22_X1 U11496 ( .A1(n10435), .A2(keyinput2), .B1(keyinput121), .B2(n10434), 
        .ZN(n10433) );
  OAI221_X1 U11497 ( .B1(n10435), .B2(keyinput2), .C1(n10434), .C2(keyinput121), .A(n10433), .ZN(n10444) );
  INV_X1 U11498 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U11499 ( .A1(n10438), .A2(keyinput19), .B1(keyinput0), .B2(n10437), 
        .ZN(n10436) );
  OAI221_X1 U11500 ( .B1(n10438), .B2(keyinput19), .C1(n10437), .C2(keyinput0), 
        .A(n10436), .ZN(n10443) );
  AOI22_X1 U11501 ( .A1(n10441), .A2(keyinput5), .B1(n10440), .B2(keyinput103), 
        .ZN(n10439) );
  OAI221_X1 U11502 ( .B1(n10441), .B2(keyinput5), .C1(n10440), .C2(keyinput103), .A(n10439), .ZN(n10442) );
  NOR4_X1 U11503 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10495) );
  AOI22_X1 U11504 ( .A1(n10448), .A2(keyinput53), .B1(keyinput67), .B2(n10447), 
        .ZN(n10446) );
  OAI221_X1 U11505 ( .B1(n10448), .B2(keyinput53), .C1(n10447), .C2(keyinput67), .A(n10446), .ZN(n10461) );
  AOI22_X1 U11506 ( .A1(n10451), .A2(keyinput95), .B1(n10450), .B2(keyinput119), .ZN(n10449) );
  OAI221_X1 U11507 ( .B1(n10451), .B2(keyinput95), .C1(n10450), .C2(
        keyinput119), .A(n10449), .ZN(n10460) );
  AOI22_X1 U11508 ( .A1(n10454), .A2(keyinput17), .B1(n10453), .B2(keyinput88), 
        .ZN(n10452) );
  OAI221_X1 U11509 ( .B1(n10454), .B2(keyinput17), .C1(n10453), .C2(keyinput88), .A(n10452), .ZN(n10459) );
  XOR2_X1 U11510 ( .A(n10455), .B(keyinput71), .Z(n10457) );
  XNOR2_X1 U11511 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput54), .ZN(n10456) );
  NAND2_X1 U11512 ( .A1(n10457), .A2(n10456), .ZN(n10458) );
  NOR4_X1 U11513 ( .A1(n10461), .A2(n10460), .A3(n10459), .A4(n10458), .ZN(
        n10494) );
  AOI22_X1 U11514 ( .A1(n10464), .A2(keyinput37), .B1(n10463), .B2(keyinput48), 
        .ZN(n10462) );
  OAI221_X1 U11515 ( .B1(n10464), .B2(keyinput37), .C1(n10463), .C2(keyinput48), .A(n10462), .ZN(n10476) );
  AOI22_X1 U11516 ( .A1(n10467), .A2(keyinput109), .B1(keyinput8), .B2(n10466), 
        .ZN(n10465) );
  OAI221_X1 U11517 ( .B1(n10467), .B2(keyinput109), .C1(n10466), .C2(keyinput8), .A(n10465), .ZN(n10475) );
  AOI22_X1 U11518 ( .A1(n10470), .A2(keyinput116), .B1(n10469), .B2(keyinput85), .ZN(n10468) );
  OAI221_X1 U11519 ( .B1(n10470), .B2(keyinput116), .C1(n10469), .C2(
        keyinput85), .A(n10468), .ZN(n10474) );
  XOR2_X1 U11520 ( .A(n9392), .B(keyinput64), .Z(n10472) );
  XNOR2_X1 U11521 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput39), .ZN(n10471)
         );
  NAND2_X1 U11522 ( .A1(n10472), .A2(n10471), .ZN(n10473) );
  NOR4_X1 U11523 ( .A1(n10476), .A2(n10475), .A3(n10474), .A4(n10473), .ZN(
        n10493) );
  AOI22_X1 U11524 ( .A1(n10479), .A2(keyinput55), .B1(n10478), .B2(keyinput70), 
        .ZN(n10477) );
  OAI221_X1 U11525 ( .B1(n10479), .B2(keyinput55), .C1(n10478), .C2(keyinput70), .A(n10477), .ZN(n10491) );
  INV_X1 U11526 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U11527 ( .A1(n10482), .A2(keyinput75), .B1(keyinput59), .B2(n10481), 
        .ZN(n10480) );
  OAI221_X1 U11528 ( .B1(n10482), .B2(keyinput75), .C1(n10481), .C2(keyinput59), .A(n10480), .ZN(n10490) );
  AOI22_X1 U11529 ( .A1(n10484), .A2(keyinput52), .B1(n9689), .B2(keyinput27), 
        .ZN(n10483) );
  OAI221_X1 U11530 ( .B1(n10484), .B2(keyinput52), .C1(n9689), .C2(keyinput27), 
        .A(n10483), .ZN(n10489) );
  INV_X1 U11531 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U11532 ( .A1(n10487), .A2(keyinput107), .B1(n10486), .B2(
        keyinput120), .ZN(n10485) );
  OAI221_X1 U11533 ( .B1(n10487), .B2(keyinput107), .C1(n10486), .C2(
        keyinput120), .A(n10485), .ZN(n10488) );
  NOR4_X1 U11534 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10492) );
  NAND4_X1 U11535 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(
        n10496) );
  AOI211_X1 U11536 ( .C1(keyinput108), .C2(n10498), .A(n10497), .B(n10496), 
        .ZN(n10499) );
  NAND4_X1 U11537 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10503) );
  XNOR2_X1 U11538 ( .A(n10504), .B(n10503), .ZN(n10506) );
  XNOR2_X1 U11539 ( .A(n10506), .B(n10505), .ZN(ADD_1068_U59) );
  OAI21_X1 U11540 ( .B1(n10509), .B2(n10508), .A(n10507), .ZN(ADD_1068_U50) );
  OAI21_X1 U11541 ( .B1(n10512), .B2(n10511), .A(n10510), .ZN(ADD_1068_U51) );
  AOI21_X1 U11542 ( .B1(n10515), .B2(n10514), .A(n10513), .ZN(ADD_1068_U54) );
  OAI21_X1 U11543 ( .B1(n10518), .B2(n10517), .A(n10516), .ZN(ADD_1068_U47) );
  OAI21_X1 U11544 ( .B1(n10521), .B2(n10520), .A(n10519), .ZN(ADD_1068_U48) );
  OAI21_X1 U11545 ( .B1(n10524), .B2(n10523), .A(n10522), .ZN(ADD_1068_U49) );
  AOI21_X1 U11546 ( .B1(n10527), .B2(n10526), .A(n10525), .ZN(ADD_1068_U53) );
  OAI21_X1 U11547 ( .B1(n10530), .B2(n10529), .A(n10528), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4911 ( .A(n9183), .Z(n4647) );
  CLKBUF_X1 U4924 ( .A(n5934), .Z(n9610) );
  CLKBUF_X1 U5068 ( .A(n6048), .Z(n9004) );
  CLKBUF_X1 U5629 ( .A(n9125), .Z(n4705) );
  CLKBUF_X1 U6423 ( .A(n8329), .Z(n4648) );
endmodule

