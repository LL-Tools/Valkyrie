

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9720, n9721, n9722, n9723, n9724, n9725, n9727, n9728, n9729, n9731,
         n9732, n9733, n9734, n9735, n9737, n9738, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501;

  INV_X2 U11164 ( .A(n20344), .ZN(n20330) );
  NOR2_X1 U11165 ( .A1(n11846), .A2(n10342), .ZN(n16083) );
  AND2_X1 U11166 ( .A1(n14510), .A2(n14335), .ZN(n20344) );
  INV_X1 U11168 ( .A(n19903), .ZN(n19907) );
  INV_X1 U11169 ( .A(n19767), .ZN(n19769) );
  OR2_X1 U11170 ( .A1(n19974), .A2(n20028), .ZN(n20086) );
  OR2_X1 U11171 ( .A1(n19944), .A2(n19949), .ZN(n20021) );
  NAND2_X1 U11173 ( .A1(n9780), .A2(n19064), .ZN(n18502) );
  AND2_X1 U11174 ( .A1(n16616), .A2(n16554), .ZN(n16570) );
  OR2_X1 U11175 ( .A1(n13328), .A2(n13322), .ZN(n13324) );
  AND3_X1 U11176 ( .A1(n19479), .A2(n10841), .A3(n13436), .ZN(n19686) );
  BUF_X1 U11177 ( .A(n11412), .Z(n11737) );
  CLKBUF_X2 U11178 ( .A(n11970), .Z(n17602) );
  BUF_X1 U11179 ( .A(n11892), .Z(n9724) );
  CLKBUF_X3 U11180 ( .A(n17457), .Z(n17613) );
  AND2_X1 U11181 ( .A1(n12988), .A2(n12920), .ZN(n10427) );
  CLKBUF_X2 U11182 ( .A(n10802), .Z(n11293) );
  CLKBUF_X2 U11183 ( .A(n11970), .Z(n16668) );
  INV_X1 U11184 ( .A(n11441), .ZN(n9742) );
  BUF_X1 U11185 ( .A(n11892), .Z(n9725) );
  AND2_X2 U11186 ( .A1(n10850), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10912) );
  BUF_X2 U11188 ( .A(n16669), .Z(n9721) );
  AND2_X2 U11189 ( .A1(n10749), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11246) );
  AND2_X1 U11190 ( .A1(n12691), .A2(n12816), .ZN(n14381) );
  AND2_X1 U11192 ( .A1(n10182), .A2(n10181), .ZN(n16669) );
  CLKBUF_X1 U11193 ( .A(n14485), .Z(n14450) );
  INV_X2 U11194 ( .A(n12146), .ZN(n19513) );
  CLKBUF_X2 U11195 ( .A(n12994), .Z(n14487) );
  CLKBUF_X2 U11196 ( .A(n14235), .Z(n14473) );
  CLKBUF_X2 U11197 ( .A(n14483), .Z(n14099) );
  CLKBUF_X2 U11198 ( .A(n12993), .Z(n14476) );
  NAND2_X1 U11199 ( .A1(n12141), .A2(n11397), .ZN(n10783) );
  CLKBUF_X1 U11200 ( .A(n12814), .Z(n20506) );
  NAND2_X1 U11201 ( .A1(n19234), .A2(n17332), .ZN(n17361) );
  INV_X2 U11202 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19234) );
  AND2_X1 U11204 ( .A1(n13018), .A2(n12813), .ZN(n12871) );
  AND2_X1 U11205 ( .A1(n10675), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13655) );
  AND2_X1 U11206 ( .A1(n13097), .A2(n21091), .ZN(n10158) );
  NAND2_X1 U11208 ( .A1(n10769), .A2(n13697), .ZN(n10792) );
  AND2_X1 U11210 ( .A1(n12662), .A2(n13451), .ZN(n12993) );
  NAND2_X1 U11211 ( .A1(n11121), .A2(n11744), .ZN(n11132) );
  INV_X1 U11212 ( .A(n11349), .ZN(n11352) );
  BUF_X1 U11213 ( .A(n10801), .Z(n11703) );
  NOR2_X1 U11214 ( .A1(n9938), .A2(n10830), .ZN(n19588) );
  OR2_X1 U11215 ( .A1(n18067), .A2(n18090), .ZN(n18027) );
  OR2_X1 U11216 ( .A1(n11864), .A2(n17361), .ZN(n9784) );
  AND2_X1 U11217 ( .A1(n13345), .A2(n14537), .ZN(n15339) );
  AND2_X1 U11218 ( .A1(n11671), .A2(n9906), .ZN(n11678) );
  INV_X1 U11219 ( .A(n11703), .ZN(n11715) );
  CLKBUF_X3 U11220 ( .A(n11397), .Z(n11789) );
  MUX2_X1 U11221 ( .A(n17970), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .S(
        n18199), .Z(n12126) );
  INV_X1 U11222 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10007) );
  INV_X1 U11223 ( .A(n11664), .ZN(n15742) );
  NAND2_X1 U11224 ( .A1(n16183), .A2(n11844), .ZN(n12450) );
  NAND2_X1 U11225 ( .A1(n11209), .A2(n11208), .ZN(n13765) );
  AND3_X1 U11226 ( .A1(n19479), .A2(n10836), .A3(n13436), .ZN(n19752) );
  INV_X1 U11227 ( .A(n17353), .ZN(n17366) );
  CLKBUF_X3 U11228 ( .A(n16669), .Z(n9722) );
  NOR2_X1 U11229 ( .A1(n16704), .A2(n18307), .ZN(n17939) );
  INV_X1 U11230 ( .A(n18117), .ZN(n18199) );
  NAND2_X1 U11231 ( .A1(n18621), .A2(n18584), .ZN(n18574) );
  INV_X1 U11232 ( .A(n20305), .ZN(n20334) );
  NOR2_X2 U11233 ( .A1(n13476), .A2(n13475), .ZN(n13577) );
  INV_X1 U11234 ( .A(n20604), .ZN(n20570) );
  NOR2_X1 U11235 ( .A1(n19808), .A2(n19742), .ZN(n19614) );
  INV_X1 U11236 ( .A(n19644), .ZN(n19676) );
  OAI21_X1 U11237 ( .B1(n19776), .B2(n19797), .A(n20033), .ZN(n19801) );
  INV_X1 U11238 ( .A(n19837), .ZN(n19872) );
  NOR2_X1 U11239 ( .A1(n19944), .A2(n19882), .ZN(n19940) );
  INV_X1 U11240 ( .A(n18164), .ZN(n18200) );
  INV_X1 U11241 ( .A(n18272), .ZN(n18281) );
  INV_X1 U11242 ( .A(n19260), .ZN(n18621) );
  AOI211_X1 U11243 ( .C1(n16311), .C2(n16640), .A(n16310), .B(n16309), .ZN(
        n16312) );
  INV_X1 U11244 ( .A(n16556), .ZN(n16846) );
  AOI211_X1 U11245 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17063), .A(n17062), 
        .B(n17061), .ZN(n17064) );
  NAND2_X1 U11246 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17372), .ZN(n17363) );
  NOR2_X1 U11247 ( .A1(n17992), .A2(n18145), .ZN(n18272) );
  NOR2_X1 U11248 ( .A1(n18502), .A2(n19060), .ZN(n18584) );
  OR2_X1 U11249 ( .A1(n11862), .A2(n19081), .ZN(n9720) );
  OAI21_X1 U11250 ( .B1(n13400), .B2(n12691), .A(n13405), .ZN(n10159) );
  NOR2_X4 U11251 ( .A1(n9747), .A2(n11647), .ZN(n11644) );
  NAND2_X2 U11252 ( .A1(n20460), .A2(n20452), .ZN(n20475) );
  NOR2_X2 U11253 ( .A1(n13274), .A2(n13356), .ZN(n13355) );
  AOI21_X2 U11254 ( .B1(n13663), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10035), 
        .ZN(n10034) );
  NOR2_X4 U11255 ( .A1(n15873), .A2(n15874), .ZN(n15868) );
  NOR2_X2 U11256 ( .A1(n15718), .A2(n16234), .ZN(n15708) );
  AND2_X4 U11257 ( .A1(n13441), .A2(n12958), .ZN(n14484) );
  NOR2_X1 U11258 ( .A1(n11863), .A2(n11861), .ZN(n11892) );
  OR2_X2 U11259 ( .A1(n17805), .A2(n10255), .ZN(n17779) );
  NOR2_X1 U11262 ( .A1(n11861), .A2(n19081), .ZN(n17457) );
  AOI21_X2 U11263 ( .B1(n16355), .B2(n16344), .A(n11800), .ZN(n16327) );
  NAND2_X4 U11264 ( .A1(n10107), .A2(n10271), .ZN(n13069) );
  NOR2_X1 U11265 ( .A1(n12129), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16850) );
  NOR2_X2 U11266 ( .A1(n11697), .A2(n15863), .ZN(n15862) );
  INV_X2 U11267 ( .A(n17505), .ZN(n9728) );
  INV_X1 U11268 ( .A(n17505), .ZN(n9729) );
  AND2_X1 U11269 ( .A1(n10307), .A2(n9858), .ZN(n10438) );
  AND2_X1 U11270 ( .A1(n10626), .A2(n9856), .ZN(n10166) );
  OAI21_X1 U11271 ( .B1(n14397), .B2(n10423), .A(n10422), .ZN(n15106) );
  INV_X1 U11272 ( .A(n12450), .ZN(n9731) );
  NOR2_X1 U11273 ( .A1(n14514), .A2(n10657), .ZN(n15821) );
  XNOR2_X1 U11274 ( .A(n11799), .B(n11741), .ZN(n15910) );
  AOI21_X1 U11275 ( .B1(n16848), .B2(n18117), .A(n16847), .ZN(n12129) );
  NAND2_X1 U11276 ( .A1(n16799), .A2(n14373), .ZN(n10395) );
  NOR2_X1 U11277 ( .A1(n15160), .A2(n10645), .ZN(n15125) );
  BUF_X2 U11278 ( .A(n10120), .Z(n15210) );
  INV_X1 U11279 ( .A(n14392), .ZN(n10420) );
  NAND2_X1 U11280 ( .A1(n9809), .A2(n10930), .ZN(n10148) );
  NOR2_X2 U11281 ( .A1(n19221), .A2(n18218), .ZN(n18145) );
  INV_X1 U11282 ( .A(n10601), .ZN(n10403) );
  INV_X2 U11283 ( .A(n18122), .ZN(n18202) );
  NAND2_X1 U11284 ( .A1(n13102), .A2(n13101), .ZN(n20568) );
  NOR2_X2 U11285 ( .A1(n9938), .A2(n19494), .ZN(n10950) );
  CLKBUF_X1 U11286 ( .A(n13370), .Z(n13102) );
  CLKBUF_X1 U11287 ( .A(n10945), .Z(n19982) );
  OR2_X1 U11288 ( .A1(n10837), .A2(n13436), .ZN(n19811) );
  NAND2_X1 U11289 ( .A1(n10389), .A2(n10388), .ZN(n13370) );
  OR2_X1 U11290 ( .A1(n10839), .A2(n13436), .ZN(n19884) );
  AND2_X1 U11291 ( .A1(n10831), .A2(n9810), .ZN(n19717) );
  NAND2_X1 U11292 ( .A1(n10157), .A2(n13099), .ZN(n13400) );
  CLKBUF_X1 U11293 ( .A(n18584), .Z(n9743) );
  NOR2_X1 U11294 ( .A1(n17779), .A2(n17901), .ZN(n17773) );
  OAI21_X1 U11295 ( .B1(n13020), .B2(n9961), .A(n9748), .ZN(n13237) );
  XNOR2_X1 U11296 ( .A(n10818), .B(n10813), .ZN(n10821) );
  AND2_X1 U11297 ( .A1(n10773), .A2(n10772), .ZN(n10818) );
  NAND2_X1 U11298 ( .A1(n12623), .A2(n9832), .ZN(n12088) );
  NOR2_X1 U11299 ( .A1(n18621), .A2(n17908), .ZN(n17909) );
  NAND2_X1 U11300 ( .A1(n10442), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10800) );
  CLKBUF_X2 U11301 ( .A(n10787), .Z(n13663) );
  NAND2_X1 U11302 ( .A1(n10223), .A2(n10225), .ZN(n10548) );
  NAND2_X1 U11303 ( .A1(n11574), .A2(n11352), .ZN(n13632) );
  OR2_X1 U11304 ( .A1(n11240), .A2(n10780), .ZN(n10781) );
  NOR2_X1 U11305 ( .A1(n17797), .A2(n12101), .ZN(n12103) );
  NOR2_X1 U11306 ( .A1(n11349), .A2(n11722), .ZN(n10794) );
  CLKBUF_X1 U11307 ( .A(n10766), .Z(n19523) );
  AND2_X1 U11309 ( .A1(n12864), .A2(n10008), .ZN(n12825) );
  CLKBUF_X2 U11311 ( .A(n12882), .Z(n15472) );
  AND4_X1 U11312 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n10661) );
  AND2_X1 U11313 ( .A1(n10282), .A2(n10283), .ZN(n12169) );
  NAND2_X2 U11315 ( .A1(n9782), .A2(n10674), .ZN(n12888) );
  NAND2_X2 U11316 ( .A1(n12670), .A2(n12669), .ZN(n12812) );
  AND4_X1 U11317 ( .A1(n12779), .A2(n12778), .A3(n12777), .A4(n12776), .ZN(
        n12785) );
  INV_X2 U11318 ( .A(n12532), .ZN(n12500) );
  CLKBUF_X2 U11319 ( .A(n14486), .Z(n14230) );
  BUF_X2 U11320 ( .A(n14119), .Z(n14477) );
  BUF_X2 U11321 ( .A(n14482), .Z(n9740) );
  BUF_X2 U11322 ( .A(n14488), .Z(n14171) );
  INV_X4 U11323 ( .A(n18481), .ZN(n9732) );
  CLKBUF_X2 U11324 ( .A(n12001), .Z(n17563) );
  AND2_X2 U11325 ( .A1(n10749), .A2(n11030), .ZN(n10882) );
  CLKBUF_X2 U11326 ( .A(n11903), .Z(n17595) );
  CLKBUF_X3 U11327 ( .A(n11963), .Z(n9737) );
  BUF_X2 U11328 ( .A(n14449), .Z(n14472) );
  NOR2_X1 U11329 ( .A1(n11864), .A2(n11860), .ZN(n11963) );
  INV_X2 U11331 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n13022) );
  INV_X4 U11333 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19226) );
  NAND2_X1 U11334 ( .A1(n10166), .A2(n10167), .ZN(n10165) );
  AND2_X1 U11335 ( .A1(n9985), .A2(n16150), .ZN(n16469) );
  NAND2_X1 U11336 ( .A1(n9731), .A2(n9919), .ZN(n9935) );
  AOI21_X1 U11337 ( .B1(n10343), .B2(n9777), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16068) );
  NOR2_X1 U11338 ( .A1(n16212), .A2(n16205), .ZN(n16204) );
  NOR2_X1 U11339 ( .A1(n15159), .A2(n15126), .ZN(n15148) );
  NAND3_X1 U11340 ( .A1(n11775), .A2(n9799), .A3(n11774), .ZN(n10600) );
  NAND2_X1 U11341 ( .A1(n10371), .A2(n10220), .ZN(n10115) );
  AND2_X1 U11342 ( .A1(n16183), .A2(n9778), .ZN(n16032) );
  NAND2_X1 U11343 ( .A1(n14397), .A2(n10114), .ZN(n10021) );
  OR2_X1 U11344 ( .A1(n14599), .A2(n14246), .ZN(n9989) );
  NAND2_X1 U11345 ( .A1(n15821), .A2(n15820), .ZN(n15819) );
  NAND2_X1 U11346 ( .A1(n15493), .A2(n15492), .ZN(n16300) );
  NAND3_X1 U11347 ( .A1(n10378), .A2(n14391), .A3(n10376), .ZN(n15209) );
  NAND2_X1 U11348 ( .A1(n10395), .A2(n10379), .ZN(n10378) );
  OAI21_X1 U11349 ( .B1(n17939), .B2(n18117), .A(n16907), .ZN(n17935) );
  NOR2_X1 U11350 ( .A1(n16706), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16848) );
  NAND2_X1 U11351 ( .A1(n16265), .A2(n16266), .ZN(n11597) );
  INV_X1 U11352 ( .A(n10370), .ZN(n10369) );
  AND2_X1 U11353 ( .A1(n15125), .A2(n14361), .ZN(n14395) );
  AND2_X1 U11354 ( .A1(n16704), .A2(n18307), .ZN(n17940) );
  AND2_X1 U11355 ( .A1(n11607), .A2(n11606), .ZN(n16235) );
  NAND2_X1 U11356 ( .A1(n11602), .A2(n16569), .ZN(n16246) );
  AND2_X1 U11357 ( .A1(n10630), .A2(n9916), .ZN(n10220) );
  OR2_X1 U11358 ( .A1(n11605), .A2(n11604), .ZN(n11607) );
  NAND2_X1 U11359 ( .A1(n14385), .A2(n16811), .ZN(n16793) );
  XNOR2_X1 U11360 ( .A(n11605), .B(n11792), .ZN(n11602) );
  AND2_X1 U11361 ( .A1(n10134), .A2(n10133), .ZN(n16226) );
  OR3_X1 U11362 ( .A1(n19980), .A2(n19979), .A3(n19978), .ZN(n20018) );
  NAND2_X1 U11363 ( .A1(n10125), .A2(n10124), .ZN(n16225) );
  NAND2_X1 U11364 ( .A1(n11596), .A2(n11792), .ZN(n10129) );
  NAND2_X1 U11365 ( .A1(n10056), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16268) );
  XNOR2_X1 U11366 ( .A(n11791), .B(n11790), .ZN(n12467) );
  INV_X1 U11367 ( .A(n10028), .ZN(n10582) );
  INV_X1 U11368 ( .A(n11595), .ZN(n10056) );
  NAND2_X1 U11369 ( .A1(n10142), .A2(n10148), .ZN(n10028) );
  NAND2_X1 U11370 ( .A1(n13903), .A2(n13902), .ZN(n15005) );
  XNOR2_X1 U11371 ( .A(n10420), .B(n15344), .ZN(n15175) );
  AND2_X1 U11372 ( .A1(n17971), .A2(n9886), .ZN(n10221) );
  NAND2_X1 U11373 ( .A1(n13584), .A2(n13583), .ZN(n13891) );
  OAI21_X1 U11374 ( .B1(n13617), .B2(n13874), .A(n13616), .ZN(n13905) );
  XNOR2_X1 U11375 ( .A(n10972), .B(n10148), .ZN(n11595) );
  NOR2_X1 U11376 ( .A1(n18317), .A2(n17961), .ZN(n18302) );
  INV_X2 U11377 ( .A(n14392), .ZN(n15189) );
  NAND2_X1 U11378 ( .A1(n13574), .A2(n10628), .ZN(n10627) );
  NAND2_X2 U11379 ( .A1(n14366), .A2(n14358), .ZN(n14392) );
  NAND2_X1 U11380 ( .A1(n10443), .A2(n10971), .ZN(n10972) );
  INV_X1 U11381 ( .A(n20021), .ZN(n20010) );
  INV_X1 U11382 ( .A(n17975), .ZN(n17970) );
  INV_X1 U11383 ( .A(n18428), .ZN(n18016) );
  NAND2_X1 U11384 ( .A1(n9817), .A2(n9756), .ZN(n10443) );
  NOR2_X2 U11385 ( .A1(n19742), .A2(n19949), .ZN(n19738) );
  OR2_X1 U11386 ( .A1(n11164), .A2(n16394), .ZN(n16112) );
  NAND2_X1 U11387 ( .A1(n9841), .A2(n10403), .ZN(n14366) );
  NOR2_X2 U11388 ( .A1(n19742), .A2(n20028), .ZN(n19794) );
  NAND2_X1 U11389 ( .A1(n9753), .A2(n10014), .ZN(n13576) );
  NAND2_X1 U11390 ( .A1(n10403), .A2(n10404), .ZN(n13574) );
  NAND2_X1 U11391 ( .A1(n18282), .A2(n12582), .ZN(n18164) );
  NAND2_X1 U11392 ( .A1(n18475), .A2(n18415), .ZN(n18109) );
  NAND2_X1 U11393 ( .A1(n16901), .A2(n10386), .ZN(n18428) );
  NAND2_X1 U11394 ( .A1(n18076), .A2(n18396), .ZN(n18075) );
  OR2_X1 U11395 ( .A1(n18292), .A2(n12582), .ZN(n18122) );
  AND4_X1 U11396 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n10849) );
  NAND2_X1 U11397 ( .A1(n13385), .A2(n9980), .ZN(n13386) );
  INV_X1 U11398 ( .A(n18261), .ZN(n18293) );
  NAND2_X1 U11399 ( .A1(n18051), .A2(n18289), .ZN(n18008) );
  INV_X1 U11400 ( .A(n18292), .ZN(n18282) );
  INV_X1 U11401 ( .A(n14423), .ZN(n20459) );
  INV_X1 U11402 ( .A(n13385), .ZN(n9979) );
  OAI22_X1 U11403 ( .A1(n21480), .A2(n19559), .B1(n10834), .B2(n10833), .ZN(
        n10835) );
  AND2_X1 U11404 ( .A1(n18027), .A2(n10240), .ZN(n10239) );
  NOR2_X2 U11406 ( .A1(n19260), .A2(n17005), .ZN(n18261) );
  AOI21_X1 U11407 ( .B1(n18027), .B2(n9757), .A(n9904), .ZN(n10236) );
  OR2_X1 U11408 ( .A1(n9994), .A2(P3_EBX_REG_27__SCAN_IN), .ZN(n17073) );
  CLKBUF_X1 U11409 ( .A(n10944), .Z(n19915) );
  AND2_X1 U11410 ( .A1(n10365), .A2(n10830), .ZN(n19779) );
  NAND2_X1 U11411 ( .A1(n18165), .A2(n18116), .ZN(n18509) );
  AND2_X1 U11412 ( .A1(n10365), .A2(n19494), .ZN(n19851) );
  AOI22_X1 U11413 ( .A1(n19654), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n20023), .ZN(n10825) );
  AOI22_X1 U11414 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19717), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U11415 ( .A1(n13370), .A2(n13369), .ZN(n13385) );
  AND2_X1 U11416 ( .A1(n13289), .A2(n12157), .ZN(n13312) );
  NOR2_X1 U11417 ( .A1(n13749), .A2(n13761), .ZN(n13760) );
  NAND2_X1 U11418 ( .A1(n10012), .A2(n13474), .ZN(n20750) );
  AND2_X1 U11419 ( .A1(n10824), .A2(n10832), .ZN(n10944) );
  AND2_X1 U11420 ( .A1(n10832), .A2(n10831), .ZN(n10945) );
  OR2_X1 U11421 ( .A1(n10839), .A2(n15771), .ZN(n19620) );
  OR2_X1 U11422 ( .A1(n10837), .A2(n15771), .ZN(n19559) );
  NAND2_X1 U11423 ( .A1(n12172), .A2(n12148), .ZN(n13492) );
  AND3_X1 U11424 ( .A1(n19479), .A2(n15771), .A3(n10836), .ZN(n20023) );
  AND3_X1 U11425 ( .A1(n19479), .A2(n15771), .A3(n10841), .ZN(n19946) );
  CLKBUF_X1 U11426 ( .A(n13463), .Z(n20775) );
  AND2_X1 U11427 ( .A1(n10830), .A2(n19479), .ZN(n10824) );
  NOR2_X1 U11428 ( .A1(n12115), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10242) );
  AND2_X1 U11429 ( .A1(n15813), .A2(n10822), .ZN(n10841) );
  NAND2_X1 U11430 ( .A1(n17773), .A2(n17661), .ZN(n17751) );
  INV_X1 U11431 ( .A(n15773), .ZN(n11425) );
  NOR2_X1 U11432 ( .A1(n16835), .A2(n10822), .ZN(n10836) );
  NAND2_X1 U11433 ( .A1(n20541), .A2(n10158), .ZN(n10157) );
  AND2_X1 U11434 ( .A1(n12947), .A2(n21091), .ZN(n9984) );
  NAND2_X1 U11435 ( .A1(n10155), .A2(n13011), .ZN(n13229) );
  NAND2_X2 U11436 ( .A1(n12753), .A2(n12752), .ZN(n13328) );
  XNOR2_X1 U11437 ( .A(n11618), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U11438 ( .A1(n20608), .A2(n10113), .ZN(n20541) );
  NAND3_X1 U11439 ( .A1(n10184), .A2(n10815), .A3(n10183), .ZN(n10112) );
  INV_X2 U11440 ( .A(n15887), .ZN(n9733) );
  NAND2_X1 U11441 ( .A1(n13237), .A2(n13096), .ZN(n13369) );
  NAND2_X1 U11443 ( .A1(n12751), .A2(n12750), .ZN(n12753) );
  INV_X2 U11444 ( .A(n13154), .ZN(n9734) );
  OR2_X2 U11445 ( .A1(n11074), .A2(n19534), .ZN(n11744) );
  BUF_X1 U11446 ( .A(n10814), .Z(n10817) );
  OAI21_X1 U11447 ( .B1(n16777), .B2(n16776), .A(n19258), .ZN(n17805) );
  OR2_X1 U11448 ( .A1(n10801), .A2(n16617), .ZN(n10807) );
  NAND2_X1 U11449 ( .A1(n10033), .A2(n10795), .ZN(n10811) );
  NAND3_X1 U11450 ( .A1(n10029), .A2(n10800), .A3(n10198), .ZN(n10810) );
  INV_X1 U11451 ( .A(n10819), .ZN(n10813) );
  INV_X2 U11452 ( .A(n17658), .ZN(n9735) );
  OAI22_X1 U11453 ( .A1(n10800), .A2(n11030), .B1(n10799), .B2(n20188), .ZN(
        n10808) );
  NAND2_X1 U11454 ( .A1(n18244), .A2(n18544), .ZN(n18243) );
  INV_X2 U11455 ( .A(n17362), .ZN(n17294) );
  OAI211_X1 U11456 ( .C1(n10548), .C2(n12104), .A(n9798), .B(n10000), .ZN(
        n18244) );
  AND3_X1 U11457 ( .A1(n12919), .A2(n10663), .A3(n12918), .ZN(n12987) );
  NAND2_X1 U11458 ( .A1(n12903), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10402) );
  AND2_X1 U11459 ( .A1(n10314), .A2(n10313), .ZN(n16691) );
  NOR3_X1 U11460 ( .A1(n12042), .A2(n12041), .A3(n12040), .ZN(n12074) );
  NAND2_X2 U11461 ( .A1(n17854), .A2(n19104), .ZN(n17919) );
  NAND3_X1 U11462 ( .A1(n10311), .A2(n10312), .A3(n11357), .ZN(n10442) );
  NAND2_X2 U11463 ( .A1(n12582), .A2(n12112), .ZN(n18117) );
  AND2_X1 U11464 ( .A1(n18234), .A2(n10560), .ZN(n10557) );
  AND3_X1 U11465 ( .A1(n12917), .A2(n10604), .A3(n10603), .ZN(n10663) );
  NAND2_X1 U11466 ( .A1(n12035), .A2(n10060), .ZN(n12046) );
  NAND2_X1 U11467 ( .A1(n10477), .A2(n10473), .ZN(n12639) );
  XNOR2_X1 U11468 ( .A(n17790), .B(n12108), .ZN(n18234) );
  INV_X2 U11469 ( .A(n11720), .ZN(n11711) );
  NOR2_X1 U11470 ( .A1(n10061), .A2(n10064), .ZN(n10060) );
  XNOR2_X1 U11471 ( .A(n12102), .B(n18556), .ZN(n10225) );
  AND2_X1 U11472 ( .A1(n13067), .A2(n9893), .ZN(n10195) );
  CLKBUF_X1 U11473 ( .A(n11240), .Z(n13686) );
  NOR2_X1 U11474 ( .A1(n12087), .A2(n12069), .ZN(n12478) );
  AND2_X1 U11475 ( .A1(n11215), .A2(n9944), .ZN(n10123) );
  NAND2_X1 U11476 ( .A1(n9795), .A2(n10794), .ZN(n11720) );
  NOR2_X1 U11477 ( .A1(n17929), .A2(n17922), .ZN(n12592) );
  AND2_X1 U11478 ( .A1(n10794), .A2(n12412), .ZN(n13067) );
  AND2_X1 U11479 ( .A1(n12890), .A2(n12889), .ZN(n12956) );
  INV_X1 U11480 ( .A(n12038), .ZN(n10061) );
  NAND2_X1 U11481 ( .A1(n10763), .A2(n11352), .ZN(n12411) );
  XNOR2_X1 U11482 ( .A(n10180), .B(n17797), .ZN(n12102) );
  NOR2_X1 U11483 ( .A1(n11434), .A2(n11534), .ZN(n10533) );
  NOR2_X1 U11484 ( .A1(n18640), .A2(n18636), .ZN(n12038) );
  CLKBUF_X1 U11485 ( .A(n12979), .Z(n14418) );
  NAND2_X1 U11486 ( .A1(n10412), .A2(n12799), .ZN(n12935) );
  INV_X2 U11487 ( .A(n11441), .ZN(n11736) );
  INV_X1 U11488 ( .A(n12077), .ZN(n18625) );
  NOR2_X1 U11489 ( .A1(n18636), .A2(n12077), .ZN(n12086) );
  AND2_X1 U11490 ( .A1(n10784), .A2(n10270), .ZN(n12412) );
  INV_X2 U11491 ( .A(n10840), .ZN(n13063) );
  NOR2_X1 U11492 ( .A1(n9991), .A2(n19518), .ZN(n9990) );
  NAND2_X1 U11493 ( .A1(n10762), .A2(n19518), .ZN(n11349) );
  INV_X1 U11494 ( .A(n10767), .ZN(n10763) );
  NAND2_X2 U11495 ( .A1(n13381), .A2(n13382), .ZN(n13833) );
  NAND2_X1 U11496 ( .A1(n10002), .A2(n17808), .ZN(n12101) );
  AND2_X1 U11497 ( .A1(n12982), .A2(n12900), .ZN(n12953) );
  NAND2_X1 U11498 ( .A1(n10708), .A2(n10707), .ZN(n10762) );
  CLKBUF_X3 U11499 ( .A(n10765), .Z(n13685) );
  NAND2_X2 U11500 ( .A1(n10765), .A2(n12146), .ZN(n11722) );
  INV_X1 U11501 ( .A(n17800), .ZN(n10002) );
  AND2_X2 U11502 ( .A1(n12711), .A2(n12812), .ZN(n13830) );
  OR3_X2 U11503 ( .A1(n10250), .A2(n10248), .A3(n10249), .ZN(n19260) );
  CLKBUF_X1 U11504 ( .A(n12899), .Z(n12914) );
  AND2_X1 U11505 ( .A1(n12798), .A2(n12691), .ZN(n10412) );
  INV_X1 U11506 ( .A(n12823), .ZN(n10020) );
  CLKBUF_X1 U11507 ( .A(n12141), .Z(n19541) );
  INV_X1 U11508 ( .A(n12871), .ZN(n13205) );
  NAND3_X2 U11509 ( .A1(n9781), .A2(n10661), .A3(n10642), .ZN(n17808) );
  INV_X2 U11510 ( .A(U212), .ZN(n16947) );
  NAND2_X1 U11511 ( .A1(n10748), .A2(n10747), .ZN(n10765) );
  INV_X1 U11512 ( .A(n12891), .ZN(n13323) );
  AND3_X1 U11513 ( .A1(n11915), .A2(n9761), .A3(n9844), .ZN(n17797) );
  NAND4_X2 U11514 ( .A1(n11024), .A2(n11023), .A3(n11022), .A4(n11021), .ZN(
        n11813) );
  NAND2_X2 U11515 ( .A1(n10761), .A2(n10760), .ZN(n12146) );
  OR2_X1 U11516 ( .A1(n10861), .A2(n10860), .ZN(n11582) );
  AND2_X2 U11517 ( .A1(n10111), .A2(n10110), .ZN(n19529) );
  NAND2_X1 U11518 ( .A1(n10109), .A2(n10108), .ZN(n19518) );
  NAND2_X1 U11519 ( .A1(n11397), .A2(n12169), .ZN(n11212) );
  NAND2_X1 U11520 ( .A1(n10048), .A2(n10047), .ZN(n12891) );
  AND2_X2 U11521 ( .A1(n10285), .A2(n10284), .ZN(n11397) );
  NAND4_X1 U11522 ( .A1(n10706), .A2(n10705), .A3(n10704), .A4(n10703), .ZN(
        n10707) );
  NAND2_X2 U11523 ( .A1(n12888), .A2(n12814), .ZN(n14416) );
  AND3_X1 U11524 ( .A1(n11900), .A2(n11899), .A3(n11898), .ZN(n10642) );
  INV_X2 U11525 ( .A(n12814), .ZN(n12691) );
  AND2_X1 U11526 ( .A1(n12812), .A2(n20532), .ZN(n12880) );
  NOR2_X2 U11527 ( .A1(n20487), .A2(n20485), .ZN(n20486) );
  OR2_X2 U11528 ( .A1(n12795), .A2(n12794), .ZN(n20532) );
  NOR2_X1 U11529 ( .A1(n12772), .A2(n12771), .ZN(n12773) );
  NOR2_X1 U11530 ( .A1(n10050), .A2(n10049), .ZN(n10048) );
  INV_X2 U11531 ( .A(U214), .ZN(n16957) );
  AND4_X1 U11532 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n12670) );
  AND4_X1 U11533 ( .A1(n12761), .A2(n12760), .A3(n12756), .A4(n12757), .ZN(
        n10047) );
  AND4_X1 U11534 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10732) );
  AND4_X1 U11535 ( .A1(n12765), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12774) );
  NAND2_X2 U11536 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20158), .ZN(n20162) );
  INV_X4 U11537 ( .A(n9784), .ZN(n17615) );
  NAND2_X1 U11538 ( .A1(n10081), .A2(n10080), .ZN(n17566) );
  BUF_X2 U11539 ( .A(n17597), .Z(n17617) );
  NAND3_X2 U11540 ( .A1(n19274), .A2(n19263), .A3(n19273), .ZN(n18481) );
  INV_X2 U11541 ( .A(n10640), .ZN(n17553) );
  INV_X2 U11542 ( .A(n16990), .ZN(U215) );
  AND2_X2 U11543 ( .A1(n10850), .A2(n11030), .ZN(n10885) );
  NAND2_X2 U11544 ( .A1(n19272), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19189) );
  NOR2_X2 U11545 ( .A1(n18853), .A2(n18756), .ZN(n18843) );
  AND2_X1 U11546 ( .A1(n15798), .A2(n19477), .ZN(n15780) );
  CLKBUF_X1 U11547 ( .A(n10850), .Z(n12393) );
  BUF_X2 U11548 ( .A(n14484), .Z(n13515) );
  BUF_X2 U11549 ( .A(n12780), .Z(n14102) );
  INV_X1 U11550 ( .A(n9784), .ZN(n9738) );
  CLKBUF_X1 U11551 ( .A(n14474), .Z(n14229) );
  NAND2_X1 U11552 ( .A1(n10383), .A2(n10382), .ZN(n17505) );
  NAND2_X1 U11553 ( .A1(n11855), .A2(n11865), .ZN(n17333) );
  AND2_X2 U11554 ( .A1(n12401), .A2(n11030), .ZN(n12257) );
  AND2_X2 U11555 ( .A1(n12400), .A2(n11030), .ZN(n12256) );
  AND2_X2 U11556 ( .A1(n12265), .A2(n11030), .ZN(n10864) );
  NOR2_X1 U11557 ( .A1(n21384), .A2(n18194), .ZN(n18192) );
  NAND2_X1 U11558 ( .A1(n19234), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11863) );
  NAND3_X1 U11559 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11622), .A3(
        n9760), .ZN(n11631) );
  AND2_X1 U11560 ( .A1(n12726), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12656) );
  AND2_X1 U11561 ( .A1(n10219), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12662) );
  AND2_X1 U11562 ( .A1(n15469), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10153) );
  AND2_X2 U11563 ( .A1(n12962), .A2(n12655), .ZN(n14485) );
  NAND2_X1 U11564 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10245) );
  NAND2_X2 U11565 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19081) );
  INV_X1 U11566 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10040) );
  AND2_X2 U11567 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13629) );
  INV_X1 U11568 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13627) );
  INV_X1 U11569 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10676) );
  INV_X1 U11570 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10677) );
  INV_X2 U11571 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10789) );
  AND2_X1 U11572 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12963) );
  NOR2_X2 U11573 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17267), .ZN(n17252) );
  INV_X2 U11574 ( .A(n12819), .ZN(n13018) );
  NOR2_X2 U11575 ( .A1(n14750), .A2(n10607), .ZN(n14691) );
  INV_X1 U11576 ( .A(n10823), .ZN(n15771) );
  NOR2_X1 U11577 ( .A1(n10823), .A2(n15813), .ZN(n10832) );
  NOR2_X2 U11578 ( .A1(n12085), .A2(n18636), .ZN(n16778) );
  NOR2_X2 U11579 ( .A1(n19343), .A2(n19319), .ZN(n15631) );
  NOR2_X4 U11580 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13451) );
  NOR2_X2 U11581 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12962) );
  OAI22_X2 U11582 ( .A1(n16429), .A2(n16628), .B1(n16430), .B2(n16629), .ZN(
        n16616) );
  INV_X4 U11583 ( .A(n10640), .ZN(n9741) );
  NOR2_X2 U11584 ( .A1(n17969), .A2(n11962), .ZN(n18303) );
  NOR2_X2 U11585 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13438) );
  NAND2_X4 U11586 ( .A1(n11621), .A2(n11620), .ZN(n11664) );
  NOR2_X2 U11587 ( .A1(n17073), .A2(P3_EBX_REG_28__SCAN_IN), .ZN(n17058) );
  NOR2_X2 U11588 ( .A1(n16647), .A2(n15797), .ZN(n15798) );
  NAND2_X1 U11589 ( .A1(n12146), .A2(n19977), .ZN(n11441) );
  OR2_X2 U11590 ( .A1(n20421), .A2(n13413), .ZN(n20433) );
  AND2_X2 U11591 ( .A1(n20253), .A2(n13245), .ZN(n20421) );
  AND2_X1 U11592 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12655) );
  NOR2_X1 U11593 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12661) );
  INV_X1 U11594 ( .A(n10792), .ZN(n10802) );
  NAND2_X1 U11595 ( .A1(n10402), .A2(n12905), .ZN(n10398) );
  OAI211_X1 U11596 ( .C1(n9983), .C2(n13384), .A(n10010), .B(n9982), .ZN(n9981) );
  NAND2_X1 U11597 ( .A1(n10011), .A2(n9790), .ZN(n10010) );
  NAND2_X1 U11598 ( .A1(n9983), .A2(n10009), .ZN(n9982) );
  NAND2_X1 U11599 ( .A1(n9984), .A2(n12948), .ZN(n9983) );
  AND2_X1 U11600 ( .A1(n19529), .A2(n12169), .ZN(n10784) );
  NAND2_X1 U11601 ( .A1(n10732), .A2(n11030), .ZN(n10285) );
  NAND2_X1 U11602 ( .A1(n10099), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10098) );
  INV_X1 U11603 ( .A(n11784), .ZN(n10099) );
  AND3_X1 U11604 ( .A1(n16063), .A2(n11773), .A3(n16061), .ZN(n11774) );
  AND4_X1 U11605 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11024) );
  AND4_X1 U11606 ( .A1(n11006), .A2(n11005), .A3(n11004), .A4(n11003), .ZN(
        n11023) );
  NOR2_X1 U11607 ( .A1(n11020), .A2(n11019), .ZN(n11021) );
  AOI21_X1 U11608 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18611), .A(
        n12059), .ZN(n12065) );
  NOR2_X1 U11609 ( .A1(n16691), .A2(n17855), .ZN(n12623) );
  NAND2_X1 U11610 ( .A1(n10718), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10271) );
  NAND2_X1 U11611 ( .A1(n10713), .A2(n11030), .ZN(n10107) );
  NOR2_X1 U11612 ( .A1(n12476), .A2(n19059), .ZN(n16695) );
  AND4_X1 U11613 ( .A1(n10900), .A2(n10899), .A3(n10898), .A4(n10897), .ZN(
        n10910) );
  AOI22_X1 U11614 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19654), .B1(
        n10945), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10899) );
  NOR2_X1 U11615 ( .A1(n15127), .A2(n9749), .ZN(n14400) );
  NAND2_X1 U11616 ( .A1(n10015), .A2(n10013), .ZN(n10404) );
  OR2_X1 U11617 ( .A1(n13474), .A2(n10014), .ZN(n10013) );
  NAND2_X1 U11618 ( .A1(n13463), .A2(n10016), .ZN(n10015) );
  AND2_X1 U11619 ( .A1(n13536), .A2(n21091), .ZN(n10016) );
  NAND2_X1 U11620 ( .A1(n9840), .A2(n12825), .ZN(n10411) );
  INV_X1 U11621 ( .A(n13830), .ZN(n13835) );
  NOR2_X1 U11622 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12663), .ZN(
        n12664) );
  NAND2_X1 U11623 ( .A1(n12818), .A2(n12813), .ZN(n12823) );
  NAND2_X1 U11624 ( .A1(n10781), .A2(n10310), .ZN(n10312) );
  NAND2_X1 U11625 ( .A1(n10054), .A2(n10778), .ZN(n10311) );
  NAND2_X1 U11626 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  INV_X1 U11627 ( .A(n11353), .ZN(n10777) );
  OR2_X1 U11628 ( .A1(n15610), .A2(n11792), .ZN(n11165) );
  AND2_X1 U11629 ( .A1(n9809), .A2(n10443), .ZN(n9977) );
  AND2_X1 U11630 ( .A1(n10930), .A2(n10971), .ZN(n9978) );
  NAND2_X1 U11631 ( .A1(n10032), .A2(n9820), .ZN(n10797) );
  NAND2_X1 U11632 ( .A1(n10188), .A2(n9795), .ZN(n10189) );
  NOR2_X1 U11633 ( .A1(n12114), .A2(n12113), .ZN(n12115) );
  INV_X1 U11634 ( .A(n12084), .ZN(n10313) );
  AND2_X1 U11635 ( .A1(n17332), .A2(n19079), .ZN(n10383) );
  AND3_X1 U11636 ( .A1(n12898), .A2(n13018), .A3(n12818), .ZN(n12864) );
  OR2_X1 U11637 ( .A1(n15472), .A2(n21091), .ZN(n14465) );
  INV_X1 U11638 ( .A(n14328), .ZN(n14468) );
  INV_X1 U11639 ( .A(n14647), .ZN(n10454) );
  AND2_X1 U11640 ( .A1(n10631), .A2(n14400), .ZN(n10630) );
  NOR2_X1 U11641 ( .A1(n15199), .A2(n9749), .ZN(n15159) );
  INV_X1 U11642 ( .A(n14816), .ZN(n14277) );
  AND2_X1 U11643 ( .A1(n14409), .A2(n14318), .ZN(n14413) );
  NAND2_X1 U11644 ( .A1(n13011), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10156) );
  NAND2_X1 U11645 ( .A1(n13020), .A2(n9748), .ZN(n9960) );
  OR2_X2 U11646 ( .A1(n12690), .A2(n12689), .ZN(n12814) );
  NAND2_X1 U11647 ( .A1(n11778), .A2(n11744), .ZN(n11771) );
  INV_X1 U11648 ( .A(n13490), .ZN(n14515) );
  INV_X1 U11649 ( .A(n15772), .ZN(n11424) );
  NAND2_X1 U11650 ( .A1(n11398), .A2(n19513), .ZN(n11534) );
  INV_X1 U11651 ( .A(n13777), .ZN(n11286) );
  NAND2_X1 U11652 ( .A1(n9783), .A2(n10930), .ZN(n11593) );
  NAND2_X1 U11653 ( .A1(n10083), .A2(n10082), .ZN(n9937) );
  INV_X1 U11654 ( .A(n10930), .ZN(n10082) );
  NAND2_X1 U11655 ( .A1(n16226), .A2(n9953), .ZN(n9952) );
  NAND2_X1 U11656 ( .A1(n9954), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9953) );
  INV_X1 U11657 ( .A(n16225), .ZN(n9954) );
  INV_X1 U11658 ( .A(n13731), .ZN(n10576) );
  INV_X1 U11659 ( .A(n13058), .ZN(n10524) );
  NAND2_X1 U11660 ( .A1(n10811), .A2(n10810), .ZN(n10814) );
  NAND2_X1 U11661 ( .A1(n9946), .A2(n10818), .ZN(n9949) );
  INV_X2 U11662 ( .A(n11534), .ZN(n11545) );
  INV_X1 U11663 ( .A(n10782), .ZN(n10027) );
  NAND2_X1 U11664 ( .A1(n10025), .A2(n10024), .ZN(n10023) );
  NAND2_X1 U11665 ( .A1(n10786), .A2(n10785), .ZN(n10024) );
  NOR2_X1 U11666 ( .A1(n17790), .A2(n12108), .ZN(n12109) );
  NAND2_X1 U11667 ( .A1(n10004), .A2(n10003), .ZN(n10550) );
  INV_X1 U11668 ( .A(n12115), .ZN(n10003) );
  OAI21_X1 U11669 ( .B1(n18207), .B2(n18206), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11959) );
  XNOR2_X1 U11670 ( .A(n17786), .B(n12109), .ZN(n12110) );
  NOR2_X1 U11671 ( .A1(n18234), .A2(n10560), .ZN(n10556) );
  AND2_X1 U11672 ( .A1(n10548), .A2(n9785), .ZN(n12106) );
  AND2_X1 U11673 ( .A1(n10452), .A2(n14318), .ZN(n14570) );
  AND2_X1 U11674 ( .A1(n15034), .A2(n10409), .ZN(n10408) );
  NOR2_X1 U11675 ( .A1(n15210), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10409) );
  NAND2_X1 U11676 ( .A1(n15034), .A2(n15043), .ZN(n15033) );
  AND2_X1 U11677 ( .A1(n14631), .A2(n14617), .ZN(n14602) );
  NAND2_X1 U11678 ( .A1(n13547), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n9968) );
  NAND2_X1 U11679 ( .A1(n13544), .A2(n10051), .ZN(n13547) );
  NAND2_X1 U11680 ( .A1(n10052), .A2(n10159), .ZN(n10051) );
  INV_X1 U11681 ( .A(n13400), .ZN(n10388) );
  NAND2_X1 U11682 ( .A1(n13833), .A2(n12806), .ZN(n12752) );
  NAND2_X1 U11683 ( .A1(n9764), .A2(n9881), .ZN(n10041) );
  NAND2_X1 U11684 ( .A1(n13097), .A2(n12946), .ZN(n10022) );
  NOR2_X1 U11685 ( .A1(n20568), .A2(n20490), .ZN(n20904) );
  AND2_X1 U11686 ( .A1(n20568), .A2(n20490), .ZN(n20871) );
  AND2_X1 U11687 ( .A1(n20568), .A2(n20567), .ZN(n20986) );
  AOI21_X1 U11688 ( .B1(n11202), .B2(n11201), .A(n11200), .ZN(n11238) );
  AOI22_X1 U11689 ( .A1(n13765), .A2(n13682), .B1(n12651), .B2(n12410), .ZN(
        n12846) );
  NAND2_X1 U11690 ( .A1(n11391), .A2(n11404), .ZN(n11740) );
  NOR3_X1 U11691 ( .A1(n11787), .A2(n11792), .A3(n16303), .ZN(n16030) );
  AOI21_X1 U11692 ( .B1(n11783), .B2(n9911), .A(n10599), .ZN(n10598) );
  OAI211_X1 U11693 ( .C1(n9797), .C2(n10187), .A(n10186), .B(n11770), .ZN(
        n11775) );
  INV_X1 U11694 ( .A(n11767), .ZN(n10187) );
  OAI21_X1 U11695 ( .B1(n11834), .B2(n10515), .A(n10513), .ZN(n16114) );
  NAND2_X1 U11696 ( .A1(n10516), .A2(n9745), .ZN(n10515) );
  AND2_X1 U11697 ( .A1(n10519), .A2(n10514), .ZN(n10513) );
  INV_X1 U11698 ( .A(n10520), .ZN(n10519) );
  INV_X1 U11699 ( .A(n10363), .ZN(n10362) );
  OAI21_X1 U11700 ( .B1(n9745), .B2(n9751), .A(n16122), .ZN(n10363) );
  NAND2_X1 U11701 ( .A1(n10362), .A2(n10359), .ZN(n10358) );
  NAND2_X1 U11702 ( .A1(n9751), .A2(n10361), .ZN(n10359) );
  NAND2_X1 U11703 ( .A1(n9731), .A2(n10341), .ZN(n16118) );
  INV_X1 U11704 ( .A(n11845), .ZN(n10341) );
  INV_X1 U11705 ( .A(n10140), .ZN(n10139) );
  OAI21_X1 U11706 ( .B1(n10141), .B2(n10510), .A(n16155), .ZN(n10140) );
  NAND2_X1 U11707 ( .A1(n11603), .A2(n9791), .ZN(n10191) );
  NOR2_X2 U11708 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20180) );
  OAI21_X1 U11709 ( .B1(n10332), .B2(n12088), .A(n9839), .ZN(n16777) );
  NAND2_X1 U11710 ( .A1(n16687), .A2(n10337), .ZN(n10332) );
  NAND2_X1 U11711 ( .A1(n17855), .A2(n19260), .ZN(n16689) );
  NAND2_X1 U11712 ( .A1(n16704), .A2(n10553), .ZN(n16706) );
  AND2_X1 U11713 ( .A1(n18307), .A2(n17921), .ZN(n10553) );
  AND2_X1 U11714 ( .A1(n12109), .A2(n12096), .ZN(n12112) );
  INV_X1 U11715 ( .A(n17783), .ZN(n12582) );
  NAND2_X1 U11716 ( .A1(n10237), .A2(n10236), .ZN(n18012) );
  XNOR2_X1 U11717 ( .A(n12110), .B(n10171), .ZN(n10558) );
  INV_X1 U11718 ( .A(n17002), .ZN(n19054) );
  OAI211_X1 U11719 ( .C1(n12067), .C2(n12066), .A(n12065), .B(n12064), .ZN(
        n19059) );
  OR2_X1 U11720 ( .A1(n12652), .A2(n13775), .ZN(n14549) );
  NAND2_X1 U11721 ( .A1(n16283), .A2(n20197), .ZN(n16287) );
  NAND2_X1 U11722 ( .A1(n10214), .A2(n9898), .ZN(n17642) );
  INV_X1 U11723 ( .A(n16775), .ZN(n10214) );
  NAND2_X1 U11724 ( .A1(n10020), .A2(n10018), .ZN(n10017) );
  NAND2_X1 U11725 ( .A1(n12879), .A2(n13323), .ZN(n10019) );
  AND2_X1 U11726 ( .A1(n11592), .A2(n10928), .ZN(n10269) );
  NAND2_X1 U11729 ( .A1(n12815), .A2(n12816), .ZN(n12976) );
  NOR2_X1 U11730 ( .A1(n12915), .A2(n10605), .ZN(n10604) );
  INV_X1 U11731 ( .A(n13341), .ZN(n10605) );
  NAND2_X1 U11732 ( .A1(n13012), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U11733 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10990) );
  INV_X1 U11734 ( .A(n10917), .ZN(n10918) );
  INV_X1 U11735 ( .A(n10921), .ZN(n10922) );
  INV_X1 U11736 ( .A(n10920), .ZN(n10923) );
  INV_X1 U11737 ( .A(n15745), .ZN(n10534) );
  NAND2_X1 U11738 ( .A1(n15775), .A2(n11813), .ZN(n10130) );
  NOR2_X1 U11739 ( .A1(n11068), .A2(n10127), .ZN(n10126) );
  INV_X1 U11740 ( .A(n15775), .ZN(n10127) );
  NOR2_X1 U11741 ( .A1(n13627), .A2(n11619), .ZN(n10505) );
  AOI21_X1 U11742 ( .B1(n10803), .B2(P2_EBX_REG_1__SCAN_IN), .A(n10771), .ZN(
        n10772) );
  NAND2_X1 U11743 ( .A1(n10030), .A2(n10790), .ZN(n10796) );
  NAND2_X1 U11744 ( .A1(n10442), .A2(n10031), .ZN(n10030) );
  NOR2_X1 U11745 ( .A1(n10789), .A2(n11619), .ZN(n10031) );
  INV_X1 U11746 ( .A(n19529), .ZN(n11204) );
  NAND2_X1 U11747 ( .A1(n11204), .A2(n13069), .ZN(n10785) );
  AOI21_X1 U11748 ( .B1(n19523), .B2(n10783), .A(n10026), .ZN(n10025) );
  NAND2_X1 U11749 ( .A1(n11212), .A2(n19518), .ZN(n10026) );
  INV_X1 U11750 ( .A(n19518), .ZN(n11350) );
  INV_X1 U11751 ( .A(n10762), .ZN(n10766) );
  AOI22_X1 U11752 ( .A1(n12264), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U11753 ( .A1(n9810), .A2(n9939), .ZN(n9938) );
  INV_X1 U11754 ( .A(n19479), .ZN(n9939) );
  NAND2_X1 U11755 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19079), .ZN(
        n11864) );
  NAND2_X1 U11756 ( .A1(n17332), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11860) );
  NAND2_X1 U11757 ( .A1(n18117), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10240) );
  XOR2_X1 U11758 ( .A(n17793), .B(n12103), .Z(n12105) );
  AOI21_X1 U11759 ( .B1(n19067), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12049), .ZN(n12055) );
  NOR2_X1 U11760 ( .A1(n12061), .A2(n12056), .ZN(n12049) );
  NAND2_X1 U11761 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19066), .ZN(
        n12056) );
  NAND2_X1 U11762 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10253) );
  NAND2_X1 U11763 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10254) );
  NAND2_X1 U11764 ( .A1(n17596), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10322) );
  NAND2_X1 U11765 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10321) );
  INV_X1 U11766 ( .A(n13528), .ZN(n10628) );
  NAND2_X1 U11767 ( .A1(n10403), .A2(n10154), .ZN(n13895) );
  AND2_X1 U11768 ( .A1(n10404), .A2(n13528), .ZN(n10154) );
  NOR2_X1 U11769 ( .A1(n10618), .A2(n10616), .ZN(n10615) );
  INV_X1 U11770 ( .A(n14246), .ZN(n10618) );
  NAND2_X1 U11771 ( .A1(n10617), .A2(n14204), .ZN(n10616) );
  INV_X1 U11772 ( .A(n14598), .ZN(n10617) );
  INV_X1 U11773 ( .A(n14616), .ZN(n14204) );
  AND2_X1 U11774 ( .A1(n10620), .A2(n14643), .ZN(n10619) );
  NOR2_X1 U11775 ( .A1(n14654), .A2(n10621), .ZN(n10620) );
  INV_X1 U11776 ( .A(n10622), .ZN(n10621) );
  AND2_X1 U11777 ( .A1(n9901), .A2(n10611), .ZN(n10609) );
  AND2_X1 U11778 ( .A1(n14739), .A2(n10612), .ZN(n10611) );
  INV_X1 U11779 ( .A(n14751), .ZN(n10612) );
  INV_X1 U11780 ( .A(n14468), .ZN(n14502) );
  AND2_X1 U11781 ( .A1(n13891), .A2(n9988), .ZN(n9987) );
  AND2_X1 U11782 ( .A1(n13890), .A2(n14915), .ZN(n9988) );
  AOI21_X1 U11783 ( .B1(n9763), .B2(n14400), .A(n9914), .ZN(n10629) );
  NAND2_X1 U11784 ( .A1(n15150), .A2(n15146), .ZN(n15127) );
  NOR2_X1 U11785 ( .A1(n10447), .A2(n14282), .ZN(n10446) );
  INV_X1 U11786 ( .A(n14276), .ZN(n10447) );
  AND2_X1 U11787 ( .A1(n15208), .A2(n14393), .ZN(n14394) );
  OR2_X1 U11788 ( .A1(n14392), .A2(n15422), .ZN(n14393) );
  INV_X1 U11789 ( .A(n16793), .ZN(n10377) );
  AND2_X1 U11790 ( .A1(n16813), .A2(n14929), .ZN(n10459) );
  AND2_X1 U11791 ( .A1(n13528), .A2(n13893), .ZN(n10625) );
  NAND2_X1 U11792 ( .A1(n9965), .A2(n9964), .ZN(n9972) );
  AOI21_X1 U11793 ( .B1(n9746), .B2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U11794 ( .A1(n15462), .A2(n9877), .ZN(n9965) );
  INV_X1 U11795 ( .A(n13427), .ZN(n14319) );
  NAND2_X1 U11796 ( .A1(n13078), .A2(n13077), .ZN(n13426) );
  INV_X1 U11797 ( .A(n13208), .ZN(n13021) );
  INV_X1 U11798 ( .A(n14357), .ZN(n9959) );
  INV_X1 U11799 ( .A(n13011), .ZN(n9961) );
  NAND2_X1 U11800 ( .A1(n12929), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10042) );
  INV_X1 U11801 ( .A(n10018), .ZN(n10039) );
  INV_X1 U11802 ( .A(n20489), .ZN(n20749) );
  INV_X1 U11803 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20905) );
  NAND4_X1 U11804 ( .A1(n10766), .A2(n19529), .A3(n19518), .A4(n13069), .ZN(
        n10779) );
  AND2_X1 U11805 ( .A1(n11119), .A2(n11115), .ZN(n10540) );
  OR2_X1 U11806 ( .A1(n11071), .A2(n10100), .ZN(n11124) );
  NAND2_X1 U11807 ( .A1(n10101), .A2(n11092), .ZN(n10100) );
  INV_X1 U11808 ( .A(n10102), .ZN(n10101) );
  NOR2_X1 U11809 ( .A1(n11042), .A2(n11055), .ZN(n11045) );
  NOR2_X1 U11810 ( .A1(n12335), .A2(n10592), .ZN(n10591) );
  INV_X1 U11811 ( .A(n15870), .ZN(n10592) );
  OR2_X1 U11812 ( .A1(n10765), .A2(n12146), .ZN(n10767) );
  OR2_X1 U11813 ( .A1(n10969), .A2(n10968), .ZN(n11430) );
  NAND2_X1 U11814 ( .A1(n10105), .A2(n11599), .ZN(n11605) );
  NAND2_X1 U11815 ( .A1(n10547), .A2(n15532), .ZN(n10546) );
  INV_X1 U11816 ( .A(n14525), .ZN(n10547) );
  NAND2_X1 U11817 ( .A1(n10568), .A2(n15511), .ZN(n10567) );
  INV_X1 U11818 ( .A(n15496), .ZN(n10568) );
  INV_X1 U11819 ( .A(n16047), .ZN(n11783) );
  INV_X1 U11820 ( .A(n10355), .ZN(n10352) );
  AOI21_X1 U11821 ( .B1(n11179), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16086), .ZN(n10355) );
  NOR2_X1 U11822 ( .A1(n11179), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10354) );
  OR2_X1 U11823 ( .A1(n16712), .A2(n11792), .ZN(n11172) );
  AND2_X1 U11824 ( .A1(n9846), .A2(n16214), .ZN(n10444) );
  NAND2_X1 U11825 ( .A1(n10528), .A2(n10527), .ZN(n10526) );
  INV_X1 U11826 ( .A(n16002), .ZN(n10527) );
  OR2_X1 U11827 ( .A1(n19317), .A2(n11792), .ZN(n11151) );
  NAND2_X1 U11828 ( .A1(n10139), .A2(n10141), .ZN(n10136) );
  AND2_X1 U11829 ( .A1(n13760), .A2(n9854), .ZN(n13797) );
  INV_X1 U11830 ( .A(n13798), .ZN(n10562) );
  INV_X1 U11831 ( .A(n12450), .ZN(n9986) );
  AND2_X1 U11832 ( .A1(n11286), .A2(n11290), .ZN(n10563) );
  NAND2_X1 U11833 ( .A1(n10129), .A2(n10128), .ZN(n10131) );
  AND2_X1 U11834 ( .A1(n19357), .A2(n11267), .ZN(n10128) );
  NAND2_X1 U11835 ( .A1(n16247), .A2(n16244), .ZN(n11603) );
  NAND2_X1 U11836 ( .A1(n11597), .A2(n16268), .ZN(n11601) );
  INV_X1 U11837 ( .A(n13603), .ZN(n10577) );
  INV_X1 U11838 ( .A(n15749), .ZN(n10133) );
  NAND2_X1 U11839 ( .A1(n10796), .A2(n10797), .ZN(n10816) );
  NAND2_X1 U11840 ( .A1(n10798), .A2(n10433), .ZN(n10815) );
  INV_X1 U11841 ( .A(n10796), .ZN(n10433) );
  INV_X1 U11842 ( .A(n10797), .ZN(n10798) );
  OR2_X1 U11843 ( .A1(n10881), .A2(n10880), .ZN(n11581) );
  OR2_X1 U11844 ( .A1(n10879), .A2(n10878), .ZN(n10880) );
  AND2_X1 U11845 ( .A1(n13069), .A2(n19977), .ZN(n11404) );
  NAND2_X1 U11846 ( .A1(n10149), .A2(n11212), .ZN(n11213) );
  AOI22_X1 U11847 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10757) );
  AND2_X1 U11848 ( .A1(n19529), .A2(n10762), .ZN(n9992) );
  INV_X1 U11849 ( .A(n11212), .ZN(n9993) );
  AND2_X1 U11850 ( .A1(n19479), .A2(n12153), .ZN(n10831) );
  NOR2_X1 U11851 ( .A1(n10829), .A2(n19479), .ZN(n10365) );
  NAND2_X1 U11852 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10289) );
  AOI21_X1 U11853 ( .B1(n12264), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n10296), .ZN(n10295) );
  NAND2_X1 U11854 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U11855 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10298) );
  NAND2_X1 U11856 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10294) );
  AOI21_X1 U11857 ( .B1(n12264), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n10291), .ZN(n10290) );
  NAND2_X1 U11858 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10292) );
  NAND2_X1 U11859 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10293) );
  INV_X1 U11860 ( .A(n10689), .ZN(n10694) );
  INV_X1 U11861 ( .A(n12169), .ZN(n12141) );
  NOR2_X1 U11862 ( .A1(n11863), .A2(n11854), .ZN(n11970) );
  NAND2_X1 U11863 ( .A1(n19226), .A2(n19079), .ZN(n11862) );
  NAND2_X1 U11864 ( .A1(n10383), .A2(n9818), .ZN(n10384) );
  NOR2_X1 U11865 ( .A1(n17361), .A2(n11861), .ZN(n11903) );
  AOI22_X1 U11866 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10078) );
  AND2_X1 U11867 ( .A1(n10503), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10502) );
  NOR2_X1 U11868 ( .A1(n16704), .A2(n10638), .ZN(n16847) );
  NAND2_X1 U11869 ( .A1(n17982), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10179) );
  INV_X1 U11870 ( .A(n16693), .ZN(n10336) );
  OAI21_X1 U11871 ( .B1(n18629), .B2(n12043), .A(n12074), .ZN(n12089) );
  NAND2_X1 U11872 ( .A1(n18632), .A2(n18629), .ZN(n10064) );
  NAND2_X1 U11873 ( .A1(n10315), .A2(n12045), .ZN(n16690) );
  NAND2_X1 U11874 ( .A1(n17815), .A2(n18636), .ZN(n10316) );
  NOR2_X1 U11875 ( .A1(n12862), .A2(n12797), .ZN(n10008) );
  AND2_X1 U11876 ( .A1(n13327), .A2(n13340), .ZN(n13339) );
  NAND2_X1 U11877 ( .A1(n14184), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14206) );
  AND2_X2 U11878 ( .A1(n14040), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14041) );
  INV_X1 U11879 ( .A(n14039), .ZN(n14040) );
  OR2_X1 U11880 ( .A1(n15112), .A2(n14468), .ZN(n14060) );
  NAND2_X1 U11881 ( .A1(n13949), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13962) );
  INV_X1 U11882 ( .A(n13948), .ZN(n13949) );
  NAND2_X1 U11883 ( .A1(n13577), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13611) );
  AND2_X1 U11884 ( .A1(n10646), .A2(n14422), .ZN(n10406) );
  NAND2_X1 U11885 ( .A1(n14603), .A2(n14322), .ZN(n14587) );
  AND2_X1 U11886 ( .A1(n10450), .A2(n14601), .ZN(n10449) );
  AND2_X1 U11887 ( .A1(n10451), .A2(n14322), .ZN(n10450) );
  INV_X1 U11888 ( .A(n14588), .ZN(n10451) );
  NAND2_X1 U11889 ( .A1(n10429), .A2(n10164), .ZN(n10163) );
  NAND2_X1 U11890 ( .A1(n10429), .A2(n15210), .ZN(n10162) );
  NAND2_X1 U11891 ( .A1(n15026), .A2(n9918), .ZN(n10375) );
  NAND3_X1 U11892 ( .A1(n10626), .A2(n10045), .A3(n10043), .ZN(n15034) );
  NAND2_X1 U11893 ( .A1(n10044), .A2(n15259), .ZN(n10043) );
  INV_X1 U11894 ( .A(n14404), .ZN(n10044) );
  NAND2_X1 U11895 ( .A1(n10160), .A2(n15189), .ZN(n15043) );
  AND2_X1 U11896 ( .A1(n14695), .A2(n9889), .ZN(n14631) );
  INV_X1 U11897 ( .A(n14632), .ZN(n10453) );
  NAND2_X1 U11898 ( .A1(n14695), .A2(n9871), .ZN(n14649) );
  NAND2_X1 U11899 ( .A1(n14695), .A2(n9869), .ZN(n14656) );
  NAND2_X1 U11900 ( .A1(n14695), .A2(n14302), .ZN(n14675) );
  NAND2_X1 U11901 ( .A1(n10400), .A2(n10629), .ZN(n10372) );
  NAND2_X1 U11902 ( .A1(n14397), .A2(n10630), .ZN(n10400) );
  OAI21_X1 U11903 ( .B1(n9830), .B2(n15189), .A(n10419), .ZN(n15099) );
  NAND2_X1 U11904 ( .A1(n15089), .A2(n15189), .ZN(n10419) );
  NOR2_X1 U11905 ( .A1(n14741), .A2(n14290), .ZN(n14733) );
  NAND2_X1 U11906 ( .A1(n10371), .A2(n10630), .ZN(n15087) );
  NAND2_X1 U11907 ( .A1(n9975), .A2(n13542), .ZN(n9974) );
  NAND2_X1 U11908 ( .A1(n13564), .A2(n10650), .ZN(n13590) );
  INV_X1 U11909 ( .A(n13589), .ZN(n13564) );
  NAND2_X1 U11910 ( .A1(n10117), .A2(n13397), .ZN(n13411) );
  NAND2_X1 U11911 ( .A1(n13017), .A2(n13016), .ZN(n13232) );
  AND2_X1 U11912 ( .A1(n13015), .A2(n13014), .ZN(n13016) );
  INV_X1 U11913 ( .A(n10427), .ZN(n10113) );
  INV_X1 U11914 ( .A(n14871), .ZN(n20988) );
  AOI21_X1 U11915 ( .B1(n20571), .B2(n20646), .A(n20705), .ZN(n20577) );
  NAND2_X1 U11916 ( .A1(n13463), .A2(n21091), .ZN(n10012) );
  NOR2_X1 U11917 ( .A1(n20653), .A2(n20647), .ZN(n20836) );
  AND4_X1 U11918 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        n12669) );
  NOR2_X1 U11919 ( .A1(n20654), .A2(n20653), .ZN(n20994) );
  AOI21_X1 U11920 ( .B1(n20953), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20653), 
        .ZN(n21035) );
  NAND2_X1 U11921 ( .A1(n10200), .A2(n10199), .ZN(n11742) );
  INV_X1 U11922 ( .A(n10779), .ZN(n10199) );
  NOR2_X1 U11923 ( .A1(n10201), .A2(n10149), .ZN(n10200) );
  INV_X1 U11924 ( .A(n13685), .ZN(n10201) );
  NAND2_X1 U11925 ( .A1(n10767), .A2(n11722), .ZN(n9944) );
  AND2_X1 U11926 ( .A1(n11367), .A2(n11366), .ZN(n13682) );
  NAND2_X1 U11927 ( .A1(n11039), .A2(n11038), .ZN(n11232) );
  NAND2_X1 U11928 ( .A1(n11586), .A2(n11751), .ZN(n11039) );
  NAND2_X1 U11929 ( .A1(n11747), .A2(n11746), .ZN(n11786) );
  INV_X1 U11930 ( .A(n11780), .ZN(n11747) );
  AND2_X1 U11931 ( .A1(n11180), .A2(n15552), .ZN(n10542) );
  OAI21_X1 U11932 ( .B1(n11111), .B2(n10095), .A(n9762), .ZN(n10097) );
  NAND2_X1 U11933 ( .A1(n11098), .A2(n10094), .ZN(n10093) );
  NAND2_X1 U11934 ( .A1(n11077), .A2(n11078), .ZN(n11074) );
  AND2_X1 U11935 ( .A1(n11423), .A2(n11422), .ZN(n15772) );
  NAND2_X1 U11937 ( .A1(n13491), .A2(n9875), .ZN(n13743) );
  AOI22_X1 U11938 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11246), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11445) );
  INV_X1 U11939 ( .A(n16650), .ZN(n13066) );
  INV_X1 U11940 ( .A(n10783), .ZN(n12415) );
  INV_X1 U11941 ( .A(n13719), .ZN(n10525) );
  NOR2_X1 U11942 ( .A1(n13719), .A2(n10530), .ZN(n13620) );
  AND3_X1 U11943 ( .A1(n11506), .A2(n11505), .A3(n11504), .ZN(n13488) );
  NOR2_X1 U11944 ( .A1(n11397), .A2(n13069), .ZN(n10270) );
  AND3_X1 U11945 ( .A1(n11428), .A2(n11427), .A3(n11426), .ZN(n15757) );
  INV_X1 U11946 ( .A(n16295), .ZN(n10580) );
  NOR2_X1 U11947 ( .A1(n10793), .A2(n10195), .ZN(n10198) );
  NAND2_X1 U11948 ( .A1(n10036), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10029) );
  NAND2_X1 U11949 ( .A1(n10272), .A2(n13632), .ZN(n10055) );
  NOR2_X2 U11950 ( .A1(n15490), .A2(n15491), .ZN(n15489) );
  NAND2_X1 U11951 ( .A1(n14530), .A2(n15511), .ZN(n15495) );
  NAND2_X1 U11952 ( .A1(n16048), .A2(n10440), .ZN(n10439) );
  NOR2_X1 U11953 ( .A1(n11696), .A2(n10570), .ZN(n10569) );
  INV_X1 U11954 ( .A(n10571), .ZN(n10570) );
  OR2_X1 U11955 ( .A1(n15556), .A2(n11184), .ZN(n16064) );
  INV_X1 U11956 ( .A(n10344), .ZN(n10342) );
  AND2_X1 U11957 ( .A1(n16106), .A2(n11766), .ZN(n16095) );
  NAND2_X1 U11958 ( .A1(n16102), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16100) );
  NOR2_X1 U11959 ( .A1(n9768), .A2(n15592), .ZN(n10511) );
  OR3_X1 U11960 ( .A1(n15645), .A2(n11792), .A3(n16461), .ZN(n16145) );
  INV_X1 U11961 ( .A(n10508), .ZN(n10141) );
  NAND2_X1 U11962 ( .A1(n9986), .A2(n10585), .ZN(n16150) );
  AND2_X1 U11963 ( .A1(n10672), .A2(n16171), .ZN(n10510) );
  NAND2_X1 U11964 ( .A1(n10509), .A2(n16171), .ZN(n10508) );
  INV_X1 U11965 ( .A(n11833), .ZN(n10509) );
  NAND2_X1 U11966 ( .A1(n9986), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16165) );
  AND3_X1 U11967 ( .A1(n11467), .A2(n11466), .A3(n11465), .ZN(n13275) );
  NAND2_X1 U11968 ( .A1(n16213), .A2(n16214), .ZN(n16166) );
  AND3_X1 U11969 ( .A1(n11454), .A2(n11453), .A3(n11452), .ZN(n13058) );
  AND2_X1 U11970 ( .A1(n19807), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19748) );
  NAND2_X1 U11971 ( .A1(n11828), .A2(n11619), .ZN(n11621) );
  NAND2_X1 U11972 ( .A1(n11207), .A2(n19411), .ZN(n11208) );
  AND2_X1 U11973 ( .A1(n19807), .A2(n19501), .ZN(n19715) );
  NAND2_X1 U11974 ( .A1(n19807), .A2(n20211), .ZN(n19742) );
  INV_X1 U11975 ( .A(n20178), .ZN(n19882) );
  NOR3_X1 U11976 ( .A1(n19915), .A2(n19937), .A3(n20207), .ZN(n19917) );
  INV_X1 U11977 ( .A(n19949), .ZN(n19912) );
  OR2_X1 U11978 ( .A1(n20190), .A2(n20199), .ZN(n19949) );
  OR2_X1 U11979 ( .A1(n19807), .A2(n19501), .ZN(n19944) );
  NAND2_X1 U11980 ( .A1(n20184), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20029) );
  INV_X1 U11981 ( .A(n17968), .ZN(n10463) );
  INV_X1 U11982 ( .A(n17381), .ZN(n10216) );
  INV_X1 U11983 ( .A(n17782), .ZN(n10257) );
  OR2_X1 U11984 ( .A1(n12592), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10477) );
  NOR2_X1 U11985 ( .A1(n10476), .A2(n10482), .ZN(n10475) );
  INV_X1 U11986 ( .A(n16859), .ZN(n16866) );
  OAI21_X1 U11987 ( .B1(n16866), .B2(n18593), .A(n10387), .ZN(n16702) );
  AOI21_X1 U11988 ( .B1(n16865), .B2(n18318), .A(n18588), .ZN(n10387) );
  NAND2_X1 U11989 ( .A1(n18016), .A2(n18321), .ZN(n17969) );
  NAND2_X1 U11990 ( .A1(n17989), .A2(n10561), .ZN(n17975) );
  AND2_X1 U11991 ( .A1(n12125), .A2(n18296), .ZN(n10561) );
  NAND2_X1 U11992 ( .A1(n18090), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12123) );
  INV_X1 U11993 ( .A(n11959), .ZN(n11957) );
  AND2_X1 U11994 ( .A1(n18480), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18436) );
  NAND2_X1 U11995 ( .A1(n10555), .A2(n10168), .ZN(n18219) );
  NAND2_X1 U11996 ( .A1(n10558), .A2(n10556), .ZN(n10555) );
  NOR2_X1 U11997 ( .A1(n10170), .A2(n10557), .ZN(n10169) );
  INV_X1 U11998 ( .A(n10556), .ZN(n10554) );
  NAND2_X1 U11999 ( .A1(n18243), .A2(n12107), .ZN(n18232) );
  INV_X1 U12000 ( .A(n12100), .ZN(n10224) );
  XNOR2_X1 U12001 ( .A(n12099), .B(n18580), .ZN(n18266) );
  NOR2_X1 U12002 ( .A1(n18266), .A2(n18267), .ZN(n18265) );
  INV_X1 U12003 ( .A(n11965), .ZN(n10249) );
  NAND2_X1 U12004 ( .A1(n10251), .A2(n11969), .ZN(n10250) );
  INV_X1 U12005 ( .A(n17815), .ZN(n18617) );
  OR2_X1 U12006 ( .A1(n13202), .A2(n13201), .ZN(n13204) );
  INV_X1 U12007 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20953) );
  XNOR2_X1 U12008 ( .A(n13229), .B(n13232), .ZN(n20567) );
  NAND2_X1 U12009 ( .A1(n12948), .A2(n12947), .ZN(n12949) );
  AND2_X1 U12010 ( .A1(n20568), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20748) );
  XNOR2_X1 U12011 ( .A(n11786), .B(n11785), .ZN(n15501) );
  OR2_X1 U12012 ( .A1(n14549), .A2(n11752), .ZN(n19356) );
  NOR2_X2 U12013 ( .A1(n11664), .A2(n19364), .ZN(n19320) );
  OR2_X1 U12014 ( .A1(n11796), .A2(n10564), .ZN(n14544) );
  AND2_X1 U12015 ( .A1(n15498), .A2(n11795), .ZN(n10564) );
  INV_X1 U12016 ( .A(n19408), .ZN(n13177) );
  XNOR2_X1 U12017 ( .A(n11820), .B(n11819), .ZN(n12576) );
  NAND2_X1 U12018 ( .A1(n16032), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U12019 ( .A1(n16183), .A2(n10366), .ZN(n16039) );
  OR2_X1 U12020 ( .A1(n15578), .A2(n15577), .ZN(n16372) );
  AOI21_X1 U12021 ( .B1(n16411), .B2(n19493), .A(n12458), .ZN(n12459) );
  INV_X1 U12022 ( .A(n19487), .ZN(n19476) );
  CLKBUF_X1 U12023 ( .A(n12153), .Z(n19494) );
  INV_X1 U12024 ( .A(n16287), .ZN(n19493) );
  NAND2_X1 U12025 ( .A1(n12653), .A2(n11822), .ZN(n16283) );
  AND2_X1 U12026 ( .A1(n11821), .A2(n13063), .ZN(n19484) );
  NAND2_X1 U12027 ( .A1(n10088), .A2(n10281), .ZN(n10087) );
  XNOR2_X1 U12028 ( .A(n11794), .B(n11793), .ZN(n12597) );
  NOR2_X1 U12029 ( .A1(n11812), .A2(n16030), .ZN(n11794) );
  NAND2_X1 U12030 ( .A1(n10436), .A2(n16054), .ZN(n10435) );
  INV_X1 U12031 ( .A(n10437), .ZN(n10436) );
  OR2_X1 U12032 ( .A1(n16338), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10146) );
  NAND2_X1 U12033 ( .A1(n16100), .A2(n10267), .ZN(n16379) );
  NAND2_X1 U12034 ( .A1(n10268), .A2(n16371), .ZN(n10267) );
  OAI21_X1 U12035 ( .B1(n16114), .B2(n11839), .A(n16112), .ZN(n11843) );
  NAND2_X1 U12036 ( .A1(n10340), .A2(n9822), .ZN(n12439) );
  NAND2_X1 U12037 ( .A1(n16118), .A2(n11371), .ZN(n10340) );
  NAND2_X1 U12038 ( .A1(n16394), .A2(n11371), .ZN(n10339) );
  OAI211_X1 U12039 ( .C1(n10523), .C2(n9843), .A(n10360), .B(n10357), .ZN(
        n16416) );
  OAI21_X1 U12040 ( .B1(n10362), .B2(n9792), .A(n10358), .ZN(n10357) );
  NAND2_X1 U12041 ( .A1(n9943), .A2(n16118), .ZN(n16415) );
  NAND2_X1 U12042 ( .A1(n9935), .A2(n16409), .ZN(n9943) );
  AND2_X1 U12043 ( .A1(n16496), .A2(n11381), .ZN(n16462) );
  INV_X1 U12044 ( .A(n16838), .ZN(n16590) );
  INV_X1 U12045 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12154) );
  INV_X1 U12046 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20205) );
  INV_X1 U12047 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20196) );
  NAND2_X1 U12048 ( .A1(n13765), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16771) );
  NAND2_X1 U12049 ( .A1(n19258), .A2(n19054), .ZN(n17853) );
  INV_X1 U12050 ( .A(n17373), .ZN(n17372) );
  NAND2_X1 U12051 ( .A1(n17410), .A2(n9899), .ZN(n13817) );
  NAND2_X1 U12052 ( .A1(n17412), .A2(n9735), .ZN(n17410) );
  NOR2_X1 U12053 ( .A1(n17440), .A2(n17124), .ZN(n17452) );
  AOI21_X1 U12054 ( .B1(n12478), .B2(n12477), .A(n16695), .ZN(n16775) );
  INV_X1 U12055 ( .A(n17673), .ZN(n17666) );
  NAND2_X1 U12056 ( .A1(n17666), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17668) );
  INV_X1 U12057 ( .A(n17743), .ZN(n17732) );
  NOR2_X1 U12058 ( .A1(n18645), .A2(n17805), .ZN(n17774) );
  NOR2_X1 U12059 ( .A1(n11881), .A2(n11880), .ZN(n17790) );
  INV_X1 U12060 ( .A(n17774), .ZN(n17806) );
  NAND2_X1 U12061 ( .A1(n12128), .A2(n18302), .ZN(n16896) );
  NAND2_X1 U12062 ( .A1(n17156), .A2(n10503), .ZN(n17994) );
  OR2_X1 U12063 ( .A1(n18058), .A2(n18374), .ZN(n9932) );
  AOI21_X1 U12064 ( .B1(n18200), .B2(n18367), .A(n9931), .ZN(n9930) );
  NOR2_X1 U12065 ( .A1(n18140), .A2(n18034), .ZN(n9931) );
  OR2_X1 U12066 ( .A1(n18092), .A2(n9928), .ZN(n9927) );
  AND2_X1 U12067 ( .A1(n18039), .A2(n18354), .ZN(n9928) );
  NAND2_X1 U12068 ( .A1(n18068), .A2(n18366), .ZN(n18058) );
  AND2_X1 U12069 ( .A1(n16901), .A2(n9773), .ZN(n18429) );
  NAND2_X1 U12070 ( .A1(n16701), .A2(n16884), .ZN(n12138) );
  INV_X1 U12071 ( .A(n16702), .ZN(n16701) );
  XNOR2_X1 U12072 ( .A(n10227), .B(n16878), .ZN(n10006) );
  AOI21_X1 U12073 ( .B1(n16897), .B2(n16706), .A(n16705), .ZN(n10227) );
  OAI21_X1 U12074 ( .B1(n16708), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n10230), .ZN(n10229) );
  NAND2_X1 U12075 ( .A1(n9732), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n10230) );
  AOI211_X1 U12076 ( .C1(n12094), .C2(n19056), .A(n12076), .B(n16693), .ZN(
        n12082) );
  AND2_X1 U12077 ( .A1(n19252), .A2(n19099), .ZN(n10331) );
  OR2_X1 U12078 ( .A1(n19209), .A2(n19112), .ZN(n10328) );
  NOR2_X1 U12079 ( .A1(n19109), .A2(n10329), .ZN(n19209) );
  NAND2_X1 U12080 ( .A1(n10330), .A2(n19258), .ZN(n10329) );
  NAND2_X1 U12081 ( .A1(n19103), .A2(n19104), .ZN(n10330) );
  AND2_X1 U12082 ( .A1(n12714), .A2(n12713), .ZN(n12721) );
  INV_X1 U12083 ( .A(n12896), .ZN(n10415) );
  AOI21_X1 U12084 ( .B1(n12707), .B2(n12732), .A(n12800), .ZN(n12735) );
  NAND2_X1 U12085 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12267) );
  NAND2_X1 U12086 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12275) );
  NAND4_X1 U12087 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(
        n10929) );
  AND4_X1 U12088 ( .A1(n10976), .A2(n10975), .A3(n10974), .A4(n10973), .ZN(
        n10986) );
  AND2_X1 U12089 ( .A1(n13698), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10035) );
  AOI22_X1 U12090 ( .A1(n10802), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10770) );
  AND2_X1 U12091 ( .A1(n10794), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10188) );
  INV_X1 U12092 ( .A(n12256), .ZN(n11012) );
  OAI21_X1 U12093 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19226), .A(
        n12050), .ZN(n12051) );
  OR2_X1 U12094 ( .A1(n12054), .A2(n12055), .ZN(n12050) );
  AND2_X1 U12095 ( .A1(n10630), .A2(n15210), .ZN(n10114) );
  INV_X1 U12096 ( .A(n14398), .ZN(n10632) );
  NAND2_X1 U12097 ( .A1(n13832), .A2(n13831), .ZN(n13893) );
  INV_X1 U12098 ( .A(n13229), .ZN(n13235) );
  OR2_X1 U12099 ( .A1(n13000), .A2(n12999), .ZN(n14380) );
  AND2_X1 U12100 ( .A1(n12816), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U12101 ( .A1(n10019), .A2(n10017), .ZN(n12884) );
  NOR2_X1 U12102 ( .A1(n10011), .A2(n9790), .ZN(n10009) );
  NAND2_X1 U12103 ( .A1(n13333), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U12104 ( .A1(n13830), .A2(n14376), .ZN(n12730) );
  AOI22_X1 U12105 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12994), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U12106 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12755) );
  INV_X1 U12107 ( .A(n12759), .ZN(n10050) );
  OR2_X1 U12108 ( .A1(n13473), .A2(n13472), .ZN(n13537) );
  AOI22_X1 U12109 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U12110 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12780), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U12111 ( .A1(n12775), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12994), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U12112 ( .A1(n11029), .A2(n11034), .ZN(n11044) );
  AND2_X1 U12113 ( .A1(n9842), .A2(n15877), .ZN(n10537) );
  INV_X1 U12114 ( .A(n11144), .ZN(n10538) );
  AOI22_X1 U12115 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12401), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U12116 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12401), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U12117 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12401), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U12118 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12354) );
  NAND2_X1 U12119 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12326) );
  NAND2_X1 U12120 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12319) );
  AOI22_X1 U12121 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12401), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U12122 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12401), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U12123 ( .A1(n10089), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10882), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U12124 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__5__SCAN_IN), .B2(n10884), .ZN(n10963) );
  AOI21_X1 U12125 ( .B1(n10935), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n10090), .ZN(n10941) );
  AND2_X1 U12126 ( .A1(n10872), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10090) );
  INV_X1 U12127 ( .A(n11720), .ZN(n10803) );
  AND4_X1 U12128 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11022) );
  INV_X1 U12129 ( .A(n10785), .ZN(n11215) );
  INV_X1 U12130 ( .A(n13069), .ZN(n9991) );
  NAND2_X1 U12131 ( .A1(n20205), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11026) );
  OR2_X1 U12132 ( .A1(n11189), .A2(n11185), .ZN(n11186) );
  NOR2_X1 U12133 ( .A1(n10479), .A2(n10483), .ZN(n10478) );
  INV_X1 U12134 ( .A(n10480), .ZN(n10479) );
  NOR2_X1 U12135 ( .A1(n18285), .A2(n10481), .ZN(n10480) );
  NOR2_X1 U12136 ( .A1(n12038), .A2(n18645), .ZN(n12039) );
  NOR2_X1 U12137 ( .A1(n14666), .A2(n10623), .ZN(n10622) );
  INV_X1 U12138 ( .A(n14682), .ZN(n10623) );
  INV_X1 U12139 ( .A(n14750), .ZN(n10610) );
  NOR2_X1 U12140 ( .A1(n13885), .A2(n13868), .ZN(n13869) );
  NAND2_X1 U12141 ( .A1(n15189), .A2(n10430), .ZN(n10429) );
  INV_X1 U12142 ( .A(n14405), .ZN(n10430) );
  INV_X1 U12143 ( .A(n14658), .ZN(n10455) );
  INV_X1 U12144 ( .A(n14402), .ZN(n10431) );
  NAND2_X1 U12145 ( .A1(n14392), .A2(n14359), .ZN(n15171) );
  INV_X1 U12146 ( .A(n14844), .ZN(n10458) );
  AND2_X1 U12147 ( .A1(n16792), .A2(n14374), .ZN(n10379) );
  NAND2_X1 U12148 ( .A1(n10410), .A2(n13533), .ZN(n14362) );
  NOR2_X1 U12149 ( .A1(n13380), .A2(n13379), .ZN(n13529) );
  AND2_X1 U12150 ( .A1(n10606), .A2(n10037), .ZN(n13341) );
  OR2_X1 U12151 ( .A1(n13010), .A2(n13009), .ZN(n13402) );
  AND2_X1 U12152 ( .A1(n13333), .A2(n14380), .ZN(n13012) );
  OR2_X1 U12153 ( .A1(n13089), .A2(n13088), .ZN(n13401) );
  AOI21_X1 U12154 ( .B1(n10020), .B2(n14318), .A(n12913), .ZN(n12890) );
  INV_X1 U12155 ( .A(n12730), .ZN(n12749) );
  OR2_X1 U12156 ( .A1(n12745), .A2(n12744), .ZN(n12748) );
  AOI22_X1 U12157 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U12158 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U12159 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U12160 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U12161 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12792) );
  OR2_X1 U12162 ( .A1(n11786), .A2(n11748), .ZN(n11791) );
  OAI21_X1 U12163 ( .B1(n19310), .B2(n15742), .A(n16715), .ZN(n15580) );
  NAND2_X1 U12164 ( .A1(n11111), .A2(n11744), .ZN(n11108) );
  NOR2_X1 U12165 ( .A1(n11124), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U12166 ( .A1(n10536), .A2(n10103), .ZN(n10102) );
  INV_X1 U12167 ( .A(n11070), .ZN(n10103) );
  INV_X1 U12168 ( .A(n11075), .ZN(n11073) );
  MUX2_X1 U12169 ( .A(n13734), .B(n11813), .S(n11789), .Z(n11078) );
  NOR2_X1 U12170 ( .A1(n10996), .A2(n10995), .ZN(n11434) );
  NOR2_X1 U12171 ( .A1(n10919), .A2(n10918), .ZN(n10926) );
  MUX2_X1 U12172 ( .A(n11032), .B(n11235), .S(n11789), .Z(n11046) );
  AOI21_X1 U12173 ( .B1(n10089), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n10092), .ZN(n11529) );
  AND2_X1 U12174 ( .A1(n10872), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10092) );
  CLKBUF_X1 U12175 ( .A(n10749), .Z(n12394) );
  CLKBUF_X1 U12176 ( .A(n10648), .Z(n12398) );
  CLKBUF_X1 U12177 ( .A(n12264), .Z(n12368) );
  AOI22_X1 U12178 ( .A1(n10089), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U12179 ( .A1(n10089), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__3__SCAN_IN), .B2(n10884), .ZN(n12214) );
  AOI22_X1 U12180 ( .A1(n10089), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12193) );
  NAND2_X1 U12181 ( .A1(n13801), .A2(n9882), .ZN(n15883) );
  AOI22_X1 U12182 ( .A1(n10089), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12183) );
  AND2_X1 U12183 ( .A1(n10594), .A2(n15900), .ZN(n10593) );
  NOR2_X1 U12184 ( .A1(n10530), .A2(n10529), .ZN(n10528) );
  INV_X1 U12185 ( .A(n13738), .ZN(n10529) );
  NAND2_X1 U12186 ( .A1(n10531), .A2(n13622), .ZN(n10530) );
  INV_X1 U12187 ( .A(n13718), .ZN(n10531) );
  NOR2_X1 U12188 ( .A1(n15541), .A2(n10490), .ZN(n10489) );
  INV_X1 U12189 ( .A(n11630), .ZN(n10498) );
  NOR2_X1 U12190 ( .A1(n10501), .A2(n10500), .ZN(n10499) );
  NAND2_X1 U12191 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10501) );
  NOR2_X1 U12192 ( .A1(n10895), .A2(n10894), .ZN(n11586) );
  NAND2_X1 U12193 ( .A1(n11574), .A2(n9827), .ZN(n10196) );
  NAND2_X1 U12194 ( .A1(n10787), .A2(n9821), .ZN(n10197) );
  NOR2_X1 U12195 ( .A1(n13067), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10272) );
  INV_X1 U12196 ( .A(n10794), .ZN(n10273) );
  INV_X1 U12197 ( .A(n16030), .ZN(n11809) );
  OR2_X1 U12198 ( .A1(n10279), .A2(n10278), .ZN(n10086) );
  AND2_X1 U12199 ( .A1(n10444), .A2(n11767), .ZN(n10185) );
  INV_X1 U12200 ( .A(n16045), .ZN(n10440) );
  NOR2_X1 U12201 ( .A1(n10441), .A2(n16315), .ZN(n10308) );
  AOI21_X1 U12202 ( .B1(n10302), .B2(n10304), .A(n10599), .ZN(n10300) );
  AND2_X1 U12203 ( .A1(n11343), .A2(n11344), .ZN(n11693) );
  OR2_X1 U12204 ( .A1(n11771), .A2(n11792), .ZN(n11784) );
  AND2_X1 U12205 ( .A1(n10572), .A2(n10573), .ZN(n10571) );
  INV_X1 U12206 ( .A(n11848), .ZN(n10572) );
  NOR2_X1 U12207 ( .A1(n10574), .A2(n15594), .ZN(n10573) );
  INV_X1 U12208 ( .A(n12455), .ZN(n10574) );
  INV_X1 U12209 ( .A(n11838), .ZN(n10516) );
  OAI21_X1 U12210 ( .B1(n11838), .B2(n10522), .A(n10521), .ZN(n10520) );
  AND2_X1 U12211 ( .A1(n12451), .A2(n16121), .ZN(n10521) );
  OR2_X1 U12212 ( .A1(n15596), .A2(n11792), .ZN(n11164) );
  NOR2_X1 U12213 ( .A1(n16441), .A2(n16392), .ZN(n16391) );
  NOR2_X1 U12214 ( .A1(n15892), .A2(n15893), .ZN(n15621) );
  NOR2_X1 U12215 ( .A1(n16474), .A2(n21372), .ZN(n10585) );
  AND2_X1 U12216 ( .A1(n16246), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U12217 ( .A1(n16269), .A2(n10194), .ZN(n10193) );
  NAND2_X1 U12218 ( .A1(n10135), .A2(n9834), .ZN(n10124) );
  NAND2_X1 U12219 ( .A1(n9945), .A2(n10126), .ZN(n10125) );
  OAI211_X1 U12220 ( .C1(n10813), .C2(n10818), .A(n10814), .B(n10816), .ZN(
        n10184) );
  NAND2_X1 U12221 ( .A1(n11593), .A2(n10306), .ZN(n10142) );
  NAND2_X1 U12222 ( .A1(n10066), .A2(n10065), .ZN(n11209) );
  NAND2_X1 U12223 ( .A1(n11619), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10065) );
  NAND2_X1 U12224 ( .A1(n10067), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U12225 ( .A1(n11203), .A2(n11238), .ZN(n10067) );
  AND2_X1 U12226 ( .A1(n10702), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10706) );
  NAND2_X1 U12227 ( .A1(n11186), .A2(n11026), .ZN(n11036) );
  OR2_X2 U12228 ( .A1(n11863), .A2(n11862), .ZN(n10640) );
  NAND2_X1 U12229 ( .A1(n10182), .A2(n11855), .ZN(n12532) );
  INV_X1 U12230 ( .A(n11860), .ZN(n10081) );
  INV_X1 U12231 ( .A(n11861), .ZN(n10080) );
  INV_X1 U12232 ( .A(n10478), .ZN(n10476) );
  NOR2_X1 U12233 ( .A1(n10478), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10474) );
  NOR2_X1 U12234 ( .A1(n11946), .A2(n10002), .ZN(n11944) );
  AND2_X1 U12235 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12110), .ZN(
        n12111) );
  OAI21_X1 U12236 ( .B1(n12112), .B2(n12582), .A(n18117), .ZN(n12113) );
  OAI21_X1 U12237 ( .B1(n12060), .B2(n12064), .A(n12065), .ZN(n17002) );
  OAI22_X1 U12238 ( .A1(n19234), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n19067), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12061) );
  NOR2_X1 U12239 ( .A1(n10064), .A2(n18625), .ZN(n10062) );
  AND3_X1 U12240 ( .A1(n10252), .A2(n11967), .A3(n11966), .ZN(n10251) );
  AND3_X1 U12241 ( .A1(n11968), .A2(n10254), .A3(n10253), .ZN(n10252) );
  AOI22_X1 U12242 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10247) );
  AOI21_X1 U12243 ( .B1(n17613), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n10325), .ZN(n10324) );
  NAND2_X1 U12244 ( .A1(n11985), .A2(n9933), .ZN(n10325) );
  NOR2_X1 U12245 ( .A1(n10323), .A2(n10320), .ZN(n10319) );
  INV_X1 U12246 ( .A(n11986), .ZN(n10323) );
  AND2_X1 U12247 ( .A1(n19226), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10382) );
  OR2_X1 U12248 ( .A1(n19235), .A2(n19119), .ZN(n18615) );
  INV_X1 U12249 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n21397) );
  NAND2_X1 U12250 ( .A1(n12797), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13382) );
  AND2_X1 U12251 ( .A1(n14872), .A2(n14332), .ZN(n14350) );
  MUX2_X1 U12252 ( .A(n14319), .B(n14318), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13429) );
  NOR2_X1 U12253 ( .A1(n13426), .A2(n10448), .ZN(n13431) );
  NAND2_X1 U12254 ( .A1(n10627), .A2(n13895), .ZN(n13617) );
  NOR2_X1 U12255 ( .A1(n13610), .A2(n13609), .ZN(n13618) );
  INV_X1 U12256 ( .A(n20384), .ZN(n13033) );
  INV_X1 U12257 ( .A(n13899), .ZN(n14503) );
  AOI21_X1 U12258 ( .B1(n14576), .B2(n14502), .A(n14501), .ZN(n14569) );
  NAND2_X1 U12259 ( .A1(n14448), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14469) );
  INV_X1 U12260 ( .A(n14585), .ZN(n10613) );
  OR2_X1 U12261 ( .A1(n15038), .A2(n14468), .ZN(n14225) );
  AND2_X1 U12262 ( .A1(n14614), .A2(n10614), .ZN(n14599) );
  INV_X1 U12263 ( .A(n10616), .ZN(n10614) );
  OR2_X1 U12264 ( .A1(n15047), .A2(n14468), .ZN(n14203) );
  CLKBUF_X1 U12265 ( .A(n14627), .Z(n14628) );
  AND2_X1 U12266 ( .A1(n14115), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14116) );
  OR2_X1 U12267 ( .A1(n15074), .A2(n14468), .ZN(n14145) );
  AND2_X1 U12268 ( .A1(n14077), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14078) );
  INV_X1 U12269 ( .A(n14076), .ZN(n14077) );
  NAND2_X1 U12270 ( .A1(n14078), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14114) );
  OR2_X1 U12271 ( .A1(n14706), .A2(n10608), .ZN(n10607) );
  INV_X1 U12272 ( .A(n10609), .ZN(n10608) );
  NAND2_X1 U12273 ( .A1(n14021), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14039) );
  NAND2_X1 U12274 ( .A1(n14015), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14020) );
  INV_X1 U12275 ( .A(n14014), .ZN(n14015) );
  INV_X1 U12276 ( .A(n13970), .ZN(n13931) );
  OR2_X2 U12277 ( .A1(n13968), .A2(n13967), .ZN(n13970) );
  INV_X1 U12278 ( .A(n14765), .ZN(n14911) );
  INV_X1 U12279 ( .A(n13896), .ZN(n13839) );
  NAND2_X1 U12280 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n13839), .ZN(
        n13885) );
  INV_X1 U12281 ( .A(n13838), .ZN(n13897) );
  NAND2_X1 U12282 ( .A1(n13897), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13896) );
  NAND2_X1 U12283 ( .A1(n14365), .A2(n13984), .ZN(n13903) );
  INV_X1 U12284 ( .A(n13611), .ZN(n13612) );
  INV_X1 U12285 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13475) );
  NAND2_X1 U12286 ( .A1(n9808), .A2(n13394), .ZN(n13462) );
  INV_X1 U12287 ( .A(n15099), .ZN(n10418) );
  AND2_X1 U12288 ( .A1(n14733), .A2(n14296), .ZN(n14695) );
  NAND2_X1 U12289 ( .A1(n14398), .A2(n10424), .ZN(n10423) );
  OR2_X1 U12290 ( .A1(n10630), .A2(n15116), .ZN(n10422) );
  NAND2_X1 U12291 ( .A1(n14277), .A2(n9883), .ZN(n14741) );
  INV_X1 U12292 ( .A(n14754), .ZN(n10445) );
  INV_X1 U12293 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10393) );
  NOR2_X1 U12294 ( .A1(n15136), .A2(n15135), .ZN(n10394) );
  NAND2_X1 U12295 ( .A1(n14277), .A2(n9870), .ZN(n14772) );
  OR2_X1 U12296 ( .A1(n14392), .A2(n21351), .ZN(n15150) );
  OR2_X1 U12297 ( .A1(n14392), .A2(n14399), .ZN(n15146) );
  AND2_X1 U12298 ( .A1(n14277), .A2(n10446), .ZN(n14787) );
  NAND2_X1 U12299 ( .A1(n14277), .A2(n14276), .ZN(n14818) );
  AND2_X1 U12300 ( .A1(n14275), .A2(n14274), .ZN(n14828) );
  NAND2_X1 U12301 ( .A1(n14919), .A2(n14913), .ZN(n14816) );
  NAND2_X1 U12302 ( .A1(n15210), .A2(n15422), .ZN(n10396) );
  AND2_X1 U12303 ( .A1(n14265), .A2(n14264), .ZN(n14917) );
  NAND2_X1 U12304 ( .A1(n14256), .A2(n9873), .ZN(n14918) );
  AND2_X1 U12305 ( .A1(n14256), .A2(n10456), .ZN(n14919) );
  AND2_X1 U12306 ( .A1(n9873), .A2(n10457), .ZN(n10456) );
  INV_X1 U12307 ( .A(n14917), .ZN(n10457) );
  NAND2_X1 U12308 ( .A1(n14256), .A2(n10459), .ZN(n14928) );
  INV_X1 U12309 ( .A(n14386), .ZN(n14385) );
  NAND2_X1 U12310 ( .A1(n14386), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16792) );
  AND2_X1 U12311 ( .A1(n14255), .A2(n14254), .ZN(n16813) );
  NAND3_X1 U12312 ( .A1(n9971), .A2(n13549), .A3(n9967), .ZN(n13550) );
  NAND2_X1 U12313 ( .A1(n9974), .A2(n9972), .ZN(n9971) );
  NAND3_X1 U12314 ( .A1(n9970), .A2(n9969), .A3(n20423), .ZN(n9967) );
  XNOR2_X1 U12315 ( .A(n14362), .B(n13555), .ZN(n13551) );
  AND2_X1 U12316 ( .A1(n13558), .A2(n13557), .ZN(n13565) );
  AND2_X1 U12317 ( .A1(n13563), .A2(n13562), .ZN(n13586) );
  OR2_X1 U12318 ( .A1(n15339), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20474) );
  NAND2_X1 U12319 ( .A1(n10414), .A2(n14409), .ZN(n13196) );
  NAND2_X1 U12320 ( .A1(n9962), .A2(n13369), .ZN(n13100) );
  NAND2_X1 U12321 ( .A1(n9960), .A2(n9958), .ZN(n9963) );
  AOI21_X1 U12322 ( .B1(n9961), .B2(n9748), .A(n9959), .ZN(n9958) );
  NAND2_X1 U12323 ( .A1(n13097), .A2(n10426), .ZN(n12947) );
  AND2_X1 U12324 ( .A1(n9764), .A2(n9852), .ZN(n10426) );
  INV_X1 U12325 ( .A(n9981), .ZN(n9980) );
  INV_X1 U12326 ( .A(n12914), .ZN(n13442) );
  NOR2_X1 U12327 ( .A1(n13440), .A2(n9902), .ZN(n13444) );
  AND3_X1 U12328 ( .A1(n12797), .A2(n12891), .A3(n12818), .ZN(n12798) );
  NAND2_X1 U12329 ( .A1(n12874), .A2(n10038), .ZN(n12875) );
  NAND2_X1 U12330 ( .A1(n12817), .A2(n10039), .ZN(n10038) );
  OAI21_X1 U12331 ( .B1(n20613), .B2(n20612), .A(n20908), .ZN(n20618) );
  INV_X1 U12332 ( .A(n20750), .ZN(n21033) );
  NAND2_X1 U12333 ( .A1(n12869), .A2(n10020), .ZN(n16744) );
  OR2_X1 U12334 ( .A1(n20221), .A2(n11612), .ZN(n11253) );
  AND2_X1 U12335 ( .A1(n10542), .A2(n15839), .ZN(n10541) );
  AOI21_X1 U12336 ( .B1(n15580), .B2(n11664), .A(n16098), .ZN(n15582) );
  AND2_X1 U12337 ( .A1(n10540), .A2(n11093), .ZN(n10539) );
  AND2_X1 U12338 ( .A1(n11136), .A2(n11139), .ZN(n15656) );
  AND2_X1 U12339 ( .A1(n11133), .A2(n11117), .ZN(n15667) );
  AND2_X1 U12340 ( .A1(n11061), .A2(n11082), .ZN(n10504) );
  MUX2_X1 U12341 ( .A(n11581), .B(n11033), .S(n19534), .Z(n11056) );
  NAND2_X1 U12342 ( .A1(n19534), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11040) );
  AND2_X1 U12343 ( .A1(n14530), .A2(n10566), .ZN(n11796) );
  NOR2_X1 U12344 ( .A1(n10567), .A2(n11795), .ZN(n10566) );
  AND2_X1 U12345 ( .A1(n13808), .A2(n15640), .ZN(n15639) );
  AND2_X1 U12346 ( .A1(n15905), .A2(n12179), .ZN(n10594) );
  AOI22_X1 U12347 ( .A1(n10089), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11512) );
  AOI21_X1 U12348 ( .B1(n10089), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n10091), .ZN(n11495) );
  AND2_X1 U12349 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10091) );
  AOI22_X1 U12350 ( .A1(n10089), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11485) );
  AND2_X1 U12351 ( .A1(n11285), .A2(n11284), .ZN(n13777) );
  AOI22_X1 U12352 ( .A1(n10089), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11472) );
  AND2_X1 U12353 ( .A1(n12172), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12173) );
  INV_X1 U12354 ( .A(n10546), .ZN(n10544) );
  NAND2_X1 U12355 ( .A1(n9766), .A2(n10590), .ZN(n10589) );
  INV_X1 U12356 ( .A(n12335), .ZN(n10590) );
  AND2_X1 U12357 ( .A1(n11554), .A2(n11553), .ZN(n15618) );
  AND2_X1 U12358 ( .A1(n11551), .A2(n11550), .ZN(n15995) );
  CLKBUF_X1 U12359 ( .A(n15883), .Z(n15890) );
  AND2_X1 U12360 ( .A1(n11549), .A2(n11548), .ZN(n16002) );
  AND3_X1 U12361 ( .A1(n11433), .A2(n11432), .A3(n11431), .ZN(n15745) );
  AND2_X1 U12362 ( .A1(n11424), .A2(n11429), .ZN(n10535) );
  OAI211_X1 U12363 ( .C1(n11534), .C2(n11401), .A(n11411), .B(n11400), .ZN(
        n13706) );
  INV_X1 U12364 ( .A(n11206), .ZN(n19411) );
  AOI21_X1 U12365 ( .B1(n19409), .B2(n19408), .A(n20228), .ZN(n19439) );
  AND2_X1 U12366 ( .A1(n9909), .A2(n16316), .ZN(n10366) );
  NAND2_X1 U12367 ( .A1(n11671), .A2(n10489), .ZN(n11679) );
  NAND2_X1 U12368 ( .A1(n11644), .A2(n9769), .ZN(n11657) );
  NAND2_X1 U12369 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10471) );
  AOI21_X1 U12370 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11289), .ZN(n13741) );
  NAND2_X1 U12371 ( .A1(n10578), .A2(n10579), .ZN(n16236) );
  NAND2_X1 U12372 ( .A1(n11603), .A2(n16246), .ZN(n10579) );
  NAND2_X1 U12373 ( .A1(n16243), .A2(n11600), .ZN(n10578) );
  AOI21_X1 U12374 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11274), .ZN(n13731) );
  NOR2_X1 U12375 ( .A1(n16282), .A2(n11623), .ZN(n10472) );
  NAND2_X1 U12376 ( .A1(n11622), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11626) );
  AND3_X1 U12377 ( .A1(n10086), .A2(n9807), .A3(n11816), .ZN(n10085) );
  NOR2_X1 U12378 ( .A1(n10600), .A2(n11816), .ZN(n10275) );
  NAND2_X1 U12379 ( .A1(n10086), .A2(n9807), .ZN(n10088) );
  OR2_X1 U12380 ( .A1(n10598), .A2(n16029), .ZN(n10279) );
  OR2_X1 U12381 ( .A1(n9754), .A2(n16029), .ZN(n10280) );
  AND2_X1 U12382 ( .A1(n11572), .A2(n10545), .ZN(n10543) );
  NOR2_X1 U12383 ( .A1(n15507), .A2(n10546), .ZN(n10545) );
  INV_X1 U12384 ( .A(n10567), .ZN(n10565) );
  OR2_X1 U12385 ( .A1(n15525), .A2(n11792), .ZN(n16045) );
  NAND2_X1 U12386 ( .A1(n16053), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16054) );
  NOR2_X1 U12387 ( .A1(n9910), .A2(n16383), .ZN(n10344) );
  AOI21_X1 U12388 ( .B1(n9744), .B2(n10353), .A(n10347), .ZN(n10346) );
  NAND2_X1 U12389 ( .A1(n16095), .A2(n9744), .ZN(n10345) );
  INV_X1 U12390 ( .A(n16064), .ZN(n10347) );
  XNOR2_X1 U12391 ( .A(n11784), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16063) );
  AND2_X1 U12392 ( .A1(n10303), .A2(n11774), .ZN(n10302) );
  OR2_X1 U12393 ( .A1(n11767), .A2(n10304), .ZN(n10303) );
  AND2_X1 U12394 ( .A1(n10351), .A2(n10349), .ZN(n10348) );
  NAND2_X1 U12395 ( .A1(n10354), .A2(n10350), .ZN(n10349) );
  OR2_X1 U12396 ( .A1(n9814), .A2(n10352), .ZN(n10351) );
  AND2_X1 U12397 ( .A1(n16381), .A2(n11386), .ZN(n16355) );
  OR2_X1 U12398 ( .A1(n12442), .A2(n11371), .ZN(n16367) );
  AND2_X1 U12399 ( .A1(n11330), .A2(n11329), .ZN(n15863) );
  NAND2_X1 U12400 ( .A1(n12454), .A2(n10571), .ZN(n11697) );
  NAND2_X1 U12401 ( .A1(n16391), .A2(n11382), .ZN(n12442) );
  NAND2_X1 U12402 ( .A1(n12454), .A2(n12455), .ZN(n12453) );
  INV_X1 U12403 ( .A(n16121), .ZN(n10364) );
  INV_X1 U12404 ( .A(n9792), .ZN(n10361) );
  NOR2_X1 U12405 ( .A1(n11836), .A2(n11837), .ZN(n16131) );
  AND2_X1 U12406 ( .A1(n11113), .A2(n11835), .ZN(n16139) );
  NAND2_X1 U12407 ( .A1(n10137), .A2(n9833), .ZN(n11834) );
  NAND2_X1 U12408 ( .A1(n16213), .A2(n10139), .ZN(n10137) );
  AND2_X1 U12409 ( .A1(n16156), .A2(n16145), .ZN(n10356) );
  AND2_X1 U12410 ( .A1(n11297), .A2(n11296), .ZN(n13798) );
  INV_X1 U12411 ( .A(n13488), .ZN(n11507) );
  AND2_X1 U12412 ( .A1(n16538), .A2(n11376), .ZN(n16482) );
  NAND2_X1 U12413 ( .A1(n13760), .A2(n9793), .ZN(n13799) );
  AND2_X1 U12414 ( .A1(n13760), .A2(n10563), .ZN(n13787) );
  AND3_X1 U12415 ( .A1(n11481), .A2(n11480), .A3(n11479), .ZN(n13356) );
  INV_X1 U12416 ( .A(n13275), .ZN(n11468) );
  AND2_X1 U12417 ( .A1(n13497), .A2(n9758), .ZN(n13751) );
  NAND2_X1 U12418 ( .A1(n9976), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16247) );
  NAND2_X1 U12419 ( .A1(n11601), .A2(n11596), .ZN(n16244) );
  AND2_X1 U12420 ( .A1(n11271), .A2(n11270), .ZN(n13603) );
  NAND2_X1 U12421 ( .A1(n13497), .A2(n9796), .ZN(n13732) );
  CLKBUF_X1 U12422 ( .A(n16243), .Z(n16258) );
  INV_X1 U12423 ( .A(n11597), .ZN(n16269) );
  NAND2_X1 U12424 ( .A1(n16296), .A2(n11591), .ZN(n11594) );
  NAND2_X1 U12425 ( .A1(n10816), .A2(n10815), .ZN(n10432) );
  AND2_X1 U12426 ( .A1(n11406), .A2(n11405), .ZN(n13188) );
  NAND2_X1 U12427 ( .A1(n13189), .A2(n13188), .ZN(n13191) );
  AND2_X1 U12428 ( .A1(n11415), .A2(n11414), .ZN(n13702) );
  NAND2_X1 U12429 ( .A1(n13703), .A2(n13702), .ZN(n13705) );
  XNOR2_X1 U12430 ( .A(n16650), .B(n12156), .ZN(n13291) );
  AOI21_X1 U12431 ( .B1(n12153), .B2(n12152), .A(n12151), .ZN(n13290) );
  AND2_X2 U12432 ( .A1(n10679), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13656) );
  NAND2_X1 U12433 ( .A1(n10122), .A2(n13654), .ZN(n13662) );
  INV_X1 U12434 ( .A(n11574), .ZN(n10122) );
  XNOR2_X1 U12435 ( .A(n12167), .B(n12165), .ZN(n13313) );
  AND2_X1 U12436 ( .A1(n11362), .A2(n11361), .ZN(n13661) );
  NAND2_X1 U12437 ( .A1(n10754), .A2(n11030), .ZN(n10761) );
  AND2_X1 U12438 ( .A1(n20190), .A2(n19502), .ZN(n19557) );
  INV_X1 U12439 ( .A(n19974), .ZN(n19913) );
  NAND2_X1 U12440 ( .A1(n10290), .A2(n9816), .ZN(n10109) );
  NAND2_X1 U12441 ( .A1(n10295), .A2(n9815), .ZN(n10108) );
  OAI21_X1 U12442 ( .B1(n10693), .B2(n10694), .A(n11030), .ZN(n10111) );
  NAND2_X1 U12443 ( .A1(n10688), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10110) );
  INV_X1 U12444 ( .A(n19546), .ZN(n19538) );
  INV_X1 U12445 ( .A(n19547), .ZN(n19539) );
  NAND2_X1 U12446 ( .A1(n20033), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19549) );
  NOR2_X2 U12447 ( .A1(n19497), .A2(n19498), .ZN(n19547) );
  OR2_X1 U12448 ( .A1(n19807), .A2(n20211), .ZN(n19974) );
  OR2_X1 U12449 ( .A1(n20190), .A2(n19502), .ZN(n20028) );
  NAND2_X1 U12450 ( .A1(n18617), .A2(n19260), .ZN(n12084) );
  NOR2_X1 U12451 ( .A1(n17045), .A2(n17294), .ZN(n17040) );
  OR2_X1 U12452 ( .A1(n17084), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n9994) );
  INV_X1 U12453 ( .A(n18009), .ZN(n10487) );
  NAND2_X1 U12454 ( .A1(n17295), .A2(n17631), .ZN(n17287) );
  NOR2_X1 U12455 ( .A1(n17312), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n17295) );
  NOR2_X1 U12456 ( .A1(n17749), .A2(n17382), .ZN(n10217) );
  NAND2_X1 U12457 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_18__SCAN_IN), 
        .ZN(n10208) );
  NOR2_X1 U12458 ( .A1(n17243), .A2(n10211), .ZN(n10210) );
  INV_X1 U12459 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U12460 ( .A1(n17876), .A2(n17874), .ZN(n10264) );
  NOR2_X1 U12461 ( .A1(n17707), .A2(n10262), .ZN(n10261) );
  NAND2_X1 U12462 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_16__SCAN_IN), 
        .ZN(n10262) );
  INV_X1 U12463 ( .A(n11862), .ZN(n10181) );
  INV_X1 U12464 ( .A(n11902), .ZN(n10381) );
  AND2_X1 U12465 ( .A1(n10385), .A2(n10384), .ZN(n11901) );
  NAND2_X1 U12466 ( .A1(n9819), .A2(n11855), .ZN(n10385) );
  NAND2_X1 U12467 ( .A1(n17332), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10246) );
  AOI22_X1 U12468 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17567), .B1(
        n11903), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11899) );
  NAND2_X1 U12469 ( .A1(n11970), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11898) );
  NAND2_X1 U12470 ( .A1(n17457), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10234) );
  NAND2_X1 U12471 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11884) );
  NOR2_X1 U12472 ( .A1(n10079), .A2(n10077), .ZN(n10076) );
  INV_X1 U12473 ( .A(n12014), .ZN(n10079) );
  NOR2_X1 U12474 ( .A1(n17853), .A2(n17814), .ZN(n17832) );
  INV_X1 U12475 ( .A(n16690), .ZN(n17855) );
  NAND2_X1 U12476 ( .A1(n12628), .A2(n10652), .ZN(n17951) );
  AND2_X1 U12477 ( .A1(n9876), .A2(n12587), .ZN(n10503) );
  AND2_X1 U12478 ( .A1(n17156), .A2(n9876), .ZN(n18005) );
  INV_X1 U12479 ( .A(n17198), .ZN(n10496) );
  NAND4_X1 U12480 ( .A1(n18192), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18123) );
  INV_X1 U12481 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18130) );
  NOR2_X1 U12482 ( .A1(n17198), .A2(n18123), .ZN(n17200) );
  INV_X1 U12483 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18194) );
  NOR2_X1 U12484 ( .A1(n18237), .A2(n18238), .ZN(n18209) );
  AND2_X1 U12485 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18252) );
  NOR2_X1 U12486 ( .A1(n18304), .A2(n9880), .ZN(n18314) );
  NOR2_X1 U12487 ( .A1(n18109), .A2(n9900), .ZN(n17962) );
  NAND2_X1 U12488 ( .A1(n17962), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17961) );
  OR2_X1 U12489 ( .A1(n18109), .A2(n10179), .ZN(n18334) );
  NOR2_X1 U12490 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18029), .ZN(
        n18010) );
  INV_X1 U12491 ( .A(n17989), .ZN(n18011) );
  NOR2_X1 U12492 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18065), .ZN(
        n18037) );
  OR2_X1 U12493 ( .A1(n18076), .A2(n18199), .ZN(n10238) );
  NOR2_X1 U12494 ( .A1(n18400), .A2(n12116), .ZN(n10549) );
  NAND2_X1 U12495 ( .A1(n10242), .A2(n9903), .ZN(n10241) );
  NAND2_X1 U12496 ( .A1(n18480), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10551) );
  NAND2_X1 U12497 ( .A1(n16901), .A2(n18436), .ZN(n18453) );
  NAND2_X1 U12498 ( .A1(n10004), .A2(n10242), .ZN(n18165) );
  NAND2_X1 U12499 ( .A1(n18223), .A2(n11956), .ZN(n18207) );
  NAND2_X1 U12500 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18224), .ZN(
        n18223) );
  NAND2_X1 U12501 ( .A1(n10548), .A2(n10001), .ZN(n10000) );
  AND2_X1 U12502 ( .A1(n12104), .A2(n9785), .ZN(n10001) );
  NOR2_X1 U12503 ( .A1(n19275), .A2(n12476), .ZN(n19060) );
  XNOR2_X1 U12504 ( .A(n17808), .B(n21317), .ZN(n18280) );
  NAND2_X1 U12505 ( .A1(n18288), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18287) );
  INV_X1 U12506 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19067) );
  NAND2_X1 U12507 ( .A1(n10336), .A2(n10335), .ZN(n10334) );
  NAND2_X1 U12508 ( .A1(n10244), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16698) );
  INV_X1 U12509 ( .A(n10245), .ZN(n10244) );
  NOR2_X2 U12510 ( .A1(n11996), .A2(n11995), .ZN(n18632) );
  NOR2_X2 U12511 ( .A1(n11980), .A2(n11979), .ZN(n18636) );
  INV_X1 U12512 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19066) );
  NAND2_X1 U12513 ( .A1(n19263), .A2(n18615), .ZN(n18690) );
  OAI21_X1 U12514 ( .B1(n18574), .B2(n19059), .A(n10662), .ZN(n19061) );
  OR3_X1 U12515 ( .A1(n13328), .A2(n12897), .A3(n20246), .ZN(n13073) );
  OR2_X1 U12516 ( .A1(n12868), .A2(n20246), .ZN(n12832) );
  NAND2_X1 U12517 ( .A1(n13073), .A2(n12832), .ZN(n14557) );
  INV_X1 U12518 ( .A(n20335), .ZN(n16781) );
  INV_X1 U12519 ( .A(n20327), .ZN(n20341) );
  AND2_X1 U12520 ( .A1(n20355), .A2(n14551), .ZN(n20350) );
  INV_X1 U12521 ( .A(n20350), .ZN(n14930) );
  INV_X1 U12522 ( .A(n14556), .ZN(n14988) );
  NOR2_X2 U12523 ( .A1(n13210), .A2(n13209), .ZN(n15006) );
  NOR2_X1 U12524 ( .A1(n13033), .A2(n20382), .ZN(n16767) );
  BUF_X1 U12525 ( .A(n16767), .Z(n20381) );
  CLKBUF_X1 U12526 ( .A(n20372), .Z(n20382) );
  INV_X1 U12527 ( .A(n20487), .ZN(n20428) );
  INV_X1 U12528 ( .A(n20421), .ZN(n15138) );
  INV_X1 U12529 ( .A(n20253), .ZN(n20429) );
  NOR2_X1 U12530 ( .A1(n14570), .A2(n14421), .ZN(n14889) );
  OR2_X1 U12531 ( .A1(n10161), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9957) );
  XNOR2_X1 U12532 ( .A(n14575), .B(n14574), .ZN(n15232) );
  AOI21_X1 U12533 ( .B1(n14572), .B2(n14571), .A(n14570), .ZN(n14575) );
  NAND2_X1 U12534 ( .A1(n10407), .A2(n10405), .ZN(n15010) );
  NAND2_X1 U12535 ( .A1(n15033), .A2(n10406), .ZN(n10405) );
  NAND2_X1 U12536 ( .A1(n10428), .A2(n10408), .ZN(n10407) );
  XNOR2_X1 U12537 ( .A(n10374), .B(n10373), .ZN(n10057) );
  INV_X1 U12538 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10373) );
  OAI211_X1 U12539 ( .C1(n15026), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10375), .B(n15025), .ZN(n10374) );
  XNOR2_X1 U12540 ( .A(n10118), .B(n15035), .ZN(n15257) );
  NAND2_X1 U12541 ( .A1(n10121), .A2(n10119), .ZN(n10118) );
  NAND2_X1 U12542 ( .A1(n15034), .A2(n10120), .ZN(n10119) );
  NAND2_X1 U12543 ( .A1(n15033), .A2(n15189), .ZN(n10121) );
  NAND2_X1 U12544 ( .A1(n10372), .A2(n15210), .ZN(n15079) );
  XNOR2_X1 U12545 ( .A(n10416), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15308) );
  NAND2_X1 U12546 ( .A1(n10421), .A2(n10417), .ZN(n10416) );
  NAND2_X1 U12547 ( .A1(n15090), .A2(n10120), .ZN(n10421) );
  NAND2_X1 U12548 ( .A1(n10418), .A2(n9878), .ZN(n10417) );
  INV_X1 U12549 ( .A(n15087), .ZN(n15117) );
  XNOR2_X1 U12550 ( .A(n10390), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15360) );
  OAI21_X1 U12551 ( .B1(n10394), .B2(n10392), .A(n10391), .ZN(n10390) );
  NAND2_X1 U12552 ( .A1(n15189), .A2(n10393), .ZN(n10392) );
  NAND2_X1 U12553 ( .A1(n10394), .A2(n10120), .ZN(n10391) );
  AND2_X1 U12554 ( .A1(n15407), .A2(n15406), .ZN(n15449) );
  INV_X1 U12555 ( .A(n9974), .ZN(n20424) );
  AND2_X1 U12556 ( .A1(n13345), .A2(n13338), .ZN(n20454) );
  OAI21_X1 U12557 ( .B1(n13456), .B2(n16829), .A(n20653), .ZN(n20483) );
  NAND2_X1 U12558 ( .A1(n12972), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16754) );
  INV_X1 U12559 ( .A(n13328), .ZN(n12972) );
  NAND2_X1 U12560 ( .A1(n10401), .A2(n20648), .ZN(n12934) );
  INV_X1 U12561 ( .A(n12948), .ZN(n10401) );
  OAI211_X1 U12562 ( .C1(n20503), .C2(n20500), .A(n20498), .B(n20836), .ZN(
        n20538) );
  OAI221_X1 U12563 ( .B1(n20908), .B2(n20546), .C1(n21030), .C2(n20545), .A(
        n21035), .ZN(n20563) );
  OAI21_X1 U12564 ( .B1(n20577), .B2(n20575), .A(n20574), .ZN(n20601) );
  OAI21_X1 U12565 ( .B1(n20672), .B2(n20655), .A(n20994), .ZN(n20673) );
  INV_X1 U12566 ( .A(n20703), .ZN(n20692) );
  OAI211_X1 U12567 ( .C1(n20710), .C2(n20913), .A(n20994), .B(n20709), .ZN(
        n20738) );
  OAI21_X1 U12568 ( .B1(n20752), .B2(n20751), .A(n21035), .ZN(n20771) );
  OAI211_X1 U12569 ( .C1(n20796), .C2(n20913), .A(n20836), .B(n20780), .ZN(
        n20798) );
  AND2_X1 U12570 ( .A1(n20742), .A2(n20871), .ZN(n20797) );
  OAI22_X1 U12571 ( .A1(n20843), .A2(n20842), .B1(n20841), .B2(n20990), .ZN(
        n20867) );
  INV_X1 U12572 ( .A(n20839), .ZN(n20868) );
  OR2_X1 U12573 ( .A1(n20873), .A2(n20829), .ZN(n20891) );
  NAND2_X1 U12574 ( .A1(n20533), .A2(n10018), .ZN(n20925) );
  OAI211_X1 U12575 ( .C1(n20914), .C2(n20913), .A(n20994), .B(n20912), .ZN(
        n20949) );
  OAI211_X1 U12576 ( .C1(n21018), .C2(n20995), .A(n20994), .B(n20993), .ZN(
        n21021) );
  INV_X1 U12577 ( .A(n20906), .ZN(n21032) );
  INV_X1 U12578 ( .A(n20921), .ZN(n21043) );
  INV_X1 U12579 ( .A(n20925), .ZN(n21049) );
  INV_X1 U12580 ( .A(n20929), .ZN(n21055) );
  INV_X1 U12581 ( .A(n20933), .ZN(n21061) );
  INV_X1 U12582 ( .A(n21088), .ZN(n21068) );
  INV_X1 U12583 ( .A(n20937), .ZN(n21067) );
  INV_X1 U12584 ( .A(n20941), .ZN(n21074) );
  NAND2_X1 U12585 ( .A1(n20987), .A2(n20986), .ZN(n21088) );
  INV_X1 U12586 ( .A(n21071), .ZN(n21084) );
  INV_X1 U12587 ( .A(n20946), .ZN(n21082) );
  AND2_X1 U12588 ( .A1(n11786), .A2(n11782), .ZN(n15515) );
  AND2_X1 U12589 ( .A1(n11181), .A2(n10542), .ZN(n15538) );
  MUX2_X1 U12590 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n11182), .S(n9802), .Z(
        n11183) );
  AND2_X1 U12591 ( .A1(n15563), .A2(n11176), .ZN(n15586) );
  AOI21_X1 U12592 ( .B1(n19307), .B2(n11664), .A(n19306), .ZN(n19310) );
  NAND2_X1 U12593 ( .A1(n14549), .A2(n11755), .ZN(n19355) );
  INV_X1 U12594 ( .A(n19320), .ZN(n16718) );
  AND2_X1 U12595 ( .A1(n19355), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19337) );
  INV_X1 U12596 ( .A(n19368), .ZN(n19324) );
  NAND2_X1 U12597 ( .A1(n11664), .A2(n19344), .ZN(n15816) );
  OR2_X1 U12598 ( .A1(n11451), .A2(n11450), .ZN(n13755) );
  OR2_X1 U12599 ( .A1(n13601), .A2(n13600), .ZN(n13754) );
  INV_X1 U12600 ( .A(n15897), .ZN(n15904) );
  INV_X1 U12601 ( .A(n20199), .ZN(n19502) );
  NAND2_X1 U12602 ( .A1(n13066), .A2(n13065), .ZN(n19501) );
  XNOR2_X1 U12603 ( .A(n10587), .B(n10586), .ZN(n10670) );
  INV_X1 U12604 ( .A(n12409), .ZN(n10586) );
  NAND2_X1 U12605 ( .A1(n15819), .A2(n12387), .ZN(n10587) );
  XNOR2_X1 U12606 ( .A(n14520), .B(n10665), .ZN(n14536) );
  INV_X1 U12607 ( .A(n15985), .ZN(n16008) );
  AND2_X1 U12608 ( .A1(n12941), .A2(n19499), .ZN(n16011) );
  AOI21_X2 U12609 ( .B1(n12846), .B2(n12414), .A(n13775), .ZN(n16017) );
  INV_X1 U12610 ( .A(n16017), .ZN(n19396) );
  INV_X1 U12611 ( .A(n16014), .ZN(n19397) );
  BUF_X1 U12612 ( .A(n19460), .Z(n20237) );
  NOR2_X1 U12614 ( .A1(n13114), .A2(n13063), .ZN(n13136) );
  OR2_X1 U12615 ( .A1(n13177), .A2(n13115), .ZN(n13154) );
  NAND2_X1 U12616 ( .A1(n16236), .A2(n16235), .ZN(n16546) );
  INV_X1 U12617 ( .A(n16283), .ZN(n19483) );
  XNOR2_X1 U12618 ( .A(n10190), .B(n16031), .ZN(n16313) );
  OAI21_X1 U12619 ( .B1(n10600), .B2(n9754), .A(n10598), .ZN(n10190) );
  NAND2_X1 U12620 ( .A1(n16322), .A2(n16838), .ZN(n10070) );
  NOR2_X1 U12621 ( .A1(n16068), .A2(n10147), .ZN(n16352) );
  AND2_X1 U12622 ( .A1(n16462), .A2(n11384), .ZN(n16381) );
  NOR2_X1 U12623 ( .A1(n10069), .A2(n10068), .ZN(n11384) );
  AND2_X1 U12624 ( .A1(n16556), .A2(n11383), .ZN(n10068) );
  NOR2_X1 U12625 ( .A1(n12442), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10069) );
  AND2_X1 U12626 ( .A1(n15589), .A2(n15588), .ZN(n16375) );
  AND2_X1 U12627 ( .A1(n10597), .A2(n11168), .ZN(n16108) );
  XNOR2_X1 U12628 ( .A(n16118), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16404) );
  INV_X1 U12629 ( .A(n9935), .ZN(n9936) );
  OAI22_X1 U12630 ( .A1(n16455), .A2(n16842), .B1(n16461), .B2(n16441), .ZN(
        n16446) );
  NOR2_X1 U12631 ( .A1(n16432), .A2(n16431), .ZN(n16433) );
  NOR2_X1 U12632 ( .A1(n16430), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16431) );
  OAI21_X1 U12634 ( .B1(n16213), .B2(n10141), .A(n10139), .ZN(n16147) );
  NAND2_X1 U12635 ( .A1(n16165), .A2(n16474), .ZN(n9985) );
  NAND2_X1 U12636 ( .A1(n10138), .A2(n10508), .ZN(n16157) );
  NAND2_X1 U12637 ( .A1(n16213), .A2(n10510), .ZN(n10138) );
  NAND2_X1 U12638 ( .A1(n16165), .A2(n9940), .ZN(n16492) );
  NAND2_X1 U12639 ( .A1(n12450), .A2(n21372), .ZN(n9940) );
  AND2_X1 U12640 ( .A1(n16535), .A2(n11378), .ZN(n16496) );
  XNOR2_X1 U12641 ( .A(n16198), .B(n16197), .ZN(n16504) );
  AND2_X1 U12642 ( .A1(n16570), .A2(n16547), .ZN(n16538) );
  NAND2_X1 U12643 ( .A1(n13054), .A2(n13053), .ZN(n13059) );
  INV_X1 U12644 ( .A(n16836), .ZN(n16633) );
  NAND2_X1 U12645 ( .A1(n13289), .A2(n13292), .ZN(n20199) );
  OR2_X1 U12646 ( .A1(n13291), .A2(n13290), .ZN(n13292) );
  NAND2_X1 U12647 ( .A1(n13311), .A2(n13314), .ZN(n20190) );
  OR2_X1 U12648 ( .A1(n13313), .A2(n13312), .ZN(n13314) );
  OAI21_X1 U12649 ( .B1(n19505), .B2(n19542), .A(n20033), .ZN(n19554) );
  AND2_X1 U12650 ( .A1(n19564), .A2(n19560), .ZN(n19582) );
  INV_X1 U12651 ( .A(n19614), .ZN(n19587) );
  OAI211_X1 U12652 ( .C1(n19612), .C2(n19597), .A(n19596), .B(n20033), .ZN(
        n19615) );
  OAI21_X1 U12653 ( .B1(n19628), .B2(n19627), .A(n19626), .ZN(n19646) );
  OAI21_X1 U12654 ( .B1(n19628), .B2(n19624), .A(n19623), .ZN(n19647) );
  INV_X1 U12655 ( .A(n19641), .ZN(n19650) );
  OAI211_X1 U12656 ( .C1(n19659), .C2(n19674), .A(n20033), .B(n19658), .ZN(
        n19677) );
  AND2_X1 U12657 ( .A1(n19683), .A2(n19682), .ZN(n19704) );
  INV_X1 U12658 ( .A(n19704), .ZN(n19711) );
  AND2_X1 U12659 ( .A1(n19715), .A2(n19912), .ZN(n19709) );
  OAI21_X1 U12660 ( .B1(n19721), .B2(n19736), .A(n20033), .ZN(n19739) );
  NAND2_X1 U12661 ( .A1(n19747), .A2(n19715), .ZN(n19767) );
  OAI211_X1 U12662 ( .C1(n19815), .C2(n19810), .A(n20033), .B(n19809), .ZN(
        n19845) );
  OAI21_X1 U12663 ( .B1(n19815), .B2(n19814), .A(n19813), .ZN(n19844) );
  OAI21_X1 U12664 ( .B1(n19881), .B2(n19850), .A(n19849), .ZN(n19871) );
  NAND2_X1 U12665 ( .A1(n19913), .A2(n20178), .ZN(n19903) );
  INV_X1 U12666 ( .A(n20056), .ZN(n19928) );
  AOI21_X1 U12667 ( .B1(n20207), .B2(n19916), .A(n19917), .ZN(n19938) );
  AND2_X1 U12668 ( .A1(n19952), .A2(n19947), .ZN(n19969) );
  OAI22_X1 U12669 ( .A1(n19512), .A2(n19539), .B1(n15998), .B2(n19538), .ZN(
        n19988) );
  OAI21_X1 U12670 ( .B1(n19985), .B2(n19984), .A(n19983), .ZN(n20017) );
  AND2_X1 U12671 ( .A1(n20033), .A2(n19506), .ZN(n20026) );
  AND2_X1 U12672 ( .A1(n20033), .A2(n19515), .ZN(n20040) );
  INV_X1 U12673 ( .A(n19988), .ZN(n20044) );
  AND2_X1 U12674 ( .A1(n20033), .A2(n19520), .ZN(n20046) );
  AND2_X1 U12675 ( .A1(n20033), .A2(n19530), .ZN(n20058) );
  INV_X1 U12676 ( .A(n20086), .ZN(n20072) );
  OR2_X1 U12677 ( .A1(n19944), .A2(n20028), .ZN(n20075) );
  INV_X1 U12678 ( .A(n20075), .ZN(n20082) );
  AND2_X1 U12679 ( .A1(n20032), .A2(n20024), .ZN(n20080) );
  AND2_X1 U12680 ( .A1(n20033), .A2(n19552), .ZN(n20079) );
  INV_X1 U12681 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19977) );
  NAND2_X1 U12682 ( .A1(n19061), .A2(n19258), .ZN(n17005) );
  NOR2_X1 U12683 ( .A1(n17294), .A2(n17027), .ZN(n17035) );
  XNOR2_X1 U12684 ( .A(n17040), .B(n10469), .ZN(n10468) );
  INV_X1 U12685 ( .A(n17041), .ZN(n10469) );
  NAND2_X1 U12686 ( .A1(n9999), .A2(n9823), .ZN(n9998) );
  OAI21_X1 U12687 ( .B1(n17044), .B2(n17377), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n9999) );
  OR2_X1 U12688 ( .A1(n17362), .A2(n17954), .ZN(n10462) );
  NAND2_X1 U12689 ( .A1(n17091), .A2(n10463), .ZN(n10461) );
  INV_X1 U12690 ( .A(n17376), .ZN(n17365) );
  INV_X1 U12691 ( .A(n9994), .ZN(n17074) );
  NOR2_X1 U12692 ( .A1(n17079), .A2(n17968), .ZN(n17078) );
  NOR2_X1 U12693 ( .A1(n17091), .A2(n17294), .ZN(n17079) );
  NAND2_X1 U12694 ( .A1(n17090), .A2(n17383), .ZN(n17084) );
  NOR2_X1 U12695 ( .A1(n17123), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n17109) );
  NAND2_X1 U12696 ( .A1(n17109), .A2(n17104), .ZN(n17103) );
  NOR2_X1 U12697 ( .A1(n17111), .A2(n18009), .ZN(n17110) );
  NOR2_X1 U12698 ( .A1(n17119), .A2(n17294), .ZN(n17111) );
  NOR2_X1 U12699 ( .A1(n17148), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17131) );
  NAND2_X1 U12700 ( .A1(n17131), .A2(n17124), .ZN(n17123) );
  NOR2_X1 U12701 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17170), .ZN(n17152) );
  NOR2_X1 U12702 ( .A1(n17193), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17178) );
  NAND2_X1 U12703 ( .A1(n17178), .A2(n17171), .ZN(n17170) );
  NOR2_X1 U12704 ( .A1(n17215), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n17202) );
  NAND2_X1 U12705 ( .A1(n17202), .A2(n17194), .ZN(n17193) );
  NOR2_X1 U12706 ( .A1(n17287), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17276) );
  NAND2_X1 U12707 ( .A1(n17276), .A2(n17270), .ZN(n17267) );
  AND3_X1 U12708 ( .A1(n9997), .A2(n9996), .A3(n9995), .ZN(n17349) );
  INV_X1 U12709 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17343) );
  AOI211_X2 U12710 ( .C1(n19115), .C2(n18932), .A(n12626), .B(n19276), .ZN(
        n17373) );
  AND2_X1 U12711 ( .A1(n17452), .A2(n9775), .ZN(n17420) );
  NAND2_X1 U12712 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(P3_EBX_REG_20__SCAN_IN), 
        .ZN(n10206) );
  NOR3_X1 U12713 ( .A1(n17489), .A2(n10208), .A3(n17149), .ZN(n17476) );
  NAND2_X1 U12714 ( .A1(n17503), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17489) );
  NOR2_X1 U12715 ( .A1(n17489), .A2(n17171), .ZN(n17502) );
  NOR2_X1 U12716 ( .A1(n17528), .A2(n17194), .ZN(n17503) );
  AND2_X1 U12717 ( .A1(n17610), .A2(n10209), .ZN(n17544) );
  AND2_X1 U12718 ( .A1(n9771), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n10209) );
  NAND2_X1 U12719 ( .A1(n17610), .A2(n9771), .ZN(n17560) );
  AND2_X1 U12720 ( .A1(n17610), .A2(n10210), .ZN(n17579) );
  NAND2_X1 U12721 ( .A1(n17610), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17591) );
  NOR2_X1 U12722 ( .A1(n17593), .A2(n17270), .ZN(n17610) );
  NOR2_X1 U12723 ( .A1(n16775), .A2(n9836), .ZN(n17635) );
  NAND2_X1 U12724 ( .A1(n9774), .A2(n12479), .ZN(n10212) );
  INV_X1 U12725 ( .A(n16681), .ZN(n17660) );
  AND2_X1 U12726 ( .A1(n17696), .A2(n9779), .ZN(n17677) );
  NAND2_X1 U12727 ( .A1(n17696), .A2(n9776), .ZN(n17684) );
  NAND2_X1 U12728 ( .A1(n17696), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17692) );
  AND2_X1 U12729 ( .A1(n17698), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17696) );
  AND2_X1 U12730 ( .A1(n17744), .A2(n10258), .ZN(n17698) );
  NOR2_X1 U12731 ( .A1(n17749), .A2(n10260), .ZN(n10258) );
  NOR2_X1 U12732 ( .A1(n17861), .A2(n17733), .ZN(n17727) );
  NOR2_X1 U12733 ( .A1(n17749), .A2(n17740), .ZN(n17734) );
  NAND2_X1 U12734 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17734), .ZN(n17733) );
  INV_X1 U12735 ( .A(n17781), .ZN(n10256) );
  INV_X1 U12736 ( .A(n12096), .ZN(n17786) );
  INV_X1 U12737 ( .A(n17810), .ZN(n17804) );
  NOR2_X1 U12738 ( .A1(n17781), .A2(n17780), .ZN(n17813) );
  INV_X1 U12739 ( .A(n17801), .ZN(n17809) );
  CLKBUF_X1 U12740 ( .A(n17850), .Z(n17848) );
  CLKBUF_X1 U12741 ( .A(n17842), .Z(n19255) );
  CLKBUF_X1 U12742 ( .A(n17916), .Z(n17908) );
  OAI211_X1 U12743 ( .C1(n18621), .C2(n19254), .A(n17855), .B(n17854), .ZN(
        n17916) );
  INV_X1 U12745 ( .A(n12639), .ZN(n17362) );
  NAND2_X1 U12746 ( .A1(n18145), .A2(n17041), .ZN(n12588) );
  NOR3_X1 U12747 ( .A1(n18095), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n18354), .ZN(n10075) );
  NAND2_X1 U12748 ( .A1(n18200), .A2(n18362), .ZN(n10073) );
  AND2_X1 U12749 ( .A1(n9773), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10386) );
  NAND2_X1 U12750 ( .A1(n10496), .A2(n10494), .ZN(n18111) );
  NOR2_X1 U12751 ( .A1(n10497), .A2(n18123), .ZN(n10494) );
  INV_X1 U12752 ( .A(n18128), .ZN(n10497) );
  INV_X1 U12753 ( .A(n18145), .ZN(n18140) );
  NAND2_X1 U12754 ( .A1(n18252), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18237) );
  INV_X1 U12755 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18238) );
  INV_X1 U12756 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18275) );
  OR2_X1 U12757 ( .A1(n17005), .A2(n18621), .ZN(n18292) );
  OAI21_X1 U12758 ( .B1(n16854), .B2(n16853), .A(n16852), .ZN(n16892) );
  OR2_X1 U12759 ( .A1(n18581), .A2(n18317), .ZN(n10175) );
  INV_X1 U12760 ( .A(n18315), .ZN(n10174) );
  INV_X1 U12761 ( .A(n18313), .ZN(n10177) );
  NAND2_X1 U12762 ( .A1(n18314), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10178) );
  NOR2_X1 U12763 ( .A1(n19060), .A2(n18462), .ZN(n18587) );
  NAND2_X1 U12764 ( .A1(n16901), .A2(n9770), .ZN(n18115) );
  AND2_X1 U12765 ( .A1(n16688), .A2(n19073), .ZN(n9934) );
  INV_X1 U12766 ( .A(n12088), .ZN(n16688) );
  INV_X1 U12767 ( .A(n18452), .ZN(n18508) );
  INV_X1 U12768 ( .A(n18595), .ZN(n18586) );
  OAI21_X1 U12769 ( .B1(n18232), .B2(n10557), .A(n10554), .ZN(n10559) );
  NOR2_X1 U12770 ( .A1(n18232), .A2(n18234), .ZN(n18233) );
  INV_X1 U12771 ( .A(n10225), .ZN(n18257) );
  NOR2_X1 U12772 ( .A1(n19260), .A2(n18545), .ZN(n18598) );
  INV_X1 U12773 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18613) );
  OR2_X1 U12774 ( .A1(n10338), .A2(n12088), .ZN(n16697) );
  INV_X1 U12775 ( .A(n16687), .ZN(n10338) );
  INV_X1 U12776 ( .A(n19111), .ZN(n10327) );
  AND2_X1 U12777 ( .A1(n12617), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20488)
         );
  CLKBUF_X1 U12779 ( .A(n16995), .Z(n21188) );
  AOI211_X1 U12780 ( .C1(n16722), .C2(n12472), .A(n12471), .B(n12470), .ZN(
        n12473) );
  NAND2_X1 U12781 ( .A1(n12466), .A2(n19322), .ZN(n12474) );
  INV_X1 U12782 ( .A(n11830), .ZN(n11831) );
  NAND2_X1 U12783 ( .A1(n10637), .A2(n12603), .ZN(n12604) );
  NAND2_X1 U12784 ( .A1(n10146), .A2(n16039), .ZN(n16323) );
  OAI21_X1 U12785 ( .B1(n16379), .B2(n19490), .A(n10266), .ZN(P2_U2991) );
  AOI21_X1 U12786 ( .B1(n16376), .B2(n19484), .A(n16101), .ZN(n10266) );
  INV_X1 U12787 ( .A(n12460), .ZN(n9941) );
  OR2_X1 U12788 ( .A1(n16415), .A2(n19490), .ZN(n9942) );
  OAI21_X1 U12789 ( .B1(n16517), .B2(n19490), .A(n10150), .ZN(P2_U3003) );
  INV_X1 U12790 ( .A(n10151), .ZN(n10150) );
  OAI21_X1 U12791 ( .B1(n16504), .B2(n16299), .A(n10152), .ZN(n10151) );
  AOI21_X1 U12792 ( .B1(n16509), .B2(n19493), .A(n16199), .ZN(n10152) );
  NAND2_X1 U12793 ( .A1(n16080), .A2(n16832), .ZN(n11615) );
  OAI21_X1 U12794 ( .B1(n12439), .B2(n16842), .A(n9838), .ZN(P2_U3025) );
  OAI21_X1 U12795 ( .B1(n16415), .B2(n16842), .A(n10286), .ZN(P2_U3027) );
  AOI21_X1 U12796 ( .B1(n10288), .B2(n16832), .A(n10287), .ZN(n10286) );
  NAND2_X1 U12797 ( .A1(n16414), .A2(n16413), .ZN(n10287) );
  INV_X1 U12798 ( .A(n16416), .ZN(n10288) );
  NAND2_X1 U12799 ( .A1(n10467), .A2(n10465), .ZN(P3_U2641) );
  NOR2_X1 U12800 ( .A1(n10466), .A2(n9998), .ZN(n10465) );
  NAND2_X1 U12801 ( .A1(n10468), .A2(n17338), .ZN(n10467) );
  NOR2_X1 U12802 ( .A1(n17051), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10466) );
  NAND2_X1 U12803 ( .A1(n17676), .A2(n17658), .ZN(n10203) );
  NAND2_X1 U12804 ( .A1(n13817), .A2(P3_EBX_REG_28__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U12805 ( .A1(n17452), .A2(n18645), .ZN(n17439) );
  NOR2_X1 U12806 ( .A1(n10213), .A2(n16775), .ZN(n17643) );
  INV_X1 U12807 ( .A(n10215), .ZN(n10213) );
  OR2_X1 U12808 ( .A1(n17666), .A2(n17665), .ZN(n17667) );
  NAND2_X1 U12809 ( .A1(n17744), .A2(n10259), .ZN(n17702) );
  AOI21_X1 U12810 ( .B1(n10006), .B2(n18200), .A(n10005), .ZN(n16877) );
  OR2_X1 U12811 ( .A1(n16876), .A2(n16875), .ZN(n10005) );
  OR3_X1 U12812 ( .A1(n18344), .A2(n18095), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18003) );
  OAI21_X1 U12813 ( .B1(n18032), .B2(n21331), .A(n10071), .ZN(P3_U2808) );
  INV_X1 U12814 ( .A(n9927), .ZN(n18032) );
  NOR3_X1 U12815 ( .A1(n10075), .A2(n10074), .A3(n10072), .ZN(n10071) );
  INV_X1 U12816 ( .A(n18020), .ZN(n10074) );
  NAND2_X1 U12817 ( .A1(n9927), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9926) );
  AND2_X1 U12818 ( .A1(n9932), .A2(n9930), .ZN(n9929) );
  NAND2_X1 U12819 ( .A1(n12138), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12139) );
  INV_X1 U12820 ( .A(n10229), .ZN(n10228) );
  OR2_X1 U12821 ( .A1(n16707), .A2(n16878), .ZN(n10231) );
  NAND2_X1 U12822 ( .A1(n10006), .A2(n18496), .ZN(n10226) );
  NAND2_X1 U12823 ( .A1(n10176), .A2(n10172), .ZN(P3_U2836) );
  AOI21_X1 U12824 ( .B1(n18316), .B2(n18496), .A(n10173), .ZN(n10172) );
  NAND2_X1 U12825 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  NAND2_X1 U12826 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  NAND2_X1 U12827 ( .A1(n19110), .A2(n10326), .ZN(P3_U2996) );
  OAI21_X1 U12828 ( .B1(n10328), .B2(n10327), .A(P3_STATE2_REG_0__SCAN_IN), 
        .ZN(n10326) );
  INV_X1 U12829 ( .A(n10328), .ZN(n19114) );
  NOR2_X1 U12830 ( .A1(n11864), .A2(n19081), .ZN(n12001) );
  NAND2_X1 U12831 ( .A1(n16183), .A2(n11611), .ZN(n11846) );
  INV_X1 U12832 ( .A(n11813), .ZN(n11792) );
  NOR2_X2 U12833 ( .A1(n10246), .A2(n10245), .ZN(n11893) );
  AND2_X1 U12834 ( .A1(n10348), .A2(n16061), .ZN(n9744) );
  INV_X2 U12835 ( .A(n15189), .ZN(n10120) );
  AND2_X1 U12836 ( .A1(n16131), .A2(n11835), .ZN(n9745) );
  NAND2_X1 U12837 ( .A1(n14681), .A2(n14682), .ZN(n14665) );
  AND2_X1 U12838 ( .A1(n13535), .A2(n14381), .ZN(n9746) );
  NAND2_X1 U12839 ( .A1(n12825), .A2(n20532), .ZN(n12897) );
  INV_X1 U12840 ( .A(n12153), .ZN(n10830) );
  OR3_X1 U12841 ( .A1(n11640), .A2(n15674), .A3(n10471), .ZN(n9747) );
  INV_X1 U12842 ( .A(n9721), .ZN(n17533) );
  AND2_X1 U12843 ( .A1(n10156), .A2(n13232), .ZN(n9748) );
  AND2_X1 U12844 ( .A1(n11151), .A2(n16444), .ZN(n11837) );
  INV_X1 U12845 ( .A(n10159), .ZN(n13546) );
  AND2_X1 U12846 ( .A1(n15189), .A2(n9905), .ZN(n9749) );
  NAND2_X1 U12847 ( .A1(n11108), .A2(n9842), .ZN(n9750) );
  NAND2_X1 U12848 ( .A1(n10610), .A2(n10611), .ZN(n14725) );
  NAND2_X1 U12849 ( .A1(n13801), .A2(n12179), .ZN(n13811) );
  OR2_X1 U12850 ( .A1(n11837), .A2(n10364), .ZN(n9751) );
  NAND2_X1 U12851 ( .A1(n13801), .A2(n10594), .ZN(n9752) );
  INV_X1 U12852 ( .A(n11855), .ZN(n11854) );
  AND2_X1 U12853 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11855) );
  OR2_X1 U12854 ( .A1(n10601), .A2(n21033), .ZN(n9753) );
  INV_X1 U12855 ( .A(n12812), .ZN(n12818) );
  BUF_X1 U12856 ( .A(n12818), .Z(n13333) );
  NOR2_X1 U12857 ( .A1(n11783), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9754) );
  AND2_X1 U12858 ( .A1(n10524), .A2(n13053), .ZN(n9755) );
  INV_X1 U12859 ( .A(n11811), .ZN(n10278) );
  AND3_X1 U12860 ( .A1(n10958), .A2(n10949), .A3(n9848), .ZN(n9756) );
  AND2_X1 U12861 ( .A1(n10240), .A2(n18199), .ZN(n9757) );
  AND2_X1 U12862 ( .A1(n9796), .A2(n10576), .ZN(n9758) );
  AND2_X1 U12863 ( .A1(n14614), .A2(n9851), .ZN(n14583) );
  AND2_X1 U12864 ( .A1(n16039), .A2(n16640), .ZN(n9759) );
  AND2_X1 U12865 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n9760) );
  AND4_X1 U12866 ( .A1(n11914), .A2(n11913), .A3(n11912), .A4(n11911), .ZN(
        n9761) );
  AND2_X1 U12867 ( .A1(n11744), .A2(n10093), .ZN(n9762) );
  AND2_X1 U12868 ( .A1(n10632), .A2(n10631), .ZN(n9763) );
  AND2_X1 U12869 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  INV_X1 U12870 ( .A(n11770), .ZN(n10304) );
  AND2_X1 U12871 ( .A1(n10042), .A2(n12925), .ZN(n9764) );
  OAI21_X1 U12872 ( .B1(n15556), .B2(n11792), .A(n11389), .ZN(n16061) );
  AND2_X1 U12873 ( .A1(n9755), .A2(n11468), .ZN(n9765) );
  NOR3_X1 U12874 ( .A1(n15847), .A2(n15846), .A3(n15849), .ZN(n9766) );
  AND2_X1 U12875 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9767) );
  OR2_X1 U12876 ( .A1(n15618), .A2(n9895), .ZN(n9768) );
  AND2_X1 U12877 ( .A1(n9767), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9769) );
  AND2_X1 U12878 ( .A1(n18436), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9770) );
  AND2_X1 U12879 ( .A1(n10210), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n9771) );
  AND2_X1 U12880 ( .A1(n10217), .A2(n10216), .ZN(n9772) );
  AND2_X1 U12881 ( .A1(n9770), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9773) );
  AND2_X1 U12882 ( .A1(n13196), .A2(n12935), .ZN(n13332) );
  AND3_X1 U12883 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(P3_EBX_REG_4__SCAN_IN), .ZN(n9774) );
  AND2_X1 U12884 ( .A1(n9772), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n9775) );
  AND2_X1 U12885 ( .A1(n10264), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9776) );
  AND2_X1 U12886 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n10344), .ZN(
        n9777) );
  AND2_X1 U12887 ( .A1(n10366), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9778) );
  AND2_X1 U12888 ( .A1(n9776), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9779) );
  NOR2_X2 U12889 ( .A1(n13069), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11412) );
  AND2_X2 U12890 ( .A1(n10648), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10872) );
  NOR2_X4 U12891 ( .A1(n16687), .A2(n12088), .ZN(n9780) );
  NAND2_X1 U12892 ( .A1(n13386), .A2(n10601), .ZN(n20489) );
  AND2_X2 U12893 ( .A1(n12265), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10863) );
  NAND2_X1 U12894 ( .A1(n10238), .A2(n10239), .ZN(n18028) );
  INV_X1 U12895 ( .A(n20532), .ZN(n14551) );
  AND2_X1 U12896 ( .A1(n10235), .A2(n10232), .ZN(n9781) );
  BUF_X2 U12897 ( .A(n17597), .Z(n17521) );
  AND4_X1 U12898 ( .A1(n12674), .A2(n12673), .A3(n12672), .A4(n12671), .ZN(
        n9782) );
  INV_X1 U12899 ( .A(n10333), .ZN(n19091) );
  OR3_X1 U12900 ( .A1(n16777), .A2(n16694), .A3(n10334), .ZN(n10333) );
  AND2_X1 U12901 ( .A1(n10929), .A2(n10928), .ZN(n9783) );
  INV_X1 U12902 ( .A(n16094), .ZN(n10350) );
  NAND2_X1 U12903 ( .A1(n10512), .A2(n10511), .ZN(n12440) );
  NOR2_X1 U12904 ( .A1(n15617), .A2(n15618), .ZN(n15613) );
  AND2_X1 U12905 ( .A1(n15859), .A2(n15861), .ZN(n15845) );
  OR2_X1 U12906 ( .A1(n11071), .A2(n10102), .ZN(n11091) );
  NOR2_X1 U12907 ( .A1(n13719), .A2(n13718), .ZN(n13621) );
  NOR2_X1 U12908 ( .A1(n15571), .A2(n11567), .ZN(n11570) );
  BUF_X1 U12909 ( .A(n12888), .Z(n12816) );
  AND2_X1 U12910 ( .A1(n11132), .A2(n10540), .ZN(n11114) );
  NAND2_X1 U12911 ( .A1(n13462), .A2(n13461), .ZN(n13892) );
  NAND2_X1 U12912 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12102), .ZN(
        n9785) );
  NAND2_X1 U12913 ( .A1(n10097), .A2(n11169), .ZN(n11174) );
  NAND2_X1 U12914 ( .A1(n10498), .A2(n10499), .ZN(n11635) );
  NAND2_X1 U12915 ( .A1(n10525), .A2(n10528), .ZN(n13737) );
  NOR2_X1 U12916 ( .A1(n18219), .A2(n12111), .ZN(n12114) );
  AND4_X1 U12917 ( .A1(n12784), .A2(n12783), .A3(n12782), .A4(n12781), .ZN(
        n9786) );
  NAND2_X1 U12918 ( .A1(n11108), .A2(n10094), .ZN(n9787) );
  AND2_X1 U12919 ( .A1(n17696), .A2(n10264), .ZN(n9788) );
  OR2_X1 U12920 ( .A1(n19334), .A2(n11112), .ZN(n11835) );
  NAND2_X1 U12922 ( .A1(n11132), .A2(n11119), .ZN(n9789) );
  NOR2_X1 U12923 ( .A1(n13529), .A2(n13381), .ZN(n9790) );
  AND2_X1 U12924 ( .A1(n16246), .A2(n16235), .ZN(n9791) );
  AND2_X1 U12925 ( .A1(n12452), .A2(n12451), .ZN(n9792) );
  AND2_X1 U12926 ( .A1(n10563), .A2(n13786), .ZN(n9793) );
  AND2_X1 U12927 ( .A1(n11107), .A2(n10538), .ZN(n9794) );
  AND2_X1 U12928 ( .A1(n12412), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9795) );
  AND2_X1 U12929 ( .A1(n10577), .A2(n13569), .ZN(n9796) );
  AND2_X1 U12930 ( .A1(n11168), .A2(n16107), .ZN(n9797) );
  OR2_X1 U12931 ( .A1(n12104), .A2(n9785), .ZN(n9798) );
  AND2_X1 U12932 ( .A1(n12454), .A2(n10569), .ZN(n14531) );
  AND2_X1 U12933 ( .A1(n14681), .A2(n10620), .ZN(n14642) );
  NAND2_X1 U12934 ( .A1(n16045), .A2(n16315), .ZN(n9799) );
  AND2_X1 U12935 ( .A1(n15621), .A2(n11316), .ZN(n12454) );
  NOR2_X1 U12936 ( .A1(n14750), .A2(n14751), .ZN(n14738) );
  OR2_X1 U12937 ( .A1(n15189), .A2(n14422), .ZN(n9800) );
  NOR2_X1 U12938 ( .A1(n18645), .A2(n17815), .ZN(n12035) );
  NAND2_X1 U12939 ( .A1(n10610), .A2(n10609), .ZN(n9801) );
  NAND2_X1 U12940 ( .A1(n11181), .A2(n11180), .ZN(n9802) );
  OR2_X1 U12941 ( .A1(n11630), .A2(n16250), .ZN(n9803) );
  OR2_X1 U12942 ( .A1(n11630), .A2(n10501), .ZN(n9804) );
  NAND2_X1 U12943 ( .A1(n10472), .A2(n11622), .ZN(n9805) );
  NAND2_X1 U12944 ( .A1(n11108), .A2(n9794), .ZN(n9806) );
  AND2_X1 U12945 ( .A1(n11810), .A2(n11809), .ZN(n9807) );
  AND2_X1 U12946 ( .A1(n14531), .A2(n14532), .ZN(n14530) );
  NOR2_X1 U12947 ( .A1(n18645), .A2(n18629), .ZN(n12090) );
  INV_X1 U12948 ( .A(n12090), .ZN(n10317) );
  NAND2_X1 U12949 ( .A1(n17955), .A2(n10221), .ZN(n16704) );
  AND2_X1 U12950 ( .A1(n13392), .A2(n13461), .ZN(n9808) );
  AND2_X1 U12951 ( .A1(n10929), .A2(n10269), .ZN(n9809) );
  INV_X1 U12952 ( .A(n10413), .ZN(n12902) );
  NAND2_X1 U12953 ( .A1(n10034), .A2(n10506), .ZN(n10819) );
  XNOR2_X1 U12954 ( .A(n11796), .B(n11721), .ZN(n12574) );
  AND2_X1 U12955 ( .A1(n10823), .A2(n16835), .ZN(n9810) );
  OR2_X1 U12956 ( .A1(n16321), .A2(n16836), .ZN(n9811) );
  AND4_X1 U12957 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n9812) );
  INV_X4 U12958 ( .A(n11789), .ZN(n19534) );
  INV_X1 U12959 ( .A(n11397), .ZN(n10106) );
  AND2_X1 U12960 ( .A1(n13801), .A2(n10593), .ZN(n9813) );
  NAND2_X1 U12961 ( .A1(n17956), .A2(n18317), .ZN(n17955) );
  AND2_X1 U12962 ( .A1(n16094), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9814) );
  NAND2_X1 U12963 ( .A1(n18075), .A2(n18117), .ZN(n17989) );
  INV_X1 U12964 ( .A(n15124), .ZN(n15197) );
  AND3_X1 U12965 ( .A1(n10294), .A2(n10683), .A3(n10682), .ZN(n9815) );
  AND3_X1 U12966 ( .A1(n10289), .A2(n10681), .A3(n10680), .ZN(n9816) );
  NOR2_X1 U12967 ( .A1(n11846), .A2(n16383), .ZN(n16102) );
  INV_X1 U12968 ( .A(n16102), .ZN(n10268) );
  AND3_X1 U12969 ( .A1(n10959), .A2(n10957), .A3(n10948), .ZN(n9817) );
  AND3_X1 U12970 ( .A1(n19226), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n9818) );
  AND3_X1 U12971 ( .A1(n19234), .A2(n17332), .A3(
        P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n9819) );
  AND2_X1 U12972 ( .A1(n10788), .A2(n10189), .ZN(n9820) );
  INV_X1 U12973 ( .A(n10037), .ZN(n12913) );
  NAND2_X1 U12974 ( .A1(n12888), .A2(n12891), .ZN(n10037) );
  AND2_X1 U12975 ( .A1(n11722), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9821) );
  AND2_X1 U12976 ( .A1(n11846), .A2(n10339), .ZN(n9822) );
  NOR2_X1 U12977 ( .A1(n17042), .A2(n17043), .ZN(n9823) );
  AND2_X1 U12978 ( .A1(n12450), .A2(n16640), .ZN(n9824) );
  INV_X1 U12979 ( .A(n11068), .ZN(n10135) );
  AND3_X1 U12980 ( .A1(n10724), .A2(n11030), .A3(n10723), .ZN(n9825) );
  OR2_X1 U12981 ( .A1(n12172), .A2(n12148), .ZN(n9826) );
  AND2_X1 U12982 ( .A1(n11352), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U12983 ( .A1(n11726), .A2(n10544), .ZN(n9828) );
  AND3_X1 U12984 ( .A1(n16320), .A2(n10070), .A3(n9811), .ZN(n9829) );
  AND2_X1 U12985 ( .A1(n15106), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9830) );
  AND4_X1 U12986 ( .A1(n10381), .A2(n11906), .A3(n11904), .A4(n11905), .ZN(
        n9831) );
  OR2_X1 U12987 ( .A1(n12047), .A2(n12048), .ZN(n9832) );
  AND2_X1 U12988 ( .A1(n11078), .A2(n11073), .ZN(n10536) );
  AND2_X1 U12989 ( .A1(n10136), .A2(n10356), .ZN(n9833) );
  NAND2_X1 U12990 ( .A1(n11069), .A2(n10130), .ZN(n9834) );
  OR2_X1 U12991 ( .A1(n16268), .A2(n11599), .ZN(n9835) );
  OR2_X1 U12992 ( .A1(n10660), .A2(n10212), .ZN(n9836) );
  INV_X1 U12993 ( .A(n11816), .ZN(n10281) );
  OAI21_X1 U12994 ( .B1(n10241), .B2(n18213), .A(n18117), .ZN(n10243) );
  AND2_X1 U12995 ( .A1(n12450), .A2(n19470), .ZN(n9837) );
  INV_X1 U12996 ( .A(n16692), .ZN(n10337) );
  OAI21_X1 U12997 ( .B1(n15516), .B2(n15742), .A(n16041), .ZN(n15502) );
  NAND2_X1 U12998 ( .A1(n12454), .A2(n10573), .ZN(n10575) );
  INV_X1 U12999 ( .A(n13384), .ZN(n10011) );
  OAI22_X1 U13000 ( .A1(n13835), .A2(n13383), .B1(n13382), .B2(n13529), .ZN(
        n13384) );
  AND2_X1 U13001 ( .A1(n12449), .A2(n12448), .ZN(n9838) );
  INV_X1 U13002 ( .A(n17361), .ZN(n10182) );
  INV_X1 U13003 ( .A(n10095), .ZN(n10094) );
  NAND2_X1 U13004 ( .A1(n10537), .A2(n10096), .ZN(n10095) );
  OR2_X1 U13005 ( .A1(n16689), .A2(n16692), .ZN(n9839) );
  AND2_X1 U13006 ( .A1(n20532), .A2(n10415), .ZN(n9840) );
  AND2_X1 U13007 ( .A1(n10404), .A2(n10625), .ZN(n9841) );
  NAND2_X1 U13008 ( .A1(n11108), .A2(n10537), .ZN(n11100) );
  NAND2_X1 U13009 ( .A1(n16064), .A2(n10098), .ZN(n10599) );
  AND2_X1 U13010 ( .A1(n9794), .A2(n11097), .ZN(n9842) );
  OR2_X1 U13011 ( .A1(n9751), .A2(n10361), .ZN(n9843) );
  INV_X1 U13012 ( .A(n10004), .ZN(n18213) );
  OR2_X1 U13013 ( .A1(n18214), .A2(n18504), .ZN(n10004) );
  INV_X1 U13014 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16250) );
  NAND2_X1 U13015 ( .A1(n11726), .A2(n15532), .ZN(n14524) );
  OR2_X2 U13016 ( .A1(n12701), .A2(n12700), .ZN(n12813) );
  AND3_X1 U13017 ( .A1(n11917), .A2(n11916), .A3(n11918), .ZN(n9844) );
  AND2_X1 U13018 ( .A1(n10523), .A2(n11835), .ZN(n9845) );
  INV_X1 U13019 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16282) );
  NAND2_X1 U13020 ( .A1(n10550), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18116) );
  AND3_X1 U13021 ( .A1(n11840), .A2(n16111), .A3(n11148), .ZN(n9846) );
  INV_X1 U13022 ( .A(n15116), .ZN(n10424) );
  AND3_X1 U13023 ( .A1(n11424), .A2(n11429), .A3(n10534), .ZN(n9847) );
  AND2_X1 U13024 ( .A1(n10946), .A2(n10947), .ZN(n9848) );
  NOR2_X2 U13025 ( .A1(n16137), .A2(n16436), .ZN(n16435) );
  AND2_X1 U13026 ( .A1(n17989), .A2(n12125), .ZN(n9849) );
  AND2_X1 U13027 ( .A1(n10499), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9850) );
  AND2_X1 U13028 ( .A1(n10615), .A2(n10613), .ZN(n9851) );
  AND2_X1 U13029 ( .A1(n12946), .A2(n9881), .ZN(n9852) );
  NAND2_X1 U13030 ( .A1(n14681), .A2(n10622), .ZN(n10624) );
  OR2_X1 U13031 ( .A1(n15617), .A2(n9768), .ZN(n9853) );
  AND2_X1 U13032 ( .A1(n9793), .A2(n10562), .ZN(n9854) );
  AND2_X1 U13033 ( .A1(n10362), .A2(n10361), .ZN(n9855) );
  AND2_X1 U13034 ( .A1(n9800), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9856) );
  INV_X1 U13035 ( .A(n10277), .ZN(n10276) );
  AOI21_X1 U13036 ( .B1(n10279), .B2(n10280), .A(n10278), .ZN(n10277) );
  AND2_X1 U13037 ( .A1(n11853), .A2(n11852), .ZN(n9857) );
  OR2_X1 U13038 ( .A1(n16046), .A2(n10439), .ZN(n9858) );
  AND2_X1 U13039 ( .A1(n9800), .A2(n10162), .ZN(n9859) );
  AND2_X1 U13040 ( .A1(n10487), .A2(n10488), .ZN(n9860) );
  NOR2_X1 U13041 ( .A1(n10355), .A2(n10354), .ZN(n10353) );
  AND2_X1 U13042 ( .A1(n10312), .A2(n10273), .ZN(n9861) );
  INV_X1 U13043 ( .A(n10518), .ZN(n10517) );
  NAND2_X1 U13044 ( .A1(n16139), .A2(n16146), .ZN(n10518) );
  INV_X1 U13045 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10679) );
  OR2_X1 U13046 ( .A1(n20532), .A2(n13022), .ZN(n9862) );
  INV_X1 U13047 ( .A(n13323), .ZN(n10018) );
  INV_X1 U13048 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U13049 ( .A1(n11220), .A2(n11742), .ZN(n11573) );
  NAND2_X1 U13050 ( .A1(n11438), .A2(n11437), .ZN(n13054) );
  AND2_X1 U13051 ( .A1(n17156), .A2(n10643), .ZN(n12635) );
  NOR2_X2 U13052 ( .A1(n11577), .A2(n20217), .ZN(n16832) );
  NAND2_X1 U13053 ( .A1(n13491), .A2(n12177), .ZN(n13742) );
  AND2_X1 U13054 ( .A1(n17452), .A2(n9772), .ZN(n9863) );
  NAND2_X1 U13055 ( .A1(n13497), .A2(n13569), .ZN(n13568) );
  OR3_X1 U13056 ( .A1(n11640), .A2(n15674), .A3(n10470), .ZN(n9864) );
  NAND2_X1 U13057 ( .A1(n13760), .A2(n11286), .ZN(n9865) );
  NOR3_X1 U13058 ( .A1(n17489), .A2(n10208), .A3(n10206), .ZN(n10205) );
  NAND2_X1 U13059 ( .A1(n17452), .A2(n10217), .ZN(n10218) );
  NAND2_X1 U13060 ( .A1(n11644), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9866) );
  NAND2_X1 U13061 ( .A1(n13054), .A2(n9755), .ZN(n9867) );
  OR2_X1 U13062 ( .A1(n11640), .A2(n15674), .ZN(n9868) );
  AND2_X1 U13063 ( .A1(n14302), .A2(n10455), .ZN(n9869) );
  AND2_X1 U13064 ( .A1(n10446), .A2(n14770), .ZN(n9870) );
  AND2_X1 U13065 ( .A1(n9869), .A2(n10454), .ZN(n9871) );
  AND2_X1 U13066 ( .A1(n12300), .A2(n15861), .ZN(n9872) );
  NAND2_X1 U13067 ( .A1(n11644), .A2(n9767), .ZN(n11651) );
  NAND2_X1 U13068 ( .A1(n11671), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11674) );
  AND2_X1 U13069 ( .A1(n10459), .A2(n10458), .ZN(n9873) );
  INV_X1 U13070 ( .A(n10532), .ZN(n12938) );
  AND2_X1 U13071 ( .A1(n13499), .A2(n13498), .ZN(n13497) );
  NOR2_X1 U13072 ( .A1(n17951), .A2(n17952), .ZN(n12629) );
  NOR2_X1 U13073 ( .A1(n13590), .A2(n13565), .ZN(n14256) );
  AND4_X1 U13074 ( .A1(n14766), .A2(n14769), .A3(n14781), .A4(n13985), .ZN(
        n9874) );
  AND2_X1 U13075 ( .A1(n17156), .A2(n10502), .ZN(n12628) );
  NAND2_X1 U13076 ( .A1(n11425), .A2(n10535), .ZN(n15744) );
  AND2_X1 U13077 ( .A1(n12177), .A2(n13744), .ZN(n9875) );
  AND2_X1 U13078 ( .A1(n10643), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9876) );
  INV_X1 U13079 ( .A(n13536), .ZN(n10014) );
  NAND2_X1 U13080 ( .A1(n11425), .A2(n11424), .ZN(n15756) );
  AND2_X1 U13081 ( .A1(n14376), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9877) );
  AND2_X1 U13082 ( .A1(n15189), .A2(n15318), .ZN(n9878) );
  AND2_X1 U13083 ( .A1(n10461), .A2(n17362), .ZN(n9879) );
  OR2_X1 U13084 ( .A1(n18319), .A2(n18305), .ZN(n9880) );
  NAND2_X1 U13085 ( .A1(n12931), .A2(n20501), .ZN(n9881) );
  INV_X1 U13086 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10500) );
  NAND2_X1 U13087 ( .A1(n20532), .A2(n12819), .ZN(n13208) );
  NAND2_X1 U13088 ( .A1(n12933), .A2(n12932), .ZN(n20648) );
  AND2_X1 U13089 ( .A1(n13797), .A2(n11301), .ZN(n13808) );
  NOR2_X2 U13090 ( .A1(n12819), .A2(n13022), .ZN(n13984) );
  AND2_X1 U13091 ( .A1(n10593), .A2(n15891), .ZN(n9882) );
  AND2_X1 U13092 ( .A1(n9870), .A2(n10445), .ZN(n9883) );
  INV_X1 U13093 ( .A(n12862), .ZN(n12863) );
  NAND2_X1 U13094 ( .A1(n12797), .A2(n20506), .ZN(n14866) );
  AND2_X1 U13095 ( .A1(n17744), .A2(n10261), .ZN(n9884) );
  NAND2_X1 U13096 ( .A1(n10781), .A2(n10309), .ZN(n9885) );
  OR2_X1 U13097 ( .A1(n11071), .A2(n11070), .ZN(n10104) );
  INV_X1 U13098 ( .A(n10207), .ZN(n17487) );
  NOR2_X1 U13099 ( .A1(n17489), .A2(n10208), .ZN(n10207) );
  OR2_X1 U13100 ( .A1(n18117), .A2(n18301), .ZN(n9886) );
  INV_X2 U13101 ( .A(n14416), .ZN(n14409) );
  INV_X1 U13102 ( .A(n10368), .ZN(n20608) );
  AND2_X1 U13103 ( .A1(n13542), .A2(n13561), .ZN(n9887) );
  AND2_X1 U13104 ( .A1(n9872), .A2(n15870), .ZN(n9888) );
  AND2_X1 U13105 ( .A1(n9871), .A2(n10453), .ZN(n9889) );
  AND2_X1 U13106 ( .A1(n9769), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9890) );
  AND2_X1 U13107 ( .A1(n10463), .A2(n10464), .ZN(n9891) );
  AND2_X1 U13108 ( .A1(n9872), .A2(n10591), .ZN(n9892) );
  AND2_X1 U13109 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n9893) );
  INV_X1 U13110 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10560) );
  NOR2_X1 U13111 ( .A1(n10660), .A2(n17611), .ZN(n10215) );
  INV_X1 U13112 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n9973) );
  AND2_X1 U13113 ( .A1(n12592), .A2(n10480), .ZN(n9894) );
  INV_X1 U13114 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10596) );
  OR2_X1 U13115 ( .A1(n10943), .A2(n10942), .ZN(n11592) );
  NAND2_X1 U13116 ( .A1(n12592), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12591) );
  INV_X1 U13117 ( .A(n19081), .ZN(n11865) );
  AND2_X1 U13118 ( .A1(n11556), .A2(n11555), .ZN(n9895) );
  NAND2_X1 U13119 ( .A1(n13239), .A2(n13238), .ZN(n13545) );
  INV_X1 U13120 ( .A(n13545), .ZN(n10052) );
  AND2_X1 U13121 ( .A1(n14256), .A2(n16813), .ZN(n9896) );
  NOR2_X1 U13122 ( .A1(n18265), .A2(n12100), .ZN(n9897) );
  AND2_X1 U13123 ( .A1(n10215), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n9898) );
  INV_X1 U13124 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10470) );
  OR2_X1 U13125 ( .A1(n17660), .A2(n17386), .ZN(n9899) );
  OR2_X1 U13126 ( .A1(n10179), .A2(n18296), .ZN(n9900) );
  AND2_X1 U13127 ( .A1(n14038), .A2(n14037), .ZN(n9901) );
  OR2_X1 U13128 ( .A1(n13439), .A2(n10425), .ZN(n9902) );
  AND2_X1 U13129 ( .A1(n12121), .A2(n10639), .ZN(n9903) );
  NAND2_X1 U13130 ( .A1(n18359), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9904) );
  OR2_X1 U13131 ( .A1(n15170), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9905) );
  AND2_X1 U13132 ( .A1(n10489), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9906) );
  NAND2_X1 U13133 ( .A1(n12953), .A2(n13021), .ZN(n13331) );
  INV_X1 U13134 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21091) );
  AND2_X1 U13135 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .ZN(n9907) );
  INV_X1 U13136 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10595) );
  NOR2_X1 U13137 ( .A1(n17139), .A2(n18072), .ZN(n17156) );
  INV_X1 U13138 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10490) );
  INV_X1 U13139 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10096) );
  INV_X1 U13140 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n9995) );
  INV_X1 U13141 ( .A(n15024), .ZN(n10164) );
  AND4_X1 U13142 ( .A1(n16344), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9908) );
  INV_X1 U13143 ( .A(n19258), .ZN(n19102) );
  NOR2_X1 U13144 ( .A1(n19105), .A2(n19273), .ZN(n19258) );
  AND2_X1 U13145 ( .A1(n11611), .A2(n9908), .ZN(n9909) );
  OR2_X1 U13146 ( .A1(n21468), .A2(n16371), .ZN(n9910) );
  NAND2_X1 U13147 ( .A1(n11702), .A2(n16315), .ZN(n9911) );
  AND2_X1 U13148 ( .A1(n10585), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9912) );
  AND2_X1 U13149 ( .A1(n15318), .A2(n14403), .ZN(n9913) );
  INV_X1 U13150 ( .A(n10260), .ZN(n10259) );
  NAND2_X1 U13151 ( .A1(n10261), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n10260) );
  OR2_X1 U13152 ( .A1(n15088), .A2(n14401), .ZN(n9914) );
  AND2_X1 U13153 ( .A1(n9912), .A2(n11844), .ZN(n9915) );
  AND2_X1 U13154 ( .A1(n9913), .A2(n14402), .ZN(n9916) );
  NAND2_X1 U13155 ( .A1(n14853), .A2(n14414), .ZN(n10602) );
  AND2_X1 U13156 ( .A1(n10495), .A2(n10496), .ZN(n9917) );
  INV_X1 U13157 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10482) );
  INV_X1 U13158 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10481) );
  INV_X1 U13159 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10483) );
  INV_X1 U13160 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n9996) );
  OR2_X1 U13161 ( .A1(n15024), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9918) );
  AND2_X1 U13162 ( .A1(n16395), .A2(n10585), .ZN(n9919) );
  INV_X1 U13163 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n9997) );
  NOR2_X1 U13164 ( .A1(n19255), .A2(n17832), .ZN(n17850) );
  INV_X1 U13165 ( .A(n21072), .ZN(n9920) );
  INV_X1 U13166 ( .A(n9920), .ZN(n9921) );
  INV_X1 U13167 ( .A(n20977), .ZN(n9922) );
  INV_X1 U13168 ( .A(n9922), .ZN(n9923) );
  INV_X1 U13169 ( .A(n21078), .ZN(n9924) );
  INV_X1 U13170 ( .A(n9924), .ZN(n9925) );
  AOI22_X2 U13171 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20486), .B1(DATAI_22_), 
        .B2(n20531), .ZN(n21016) );
  AOI22_X2 U13172 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20486), .B1(DATAI_16_), 
        .B2(n20531), .ZN(n21041) );
  AOI22_X2 U13173 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20486), .B1(DATAI_28_), 
        .B2(n20531), .ZN(n21065) );
  AOI22_X2 U13174 ( .A1(DATAI_19_), .A2(n20531), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20486), .ZN(n21059) );
  AOI22_X2 U13175 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20486), .B1(DATAI_26_), 
        .B2(n20531), .ZN(n21053) );
  AOI22_X2 U13176 ( .A1(DATAI_31_), .A2(n20531), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20486), .ZN(n21089) );
  NAND2_X1 U13177 ( .A1(n18905), .A2(n18964), .ZN(n18639) );
  AOI22_X2 U13178 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19546), .ZN(n19996) );
  NOR2_X2 U13179 ( .A1(n19499), .A2(n19498), .ZN(n19546) );
  AOI22_X2 U13180 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20486), .B1(DATAI_25_), 
        .B2(n20531), .ZN(n21047) );
  NAND3_X1 U13181 ( .A1(n18033), .A2(n9929), .A3(n9926), .ZN(P3_U2809) );
  AOI22_X1 U13182 ( .A1(n11970), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9721), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9933) );
  NOR2_X2 U13183 ( .A1(n10318), .A2(n11984), .ZN(n18640) );
  NOR2_X4 U13184 ( .A1(n19072), .A2(n9934), .ZN(n19064) );
  NAND2_X1 U13185 ( .A1(n12092), .A2(n12091), .ZN(n19072) );
  INV_X2 U13186 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17332) );
  AND2_X2 U13187 ( .A1(n10824), .A2(n9810), .ZN(n19654) );
  NOR2_X1 U13188 ( .A1(n16125), .A2(n9936), .ZN(n16417) );
  NAND3_X1 U13189 ( .A1(n9937), .A2(n11593), .A3(n10580), .ZN(n16296) );
  NAND2_X1 U13190 ( .A1(n9937), .A2(n11593), .ZN(n9945) );
  NAND2_X1 U13191 ( .A1(n9942), .A2(n9941), .ZN(P2_U2995) );
  INV_X1 U13192 ( .A(n9944), .ZN(n14550) );
  NAND2_X1 U13193 ( .A1(n9945), .A2(n16295), .ZN(n16615) );
  OAI21_X1 U13194 ( .B1(n9945), .B2(n11813), .A(n15775), .ZN(n16275) );
  NAND3_X1 U13195 ( .A1(n10811), .A2(n10819), .A3(n10810), .ZN(n9946) );
  XNOR2_X2 U13196 ( .A(n10432), .B(n9947), .ZN(n12164) );
  NAND2_X1 U13197 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  NAND2_X1 U13198 ( .A1(n10814), .A2(n10813), .ZN(n9948) );
  NAND2_X2 U13199 ( .A1(n9951), .A2(n9950), .ZN(n16213) );
  AOI21_X2 U13200 ( .B1(n16227), .B2(n11089), .A(n11088), .ZN(n9950) );
  NAND2_X2 U13201 ( .A1(n10129), .A2(n19357), .ZN(n16227) );
  NAND3_X1 U13202 ( .A1(n9952), .A2(n10131), .A3(n10132), .ZN(n9951) );
  NAND2_X1 U13203 ( .A1(n10161), .A2(n10165), .ZN(n15017) );
  NAND4_X1 U13204 ( .A1(n9957), .A2(n9956), .A3(n14407), .A4(n9955), .ZN(
        n14408) );
  NAND3_X1 U13205 ( .A1(n10161), .A2(n10165), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9955) );
  OR2_X1 U13206 ( .A1(n10165), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9956) );
  NAND2_X1 U13207 ( .A1(n9963), .A2(n13094), .ZN(n9962) );
  AOI21_X2 U13208 ( .B1(n15462), .B2(n14376), .A(n9746), .ZN(n13593) );
  NAND2_X1 U13209 ( .A1(n9966), .A2(n13576), .ZN(n9975) );
  AND2_X1 U13210 ( .A1(n13574), .A2(n14376), .ZN(n9966) );
  INV_X1 U13211 ( .A(n13593), .ZN(n13543) );
  NAND2_X1 U13212 ( .A1(n9968), .A2(n13548), .ZN(n20423) );
  NAND2_X1 U13213 ( .A1(n9975), .A2(n9887), .ZN(n9969) );
  NAND2_X1 U13214 ( .A1(n13593), .A2(n9973), .ZN(n9970) );
  INV_X1 U13215 ( .A(n11602), .ZN(n9976) );
  INV_X1 U13216 ( .A(n11598), .ZN(n10105) );
  NAND2_X2 U13217 ( .A1(n9978), .A2(n9977), .ZN(n11598) );
  NAND2_X2 U13218 ( .A1(n9979), .A2(n9981), .ZN(n10601) );
  NAND4_X1 U13219 ( .A1(n10664), .A2(n14839), .A3(n9987), .A4(n13892), .ZN(
        n14765) );
  INV_X1 U13220 ( .A(n14765), .ZN(n13986) );
  NAND2_X2 U13221 ( .A1(n9989), .A2(n14584), .ZN(n15028) );
  AND3_X2 U13222 ( .A1(n9993), .A2(n9992), .A3(n9990), .ZN(n10782) );
  NOR2_X2 U13223 ( .A1(n17039), .A2(n17365), .ZN(n17044) );
  NAND3_X1 U13224 ( .A1(n10169), .A2(n10558), .A3(n18243), .ZN(n10168) );
  AND2_X2 U13225 ( .A1(n10651), .A2(n9831), .ZN(n17800) );
  NAND2_X2 U13226 ( .A1(n10550), .A2(n10549), .ZN(n18090) );
  AND2_X2 U13227 ( .A1(n10425), .A2(n12958), .ZN(n12994) );
  AND2_X2 U13228 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12958) );
  AND2_X2 U13229 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10425) );
  AND2_X2 U13230 ( .A1(n12664), .A2(n13441), .ZN(n14235) );
  NAND2_X2 U13232 ( .A1(n13323), .A2(n12892), .ZN(n12862) );
  XNOR2_X1 U13233 ( .A(n14366), .B(n13837), .ZN(n14375) );
  XNOR2_X2 U13234 ( .A(n12948), .B(n20648), .ZN(n13463) );
  INV_X1 U13235 ( .A(n10402), .ZN(n12923) );
  AND2_X2 U13236 ( .A1(n10626), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15061) );
  NAND2_X2 U13237 ( .A1(n14404), .A2(n15210), .ZN(n10626) );
  NAND2_X2 U13238 ( .A1(n10021), .A2(n10369), .ZN(n14404) );
  NAND2_X2 U13239 ( .A1(n10022), .A2(n10041), .ZN(n12948) );
  NAND2_X2 U13240 ( .A1(n10368), .A2(n10427), .ZN(n13097) );
  NAND3_X2 U13241 ( .A1(n10367), .A2(n10398), .A3(n10397), .ZN(n10368) );
  NAND3_X1 U13242 ( .A1(n10027), .A2(n20229), .A3(n10023), .ZN(n11357) );
  NAND2_X1 U13243 ( .A1(n10028), .A2(n16592), .ZN(n10584) );
  XNOR2_X1 U13244 ( .A(n10582), .B(n16592), .ZN(n16279) );
  NAND2_X1 U13245 ( .A1(n10036), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10032) );
  NAND3_X1 U13246 ( .A1(n10053), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10055), 
        .ZN(n10033) );
  NAND2_X2 U13247 ( .A1(n10197), .A2(n10196), .ZN(n10036) );
  INV_X1 U13248 ( .A(n10036), .ZN(n10801) );
  NAND2_X1 U13249 ( .A1(n10036), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10773) );
  NAND2_X2 U13250 ( .A1(n14364), .A2(n14363), .ZN(n16799) );
  NAND2_X1 U13251 ( .A1(n13550), .A2(n13551), .ZN(n14364) );
  AND4_X4 U13252 ( .A1(n10040), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12775) );
  XNOR2_X2 U13253 ( .A(n10601), .B(n20750), .ZN(n15462) );
  INV_X1 U13254 ( .A(n15078), .ZN(n10046) );
  AOI21_X1 U13255 ( .B1(n10046), .B2(n15259), .A(n14441), .ZN(n10045) );
  NAND2_X1 U13256 ( .A1(n15023), .A2(n15259), .ZN(n10167) );
  NAND2_X2 U13257 ( .A1(n14404), .A2(n15078), .ZN(n15023) );
  NAND3_X1 U13258 ( .A1(n12758), .A2(n12754), .A3(n12755), .ZN(n10049) );
  NAND2_X1 U13259 ( .A1(n13418), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13544) );
  XNOR2_X1 U13260 ( .A(n13545), .B(n10159), .ZN(n13418) );
  OAI21_X1 U13261 ( .B1(n15023), .B2(n10163), .A(n9859), .ZN(n10161) );
  NAND4_X1 U13262 ( .A1(n9861), .A2(n11357), .A3(n13632), .A4(n10311), .ZN(
        n10053) );
  NAND3_X1 U13263 ( .A1(n10775), .A2(n13685), .A3(n10774), .ZN(n10054) );
  AND2_X2 U13264 ( .A1(n10123), .A2(n10768), .ZN(n11574) );
  NAND2_X1 U13265 ( .A1(n10056), .A2(n11792), .ZN(n10134) );
  OAI21_X1 U13266 ( .B1(n10057), .B2(n20253), .A(n15032), .ZN(P1_U2971) );
  OAI21_X1 U13267 ( .B1(n10057), .B2(n15456), .A(n15249), .ZN(P1_U3003) );
  OAI211_X1 U13268 ( .C1(n19490), .C2(n16323), .A(n10058), .B(n16049), .ZN(
        P2_U2986) );
  NAND2_X1 U13269 ( .A1(n10059), .A2(n19484), .ZN(n10058) );
  NAND2_X1 U13270 ( .A1(n10438), .A2(n10435), .ZN(n10059) );
  NAND3_X1 U13271 ( .A1(n10062), .A2(n12038), .A3(n12035), .ZN(n10063) );
  NAND2_X1 U13272 ( .A1(n10063), .A2(n16690), .ZN(n10314) );
  INV_X1 U13273 ( .A(n10063), .ZN(n12075) );
  NAND2_X1 U13274 ( .A1(n13765), .A2(n13063), .ZN(n19405) );
  NAND3_X1 U13275 ( .A1(n18021), .A2(n18363), .A3(n10073), .ZN(n10072) );
  NAND2_X2 U13276 ( .A1(n9812), .A2(n10076), .ZN(n17815) );
  NAND3_X1 U13277 ( .A1(n12012), .A2(n12013), .A3(n10078), .ZN(n10077) );
  INV_X1 U13278 ( .A(n9783), .ZN(n10083) );
  NAND3_X1 U13279 ( .A1(n10274), .A2(n10087), .A3(n10084), .ZN(n12567) );
  OAI21_X1 U13280 ( .B1(n10600), .B2(n10276), .A(n10085), .ZN(n10084) );
  CLKBUF_X1 U13281 ( .A(n10935), .Z(n10089) );
  INV_X1 U13282 ( .A(n10104), .ZN(n11077) );
  NOR2_X2 U13283 ( .A1(n10779), .A2(n10149), .ZN(n13697) );
  NAND2_X2 U13284 ( .A1(n10106), .A2(n12141), .ZN(n10149) );
  XNOR2_X2 U13285 ( .A(n10112), .B(n10809), .ZN(n10823) );
  NOR2_X1 U13286 ( .A1(n10112), .A2(n11258), .ZN(n13499) );
  NAND2_X1 U13287 ( .A1(n16493), .A2(n9824), .ZN(n16502) );
  NAND2_X1 U13288 ( .A1(n16493), .A2(n9837), .ZN(n16188) );
  OAI21_X1 U13289 ( .B1(n12439), .B2(n19490), .A(n9857), .ZN(P2_U2993) );
  NAND2_X2 U13290 ( .A1(n10115), .A2(n15189), .ZN(n15078) );
  NAND2_X1 U13291 ( .A1(n15124), .A2(n10116), .ZN(n10371) );
  AND2_X1 U13292 ( .A1(n14395), .A2(n14398), .ZN(n10116) );
  NAND2_X2 U13293 ( .A1(n15124), .A2(n14395), .ZN(n14397) );
  NAND3_X1 U13294 ( .A1(n13386), .A2(n14376), .A3(n10601), .ZN(n10117) );
  OAI211_X1 U13295 ( .C1(n20489), .C2(n13874), .A(n13391), .B(n13390), .ZN(
        n13392) );
  XNOR2_X2 U13296 ( .A(n11598), .B(n11599), .ZN(n11596) );
  AOI21_X1 U13297 ( .B1(n16225), .B2(n16593), .A(n11081), .ZN(n10132) );
  AND2_X2 U13298 ( .A1(n10305), .A2(n10896), .ZN(n10930) );
  NAND2_X1 U13299 ( .A1(n9759), .A2(n10146), .ZN(n10145) );
  INV_X1 U13300 ( .A(n10438), .ZN(n10143) );
  NAND2_X1 U13301 ( .A1(n10143), .A2(n16832), .ZN(n10144) );
  NAND4_X1 U13302 ( .A1(n10434), .A2(n10145), .A3(n10144), .A4(n9829), .ZN(
        P2_U3018) );
  INV_X1 U13303 ( .A(n16055), .ZN(n10147) );
  NAND2_X1 U13304 ( .A1(n16183), .A2(n9909), .ZN(n16055) );
  NAND3_X1 U13305 ( .A1(n10149), .A2(n19529), .A3(n11212), .ZN(n11218) );
  OAI22_X1 U13306 ( .A1(n10762), .A2(n10783), .B1(n13685), .B2(n10149), .ZN(
        n10768) );
  AND2_X4 U13307 ( .A1(n10153), .A2(n10425), .ZN(n14475) );
  AND2_X2 U13308 ( .A1(n12662), .A2(n10153), .ZN(n14483) );
  NAND3_X1 U13309 ( .A1(n15171), .A2(n15175), .A3(n15173), .ZN(n15160) );
  NAND2_X1 U13310 ( .A1(n13020), .A2(n21091), .ZN(n10155) );
  XNOR2_X2 U13311 ( .A(n12988), .B(n12987), .ZN(n13020) );
  NAND2_X1 U13312 ( .A1(n20541), .A2(n13097), .ZN(n14871) );
  NAND3_X1 U13313 ( .A1(n14404), .A2(n15078), .A3(n10164), .ZN(n10160) );
  INV_X1 U13314 ( .A(n12107), .ZN(n10170) );
  INV_X1 U13315 ( .A(n10558), .ZN(n18220) );
  INV_X1 U13316 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10171) );
  NOR2_X2 U13317 ( .A1(n18109), .A2(n18423), .ZN(n18352) );
  INV_X1 U13318 ( .A(n12101), .ZN(n10180) );
  NAND2_X1 U13319 ( .A1(n16183), .A2(n9915), .ZN(n16137) );
  NAND3_X2 U13320 ( .A1(n10192), .A2(n11607), .A3(n10191), .ZN(n16183) );
  NAND3_X1 U13321 ( .A1(n10816), .A2(n10813), .A3(n10818), .ZN(n10183) );
  NAND2_X1 U13322 ( .A1(n10185), .A2(n16213), .ZN(n10186) );
  NAND2_X1 U13323 ( .A1(n16213), .A2(n10444), .ZN(n10597) );
  NAND2_X2 U13324 ( .A1(n10597), .A2(n9797), .ZN(n16106) );
  INV_X1 U13325 ( .A(n13067), .ZN(n11363) );
  INV_X2 U13326 ( .A(n12164), .ZN(n19479) );
  NAND3_X1 U13327 ( .A1(n16243), .A2(n16235), .A3(n11600), .ZN(n10192) );
  OAI211_X2 U13328 ( .C1(n11601), .C2(n10194), .A(n10193), .B(n9835), .ZN(
        n16243) );
  INV_X1 U13329 ( .A(n11596), .ZN(n10194) );
  CLKBUF_X1 U13330 ( .A(n13697), .Z(n10202) );
  INV_X1 U13331 ( .A(n10202), .ZN(n10309) );
  NOR2_X1 U13332 ( .A1(n13697), .A2(n20229), .ZN(n10310) );
  NAND2_X1 U13333 ( .A1(n12924), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10399) );
  NAND2_X1 U13334 ( .A1(n10582), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10581) );
  NAND2_X2 U13335 ( .A1(n15209), .A2(n14394), .ZN(n15124) );
  INV_X1 U13336 ( .A(n13100), .ZN(n10389) );
  OAI211_X2 U13337 ( .C1(n10764), .C2(n12411), .A(n11220), .B(n11742), .ZN(
        n10787) );
  NAND2_X1 U13338 ( .A1(n10583), .A2(n10581), .ZN(n16265) );
  NAND3_X1 U13339 ( .A1(n13819), .A2(n10204), .A3(n10203), .ZN(P3_U2675) );
  INV_X1 U13340 ( .A(n10205), .ZN(n17440) );
  NOR2_X1 U13341 ( .A1(n16775), .A2(n10660), .ZN(n17655) );
  INV_X1 U13342 ( .A(n10218), .ZN(n17423) );
  NAND2_X1 U13343 ( .A1(n12127), .A2(n18199), .ZN(n17971) );
  NAND2_X1 U13345 ( .A1(n12127), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10222) );
  OAI21_X1 U13346 ( .B1(n18267), .B2(n18266), .A(n10224), .ZN(n10223) );
  NAND3_X1 U13347 ( .A1(n10231), .A2(n10228), .A3(n10226), .ZN(P3_U2833) );
  INV_X1 U13348 ( .A(n10233), .ZN(n10232) );
  OAI21_X1 U13349 ( .B1(n17333), .B2(n17654), .A(n10234), .ZN(n10233) );
  NAND2_X1 U13350 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10235) );
  NAND2_X1 U13351 ( .A1(n18076), .A2(n10239), .ZN(n10237) );
  INV_X1 U13352 ( .A(n10243), .ZN(n18089) );
  NAND2_X1 U13353 ( .A1(n11964), .A2(n10247), .ZN(n10248) );
  NAND4_X1 U13354 ( .A1(n10257), .A2(n10256), .A3(n9907), .A4(
        P3_EAX_REG_2__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U13355 ( .A1(n17744), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17740) );
  INV_X1 U13356 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n10263) );
  OAI21_X1 U13357 ( .B1(n15257), .B2(n20253), .A(n15041), .ZN(P1_U2972) );
  NAND2_X1 U13358 ( .A1(n10265), .A2(n14398), .ZN(n10631) );
  NOR2_X1 U13359 ( .A1(n14392), .A2(n14396), .ZN(n10265) );
  OAI21_X1 U13360 ( .B1(n10600), .B2(n10280), .A(n10279), .ZN(n11812) );
  NAND2_X1 U13361 ( .A1(n10277), .A2(n10275), .ZN(n10274) );
  NAND4_X1 U13362 ( .A1(n10720), .A2(n10666), .A3(n10721), .A4(n10722), .ZN(
        n10282) );
  NAND3_X1 U13363 ( .A1(n9825), .A2(n10725), .A3(n10726), .ZN(n10283) );
  NAND4_X1 U13364 ( .A1(n10734), .A2(n10658), .A3(n10735), .A4(n10736), .ZN(
        n10284) );
  NAND3_X1 U13365 ( .A1(n10293), .A2(n11030), .A3(n10292), .ZN(n10291) );
  NAND3_X1 U13366 ( .A1(n10298), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10297), .ZN(n10296) );
  NAND2_X1 U13367 ( .A1(n10299), .A2(n10302), .ZN(n16066) );
  OR2_X1 U13368 ( .A1(n16106), .A2(n10304), .ZN(n10299) );
  NAND2_X2 U13369 ( .A1(n10301), .A2(n10300), .ZN(n16044) );
  NAND2_X1 U13370 ( .A1(n16106), .A2(n10302), .ZN(n10301) );
  NAND4_X1 U13371 ( .A1(n10848), .A2(n10849), .A3(n10846), .A4(n10847), .ZN(
        n10305) );
  INV_X1 U13372 ( .A(n11592), .ZN(n10306) );
  NAND2_X1 U13373 ( .A1(n16053), .A2(n10308), .ZN(n10307) );
  INV_X1 U13374 ( .A(n10832), .ZN(n10829) );
  XNOR2_X2 U13375 ( .A(n16044), .B(n16045), .ZN(n16053) );
  INV_X1 U13376 ( .A(n10314), .ZN(n17004) );
  NOR2_X1 U13377 ( .A1(n10317), .A2(n10316), .ZN(n10315) );
  NAND3_X1 U13378 ( .A1(n11982), .A2(n10324), .A3(n10319), .ZN(n10318) );
  NAND3_X1 U13379 ( .A1(n11983), .A2(n10322), .A3(n10321), .ZN(n10320) );
  NAND3_X1 U13380 ( .A1(n19100), .A2(n19101), .A3(n10331), .ZN(n19109) );
  INV_X1 U13381 ( .A(n16695), .ZN(n10335) );
  INV_X1 U13382 ( .A(n11846), .ZN(n10343) );
  NAND2_X1 U13383 ( .A1(n10345), .A2(n10346), .ZN(n16065) );
  OAI21_X1 U13384 ( .B1(n16095), .B2(n10353), .A(n10348), .ZN(n16062) );
  AOI21_X1 U13385 ( .B1(n16095), .B2(n16094), .A(n11179), .ZN(n16088) );
  NAND2_X1 U13386 ( .A1(n10523), .A2(n9855), .ZN(n10360) );
  AOI21_X1 U13387 ( .B1(n10523), .B2(n9745), .A(n11837), .ZN(n16123) );
  OR2_X2 U13388 ( .A1(n10399), .A2(n12923), .ZN(n10367) );
  OAI21_X1 U13389 ( .B1(n10629), .B2(n15189), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10370) );
  NAND2_X1 U13390 ( .A1(n10395), .A2(n14374), .ZN(n16791) );
  NAND2_X1 U13391 ( .A1(n10377), .A2(n16792), .ZN(n10376) );
  NAND2_X1 U13392 ( .A1(n10380), .A2(n16792), .ZN(n15218) );
  NAND2_X1 U13393 ( .A1(n16791), .A2(n16793), .ZN(n10380) );
  AND2_X2 U13394 ( .A1(n15124), .A2(n10396), .ZN(n15199) );
  NAND3_X1 U13395 ( .A1(n12923), .A2(n10399), .A3(n12906), .ZN(n10397) );
  NAND3_X1 U13396 ( .A1(n13895), .A2(n10627), .A3(n14376), .ZN(n10410) );
  NAND4_X1 U13397 ( .A1(n13196), .A2(n10411), .A3(n12935), .A4(n13331), .ZN(
        n12903) );
  INV_X1 U13398 ( .A(n12901), .ZN(n10414) );
  NAND2_X1 U13399 ( .A1(n12799), .A2(n12798), .ZN(n10413) );
  AND2_X4 U13400 ( .A1(n13451), .A2(n10425), .ZN(n14474) );
  AND2_X1 U13401 ( .A1(n15043), .A2(n14405), .ZN(n10428) );
  OR2_X1 U13402 ( .A1(n15087), .A2(n10431), .ZN(n15089) );
  OR2_X1 U13403 ( .A1(n10435), .A2(n16625), .ZN(n10434) );
  OAI21_X1 U13404 ( .B1(n16046), .B2(n16045), .A(n10441), .ZN(n10437) );
  INV_X1 U13405 ( .A(n16048), .ZN(n10441) );
  NAND2_X1 U13406 ( .A1(n10442), .A2(n10505), .ZN(n10506) );
  AND2_X2 U13407 ( .A1(n13451), .A2(n13441), .ZN(n14119) );
  NOR2_X1 U13408 ( .A1(n13079), .A2(n14416), .ZN(n10448) );
  XNOR2_X1 U13409 ( .A(n13426), .B(n13079), .ZN(n14873) );
  NAND2_X1 U13410 ( .A1(n14602), .A2(n10449), .ZN(n10452) );
  AND2_X1 U13411 ( .A1(n14602), .A2(n14601), .ZN(n14603) );
  INV_X1 U13412 ( .A(n10452), .ZN(n14586) );
  NAND3_X1 U13413 ( .A1(n12475), .A2(n12473), .A3(n12474), .ZN(P2_U2825) );
  NAND2_X1 U13414 ( .A1(n10460), .A2(n10462), .ZN(n17026) );
  NAND2_X1 U13415 ( .A1(n17091), .A2(n9891), .ZN(n10460) );
  INV_X1 U13416 ( .A(n17954), .ZN(n10464) );
  INV_X1 U13417 ( .A(n11631), .ZN(n11616) );
  AOI21_X1 U13418 ( .B1(n12592), .B2(n10475), .A(n10474), .ZN(n10473) );
  NAND2_X1 U13419 ( .A1(n10486), .A2(n10484), .ZN(n17098) );
  NAND2_X1 U13420 ( .A1(n17119), .A2(n9860), .ZN(n10484) );
  AOI21_X1 U13421 ( .B1(n17119), .B2(n10487), .A(n17294), .ZN(n10485) );
  NAND2_X1 U13422 ( .A1(n17294), .A2(n10488), .ZN(n10486) );
  INV_X1 U13423 ( .A(n17997), .ZN(n10488) );
  NOR2_X1 U13424 ( .A1(n18123), .A2(n10491), .ZN(n10495) );
  NAND2_X1 U13425 ( .A1(n18128), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10491) );
  NAND2_X1 U13426 ( .A1(n10496), .A2(n10492), .ZN(n17139) );
  NOR2_X1 U13427 ( .A1(n18123), .A2(n10493), .ZN(n10492) );
  NAND3_X1 U13428 ( .A1(n18128), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        n10649), .ZN(n10493) );
  AND2_X2 U13429 ( .A1(n11644), .A2(n9890), .ZN(n11655) );
  NAND2_X1 U13430 ( .A1(n10498), .A2(n9850), .ZN(n11638) );
  NOR2_X2 U13431 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10678) );
  NAND2_X1 U13432 ( .A1(n11045), .A2(n11061), .ZN(n11084) );
  NAND2_X1 U13433 ( .A1(n11045), .A2(n10504), .ZN(n11071) );
  CLKBUF_X1 U13434 ( .A(n12400), .Z(n10507) );
  AND2_X2 U13435 ( .A1(n12400), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10936) );
  INV_X1 U13436 ( .A(n15617), .ZN(n10512) );
  NAND2_X1 U13437 ( .A1(n11834), .A2(n10517), .ZN(n10523) );
  AND2_X1 U13438 ( .A1(n11834), .A2(n16146), .ZN(n16138) );
  NAND3_X1 U13439 ( .A1(n10516), .A2(n9745), .A3(n10518), .ZN(n10514) );
  INV_X1 U13440 ( .A(n11837), .ZN(n10522) );
  NAND2_X1 U13441 ( .A1(n13054), .A2(n9765), .ZN(n13274) );
  NOR2_X2 U13442 ( .A1(n13719), .A2(n10526), .ZN(n15993) );
  AOI21_X1 U13443 ( .B1(n11425), .B2(n9847), .A(n10533), .ZN(n10532) );
  NAND2_X1 U13444 ( .A1(n11108), .A2(n11107), .ZN(n11106) );
  NAND2_X1 U13445 ( .A1(n11132), .A2(n10539), .ZN(n11109) );
  NAND2_X1 U13446 ( .A1(n11181), .A2(n10541), .ZN(n11778) );
  AND2_X1 U13447 ( .A1(n11570), .A2(n11572), .ZN(n11726) );
  NAND2_X1 U13448 ( .A1(n11570), .A2(n10543), .ZN(n15490) );
  INV_X1 U13449 ( .A(n10548), .ZN(n18256) );
  OR2_X1 U13450 ( .A1(n18116), .A2(n10551), .ZN(n18101) );
  NAND3_X2 U13451 ( .A1(n10552), .A2(n10655), .A3(n11883), .ZN(n18288) );
  NOR2_X1 U13452 ( .A1(n11886), .A2(n11887), .ZN(n10552) );
  INV_X1 U13453 ( .A(n10559), .ZN(n18221) );
  INV_X2 U13454 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19079) );
  NAND2_X1 U13455 ( .A1(n14530), .A2(n10565), .ZN(n15498) );
  INV_X1 U13456 ( .A(n10575), .ZN(n11847) );
  NAND3_X1 U13457 ( .A1(n13497), .A2(n9758), .A3(n13750), .ZN(n13749) );
  NAND2_X1 U13458 ( .A1(n11594), .A2(n10584), .ZN(n10583) );
  INV_X1 U13459 ( .A(n11594), .ZN(n16280) );
  XNOR2_X2 U13460 ( .A(n10820), .B(n10821), .ZN(n12153) );
  NAND2_X2 U13461 ( .A1(n10782), .A2(n20229), .ZN(n11220) );
  OR2_X2 U13462 ( .A1(n13495), .A2(n12173), .ZN(n13491) );
  AND2_X1 U13463 ( .A1(n15868), .A2(n15870), .ZN(n15859) );
  AOI21_X1 U13464 ( .B1(n15868), .B2(n9888), .A(n9766), .ZN(n12336) );
  NAND2_X1 U13465 ( .A1(n10588), .A2(n10589), .ZN(n15833) );
  NAND2_X1 U13466 ( .A1(n15868), .A2(n9892), .ZN(n10588) );
  NAND3_X1 U13467 ( .A1(n14853), .A2(n12916), .A3(n14414), .ZN(n10603) );
  INV_X2 U13468 ( .A(n14318), .ZN(n14414) );
  NAND2_X1 U13469 ( .A1(n12914), .A2(n13018), .ZN(n10606) );
  NAND2_X1 U13470 ( .A1(n14614), .A2(n10615), .ZN(n14584) );
  NAND2_X1 U13471 ( .A1(n14614), .A2(n14204), .ZN(n14597) );
  NAND2_X1 U13472 ( .A1(n14681), .A2(n10619), .ZN(n14627) );
  INV_X1 U13473 ( .A(n10624), .ZN(n14653) );
  NAND2_X1 U13474 ( .A1(n11616), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11630) );
  NAND2_X1 U13475 ( .A1(n11508), .A2(n11507), .ZN(n13719) );
  INV_X1 U13476 ( .A(n13423), .ZN(n11508) );
  NAND2_X1 U13477 ( .A1(n15639), .A2(n15898), .ZN(n15892) );
  AOI21_X1 U13478 ( .B1(n15232), .B2(n20350), .A(n10654), .ZN(n14891) );
  MUX2_X1 U13479 ( .A(n16065), .B(n16064), .S(n16063), .Z(n16067) );
  AOI22_X1 U13480 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U13481 ( .A1(n12597), .A2(n19484), .ZN(n12607) );
  BUF_X1 U13482 ( .A(n16054), .Z(n16333) );
  CLKBUF_X1 U13483 ( .A(n15873), .Z(n15879) );
  NAND2_X1 U13484 ( .A1(n13895), .A2(n13894), .ZN(n14365) );
  CLKBUF_X1 U13485 ( .A(n15993), .Z(n15994) );
  NAND2_X1 U13486 ( .A1(n15993), .A2(n11552), .ZN(n15617) );
  XNOR2_X1 U13487 ( .A(n17800), .B(n12098), .ZN(n12099) );
  INV_X1 U13488 ( .A(n17808), .ZN(n12098) );
  OAI21_X1 U13489 ( .B1(n12164), .B2(n12163), .A(n12162), .ZN(n12167) );
  CLKBUF_X1 U13490 ( .A(n12164), .Z(n13315) );
  NOR2_X1 U13491 ( .A1(n10779), .A2(n11212), .ZN(n11240) );
  CLKBUF_X1 U13492 ( .A(n13743), .Z(n13789) );
  INV_X1 U13493 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U13494 ( .A1(n12882), .A2(n12892), .B1(n12881), .B2(n13208), .ZN(
        n12883) );
  AOI22_X1 U13495 ( .A1(n12264), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10758) );
  AND2_X2 U13496 ( .A1(n12264), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10862) );
  NAND2_X1 U13497 ( .A1(n15489), .A2(n11797), .ZN(n11799) );
  OR2_X1 U13498 ( .A1(n10811), .A2(n10810), .ZN(n10812) );
  NOR2_X2 U13499 ( .A1(n14627), .A2(n14630), .ZN(n14614) );
  OAI21_X2 U13500 ( .B1(n16835), .B2(n12163), .A(n12155), .ZN(n16650) );
  OR2_X1 U13501 ( .A1(n12598), .A2(n16842), .ZN(n10633) );
  NOR2_X1 U13502 ( .A1(n11804), .A2(n11803), .ZN(n10634) );
  OR2_X1 U13503 ( .A1(n14544), .A2(n16836), .ZN(n10635) );
  NOR2_X1 U13504 ( .A1(n11579), .A2(n11578), .ZN(n10636) );
  INV_X1 U13505 ( .A(n14932), .ZN(n20351) );
  INV_X1 U13506 ( .A(n13269), .ZN(n20392) );
  NAND2_X1 U13507 ( .A1(n13204), .A2(n13203), .ZN(n14552) );
  OR2_X1 U13508 ( .A1(n14544), .A2(n16287), .ZN(n10637) );
  NAND2_X1 U13509 ( .A1(n12131), .A2(n18199), .ZN(n10638) );
  AND3_X1 U13510 ( .A1(n12120), .A2(n18423), .A3(n12119), .ZN(n10639) );
  INV_X1 U13511 ( .A(n19322), .ZN(n19366) );
  AND2_X1 U13512 ( .A1(n12334), .A2(n12333), .ZN(n10641) );
  INV_X1 U13513 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14406) );
  INV_X1 U13514 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16259) );
  AND2_X1 U13515 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10643) );
  AND2_X1 U13516 ( .A1(n10738), .A2(n10737), .ZN(n10644) );
  AND2_X1 U13517 ( .A1(n14392), .A2(n15377), .ZN(n10645) );
  AND2_X1 U13518 ( .A1(n15210), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10646) );
  AND2_X1 U13519 ( .A1(n10635), .A2(n11806), .ZN(n10647) );
  AND2_X4 U13520 ( .A1(n13629), .A2(n10789), .ZN(n10648) );
  AND2_X1 U13521 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10649) );
  NAND2_X1 U13522 ( .A1(n12887), .A2(n12976), .ZN(n12979) );
  AND2_X1 U13524 ( .A1(n13586), .A2(n13585), .ZN(n10650) );
  INV_X1 U13525 ( .A(n15878), .ZN(n15884) );
  INV_X1 U13526 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11092) );
  AND4_X1 U13527 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n10651) );
  INV_X1 U13528 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11819) );
  AND2_X1 U13529 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10652) );
  AND2_X1 U13530 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .ZN(n10653) );
  AND2_X1 U13531 ( .A1(n14922), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n10654) );
  AND4_X1 U13532 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n10655) );
  NOR2_X1 U13533 ( .A1(n12595), .A2(n12594), .ZN(n10656) );
  OR2_X1 U13534 ( .A1(n12382), .A2(n14519), .ZN(n10657) );
  AND2_X1 U13535 ( .A1(n10733), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10658) );
  CLKBUF_X3 U13536 ( .A(n11963), .Z(n17564) );
  AND2_X1 U13537 ( .A1(n10743), .A2(n10742), .ZN(n10659) );
  OR3_X1 U13538 ( .A1(n18617), .A2(n18621), .A3(n19102), .ZN(n10660) );
  NAND2_X1 U13539 ( .A1(n11799), .A2(n11798), .ZN(n12465) );
  OR2_X1 U13540 ( .A1(n19055), .A2(n12581), .ZN(n10662) );
  AND3_X1 U13541 ( .A1(n13905), .A2(n15005), .A3(n13904), .ZN(n10664) );
  INV_X1 U13542 ( .A(n14614), .ZN(n14629) );
  OR2_X1 U13543 ( .A1(n13063), .A2(n14519), .ZN(n10665) );
  AND2_X1 U13544 ( .A1(n10719), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10666) );
  OAI21_X1 U13545 ( .B1(n18090), .B2(n17984), .A(n12124), .ZN(n12125) );
  AND2_X1 U13546 ( .A1(n12139), .A2(n12593), .ZN(n10667) );
  INV_X1 U13547 ( .A(n12146), .ZN(n10840) );
  AND2_X1 U13548 ( .A1(n15797), .A2(n16647), .ZN(n10668) );
  OR2_X1 U13549 ( .A1(n12463), .A2(n15816), .ZN(n10669) );
  INV_X1 U13550 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n11619) );
  AND2_X1 U13551 ( .A1(n16061), .A2(n16064), .ZN(n10671) );
  AND4_X1 U13552 ( .A1(n16195), .A2(n16180), .A3(n16214), .A4(n16201), .ZN(
        n10672) );
  OR2_X1 U13553 ( .A1(n12576), .A2(n19490), .ZN(n10673) );
  INV_X1 U13554 ( .A(n12412), .ZN(n10776) );
  AND4_X1 U13555 ( .A1(n12678), .A2(n12677), .A3(n12676), .A4(n12675), .ZN(
        n10674) );
  AND2_X1 U13556 ( .A1(n12899), .A2(n12898), .ZN(n12982) );
  AND2_X1 U13557 ( .A1(n14866), .A2(n13442), .ZN(n12894) );
  AND2_X1 U13558 ( .A1(n14853), .A2(n12702), .ZN(n12732) );
  AND2_X1 U13559 ( .A1(n13095), .A2(n14357), .ZN(n13096) );
  NOR2_X1 U13560 ( .A1(n13833), .A2(n12719), .ZN(n12731) );
  AND2_X1 U13561 ( .A1(n20953), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12708) );
  OR2_X1 U13562 ( .A1(n12412), .A2(n19523), .ZN(n10774) );
  AOI22_X1 U13563 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10692) );
  OR2_X1 U13564 ( .A1(n13512), .A2(n13511), .ZN(n13539) );
  NOR2_X1 U13565 ( .A1(n10923), .A2(n10922), .ZN(n10924) );
  NAND2_X1 U13566 ( .A1(n19518), .A2(n12146), .ZN(n10780) );
  INV_X1 U13567 ( .A(n15834), .ZN(n12333) );
  AND2_X1 U13568 ( .A1(n10805), .A2(n10804), .ZN(n10806) );
  INV_X1 U13569 ( .A(n12257), .ZN(n11017) );
  INV_X1 U13570 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10675) );
  OR2_X1 U13572 ( .A1(n14318), .A2(n14416), .ZN(n13427) );
  INV_X1 U13573 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12726) );
  NAND2_X1 U13574 ( .A1(n11232), .A2(n11789), .ZN(n11041) );
  OR2_X1 U13575 ( .A1(n11695), .A2(n15863), .ZN(n11696) );
  INV_X1 U13576 ( .A(n11219), .ZN(n11221) );
  AND2_X1 U13577 ( .A1(n10998), .A2(n10997), .ZN(n11599) );
  INV_X1 U13578 ( .A(n18019), .ZN(n12587) );
  INV_X1 U13579 ( .A(n14185), .ZN(n14184) );
  INV_X1 U13580 ( .A(n14114), .ZN(n14115) );
  NAND2_X1 U13581 ( .A1(n12979), .A2(n12862), .ZN(n12889) );
  INV_X1 U13582 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U13583 ( .A1(n11041), .A2(n11040), .ZN(n11055) );
  NOR2_X1 U13584 ( .A1(n14515), .A2(n12147), .ZN(n12148) );
  AND2_X1 U13585 ( .A1(n15833), .A2(n15836), .ZN(n12338) );
  INV_X1 U13586 ( .A(n11740), .ZN(n11413) );
  INV_X1 U13587 ( .A(n15757), .ZN(n11429) );
  INV_X1 U13588 ( .A(n15623), .ZN(n11316) );
  INV_X1 U13589 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n21268) );
  AND2_X1 U13590 ( .A1(n12748), .A2(n12747), .ZN(n12806) );
  NOR2_X1 U13591 ( .A1(n14324), .A2(n15027), .ZN(n14448) );
  INV_X1 U13592 ( .A(n14020), .ZN(n14021) );
  NAND2_X1 U13593 ( .A1(n13931), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13948) );
  NAND2_X1 U13594 ( .A1(n13869), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13968) );
  NOR2_X1 U13595 ( .A1(n14817), .A2(n14828), .ZN(n14276) );
  AND2_X1 U13596 ( .A1(n12930), .A2(n21029), .ZN(n20776) );
  AND3_X1 U13597 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21091), .A3(n20491), 
        .ZN(n20533) );
  INV_X1 U13598 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20830) );
  INV_X1 U13599 ( .A(n11781), .ZN(n11746) );
  OAI22_X1 U13600 ( .A1(n11044), .A2(n11043), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11030), .ZN(n11202) );
  INV_X1 U13601 ( .A(n13810), .ZN(n12179) );
  INV_X1 U13602 ( .A(n13806), .ZN(n11301) );
  AND3_X1 U13603 ( .A1(n19541), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12146), 
        .ZN(n13490) );
  AND2_X1 U13604 ( .A1(n11223), .A2(n11222), .ZN(n11367) );
  INV_X1 U13605 ( .A(n13741), .ZN(n11290) );
  AND3_X1 U13606 ( .A1(n11521), .A2(n11520), .A3(n11519), .ZN(n13718) );
  INV_X1 U13607 ( .A(n11722), .ZN(n11751) );
  NAND2_X1 U13608 ( .A1(n10759), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10760) );
  NAND2_X1 U13609 ( .A1(n18209), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17198) );
  NAND2_X1 U13610 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .ZN(n17381) );
  INV_X2 U13611 ( .A(n17566), .ZN(n16674) );
  INV_X1 U13612 ( .A(n12105), .ZN(n12104) );
  NAND2_X1 U13613 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  INV_X1 U13614 ( .A(n20337), .ZN(n20322) );
  OR2_X1 U13615 ( .A1(n14557), .A2(n14330), .ZN(n14872) );
  INV_X1 U13616 ( .A(n14413), .ZN(n14317) );
  OR2_X1 U13617 ( .A1(n14926), .A2(n14927), .ZN(n14924) );
  NAND2_X1 U13618 ( .A1(n15007), .A2(n13207), .ZN(n14986) );
  NAND2_X1 U13619 ( .A1(n14116), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14165) );
  NAND2_X1 U13620 ( .A1(n14041), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14076) );
  AOI21_X1 U13621 ( .B1(n14800), .B2(n14768), .A(n14767), .ZN(n14803) );
  NAND2_X1 U13622 ( .A1(n14911), .A2(n14799), .ZN(n14800) );
  INV_X1 U13623 ( .A(n13393), .ZN(n13394) );
  INV_X1 U13624 ( .A(n14573), .ZN(n14574) );
  OR2_X2 U13625 ( .A1(n15341), .A2(n15339), .ZN(n15426) );
  OAI21_X1 U13626 ( .B1(n16753), .B2(n13457), .A(n16754), .ZN(n20491) );
  OR3_X1 U13627 ( .A1(n12876), .A2(n13202), .A3(n12875), .ZN(n16730) );
  AND2_X1 U13628 ( .A1(n20611), .A2(n20640), .ZN(n20619) );
  INV_X1 U13629 ( .A(n20567), .ZN(n20490) );
  INV_X1 U13630 ( .A(n15816), .ZN(n15787) );
  AND2_X1 U13631 ( .A1(n11560), .A2(n11559), .ZN(n12441) );
  AND2_X1 U13632 ( .A1(n16017), .A2(n12427), .ZN(n15985) );
  XNOR2_X1 U13633 ( .A(n16032), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12598) );
  OAI21_X1 U13634 ( .B1(n19618), .B2(n19882), .A(n20180), .ZN(n19628) );
  OR2_X1 U13635 ( .A1(n19944), .A2(n19808), .ZN(n19837) );
  INV_X1 U13636 ( .A(n20033), .ZN(n19978) );
  NAND2_X1 U13637 ( .A1(n20033), .A2(n20201), .ZN(n19498) );
  NAND2_X1 U13638 ( .A1(n17044), .A2(n17390), .ZN(n17033) );
  NOR2_X1 U13639 ( .A1(n17098), .A2(n17294), .ZN(n17092) );
  NOR2_X1 U13640 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17242), .ZN(n17223) );
  NAND2_X1 U13641 ( .A1(n19276), .A2(n17815), .ZN(n12641) );
  NAND2_X1 U13642 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17544), .ZN(n17528) );
  AND2_X1 U13643 ( .A1(n17806), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17665) );
  AND2_X1 U13644 ( .A1(n17750), .A2(n10653), .ZN(n17661) );
  NAND2_X1 U13645 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11904) );
  INV_X1 U13646 ( .A(n12632), .ZN(n12633) );
  INV_X1 U13647 ( .A(n18005), .ZN(n18017) );
  INV_X1 U13648 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18129) );
  XNOR2_X1 U13649 ( .A(n14326), .B(n14562), .ZN(n14510) );
  INV_X1 U13650 ( .A(n14856), .ZN(n20298) );
  AND2_X1 U13651 ( .A1(n14350), .A2(n14348), .ZN(n20337) );
  INV_X1 U13652 ( .A(n20355), .ZN(n14922) );
  NOR2_X1 U13653 ( .A1(n14924), .A2(n14841), .ZN(n14916) );
  AND2_X1 U13654 ( .A1(n13618), .A2(n13905), .ZN(n15004) );
  INV_X1 U13655 ( .A(n14986), .ZN(n13210) );
  INV_X1 U13656 ( .A(n13278), .ZN(n20418) );
  INV_X1 U13657 ( .A(n20488), .ZN(n20485) );
  OR2_X1 U13658 ( .A1(n13328), .A2(n20246), .ZN(n13241) );
  NAND2_X1 U13659 ( .A1(n13612), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13838) );
  NAND2_X1 U13660 ( .A1(n13483), .A2(n13482), .ZN(n13904) );
  AND2_X1 U13661 ( .A1(n15426), .A2(n20474), .ZN(n20464) );
  INV_X1 U13662 ( .A(n15456), .ZN(n20477) );
  NAND2_X1 U13663 ( .A1(n21091), .A2(n20491), .ZN(n20653) );
  NOR2_X1 U13664 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14540) );
  OAI22_X1 U13665 ( .A1(n20503), .A2(n20502), .B1(n20841), .B2(n20650), .ZN(
        n20537) );
  OAI22_X1 U13666 ( .A1(n20577), .A2(n20576), .B1(n20712), .B2(n20841), .ZN(
        n20600) );
  OAI22_X1 U13667 ( .A1(n20619), .A2(n20618), .B1(n13022), .B2(n20617), .ZN(
        n20642) );
  OAI21_X1 U13668 ( .B1(n20616), .B2(n20618), .A(n20615), .ZN(n20643) );
  NOR2_X1 U13669 ( .A1(n15462), .A2(n20749), .ZN(n20605) );
  OAI22_X1 U13670 ( .A1(n20714), .A2(n20713), .B1(n20712), .B2(n20989), .ZN(
        n20737) );
  NOR2_X1 U13671 ( .A1(n20568), .A2(n20567), .ZN(n20807) );
  NOR2_X1 U13672 ( .A1(n20489), .A2(n20750), .ZN(n20742) );
  INV_X1 U13673 ( .A(n20865), .ZN(n20824) );
  INV_X1 U13674 ( .A(n20807), .ZN(n20959) );
  OAI21_X1 U13675 ( .B1(n20881), .B2(n20880), .A(n21035), .ZN(n20901) );
  OAI22_X1 U13676 ( .A1(n20918), .A2(n20917), .B1(n20916), .B2(n20989), .ZN(
        n20948) );
  NAND2_X1 U13677 ( .A1(n15462), .A2(n20489), .ZN(n20873) );
  OAI21_X1 U13678 ( .B1(n20958), .B2(n20957), .A(n21035), .ZN(n20982) );
  NOR2_X2 U13679 ( .A1(n20960), .A2(n20959), .ZN(n21020) );
  NOR2_X1 U13680 ( .A1(n20489), .A2(n21033), .ZN(n20987) );
  INV_X1 U13681 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21090) );
  INV_X1 U13682 ( .A(n19356), .ZN(n16722) );
  AND2_X1 U13683 ( .A1(n13177), .A2(n13696), .ZN(n19322) );
  AND2_X1 U13684 ( .A1(n11227), .A2(n11238), .ZN(n13680) );
  INV_X1 U13685 ( .A(n13801), .ZN(n13802) );
  AND2_X1 U13686 ( .A1(n16017), .A2(n12416), .ZN(n12941) );
  INV_X1 U13687 ( .A(n16023), .ZN(n19398) );
  INV_X1 U13688 ( .A(n12598), .ZN(n12605) );
  AND2_X1 U13689 ( .A1(n16283), .A2(n12853), .ZN(n19487) );
  INV_X1 U13690 ( .A(n19490), .ZN(n19470) );
  OAI21_X1 U13691 ( .B1(n16435), .B2(n16434), .A(n16433), .ZN(n16447) );
  INV_X1 U13692 ( .A(n16842), .ZN(n16640) );
  INV_X1 U13693 ( .A(n19501), .ZN(n20211) );
  NAND2_X1 U13694 ( .A1(n19509), .A2(n19508), .ZN(n19553) );
  INV_X1 U13695 ( .A(n19576), .ZN(n19583) );
  OAI21_X1 U13696 ( .B1(n19592), .B2(n20207), .A(n19594), .ZN(n19613) );
  AND2_X1 U13697 ( .A1(n19715), .A2(n20178), .ZN(n19641) );
  OAI21_X1 U13698 ( .B1(n19689), .B2(n19688), .A(n19687), .ZN(n19710) );
  NAND2_X1 U13699 ( .A1(n19781), .A2(n19780), .ZN(n19800) );
  INV_X1 U13700 ( .A(n19557), .ZN(n19808) );
  AND2_X1 U13701 ( .A1(n20190), .A2(n20199), .ZN(n20178) );
  INV_X1 U13702 ( .A(n20087), .ZN(n19939) );
  INV_X1 U13703 ( .A(n19973), .ZN(n19966) );
  INV_X1 U13704 ( .A(n19991), .ZN(n20041) );
  INV_X1 U13705 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19221) );
  NAND2_X1 U13706 ( .A1(n17033), .A2(n17032), .ZN(n17034) );
  NOR2_X1 U13707 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17339), .ZN(n17323) );
  NOR2_X2 U13708 ( .A1(n12640), .A2(n12641), .ZN(n17353) );
  NAND2_X1 U13709 ( .A1(n12564), .A2(n12563), .ZN(n12565) );
  INV_X1 U13710 ( .A(n17696), .ZN(n17697) );
  NAND2_X1 U13711 ( .A1(n12131), .A2(n18302), .ZN(n16865) );
  NAND2_X1 U13712 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18019) );
  INV_X1 U13713 ( .A(n18690), .ZN(n18905) );
  INV_X1 U13714 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19273) );
  INV_X1 U13715 ( .A(n18485), .ZN(n18496) );
  INV_X1 U13716 ( .A(n18581), .ZN(n18588) );
  AOI21_X2 U13717 ( .B1(n12082), .B2(n12081), .A(n19102), .ZN(n18595) );
  INV_X1 U13718 ( .A(n18639), .ZN(n18998) );
  AND3_X1 U13719 ( .A1(n19134), .A2(n19189), .A3(n19124), .ZN(n19259) );
  INV_X1 U13720 ( .A(n19499), .ZN(n19497) );
  INV_X1 U13721 ( .A(n20333), .ZN(n20294) );
  OR2_X2 U13722 ( .A1(n14510), .A2(n14334), .ZN(n14856) );
  AND2_X1 U13723 ( .A1(n12986), .A2(n13203), .ZN(n20355) );
  OR2_X1 U13724 ( .A1(n14916), .A2(n14842), .ZN(n15221) );
  OR2_X1 U13725 ( .A1(n15004), .A2(n13619), .ZN(n16803) );
  OR2_X1 U13726 ( .A1(n13241), .A2(n13032), .ZN(n20384) );
  NOR2_X1 U13727 ( .A1(n13073), .A2(n13072), .ZN(n13269) );
  OR2_X2 U13728 ( .A1(n13241), .A2(n16744), .ZN(n20253) );
  INV_X1 U13729 ( .A(n20454), .ZN(n20471) );
  INV_X1 U13730 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16728) );
  NAND2_X1 U13731 ( .A1(n20605), .A2(n20904), .ZN(n20566) );
  NAND2_X1 U13732 ( .A1(n20605), .A2(n20807), .ZN(n20604) );
  NAND2_X1 U13733 ( .A1(n20605), .A2(n20986), .ZN(n20646) );
  NAND2_X1 U13734 ( .A1(n20605), .A2(n20871), .ZN(n20676) );
  NAND2_X1 U13735 ( .A1(n20742), .A2(n20904), .ZN(n20703) );
  NAND2_X1 U13736 ( .A1(n20742), .A2(n20807), .ZN(n20741) );
  NAND2_X1 U13737 ( .A1(n20742), .A2(n20986), .ZN(n20774) );
  NAND2_X1 U13738 ( .A1(n20878), .A2(n20904), .ZN(n20828) );
  OR2_X1 U13739 ( .A1(n20873), .A2(n20959), .ZN(n20865) );
  OR2_X1 U13740 ( .A1(n20873), .A2(n20872), .ZN(n20952) );
  NAND2_X1 U13741 ( .A1(n20987), .A2(n20904), .ZN(n20985) );
  NAND2_X1 U13742 ( .A1(n20987), .A2(n20871), .ZN(n21071) );
  OR2_X1 U13743 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20244), .ZN(n21185) );
  OR2_X1 U13744 ( .A1(n14549), .A2(n11723), .ZN(n19368) );
  INV_X1 U13745 ( .A(n19337), .ZN(n19375) );
  INV_X1 U13746 ( .A(n15824), .ZN(n15887) );
  NOR2_X1 U13747 ( .A1(n12436), .A2(n12435), .ZN(n12437) );
  AND2_X1 U13748 ( .A1(n16023), .A2(n16014), .ZN(n16015) );
  AND2_X1 U13749 ( .A1(n16008), .A2(n12942), .ZN(n19403) );
  NOR2_X1 U13750 ( .A1(n19439), .A2(n20237), .ZN(n19435) );
  INV_X1 U13751 ( .A(n19439), .ZN(n19469) );
  INV_X1 U13752 ( .A(n13136), .ZN(n19408) );
  AOI21_X1 U13753 ( .B1(n12605), .B2(n19470), .A(n12604), .ZN(n12606) );
  INV_X1 U13754 ( .A(n19484), .ZN(n16299) );
  INV_X1 U13755 ( .A(n16832), .ZN(n16625) );
  NAND2_X1 U13756 ( .A1(n19557), .A2(n19715), .ZN(n19576) );
  OR2_X1 U13757 ( .A1(n19742), .A2(n19882), .ZN(n19644) );
  INV_X1 U13758 ( .A(n19709), .ZN(n19697) );
  INV_X1 U13759 ( .A(n19794), .ZN(n19804) );
  OR2_X1 U13760 ( .A1(n19974), .A2(n19808), .ZN(n19842) );
  INV_X1 U13761 ( .A(n19940), .ZN(n19911) );
  NAND2_X1 U13762 ( .A1(n19913), .A2(n19912), .ZN(n19973) );
  NOR2_X1 U13763 ( .A1(n13700), .A2(n13766), .ZN(n13730) );
  NOR2_X1 U13764 ( .A1(n19053), .A2(n17853), .ZN(n19276) );
  AOI21_X1 U13765 ( .B1(n17036), .B2(n17035), .A(n17034), .ZN(n17037) );
  INV_X1 U13766 ( .A(n17377), .ZN(n17334) );
  NOR2_X1 U13767 ( .A1(n17390), .A2(n17389), .ZN(n17408) );
  NOR2_X1 U13768 ( .A1(n11871), .A2(n11870), .ZN(n17783) );
  INV_X1 U13769 ( .A(n17832), .ZN(n17852) );
  NAND2_X1 U13770 ( .A1(n18481), .A2(n18586), .ZN(n18581) );
  INV_X1 U13771 ( .A(n18598), .ZN(n18593) );
  AOI211_X1 U13772 ( .C1(n19258), .C2(n10333), .A(n18616), .B(n16696), .ZN(
        n19240) );
  INV_X1 U13773 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19134) );
  INV_X1 U13774 ( .A(n16958), .ZN(n16954) );
  NAND2_X1 U13775 ( .A1(n12596), .A2(n10656), .ZN(P3_U2800) );
  AND2_X4 U13776 ( .A1(n13655), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10749) );
  AND2_X4 U13777 ( .A1(n13655), .A2(n10789), .ZN(n10850) );
  AND3_X4 U13778 ( .A1(n10677), .A2(n10676), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12401) );
  AND2_X4 U13779 ( .A1(n10678), .A2(n13627), .ZN(n12400) );
  AOI22_X1 U13780 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10681) );
  AND2_X4 U13781 ( .A1(n13656), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10855) );
  AND2_X4 U13782 ( .A1(n13629), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12265) );
  AOI22_X1 U13783 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10680) );
  AND2_X4 U13784 ( .A1(n13656), .A2(n10789), .ZN(n10727) );
  BUF_X4 U13785 ( .A(n10727), .Z(n12264) );
  AOI22_X1 U13786 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13787 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13788 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13789 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13790 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10685) );
  BUF_X4 U13791 ( .A(n10727), .Z(n12399) );
  AOI22_X1 U13792 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10684) );
  NAND4_X1 U13793 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n10688) );
  AOI22_X1 U13794 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13795 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13796 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10690) );
  NAND3_X1 U13797 ( .A1(n10692), .A2(n10691), .A3(n10690), .ZN(n10693) );
  AOI22_X1 U13798 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13799 ( .A1(n12264), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10695) );
  NAND2_X1 U13800 ( .A1(n10696), .A2(n10695), .ZN(n10700) );
  AOI22_X1 U13801 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13802 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10697) );
  NAND2_X1 U13803 ( .A1(n10698), .A2(n10697), .ZN(n10699) );
  NOR2_X1 U13804 ( .A1(n10700), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U13805 ( .A1(n10701), .A2(n11030), .ZN(n10708) );
  AOI22_X1 U13806 ( .A1(n12264), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13807 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13808 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13809 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13810 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13811 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13812 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13813 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10709) );
  NAND4_X1 U13814 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10713) );
  AOI22_X1 U13815 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13816 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13817 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13818 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10714) );
  NAND4_X1 U13819 ( .A1(n10717), .A2(n10716), .A3(n10715), .A4(n10714), .ZN(
        n10718) );
  AOI22_X1 U13820 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13821 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13822 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13823 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13824 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10724) );
  AOI22_X1 U13825 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13826 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13827 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13828 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13829 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13830 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13831 ( .A1(n10727), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13832 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13833 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13834 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13835 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13836 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10740) );
  AOI22_X1 U13837 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U13838 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13839 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10737) );
  NAND3_X1 U13840 ( .A1(n10740), .A2(n10739), .A3(n10644), .ZN(n10741) );
  NAND2_X1 U13841 ( .A1(n10741), .A2(n11030), .ZN(n10748) );
  AOI22_X1 U13842 ( .A1(n12264), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13843 ( .A1(n10749), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10850), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13844 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13845 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10742) );
  NAND3_X1 U13846 ( .A1(n10745), .A2(n10744), .A3(n10659), .ZN(n10746) );
  NAND2_X1 U13847 ( .A1(n10746), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10747) );
  AOI22_X1 U13848 ( .A1(n10850), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10749), .ZN(n10753) );
  AOI22_X1 U13849 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10751) );
  NAND4_X1 U13850 ( .A1(n10753), .A2(n10752), .A3(n10751), .A4(n10750), .ZN(
        n10754) );
  AOI22_X1 U13851 ( .A1(n10855), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12265), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13852 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10755) );
  NAND4_X1 U13853 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10759) );
  NAND3_X1 U13854 ( .A1(n10106), .A2(n12169), .A3(n13069), .ZN(n10764) );
  NOR2_X1 U13855 ( .A1(n11722), .A2(n11619), .ZN(n10769) );
  INV_X1 U13856 ( .A(n10770), .ZN(n10771) );
  NAND2_X1 U13857 ( .A1(n10783), .A2(n11204), .ZN(n11219) );
  NAND3_X1 U13858 ( .A1(n11219), .A2(n13069), .A3(n11218), .ZN(n11358) );
  NAND2_X1 U13859 ( .A1(n11358), .A2(n19523), .ZN(n10775) );
  NAND2_X1 U13860 ( .A1(n10783), .A2(n19513), .ZN(n11353) );
  INV_X1 U13861 ( .A(n10784), .ZN(n10786) );
  NOR2_X1 U13862 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U13863 ( .A1(n10802), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10788) );
  AOI21_X1 U13864 ( .B1(n11619), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10790) );
  INV_X1 U13865 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13181) );
  INV_X1 U13866 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19294) );
  INV_X1 U13867 ( .A(n13698), .ZN(n10799) );
  NAND2_X1 U13868 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10791) );
  OAI211_X1 U13869 ( .C1(n10792), .C2(n19294), .A(n10799), .B(n10791), .ZN(
        n10793) );
  NAND2_X1 U13870 ( .A1(n13698), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10795) );
  INV_X1 U13871 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20188) );
  INV_X1 U13872 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16617) );
  AOI22_X1 U13873 ( .A1(n11293), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10805) );
  NAND2_X1 U13874 ( .A1(n10803), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10804) );
  NAND2_X2 U13875 ( .A1(n10807), .A2(n10806), .ZN(n11257) );
  XNOR2_X2 U13876 ( .A(n10808), .B(n11257), .ZN(n10809) );
  NAND2_X2 U13877 ( .A1(n10817), .A2(n10812), .ZN(n16835) );
  INV_X1 U13878 ( .A(n10817), .ZN(n10820) );
  NAND2_X1 U13879 ( .A1(n10950), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10828) );
  INV_X1 U13881 ( .A(n16835), .ZN(n15813) );
  AOI22_X1 U13882 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19752), .B1(
        n19946), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10827) );
  INV_X1 U13883 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n21480) );
  NAND2_X1 U13884 ( .A1(n13315), .A2(n10841), .ZN(n10837) );
  INV_X1 U13885 ( .A(n10945), .ZN(n10834) );
  INV_X1 U13886 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10833) );
  AOI21_X1 U13887 ( .B1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n19851), .A(
        n10835), .ZN(n10848) );
  AOI22_X1 U13888 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19588), .B1(
        n19779), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10847) );
  INV_X1 U13889 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10838) );
  NAND2_X1 U13890 ( .A1(n13315), .A2(n10836), .ZN(n10839) );
  INV_X1 U13891 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10869) );
  OAI22_X1 U13892 ( .A1(n10838), .A2(n19620), .B1(n19811), .B2(n10869), .ZN(
        n10845) );
  INV_X1 U13893 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10843) );
  NAND2_X1 U13894 ( .A1(n19686), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10842) );
  OAI211_X1 U13895 ( .C1(n19884), .C2(n10843), .A(n13063), .B(n10842), .ZN(
        n10844) );
  NOR2_X1 U13896 ( .A1(n10845), .A2(n10844), .ZN(n10846) );
  AOI22_X1 U13897 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10885), .B1(
        n11246), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13898 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n10882), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10853) );
  AND2_X2 U13899 ( .A1(n12264), .A2(n11030), .ZN(n10884) );
  AOI22_X1 U13900 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n10912), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10852) );
  AND2_X2 U13901 ( .A1(n12395), .A2(n11030), .ZN(n10935) );
  AOI22_X1 U13902 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10851) );
  NAND4_X1 U13903 ( .A1(n10854), .A2(n10853), .A3(n10852), .A4(n10851), .ZN(
        n10861) );
  AND2_X2 U13904 ( .A1(n10855), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10883) );
  AOI22_X1 U13905 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10859) );
  AND2_X2 U13906 ( .A1(n10648), .A2(n11030), .ZN(n10911) );
  AOI22_X1 U13907 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10911), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n12256), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13909 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12257), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10856) );
  NAND4_X1 U13910 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10860) );
  AND2_X1 U13911 ( .A1(n19513), .A2(n11582), .ZN(n12856) );
  AOI22_X1 U13912 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13913 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13914 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U13915 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10865) );
  NAND4_X1 U13916 ( .A1(n10868), .A2(n10867), .A3(n10866), .A4(n10865), .ZN(
        n10881) );
  INV_X1 U13917 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10870) );
  INV_X1 U13918 ( .A(n10937), .ZN(n11013) );
  INV_X1 U13919 ( .A(n10936), .ZN(n11016) );
  OAI22_X1 U13920 ( .A1(n10870), .A2(n11013), .B1(n11016), .B2(n10869), .ZN(
        n10871) );
  INV_X1 U13921 ( .A(n10871), .ZN(n10876) );
  NAND2_X1 U13922 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10875) );
  NAND2_X1 U13923 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10874) );
  AOI22_X1 U13924 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10873) );
  NAND4_X1 U13925 ( .A1(n10876), .A2(n10875), .A3(n10874), .A4(n10873), .ZN(
        n10879) );
  INV_X1 U13926 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10877) );
  OAI22_X1 U13927 ( .A1(n10877), .A2(n11017), .B1(n11012), .B2(n21480), .ZN(
        n10878) );
  NAND2_X1 U13928 ( .A1(n12856), .A2(n11581), .ZN(n11587) );
  AOI22_X1 U13929 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10882), .B1(
        n10883), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13930 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10912), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U13931 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13932 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10886) );
  NAND4_X1 U13933 ( .A1(n10889), .A2(n10888), .A3(n10887), .A4(n10886), .ZN(
        n10895) );
  AOI22_X1 U13934 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13935 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10911), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13936 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12257), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13937 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12256), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10890) );
  NAND4_X1 U13938 ( .A1(n10893), .A2(n10892), .A3(n10891), .A4(n10890), .ZN(
        n10894) );
  NAND2_X1 U13939 ( .A1(n11587), .A2(n11586), .ZN(n10896) );
  AOI22_X1 U13940 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19717), .B1(
        n10944), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13941 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19752), .B1(
        n20023), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13942 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19686), .B1(
        n19946), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13943 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19588), .B1(
        n19851), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13944 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10950), .B1(
        n19779), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10908) );
  INV_X1 U13945 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10902) );
  INV_X1 U13946 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10901) );
  OAI22_X1 U13947 ( .A1(n10902), .A2(n19559), .B1(n19620), .B2(n10901), .ZN(
        n10906) );
  INV_X1 U13948 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10904) );
  INV_X1 U13949 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10903) );
  OAI22_X1 U13950 ( .A1(n10904), .A2(n19811), .B1(n19884), .B2(n10903), .ZN(
        n10905) );
  NOR2_X1 U13951 ( .A1(n10906), .A2(n10905), .ZN(n10907) );
  AOI22_X1 U13952 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13953 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13954 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U13955 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10913) );
  NAND4_X1 U13956 ( .A1(n10916), .A2(n10915), .A3(n10914), .A4(n10913), .ZN(
        n10919) );
  AOI22_X1 U13957 ( .A1(n10936), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13958 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10935), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13959 ( .A1(n12256), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13960 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10921) );
  NAND3_X1 U13961 ( .A1(n10926), .A2(n10925), .A3(n10924), .ZN(n11421) );
  INV_X1 U13962 ( .A(n11421), .ZN(n10927) );
  NAND2_X1 U13963 ( .A1(n10927), .A2(n19513), .ZN(n10928) );
  AOI22_X1 U13964 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10882), .B1(
        n11246), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13965 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10912), .B1(
        n10883), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13966 ( .A1(n10862), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13967 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10931) );
  NAND4_X1 U13968 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10943) );
  AOI22_X1 U13969 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U13970 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12256), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13971 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12257), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10938) );
  NAND4_X1 U13972 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10942) );
  AOI22_X1 U13973 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19654), .B1(
        n19915), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13974 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19717), .B1(
        n19982), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13975 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19686), .B1(
        n20023), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13976 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19752), .B1(
        n19946), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13977 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10950), .B1(
        n19588), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13978 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19779), .B1(
        n19851), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10958) );
  INV_X1 U13979 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10952) );
  INV_X1 U13980 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10951) );
  OAI22_X1 U13981 ( .A1(n10952), .A2(n19811), .B1(n19884), .B2(n10951), .ZN(
        n10956) );
  INV_X1 U13982 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10954) );
  INV_X1 U13983 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10953) );
  OAI22_X1 U13984 ( .A1(n10954), .A2(n19559), .B1(n19620), .B2(n10953), .ZN(
        n10955) );
  NOR2_X1 U13985 ( .A1(n10956), .A2(n10955), .ZN(n10957) );
  AOI22_X1 U13986 ( .A1(n10936), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U13987 ( .A1(n12256), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13988 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10960) );
  NAND4_X1 U13989 ( .A1(n10963), .A2(n10962), .A3(n10961), .A4(n10960), .ZN(
        n10969) );
  AOI22_X1 U13990 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U13991 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U13992 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U13993 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10964) );
  NAND4_X1 U13994 ( .A1(n10967), .A2(n10966), .A3(n10965), .A4(n10964), .ZN(
        n10968) );
  INV_X1 U13995 ( .A(n11430), .ZN(n10970) );
  NAND2_X1 U13996 ( .A1(n10970), .A2(n19513), .ZN(n10971) );
  AOI22_X1 U13997 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19717), .B1(
        n19915), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U13998 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19654), .B1(
        n19982), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U13999 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19946), .B1(
        n20023), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U14000 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19752), .B1(
        n19686), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U14001 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10950), .B1(
        n19851), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U14002 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19588), .B1(
        n19779), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10984) );
  INV_X1 U14003 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10978) );
  INV_X1 U14004 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10977) );
  OAI22_X1 U14005 ( .A1(n10978), .A2(n19559), .B1(n19884), .B2(n10977), .ZN(
        n10982) );
  INV_X1 U14006 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10980) );
  INV_X1 U14007 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10979) );
  OAI22_X1 U14008 ( .A1(n10980), .A2(n19620), .B1(n19811), .B2(n10979), .ZN(
        n10981) );
  NOR2_X1 U14009 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  NAND4_X1 U14010 ( .A1(n10986), .A2(n10985), .A3(n10984), .A4(n10983), .ZN(
        n10998) );
  AOI22_X1 U14011 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10936), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12256), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U14013 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10987) );
  NAND4_X1 U14014 ( .A1(n10990), .A2(n10989), .A3(n10988), .A4(n10987), .ZN(
        n10996) );
  AOI22_X1 U14015 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14016 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U14017 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U14018 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10991) );
  NAND4_X1 U14019 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n10995) );
  NAND2_X1 U14020 ( .A1(n11434), .A2(n19513), .ZN(n10997) );
  NAND2_X1 U14021 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11002) );
  NAND2_X1 U14022 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11001) );
  NAND2_X1 U14023 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11000) );
  NAND2_X1 U14024 ( .A1(n10864), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10999) );
  NAND2_X1 U14025 ( .A1(n10935), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11006) );
  NAND2_X1 U14026 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11005) );
  NAND2_X1 U14027 ( .A1(n10862), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11004) );
  NAND2_X1 U14028 ( .A1(n10872), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11003) );
  NAND2_X1 U14029 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U14030 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U14031 ( .A1(n10911), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11008) );
  NAND2_X1 U14032 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11007) );
  INV_X1 U14033 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11014) );
  INV_X1 U14034 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11011) );
  OAI22_X1 U14035 ( .A1(n11014), .A2(n11013), .B1(n11012), .B2(n11011), .ZN(
        n11020) );
  INV_X1 U14036 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11018) );
  INV_X1 U14037 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11015) );
  OAI22_X1 U14038 ( .A1(n11018), .A2(n11017), .B1(n11016), .B2(n11015), .ZN(
        n11019) );
  INV_X1 U14039 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11032) );
  NAND2_X1 U14040 ( .A1(n13627), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11025) );
  NAND2_X1 U14041 ( .A1(n11026), .A2(n11025), .ZN(n11189) );
  NAND2_X1 U14042 ( .A1(n12154), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11185) );
  INV_X1 U14043 ( .A(n11036), .ZN(n11028) );
  NAND2_X1 U14044 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20196), .ZN(
        n11027) );
  NAND2_X1 U14045 ( .A1(n11028), .A2(n11027), .ZN(n11029) );
  NAND2_X1 U14046 ( .A1(n10789), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11034) );
  XNOR2_X1 U14047 ( .A(n11030), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11043) );
  INV_X1 U14048 ( .A(n11043), .ZN(n11031) );
  XNOR2_X1 U14049 ( .A(n11044), .B(n11031), .ZN(n11196) );
  MUX2_X1 U14050 ( .A(n11421), .B(n11196), .S(n11722), .Z(n11235) );
  NOR2_X1 U14051 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n11033) );
  NAND2_X1 U14052 ( .A1(n11046), .A2(n11056), .ZN(n11042) );
  OAI21_X1 U14053 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n10789), .A(
        n11034), .ZN(n11035) );
  XNOR2_X1 U14054 ( .A(n11036), .B(n11035), .ZN(n11242) );
  INV_X1 U14055 ( .A(n11242), .ZN(n11037) );
  NAND2_X1 U14056 ( .A1(n11722), .A2(n11037), .ZN(n11038) );
  INV_X1 U14057 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11199) );
  NAND2_X1 U14058 ( .A1(n11199), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11201) );
  OR2_X1 U14059 ( .A1(n11202), .A2(n11201), .ZN(n11197) );
  MUX2_X1 U14060 ( .A(n11592), .B(n11197), .S(n11722), .Z(n11236) );
  MUX2_X1 U14061 ( .A(n11236), .B(n21249), .S(n19534), .Z(n11061) );
  INV_X1 U14062 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13571) );
  MUX2_X1 U14063 ( .A(n11430), .B(n13571), .S(n19534), .Z(n11082) );
  MUX2_X1 U14064 ( .A(n11434), .B(P2_EBX_REG_6__SCAN_IN), .S(n19534), .Z(
        n11070) );
  XNOR2_X1 U14065 ( .A(n11071), .B(n11070), .ZN(n19357) );
  INV_X1 U14066 ( .A(n11045), .ZN(n11063) );
  INV_X1 U14067 ( .A(n11056), .ZN(n11051) );
  INV_X1 U14068 ( .A(n11046), .ZN(n11047) );
  OAI21_X1 U14069 ( .B1(n11051), .B2(n11055), .A(n11047), .ZN(n11048) );
  NAND2_X1 U14070 ( .A1(n11063), .A2(n11048), .ZN(n15775) );
  INV_X1 U14071 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13070) );
  INV_X1 U14072 ( .A(n11582), .ZN(n11401) );
  NAND2_X1 U14073 ( .A1(n10679), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11049) );
  AND2_X1 U14074 ( .A1(n11185), .A2(n11049), .ZN(n11241) );
  INV_X1 U14075 ( .A(n11241), .ZN(n11190) );
  MUX2_X1 U14076 ( .A(n11401), .B(n11190), .S(n11722), .Z(n11234) );
  MUX2_X1 U14077 ( .A(n13070), .B(n11234), .S(n11789), .Z(n15809) );
  NOR2_X1 U14078 ( .A1(n15809), .A2(n13181), .ZN(n12852) );
  NAND3_X1 U14079 ( .A1(n19534), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11050) );
  NAND2_X1 U14080 ( .A1(n11051), .A2(n11050), .ZN(n11052) );
  INV_X1 U14081 ( .A(n11052), .ZN(n15800) );
  NAND2_X1 U14082 ( .A1(n12852), .A2(n15800), .ZN(n13183) );
  INV_X1 U14083 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16654) );
  NAND2_X1 U14084 ( .A1(n13183), .A2(n16654), .ZN(n11054) );
  INV_X1 U14085 ( .A(n12852), .ZN(n11053) );
  NAND2_X1 U14086 ( .A1(n11053), .A2(n11052), .ZN(n13182) );
  AND2_X1 U14087 ( .A1(n11054), .A2(n13182), .ZN(n16638) );
  INV_X1 U14088 ( .A(n11055), .ZN(n11057) );
  XNOR2_X1 U14089 ( .A(n11057), .B(n11056), .ZN(n15793) );
  XNOR2_X1 U14090 ( .A(n15793), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n16639) );
  NAND2_X1 U14091 ( .A1(n16638), .A2(n16639), .ZN(n11060) );
  INV_X1 U14092 ( .A(n15793), .ZN(n11058) );
  NAND2_X1 U14093 ( .A1(n11058), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11059) );
  AND2_X1 U14094 ( .A1(n11060), .A2(n11059), .ZN(n11064) );
  INV_X1 U14095 ( .A(n11061), .ZN(n11062) );
  XNOR2_X1 U14096 ( .A(n11063), .B(n11062), .ZN(n16276) );
  INV_X1 U14097 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16592) );
  AND2_X1 U14098 ( .A1(n16276), .A2(n16592), .ZN(n11065) );
  AOI21_X1 U14099 ( .B1(n11064), .B2(n16617), .A(n11065), .ZN(n11069) );
  INV_X1 U14100 ( .A(n11064), .ZN(n16290) );
  INV_X1 U14101 ( .A(n11065), .ZN(n11066) );
  NAND3_X1 U14102 ( .A1(n16290), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n11066), .ZN(n11067) );
  OAI21_X1 U14103 ( .B1(n16276), .B2(n16592), .A(n11067), .ZN(n11068) );
  INV_X1 U14104 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16593) );
  INV_X1 U14105 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13734) );
  INV_X1 U14106 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11072) );
  NOR2_X1 U14107 ( .A1(n11789), .A2(n11072), .ZN(n11075) );
  NAND2_X1 U14108 ( .A1(n11074), .A2(n11075), .ZN(n11076) );
  NAND2_X1 U14109 ( .A1(n11091), .A2(n11076), .ZN(n15725) );
  OR2_X1 U14110 ( .A1(n15725), .A2(n11792), .ZN(n11087) );
  INV_X1 U14111 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16558) );
  NAND2_X1 U14112 ( .A1(n11087), .A2(n16558), .ZN(n16224) );
  INV_X1 U14113 ( .A(n11078), .ZN(n11079) );
  NAND2_X1 U14114 ( .A1(n10104), .A2(n11079), .ZN(n11080) );
  NAND2_X1 U14115 ( .A1(n11074), .A2(n11080), .ZN(n15733) );
  INV_X1 U14116 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16569) );
  NAND2_X1 U14117 ( .A1(n15733), .A2(n16569), .ZN(n16239) );
  NAND2_X1 U14118 ( .A1(n16224), .A2(n16239), .ZN(n11081) );
  INV_X1 U14119 ( .A(n11082), .ZN(n11083) );
  NAND2_X1 U14120 ( .A1(n11084), .A2(n11083), .ZN(n11085) );
  AND2_X1 U14121 ( .A1(n11071), .A2(n11085), .ZN(n15749) );
  AND3_X1 U14122 ( .A1(n16224), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n16239), .ZN(n11089) );
  OR2_X1 U14123 ( .A1(n15733), .A2(n16569), .ZN(n16240) );
  NAND2_X1 U14124 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11369) );
  OR2_X1 U14125 ( .A1(n15733), .A2(n11369), .ZN(n11086) );
  NAND2_X1 U14126 ( .A1(n11813), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11604) );
  OR2_X1 U14127 ( .A1(n15725), .A2(n11604), .ZN(n16223) );
  OAI211_X1 U14128 ( .C1(n11087), .C2(n16240), .A(n11086), .B(n16223), .ZN(
        n11088) );
  NAND2_X1 U14129 ( .A1(n19534), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11090) );
  XNOR2_X1 U14130 ( .A(n11091), .B(n11090), .ZN(n15710) );
  NAND2_X1 U14131 ( .A1(n15710), .A2(n11813), .ZN(n11158) );
  INV_X1 U14132 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16537) );
  NAND2_X1 U14133 ( .A1(n11158), .A2(n16537), .ZN(n16214) );
  INV_X1 U14134 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13748) );
  NAND2_X1 U14135 ( .A1(n11129), .A2(n13748), .ZN(n11121) );
  NAND2_X1 U14136 ( .A1(n19534), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U14137 ( .A1(n19534), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11115) );
  OAI21_X1 U14138 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n19534), .ZN(n11093) );
  INV_X1 U14139 ( .A(n11109), .ZN(n11095) );
  NAND2_X1 U14140 ( .A1(n11095), .A2(n11094), .ZN(n11111) );
  NAND2_X1 U14141 ( .A1(n19534), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11107) );
  INV_X1 U14142 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15625) );
  NOR2_X1 U14143 ( .A1(n11789), .A2(n15625), .ZN(n11144) );
  INV_X1 U14144 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11096) );
  NOR2_X1 U14145 ( .A1(n11789), .A2(n11096), .ZN(n11104) );
  INV_X1 U14146 ( .A(n11104), .ZN(n11097) );
  INV_X1 U14147 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15877) );
  NOR2_X1 U14148 ( .A1(n11789), .A2(n10096), .ZN(n11099) );
  INV_X1 U14149 ( .A(n11744), .ZN(n11098) );
  AOI21_X1 U14150 ( .B1(n11100), .B2(n11099), .A(n11098), .ZN(n11101) );
  NAND2_X1 U14151 ( .A1(n11101), .A2(n9787), .ZN(n19303) );
  OR2_X1 U14152 ( .A1(n19303), .A2(n11792), .ZN(n11149) );
  INV_X1 U14153 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11371) );
  NAND2_X1 U14154 ( .A1(n11149), .A2(n11371), .ZN(n11840) );
  NAND2_X1 U14155 ( .A1(n19534), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11102) );
  MUX2_X1 U14156 ( .A(n19534), .B(n11102), .S(n9750), .Z(n11103) );
  NAND2_X1 U14157 ( .A1(n11103), .A2(n11100), .ZN(n15596) );
  INV_X1 U14158 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16394) );
  NAND2_X1 U14159 ( .A1(n11164), .A2(n16394), .ZN(n16111) );
  NAND2_X1 U14160 ( .A1(n9806), .A2(n11104), .ZN(n11105) );
  NAND2_X1 U14161 ( .A1(n9750), .A2(n11105), .ZN(n15610) );
  INV_X1 U14162 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16409) );
  NAND2_X1 U14163 ( .A1(n11165), .A2(n16409), .ZN(n12451) );
  OAI21_X1 U14164 ( .B1(n11108), .B2(n11107), .A(n11106), .ZN(n19317) );
  INV_X1 U14165 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16444) );
  NAND3_X1 U14166 ( .A1(n11109), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n19534), 
        .ZN(n11110) );
  NAND3_X1 U14167 ( .A1(n11111), .A2(n11744), .A3(n11110), .ZN(n19334) );
  INV_X1 U14168 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16436) );
  OAI21_X1 U14169 ( .B1(n19334), .B2(n11792), .A(n16436), .ZN(n11113) );
  NAND2_X1 U14170 ( .A1(n11813), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11112) );
  INV_X1 U14171 ( .A(n11114), .ZN(n11133) );
  INV_X1 U14172 ( .A(n11115), .ZN(n11116) );
  NAND2_X1 U14173 ( .A1(n9789), .A2(n11116), .ZN(n11117) );
  NAND2_X1 U14174 ( .A1(n15667), .A2(n11813), .ZN(n11118) );
  INV_X1 U14175 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21372) );
  NAND2_X1 U14176 ( .A1(n11118), .A2(n21372), .ZN(n16171) );
  INV_X1 U14177 ( .A(n11119), .ZN(n11120) );
  NAND2_X1 U14178 ( .A1(n11121), .A2(n11120), .ZN(n11122) );
  NAND2_X1 U14179 ( .A1(n9789), .A2(n11122), .ZN(n15675) );
  OR2_X1 U14180 ( .A1(n15675), .A2(n11792), .ZN(n11123) );
  INV_X1 U14181 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21438) );
  NAND2_X1 U14182 ( .A1(n11123), .A2(n21438), .ZN(n16180) );
  NAND2_X1 U14183 ( .A1(n19534), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11126) );
  INV_X1 U14184 ( .A(n11124), .ZN(n11125) );
  MUX2_X1 U14185 ( .A(n11126), .B(P2_EBX_REG_10__SCAN_IN), .S(n11125), .Z(
        n11127) );
  NAND2_X1 U14186 ( .A1(n11127), .A2(n11744), .ZN(n15700) );
  OR2_X1 U14187 ( .A1(n15700), .A2(n11792), .ZN(n11128) );
  INV_X1 U14188 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16205) );
  NAND2_X1 U14189 ( .A1(n11128), .A2(n16205), .ZN(n16201) );
  INV_X1 U14190 ( .A(n11129), .ZN(n11130) );
  AND3_X1 U14191 ( .A1(n11130), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n19534), .ZN(
        n11131) );
  NOR2_X1 U14192 ( .A1(n11132), .A2(n11131), .ZN(n15686) );
  NAND2_X1 U14193 ( .A1(n15686), .A2(n11813), .ZN(n11155) );
  INV_X1 U14194 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U14195 ( .A1(n11155), .A2(n11370), .ZN(n16195) );
  AND4_X1 U14196 ( .A1(n16171), .A2(n16180), .A3(n16201), .A4(n16195), .ZN(
        n11142) );
  NAND2_X1 U14197 ( .A1(n19534), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11134) );
  MUX2_X1 U14198 ( .A(n19534), .B(n11134), .S(n11133), .Z(n11136) );
  INV_X1 U14199 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11135) );
  NAND2_X1 U14200 ( .A1(n11114), .A2(n11135), .ZN(n11139) );
  NAND2_X1 U14201 ( .A1(n15656), .A2(n11813), .ZN(n11152) );
  INV_X1 U14202 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16474) );
  NAND2_X1 U14203 ( .A1(n11152), .A2(n16474), .ZN(n16155) );
  INV_X1 U14204 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11137) );
  NOR2_X1 U14205 ( .A1(n11789), .A2(n11137), .ZN(n11138) );
  NAND2_X1 U14206 ( .A1(n11139), .A2(n11138), .ZN(n11140) );
  NAND2_X1 U14207 ( .A1(n11140), .A2(n11109), .ZN(n15645) );
  OR2_X1 U14208 ( .A1(n15645), .A2(n11792), .ZN(n11141) );
  INV_X1 U14209 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16461) );
  NAND2_X1 U14210 ( .A1(n11141), .A2(n16461), .ZN(n16146) );
  NAND4_X1 U14211 ( .A1(n16139), .A2(n11142), .A3(n16155), .A4(n16146), .ZN(
        n11143) );
  NOR2_X1 U14212 ( .A1(n11837), .A2(n11143), .ZN(n11147) );
  NAND2_X1 U14213 ( .A1(n11106), .A2(n11144), .ZN(n11145) );
  AND2_X1 U14214 ( .A1(n9806), .A2(n11145), .ZN(n15624) );
  NAND2_X1 U14215 ( .A1(n15624), .A2(n11813), .ZN(n11161) );
  INV_X1 U14216 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U14217 ( .A1(n11161), .A2(n11146), .ZN(n16121) );
  AND3_X1 U14218 ( .A1(n12451), .A2(n11147), .A3(n16121), .ZN(n11148) );
  INV_X1 U14219 ( .A(n11149), .ZN(n11150) );
  NAND2_X1 U14220 ( .A1(n11150), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11841) );
  NOR2_X1 U14221 ( .A1(n11151), .A2(n16444), .ZN(n11836) );
  INV_X1 U14222 ( .A(n11152), .ZN(n11153) );
  NAND2_X1 U14223 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16156) );
  AND2_X1 U14224 ( .A1(n11813), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11154) );
  NAND2_X1 U14225 ( .A1(n15667), .A2(n11154), .ZN(n16170) );
  OR3_X1 U14226 ( .A1(n15675), .A2(n11792), .A3(n21438), .ZN(n16179) );
  NAND2_X1 U14227 ( .A1(n16170), .A2(n16179), .ZN(n11159) );
  INV_X1 U14228 ( .A(n11155), .ZN(n11156) );
  NAND2_X1 U14229 ( .A1(n11156), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16196) );
  NAND2_X1 U14230 ( .A1(n11813), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11157) );
  OR2_X1 U14231 ( .A1(n15700), .A2(n11157), .ZN(n16200) );
  OR2_X1 U14232 ( .A1(n11158), .A2(n16537), .ZN(n16216) );
  AND2_X1 U14233 ( .A1(n16200), .A2(n16216), .ZN(n16192) );
  NAND2_X1 U14234 ( .A1(n16196), .A2(n16192), .ZN(n16168) );
  NOR2_X1 U14235 ( .A1(n11159), .A2(n16168), .ZN(n11833) );
  NAND4_X1 U14236 ( .A1(n16156), .A2(n11833), .A3(n11835), .A4(n16145), .ZN(
        n11160) );
  NOR2_X1 U14237 ( .A1(n11836), .A2(n11160), .ZN(n11163) );
  INV_X1 U14238 ( .A(n11161), .ZN(n11162) );
  NAND2_X1 U14239 ( .A1(n11162), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16122) );
  AND2_X1 U14240 ( .A1(n11163), .A2(n16122), .ZN(n11167) );
  INV_X1 U14241 ( .A(n11165), .ZN(n11166) );
  NAND2_X1 U14242 ( .A1(n11166), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12452) );
  AND4_X1 U14243 ( .A1(n11841), .A2(n11167), .A3(n16112), .A4(n12452), .ZN(
        n11168) );
  NAND2_X1 U14244 ( .A1(n19534), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11169) );
  INV_X1 U14245 ( .A(n11169), .ZN(n11170) );
  NAND2_X1 U14246 ( .A1(n9787), .A2(n11170), .ZN(n11171) );
  NAND2_X1 U14247 ( .A1(n11174), .A2(n11171), .ZN(n16712) );
  XNOR2_X1 U14248 ( .A(n11172), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16107) );
  INV_X1 U14249 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16383) );
  NAND2_X1 U14250 ( .A1(n11172), .A2(n16383), .ZN(n11766) );
  INV_X1 U14251 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11173) );
  NOR2_X1 U14252 ( .A1(n11789), .A2(n11173), .ZN(n11175) );
  NOR2_X2 U14253 ( .A1(n11174), .A2(n11175), .ZN(n11181) );
  INV_X1 U14254 ( .A(n11181), .ZN(n15563) );
  NAND2_X1 U14255 ( .A1(n11174), .A2(n11175), .ZN(n11176) );
  NAND2_X1 U14256 ( .A1(n15586), .A2(n11813), .ZN(n11177) );
  XNOR2_X1 U14257 ( .A(n11177), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16094) );
  AND2_X1 U14258 ( .A1(n11813), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11178) );
  NAND2_X1 U14259 ( .A1(n15586), .A2(n11178), .ZN(n11769) );
  INV_X1 U14260 ( .A(n11769), .ZN(n11179) );
  INV_X1 U14261 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21468) );
  AND2_X1 U14262 ( .A1(n11744), .A2(n11813), .ZN(n16086) );
  INV_X1 U14263 ( .A(n16086), .ZN(n11772) );
  NAND2_X1 U14264 ( .A1(n19534), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11182) );
  INV_X1 U14265 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U14266 ( .A1(n11183), .A2(n11744), .ZN(n15556) );
  INV_X1 U14267 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11389) );
  NAND2_X1 U14268 ( .A1(n11813), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11184) );
  XNOR2_X1 U14269 ( .A(n16062), .B(n10671), .ZN(n16080) );
  INV_X1 U14270 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21283) );
  INV_X1 U14271 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20100) );
  INV_X1 U14272 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20089) );
  NOR2_X1 U14273 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n20099) );
  INV_X1 U14274 ( .A(n20099), .ZN(n20090) );
  OAI211_X1 U14275 ( .C1(n21283), .C2(n20100), .A(n20089), .B(n20090), .ZN(
        n20228) );
  NAND2_X1 U14276 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20238) );
  INV_X1 U14277 ( .A(n20238), .ZN(n20103) );
  NOR2_X1 U14278 ( .A1(n20228), .A2(n20103), .ZN(n12841) );
  NAND2_X1 U14279 ( .A1(n11350), .A2(n12841), .ZN(n11211) );
  NAND2_X1 U14280 ( .A1(n11189), .A2(n11185), .ZN(n11231) );
  AND2_X1 U14281 ( .A1(n11186), .A2(n11231), .ZN(n11225) );
  OAI21_X1 U14282 ( .B1(n13063), .B2(n11241), .A(n11225), .ZN(n11188) );
  NAND2_X1 U14283 ( .A1(n19513), .A2(n11242), .ZN(n11187) );
  AOI21_X1 U14284 ( .B1(n11188), .B2(n11187), .A(n13685), .ZN(n11195) );
  NOR2_X1 U14285 ( .A1(n11190), .A2(n11189), .ZN(n11191) );
  NOR2_X1 U14286 ( .A1(n11722), .A2(n11191), .ZN(n11194) );
  NAND2_X1 U14287 ( .A1(n13685), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U14288 ( .A1(n11206), .A2(n13063), .ZN(n11192) );
  MUX2_X1 U14289 ( .A(n11192), .B(n11722), .S(n11242), .Z(n11193) );
  OAI21_X1 U14290 ( .B1(n11195), .B2(n11194), .A(n11193), .ZN(n11198) );
  NAND2_X1 U14291 ( .A1(n11197), .A2(n11196), .ZN(n11224) );
  MUX2_X1 U14292 ( .A(n11198), .B(n11722), .S(n11224), .Z(n11203) );
  NOR2_X1 U14293 ( .A1(n11199), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11200) );
  INV_X1 U14294 ( .A(n11209), .ZN(n11205) );
  OAI21_X1 U14295 ( .B1(n11205), .B2(n13685), .A(n11204), .ZN(n11210) );
  INV_X1 U14296 ( .A(n11238), .ZN(n11207) );
  MUX2_X1 U14297 ( .A(n11211), .B(n11210), .S(n19405), .Z(n11256) );
  NAND2_X1 U14298 ( .A1(n11213), .A2(n13069), .ZN(n11214) );
  AND2_X1 U14299 ( .A1(n19513), .A2(n13685), .ZN(n20226) );
  NAND2_X1 U14300 ( .A1(n11214), .A2(n20226), .ZN(n11359) );
  NAND2_X1 U14301 ( .A1(n11215), .A2(n19513), .ZN(n11365) );
  AOI21_X1 U14302 ( .B1(n13685), .B2(n13069), .A(n11350), .ZN(n11216) );
  NAND2_X1 U14303 ( .A1(n11365), .A2(n11216), .ZN(n11217) );
  AND4_X1 U14304 ( .A1(n11359), .A2(n11349), .A3(n11218), .A4(n11217), .ZN(
        n11223) );
  OAI21_X1 U14305 ( .B1(n11221), .B2(n11350), .A(n11220), .ZN(n11222) );
  INV_X1 U14306 ( .A(n11224), .ZN(n11244) );
  AND2_X1 U14307 ( .A1(n11242), .A2(n11225), .ZN(n11226) );
  NAND2_X1 U14308 ( .A1(n11244), .A2(n11226), .ZN(n11227) );
  NAND3_X1 U14309 ( .A1(n13680), .A2(n10202), .A3(n12841), .ZN(n11228) );
  AND2_X1 U14310 ( .A1(n11367), .A2(n11228), .ZN(n12843) );
  MUX2_X1 U14311 ( .A(n10202), .B(n11350), .S(n19513), .Z(n11229) );
  NAND3_X1 U14312 ( .A1(n11229), .A2(n20238), .A3(n13680), .ZN(n11230) );
  NAND2_X1 U14313 ( .A1(n12843), .A2(n11230), .ZN(n11254) );
  INV_X1 U14314 ( .A(n11231), .ZN(n11233) );
  OAI21_X1 U14315 ( .B1(n11234), .B2(n11233), .A(n11232), .ZN(n11237) );
  NAND3_X1 U14316 ( .A1(n11237), .A2(n11236), .A3(n11235), .ZN(n11239) );
  NAND2_X1 U14317 ( .A1(n11239), .A2(n11238), .ZN(n20221) );
  NAND2_X1 U14318 ( .A1(n13686), .A2(n20226), .ZN(n11612) );
  AND2_X1 U14319 ( .A1(n11242), .A2(n11241), .ZN(n11243) );
  AOI21_X1 U14320 ( .B1(n11244), .B2(n11243), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n11245) );
  NAND2_X1 U14321 ( .A1(n13680), .A2(n11245), .ZN(n11251) );
  INV_X1 U14322 ( .A(n11246), .ZN(n11248) );
  NAND3_X1 U14323 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11247) );
  AND2_X1 U14324 ( .A1(n11199), .A2(n11247), .ZN(n12850) );
  NAND2_X1 U14325 ( .A1(n11248), .A2(n12850), .ZN(n11249) );
  INV_X1 U14326 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12654) );
  NAND2_X1 U14327 ( .A1(n11249), .A2(n12654), .ZN(n11250) );
  NAND2_X1 U14328 ( .A1(n11250), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20208) );
  NAND2_X1 U14329 ( .A1(n11251), .A2(n20208), .ZN(n20216) );
  NAND3_X1 U14330 ( .A1(n20216), .A2(n13686), .A3(n13063), .ZN(n11252) );
  NAND2_X1 U14331 ( .A1(n11253), .A2(n11252), .ZN(n11818) );
  NOR2_X1 U14332 ( .A1(n11254), .A2(n11818), .ZN(n11255) );
  NAND3_X1 U14333 ( .A1(n16648), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n13775) );
  AOI21_X2 U14334 ( .B1(n11256), .B2(n11255), .A(n13775), .ZN(n11613) );
  INV_X1 U14335 ( .A(n11613), .ZN(n11577) );
  NAND2_X1 U14336 ( .A1(n13686), .A2(n11751), .ZN(n20217) );
  INV_X1 U14337 ( .A(n11257), .ZN(n11258) );
  OR2_X1 U14338 ( .A1(n11703), .A2(n16592), .ZN(n11262) );
  AOI22_X1 U14339 ( .A1(n11293), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11260) );
  NAND2_X1 U14340 ( .A1(n11711), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11259) );
  AND2_X1 U14341 ( .A1(n11260), .A2(n11259), .ZN(n11261) );
  NAND2_X1 U14342 ( .A1(n11262), .A2(n11261), .ZN(n13498) );
  OR2_X1 U14343 ( .A1(n11703), .A2(n16593), .ZN(n11266) );
  AOI22_X1 U14344 ( .A1(n11293), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11264) );
  NAND2_X1 U14345 ( .A1(n11711), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11263) );
  AND2_X1 U14346 ( .A1(n11264), .A2(n11263), .ZN(n11265) );
  NAND2_X1 U14347 ( .A1(n11266), .A2(n11265), .ZN(n13569) );
  INV_X1 U14348 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11267) );
  OR2_X1 U14349 ( .A1(n11703), .A2(n11267), .ZN(n11271) );
  AOI22_X1 U14350 ( .A1(n11293), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11269) );
  NAND2_X1 U14351 ( .A1(n11711), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11268) );
  AND2_X1 U14352 ( .A1(n11269), .A2(n11268), .ZN(n11270) );
  AOI22_X1 U14353 ( .A1(n11293), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11273) );
  NAND2_X1 U14354 ( .A1(n11711), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11272) );
  NAND2_X1 U14355 ( .A1(n11273), .A2(n11272), .ZN(n11274) );
  OR2_X1 U14356 ( .A1(n11703), .A2(n16558), .ZN(n11278) );
  AOI22_X1 U14357 ( .A1(n11293), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14358 ( .A1(n11711), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11275) );
  AND2_X1 U14359 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  NAND2_X1 U14360 ( .A1(n11278), .A2(n11277), .ZN(n13750) );
  AOI22_X1 U14361 ( .A1(n11293), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11280) );
  NAND2_X1 U14362 ( .A1(n11711), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11279) );
  NAND2_X1 U14363 ( .A1(n11280), .A2(n11279), .ZN(n11281) );
  AOI21_X1 U14364 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11281), .ZN(n13761) );
  OR2_X1 U14365 ( .A1(n11703), .A2(n16205), .ZN(n11285) );
  AOI22_X1 U14366 ( .A1(n11293), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11283) );
  NAND2_X1 U14367 ( .A1(n11711), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11282) );
  AND2_X1 U14368 ( .A1(n11283), .A2(n11282), .ZN(n11284) );
  AOI22_X1 U14369 ( .A1(n11293), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11288) );
  NAND2_X1 U14370 ( .A1(n11711), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11287) );
  NAND2_X1 U14371 ( .A1(n11288), .A2(n11287), .ZN(n11289) );
  INV_X1 U14372 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n21420) );
  OR2_X1 U14373 ( .A1(n11703), .A2(n21438), .ZN(n11292) );
  AOI22_X1 U14374 ( .A1(n11293), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11291) );
  OAI211_X1 U14375 ( .C1(n11720), .C2(n21420), .A(n11292), .B(n11291), .ZN(
        n13786) );
  OR2_X1 U14376 ( .A1(n11703), .A2(n21372), .ZN(n11297) );
  AOI22_X1 U14377 ( .A1(n11716), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11295) );
  NAND2_X1 U14378 ( .A1(n11711), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11294) );
  AND2_X1 U14379 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  AOI22_X1 U14380 ( .A1(n11716), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11299) );
  NAND2_X1 U14381 ( .A1(n11711), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11298) );
  NAND2_X1 U14382 ( .A1(n11299), .A2(n11298), .ZN(n11300) );
  AOI21_X1 U14383 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11300), .ZN(n13806) );
  OR2_X1 U14384 ( .A1(n11703), .A2(n16461), .ZN(n11305) );
  AOI22_X1 U14385 ( .A1(n11716), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11303) );
  NAND2_X1 U14386 ( .A1(n11711), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11302) );
  AND2_X1 U14387 ( .A1(n11303), .A2(n11302), .ZN(n11304) );
  NAND2_X1 U14388 ( .A1(n11305), .A2(n11304), .ZN(n15640) );
  OR2_X1 U14389 ( .A1(n11703), .A2(n16436), .ZN(n11309) );
  AOI22_X1 U14390 ( .A1(n11716), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11307) );
  NAND2_X1 U14391 ( .A1(n11711), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11306) );
  AND2_X1 U14392 ( .A1(n11307), .A2(n11306), .ZN(n11308) );
  NAND2_X1 U14393 ( .A1(n11309), .A2(n11308), .ZN(n15898) );
  AOI22_X1 U14394 ( .A1(n11716), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11311) );
  NAND2_X1 U14395 ( .A1(n11711), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U14396 ( .A1(n11311), .A2(n11310), .ZN(n11312) );
  AOI21_X1 U14397 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11312), .ZN(n15893) );
  AOI22_X1 U14398 ( .A1(n11716), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11314) );
  NAND2_X1 U14399 ( .A1(n11711), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U14400 ( .A1(n11314), .A2(n11313), .ZN(n11315) );
  AOI21_X1 U14401 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11315), .ZN(n15623) );
  OR2_X1 U14402 ( .A1(n11703), .A2(n16409), .ZN(n11320) );
  AOI22_X1 U14403 ( .A1(n11716), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11318) );
  NAND2_X1 U14404 ( .A1(n11711), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11317) );
  AND2_X1 U14405 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  NAND2_X1 U14406 ( .A1(n11320), .A2(n11319), .ZN(n12455) );
  AOI22_X1 U14407 ( .A1(n11716), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11322) );
  NAND2_X1 U14408 ( .A1(n11711), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11321) );
  NAND2_X1 U14409 ( .A1(n11322), .A2(n11321), .ZN(n11323) );
  AOI21_X1 U14410 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11323), .ZN(n15594) );
  AOI22_X1 U14411 ( .A1(n11716), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11325) );
  NAND2_X1 U14412 ( .A1(n11711), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14413 ( .A1(n11325), .A2(n11324), .ZN(n11326) );
  AOI21_X1 U14414 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11326), .ZN(n11848) );
  OR2_X1 U14415 ( .A1(n11703), .A2(n16383), .ZN(n11330) );
  AOI22_X1 U14416 ( .A1(n11716), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11328) );
  NAND2_X1 U14417 ( .A1(n11711), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11327) );
  AND2_X1 U14418 ( .A1(n11328), .A2(n11327), .ZN(n11329) );
  OR2_X1 U14419 ( .A1(n11703), .A2(n11389), .ZN(n11334) );
  AOI22_X1 U14420 ( .A1(n11716), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11332) );
  NAND2_X1 U14421 ( .A1(n11711), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11331) );
  AND2_X1 U14422 ( .A1(n11332), .A2(n11331), .ZN(n11333) );
  AND2_X1 U14423 ( .A1(n11334), .A2(n11333), .ZN(n11345) );
  INV_X1 U14424 ( .A(n11345), .ZN(n11343) );
  OR2_X1 U14425 ( .A1(n11703), .A2(n21468), .ZN(n11338) );
  AOI22_X1 U14426 ( .A1(n11716), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11336) );
  NAND2_X1 U14427 ( .A1(n11711), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11335) );
  AND2_X1 U14428 ( .A1(n11336), .A2(n11335), .ZN(n11337) );
  NAND2_X1 U14429 ( .A1(n11338), .A2(n11337), .ZN(n15560) );
  INV_X1 U14430 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16371) );
  OR2_X1 U14431 ( .A1(n11703), .A2(n16371), .ZN(n11342) );
  AOI22_X1 U14432 ( .A1(n11716), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11340) );
  NAND2_X1 U14433 ( .A1(n11711), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11339) );
  AND2_X1 U14434 ( .A1(n11340), .A2(n11339), .ZN(n11341) );
  NAND2_X1 U14435 ( .A1(n11342), .A2(n11341), .ZN(n15576) );
  AND2_X1 U14436 ( .A1(n15560), .A2(n15576), .ZN(n11344) );
  NAND2_X1 U14437 ( .A1(n15862), .A2(n11693), .ZN(n15535) );
  NAND2_X1 U14438 ( .A1(n15862), .A2(n11344), .ZN(n15562) );
  NAND2_X1 U14439 ( .A1(n15562), .A2(n11345), .ZN(n11346) );
  NAND2_X1 U14440 ( .A1(n15535), .A2(n11346), .ZN(n16078) );
  NAND2_X1 U14441 ( .A1(n13663), .A2(n19513), .ZN(n11347) );
  NAND2_X1 U14442 ( .A1(n11347), .A2(n13632), .ZN(n11348) );
  NAND2_X1 U14443 ( .A1(n11613), .A2(n11348), .ZN(n16836) );
  NOR2_X1 U14444 ( .A1(n13181), .A2(n16654), .ZN(n13180) );
  NAND2_X1 U14445 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13180), .ZN(
        n16629) );
  NAND2_X1 U14446 ( .A1(n11349), .A2(n19529), .ZN(n11351) );
  AOI22_X1 U14447 ( .A1(n14550), .A2(n11351), .B1(n11350), .B2(n13685), .ZN(
        n11356) );
  NAND2_X1 U14448 ( .A1(n11353), .A2(n11352), .ZN(n11354) );
  MUX2_X1 U14449 ( .A(n12411), .B(n11354), .S(n10776), .Z(n11355) );
  AND3_X1 U14450 ( .A1(n11357), .A2(n11356), .A3(n11355), .ZN(n11362) );
  NAND2_X1 U14451 ( .A1(n11358), .A2(n12146), .ZN(n13654) );
  NAND2_X1 U14452 ( .A1(n13654), .A2(n11359), .ZN(n11360) );
  NAND2_X1 U14453 ( .A1(n11360), .A2(n19523), .ZN(n11361) );
  NAND2_X1 U14454 ( .A1(n13661), .A2(n11363), .ZN(n11364) );
  NAND2_X1 U14455 ( .A1(n11613), .A2(n11364), .ZN(n16430) );
  INV_X1 U14456 ( .A(n11365), .ZN(n11366) );
  NAND2_X1 U14457 ( .A1(n11613), .A2(n13682), .ZN(n16429) );
  NOR2_X1 U14458 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13180), .ZN(
        n16628) );
  AND2_X1 U14459 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16591) );
  AND2_X1 U14460 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11368) );
  AND2_X1 U14461 ( .A1(n16591), .A2(n11368), .ZN(n16554) );
  INV_X1 U14462 ( .A(n11369), .ZN(n16547) );
  NAND2_X1 U14463 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16506) );
  NOR2_X1 U14464 ( .A1(n16506), .A2(n11370), .ZN(n11376) );
  NAND2_X1 U14465 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21214) );
  NOR2_X1 U14466 ( .A1(n21214), .A2(n16474), .ZN(n11379) );
  NAND2_X1 U14467 ( .A1(n16482), .A2(n11379), .ZN(n16441) );
  AND3_X1 U14468 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16418) );
  NAND2_X1 U14469 ( .A1(n16418), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16392) );
  AND2_X1 U14470 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11382) );
  NOR2_X1 U14471 ( .A1(n16371), .A2(n16383), .ZN(n11385) );
  NAND2_X1 U14472 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n11385), .ZN(
        n11372) );
  NOR2_X1 U14473 ( .A1(n16367), .A2(n11372), .ZN(n16346) );
  NAND2_X1 U14474 ( .A1(n16430), .A2(n16429), .ZN(n16556) );
  NOR2_X1 U14475 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20179) );
  NOR2_X1 U14476 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11688) );
  NAND2_X1 U14477 ( .A1(n20179), .A2(n11688), .ZN(n19333) );
  NAND2_X1 U14478 ( .A1(n11577), .A2(n19333), .ZN(n16627) );
  NAND2_X1 U14479 ( .A1(n16846), .A2(n16627), .ZN(n16340) );
  INV_X1 U14480 ( .A(n16430), .ZN(n16632) );
  NAND2_X1 U14481 ( .A1(n16632), .A2(n16629), .ZN(n16553) );
  NAND2_X1 U14482 ( .A1(n16554), .A2(n16547), .ZN(n11373) );
  NOR2_X1 U14483 ( .A1(n16628), .A2(n11373), .ZN(n11374) );
  NAND3_X1 U14484 ( .A1(n16553), .A2(n11374), .A3(n16627), .ZN(n11375) );
  NAND2_X1 U14485 ( .A1(n16340), .A2(n11375), .ZN(n16535) );
  INV_X1 U14486 ( .A(n11376), .ZN(n11377) );
  NAND2_X1 U14487 ( .A1(n16556), .A2(n11377), .ZN(n11378) );
  INV_X1 U14488 ( .A(n11379), .ZN(n11380) );
  NAND2_X1 U14489 ( .A1(n16556), .A2(n11380), .ZN(n11381) );
  INV_X1 U14490 ( .A(n16392), .ZN(n16395) );
  NAND2_X1 U14491 ( .A1(n16395), .A2(n11382), .ZN(n11383) );
  INV_X1 U14492 ( .A(n11385), .ZN(n16368) );
  AOI21_X1 U14493 ( .B1(n16556), .B2(n16368), .A(n21468), .ZN(n11386) );
  INV_X1 U14494 ( .A(n16340), .ZN(n11800) );
  NOR3_X1 U14495 ( .A1(n16355), .A2(n11800), .A3(n11389), .ZN(n11388) );
  INV_X1 U14496 ( .A(n19333), .ZN(n16281) );
  NAND2_X1 U14497 ( .A1(n16281), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16074) );
  INV_X1 U14498 ( .A(n16074), .ZN(n11387) );
  AOI211_X1 U14499 ( .C1(n16346), .C2(n11389), .A(n11388), .B(n11387), .ZN(
        n11390) );
  OAI21_X1 U14500 ( .B1(n16078), .B2(n16836), .A(n11390), .ZN(n11579) );
  NOR2_X1 U14501 ( .A1(n12146), .A2(n11397), .ZN(n11391) );
  NAND2_X1 U14502 ( .A1(n11413), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11396) );
  INV_X1 U14503 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11393) );
  NAND2_X1 U14504 ( .A1(n13063), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11392) );
  OAI211_X1 U14505 ( .C1(n13069), .C2(n11393), .A(n11392), .B(n19977), .ZN(
        n11394) );
  INV_X1 U14506 ( .A(n11394), .ZN(n11395) );
  NAND2_X1 U14507 ( .A1(n11396), .A2(n11395), .ZN(n13707) );
  AND2_X1 U14508 ( .A1(n11397), .A2(n19977), .ZN(n11398) );
  NAND2_X1 U14509 ( .A1(n12415), .A2(n9742), .ZN(n11411) );
  INV_X1 U14510 ( .A(n11404), .ZN(n11399) );
  NAND2_X1 U14511 ( .A1(n12154), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20206) );
  NAND2_X1 U14512 ( .A1(n11399), .A2(n20206), .ZN(n11400) );
  NAND2_X1 U14513 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  AOI22_X1 U14514 ( .A1(n11412), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11736), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11403) );
  NAND2_X1 U14515 ( .A1(n11413), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11402) );
  NAND2_X1 U14516 ( .A1(n11403), .A2(n11402), .ZN(n11407) );
  XNOR2_X1 U14517 ( .A(n13708), .B(n11407), .ZN(n13189) );
  AOI22_X1 U14518 ( .A1(n10783), .A2(n11404), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11406) );
  NAND2_X1 U14519 ( .A1(n11545), .A2(n11581), .ZN(n11405) );
  INV_X1 U14520 ( .A(n11407), .ZN(n11408) );
  NAND2_X1 U14521 ( .A1(n13708), .A2(n11408), .ZN(n11409) );
  NAND2_X1 U14522 ( .A1(n13191), .A2(n11409), .ZN(n11416) );
  NAND2_X1 U14523 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11410) );
  OAI211_X1 U14524 ( .C1(n11534), .C2(n11586), .A(n11411), .B(n11410), .ZN(
        n11417) );
  XNOR2_X1 U14525 ( .A(n11416), .B(n11417), .ZN(n13703) );
  AOI22_X1 U14526 ( .A1(n11737), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11736), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11415) );
  NAND2_X1 U14527 ( .A1(n11733), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11414) );
  INV_X1 U14528 ( .A(n11417), .ZN(n11418) );
  NAND2_X1 U14529 ( .A1(n11416), .A2(n11418), .ZN(n11419) );
  NAND2_X1 U14530 ( .A1(n13705), .A2(n11419), .ZN(n15773) );
  OAI22_X1 U14531 ( .A1(n11441), .A2(n16617), .B1(n20188), .B2(n19977), .ZN(
        n11420) );
  AOI21_X1 U14532 ( .B1(P2_REIP_REG_3__SCAN_IN), .B2(n11733), .A(n11420), .ZN(
        n11423) );
  AOI22_X1 U14533 ( .A1(n11545), .A2(n11421), .B1(n11737), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14534 ( .A1(n11737), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11736), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U14535 ( .A1(n11733), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11427) );
  NAND2_X1 U14536 ( .A1(n11545), .A2(n11592), .ZN(n11426) );
  AOI22_X1 U14537 ( .A1(n11737), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11736), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11433) );
  NAND2_X1 U14538 ( .A1(n11733), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11432) );
  NAND2_X1 U14539 ( .A1(n11545), .A2(n11430), .ZN(n11431) );
  AOI22_X1 U14540 ( .A1(n11737), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11736), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11436) );
  NAND2_X1 U14541 ( .A1(n11733), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U14542 ( .A1(n11436), .A2(n11435), .ZN(n12939) );
  NAND2_X1 U14543 ( .A1(n12938), .A2(n12939), .ZN(n11438) );
  NAND2_X1 U14544 ( .A1(n11545), .A2(n11813), .ZN(n11437) );
  AOI22_X1 U14545 ( .A1(n11737), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11736), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U14546 ( .A1(n11733), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11439) );
  NAND2_X1 U14547 ( .A1(n11440), .A2(n11439), .ZN(n13053) );
  AOI22_X1 U14548 ( .A1(n11737), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11736), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U14549 ( .A1(n11733), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14550 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14551 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14552 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11442) );
  NAND4_X1 U14553 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11451) );
  AOI22_X1 U14554 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n10882), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14555 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n10936), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14556 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n12256), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14557 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10911), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11446) );
  NAND4_X1 U14558 ( .A1(n11449), .A2(n11448), .A3(n11447), .A4(n11446), .ZN(
        n11450) );
  NAND2_X1 U14559 ( .A1(n11545), .A2(n13755), .ZN(n11452) );
  AOI22_X1 U14560 ( .A1(n11737), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11736), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U14561 ( .A1(n11733), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14562 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10884), .B1(
        n10089), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14563 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10937), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14564 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12257), .B1(
        n12256), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14565 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11455) );
  NAND4_X1 U14566 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(
        n11464) );
  AOI22_X1 U14567 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14568 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14569 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14570 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11459) );
  NAND4_X1 U14571 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n11463) );
  OR2_X1 U14572 ( .A1(n11464), .A2(n11463), .ZN(n13759) );
  NAND2_X1 U14573 ( .A1(n11545), .A2(n13759), .ZN(n11465) );
  AOI22_X1 U14574 ( .A1(n11737), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14575 ( .A1(n11733), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14576 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12257), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14577 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12256), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14578 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11469) );
  NAND4_X1 U14579 ( .A1(n11472), .A2(n11471), .A3(n11470), .A4(n11469), .ZN(
        n11478) );
  AOI22_X1 U14580 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n11246), .B1(
        n10883), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14581 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14582 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14583 ( .A1(n10862), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11473) );
  NAND4_X1 U14584 ( .A1(n11476), .A2(n11475), .A3(n11474), .A4(n11473), .ZN(
        n11477) );
  OR2_X1 U14585 ( .A1(n11478), .A2(n11477), .ZN(n13782) );
  NAND2_X1 U14586 ( .A1(n11545), .A2(n13782), .ZN(n11479) );
  INV_X1 U14587 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20127) );
  AOI22_X1 U14588 ( .A1(n11737), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14589 ( .A1(n10936), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14590 ( .A1(n12256), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14591 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14592 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11491) );
  AOI22_X1 U14593 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14594 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14595 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14596 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14597 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  OR2_X1 U14598 ( .A1(n11491), .A2(n11490), .ZN(n13744) );
  NAND2_X1 U14599 ( .A1(n11545), .A2(n13744), .ZN(n11492) );
  OAI211_X1 U14600 ( .C1(n11740), .C2(n20127), .A(n11493), .B(n11492), .ZN(
        n13424) );
  NAND2_X1 U14601 ( .A1(n13355), .A2(n13424), .ZN(n13423) );
  AOI22_X1 U14602 ( .A1(n11737), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11506) );
  INV_X2 U14603 ( .A(n11740), .ZN(n11733) );
  NAND2_X1 U14604 ( .A1(n11733), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14605 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10882), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U14606 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11246), .B1(
        n10883), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14607 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11494) );
  NAND4_X1 U14608 ( .A1(n11497), .A2(n11496), .A3(n11495), .A4(n11494), .ZN(
        n11503) );
  AOI22_X1 U14609 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14610 ( .A1(n10862), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14611 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10937), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14612 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12257), .B1(
        n12256), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11498) );
  NAND4_X1 U14613 ( .A1(n11501), .A2(n11500), .A3(n11499), .A4(n11498), .ZN(
        n11502) );
  OR2_X1 U14614 ( .A1(n11503), .A2(n11502), .ZN(n13792) );
  NAND2_X1 U14615 ( .A1(n11545), .A2(n13792), .ZN(n11504) );
  AOI22_X1 U14616 ( .A1(n11737), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11521) );
  NAND2_X1 U14617 ( .A1(n11733), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14618 ( .A1(n10936), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14619 ( .A1(n12256), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14620 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11509) );
  NAND4_X1 U14621 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11518) );
  AOI22_X1 U14622 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14623 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14624 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14625 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11513) );
  NAND4_X1 U14626 ( .A1(n11516), .A2(n11515), .A3(n11514), .A4(n11513), .ZN(
        n11517) );
  OR2_X1 U14627 ( .A1(n11518), .A2(n11517), .ZN(n13803) );
  NAND2_X1 U14628 ( .A1(n11545), .A2(n13803), .ZN(n11519) );
  AOI22_X1 U14629 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10882), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14630 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10883), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14631 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14632 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U14633 ( .A1(n11525), .A2(n11524), .A3(n11523), .A4(n11522), .ZN(
        n11531) );
  AOI22_X1 U14634 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10863), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14635 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10937), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14636 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12256), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11526) );
  NAND4_X1 U14637 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11530) );
  NOR2_X1 U14638 ( .A1(n11531), .A2(n11530), .ZN(n13810) );
  AOI22_X1 U14639 ( .A1(n11737), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14640 ( .A1(n11733), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11532) );
  OAI211_X1 U14641 ( .C1(n13810), .C2(n11534), .A(n11533), .B(n11532), .ZN(
        n13622) );
  INV_X1 U14642 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20134) );
  AOI22_X1 U14643 ( .A1(n11737), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14644 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10884), .B1(
        n10089), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14645 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10936), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14646 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12257), .B1(
        n12256), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14647 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11535) );
  NAND4_X1 U14648 ( .A1(n11538), .A2(n11537), .A3(n11536), .A4(n11535), .ZN(
        n11544) );
  AOI22_X1 U14649 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14650 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14651 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14652 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11539) );
  NAND4_X1 U14653 ( .A1(n11542), .A2(n11541), .A3(n11540), .A4(n11539), .ZN(
        n11543) );
  OR2_X1 U14654 ( .A1(n11544), .A2(n11543), .ZN(n15905) );
  NAND2_X1 U14655 ( .A1(n11545), .A2(n15905), .ZN(n11546) );
  OAI211_X1 U14656 ( .C1(n11740), .C2(n20134), .A(n11547), .B(n11546), .ZN(
        n13738) );
  AOI22_X1 U14657 ( .A1(n11737), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n9742), .B2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U14658 ( .A1(n11733), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14659 ( .A1(n11737), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U14660 ( .A1(n11733), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11550) );
  INV_X1 U14661 ( .A(n15995), .ZN(n11552) );
  AOI22_X1 U14662 ( .A1(n11737), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n9742), .B2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U14663 ( .A1(n11733), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14664 ( .A1(n11412), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U14665 ( .A1(n11733), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14666 ( .A1(n11412), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n9742), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U14667 ( .A1(n11733), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11557) );
  AND2_X1 U14668 ( .A1(n11558), .A2(n11557), .ZN(n15592) );
  AOI22_X1 U14669 ( .A1(n11412), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11560) );
  NAND2_X1 U14670 ( .A1(n11733), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11559) );
  NOR2_X2 U14671 ( .A1(n12440), .A2(n12441), .ZN(n15959) );
  AOI22_X1 U14672 ( .A1(n11412), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n9742), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11562) );
  NAND2_X1 U14673 ( .A1(n11733), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14674 ( .A1(n11562), .A2(n11561), .ZN(n15958) );
  NAND2_X1 U14675 ( .A1(n15959), .A2(n15958), .ZN(n15571) );
  AOI22_X1 U14676 ( .A1(n11412), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11564) );
  NAND2_X1 U14677 ( .A1(n11733), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11563) );
  AND2_X1 U14678 ( .A1(n11564), .A2(n11563), .ZN(n15572) );
  AOI22_X1 U14679 ( .A1(n11412), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n9742), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U14680 ( .A1(n11733), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11565) );
  AND2_X1 U14681 ( .A1(n11566), .A2(n11565), .ZN(n15587) );
  OR2_X1 U14682 ( .A1(n15572), .A2(n15587), .ZN(n11567) );
  AOI22_X1 U14683 ( .A1(n11737), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n9742), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14684 ( .A1(n11733), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U14685 ( .A1(n11569), .A2(n11568), .ZN(n11572) );
  INV_X1 U14686 ( .A(n11726), .ZN(n11571) );
  OAI21_X1 U14687 ( .B1(n11570), .B2(n11572), .A(n11571), .ZN(n15944) );
  NAND2_X1 U14688 ( .A1(n11573), .A2(n13063), .ZN(n11575) );
  NAND2_X1 U14689 ( .A1(n9885), .A2(n11574), .ZN(n13630) );
  AND2_X1 U14690 ( .A1(n11575), .A2(n13630), .ZN(n11576) );
  NOR2_X2 U14691 ( .A1(n11577), .A2(n11576), .ZN(n16838) );
  NOR2_X1 U14692 ( .A1(n15944), .A2(n16590), .ZN(n11578) );
  INV_X1 U14693 ( .A(n12856), .ZN(n11580) );
  NAND2_X1 U14694 ( .A1(n11580), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12858) );
  XNOR2_X1 U14695 ( .A(n11582), .B(n11581), .ZN(n11583) );
  NOR2_X1 U14696 ( .A1(n12858), .A2(n11583), .ZN(n11585) );
  AOI21_X1 U14697 ( .B1(n12858), .B2(n11583), .A(n11585), .ZN(n13187) );
  INV_X1 U14698 ( .A(n13187), .ZN(n11584) );
  NOR2_X1 U14699 ( .A1(n16654), .A2(n11584), .ZN(n13185) );
  NOR2_X1 U14700 ( .A1(n11585), .A2(n13185), .ZN(n11588) );
  XOR2_X1 U14701 ( .A(n10596), .B(n11588), .Z(n16636) );
  XNOR2_X1 U14702 ( .A(n11587), .B(n11586), .ZN(n16635) );
  NAND2_X1 U14703 ( .A1(n16636), .A2(n16635), .ZN(n16634) );
  OR2_X1 U14704 ( .A1(n11588), .A2(n10596), .ZN(n11589) );
  NAND2_X1 U14705 ( .A1(n16634), .A2(n11589), .ZN(n11590) );
  XNOR2_X1 U14706 ( .A(n11590), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16295) );
  NAND2_X1 U14707 ( .A1(n11590), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11591) );
  NAND2_X1 U14708 ( .A1(n11595), .A2(n16593), .ZN(n16266) );
  OAI21_X1 U14709 ( .B1(n11605), .B2(n11792), .A(n16558), .ZN(n11606) );
  AND3_X1 U14710 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11608) );
  NAND2_X1 U14711 ( .A1(n16395), .A2(n11608), .ZN(n11845) );
  NAND2_X1 U14712 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11609) );
  NOR2_X1 U14713 ( .A1(n16506), .A2(n11609), .ZN(n11844) );
  NAND3_X1 U14714 ( .A1(n11844), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11610) );
  NOR2_X1 U14715 ( .A1(n11845), .A2(n11610), .ZN(n11611) );
  XNOR2_X1 U14716 ( .A(n16083), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16082) );
  INV_X1 U14717 ( .A(n11612), .ZN(n20220) );
  NAND2_X1 U14718 ( .A1(n11613), .A2(n20220), .ZN(n16842) );
  OR2_X1 U14719 ( .A1(n16082), .A2(n16842), .ZN(n11614) );
  NAND3_X1 U14720 ( .A1(n11615), .A2(n10636), .A3(n11614), .ZN(P2_U3021) );
  AND2_X2 U14721 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11622) );
  INV_X1 U14722 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16206) );
  INV_X1 U14723 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n21400) );
  OR2_X2 U14724 ( .A1(n11638), .A2(n21400), .ZN(n11640) );
  INV_X1 U14725 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15674) );
  INV_X1 U14726 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16159) );
  INV_X1 U14727 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11647) );
  INV_X1 U14728 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15629) );
  INV_X1 U14729 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11656) );
  AND2_X2 U14730 ( .A1(n11655), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11660) );
  NAND2_X1 U14731 ( .A1(n11660), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11665) );
  INV_X1 U14732 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16714) );
  OR2_X2 U14733 ( .A1(n11665), .A2(n16714), .ZN(n11669) );
  INV_X1 U14734 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16096) );
  OR2_X2 U14735 ( .A1(n11669), .A2(n16096), .ZN(n11672) );
  INV_X1 U14736 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15565) );
  NOR2_X2 U14737 ( .A1(n11672), .A2(n15565), .ZN(n11671) );
  INV_X1 U14738 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15541) );
  INV_X1 U14739 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16050) );
  AND2_X2 U14740 ( .A1(n11678), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11681) );
  NAND2_X1 U14741 ( .A1(n11681), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11685) );
  INV_X1 U14742 ( .A(n11685), .ZN(n11617) );
  NAND2_X1 U14743 ( .A1(n11617), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U14744 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11620) );
  MUX2_X1 U14745 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n16647) );
  INV_X1 U14746 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19486) );
  MUX2_X1 U14747 ( .A(n19486), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n15797) );
  INV_X1 U14748 ( .A(n11622), .ZN(n11624) );
  OAI21_X1 U14749 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n11624), .ZN(n19477) );
  INV_X1 U14750 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11623) );
  NAND2_X1 U14751 ( .A1(n11624), .A2(n11623), .ZN(n11625) );
  NAND2_X1 U14752 ( .A1(n11626), .A2(n11625), .ZN(n16293) );
  NAND2_X1 U14753 ( .A1(n15780), .A2(n16293), .ZN(n15765) );
  NAND2_X1 U14754 ( .A1(n11626), .A2(n16282), .ZN(n11627) );
  AND2_X1 U14755 ( .A1(n9805), .A2(n11627), .ZN(n16285) );
  NOR2_X1 U14756 ( .A1(n15765), .A2(n16285), .ZN(n15741) );
  INV_X1 U14757 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U14758 ( .A1(n9805), .A2(n11628), .ZN(n11629) );
  NAND2_X1 U14759 ( .A1(n11631), .A2(n11629), .ZN(n16271) );
  NAND2_X1 U14760 ( .A1(n15741), .A2(n16271), .ZN(n19361) );
  NAND2_X1 U14761 ( .A1(n11631), .A2(n16259), .ZN(n11632) );
  AND2_X1 U14762 ( .A1(n11630), .A2(n11632), .ZN(n19363) );
  OR2_X1 U14763 ( .A1(n19361), .A2(n19363), .ZN(n15730) );
  NAND2_X1 U14764 ( .A1(n11630), .A2(n16250), .ZN(n11633) );
  AND2_X1 U14765 ( .A1(n9803), .A2(n11633), .ZN(n16252) );
  OR2_X1 U14766 ( .A1(n15730), .A2(n16252), .ZN(n15718) );
  INV_X1 U14767 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16231) );
  NAND2_X1 U14768 ( .A1(n9803), .A2(n16231), .ZN(n11634) );
  AND2_X1 U14769 ( .A1(n9804), .A2(n11634), .ZN(n16234) );
  NAND2_X1 U14770 ( .A1(n9804), .A2(n10500), .ZN(n11636) );
  NAND2_X1 U14771 ( .A1(n11635), .A2(n11636), .ZN(n16218) );
  NAND2_X1 U14772 ( .A1(n15708), .A2(n16218), .ZN(n15696) );
  NAND2_X1 U14773 ( .A1(n11635), .A2(n16206), .ZN(n11637) );
  AND2_X1 U14774 ( .A1(n11638), .A2(n11637), .ZN(n16209) );
  OR2_X1 U14775 ( .A1(n15696), .A2(n16209), .ZN(n15690) );
  NAND2_X1 U14776 ( .A1(n11638), .A2(n21400), .ZN(n11639) );
  AND2_X1 U14777 ( .A1(n11640), .A2(n11639), .ZN(n16190) );
  NOR2_X1 U14778 ( .A1(n15690), .A2(n16190), .ZN(n15672) );
  NAND2_X1 U14779 ( .A1(n11640), .A2(n15674), .ZN(n11641) );
  NAND2_X1 U14780 ( .A1(n9868), .A2(n11641), .ZN(n16185) );
  AND2_X1 U14781 ( .A1(n15672), .A2(n16185), .ZN(n15661) );
  NAND2_X1 U14782 ( .A1(n9868), .A2(n10470), .ZN(n11642) );
  NAND2_X1 U14783 ( .A1(n9864), .A2(n11642), .ZN(n16175) );
  NAND2_X1 U14784 ( .A1(n15661), .A2(n16175), .ZN(n15649) );
  NAND2_X1 U14785 ( .A1(n9864), .A2(n16159), .ZN(n11643) );
  AND2_X1 U14786 ( .A1(n9747), .A2(n11643), .ZN(n16162) );
  OR2_X1 U14787 ( .A1(n15649), .A2(n16162), .ZN(n19341) );
  INV_X1 U14788 ( .A(n11644), .ZN(n11649) );
  INV_X1 U14789 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11645) );
  NAND2_X1 U14790 ( .A1(n11649), .A2(n11645), .ZN(n11646) );
  NAND2_X1 U14791 ( .A1(n9866), .A2(n11646), .ZN(n19340) );
  NAND2_X1 U14792 ( .A1(n9747), .A2(n11647), .ZN(n11648) );
  NAND2_X1 U14793 ( .A1(n11649), .A2(n11648), .ZN(n19338) );
  NAND2_X1 U14794 ( .A1(n19340), .A2(n19338), .ZN(n11650) );
  OR2_X1 U14795 ( .A1(n19341), .A2(n11650), .ZN(n19343) );
  INV_X1 U14796 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11652) );
  NAND2_X1 U14797 ( .A1(n9866), .A2(n11652), .ZN(n11653) );
  AND2_X1 U14798 ( .A1(n11651), .A2(n11653), .ZN(n19319) );
  NAND2_X1 U14799 ( .A1(n11651), .A2(n15629), .ZN(n11654) );
  NAND2_X1 U14800 ( .A1(n11657), .A2(n11654), .ZN(n16127) );
  AND2_X1 U14801 ( .A1(n15631), .A2(n16127), .ZN(n15604) );
  INV_X1 U14802 ( .A(n11655), .ZN(n11662) );
  NAND2_X1 U14803 ( .A1(n11657), .A2(n11656), .ZN(n11658) );
  NAND2_X1 U14804 ( .A1(n11662), .A2(n11658), .ZN(n15605) );
  NAND2_X1 U14805 ( .A1(n15604), .A2(n15605), .ZN(n11659) );
  NAND2_X1 U14806 ( .A1(n11664), .A2(n11659), .ZN(n15595) );
  INV_X1 U14807 ( .A(n11660), .ZN(n11666) );
  INV_X1 U14808 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11661) );
  NAND2_X1 U14809 ( .A1(n11662), .A2(n11661), .ZN(n11663) );
  NAND2_X1 U14810 ( .A1(n11666), .A2(n11663), .ZN(n16116) );
  NAND2_X1 U14811 ( .A1(n15595), .A2(n16116), .ZN(n19307) );
  INV_X1 U14812 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21415) );
  NAND2_X1 U14813 ( .A1(n11666), .A2(n21415), .ZN(n11667) );
  AND2_X1 U14814 ( .A1(n11665), .A2(n11667), .ZN(n19306) );
  NAND2_X1 U14815 ( .A1(n11665), .A2(n16714), .ZN(n11668) );
  NAND2_X1 U14816 ( .A1(n11669), .A2(n11668), .ZN(n16715) );
  NAND2_X1 U14817 ( .A1(n11669), .A2(n16096), .ZN(n11670) );
  AND2_X1 U14818 ( .A1(n11672), .A2(n11670), .ZN(n16098) );
  INV_X1 U14819 ( .A(n11671), .ZN(n11675) );
  NAND2_X1 U14820 ( .A1(n11672), .A2(n15565), .ZN(n11673) );
  NAND2_X1 U14821 ( .A1(n11675), .A2(n11673), .ZN(n16089) );
  OAI21_X1 U14822 ( .B1(n15582), .B2(n15742), .A(n16089), .ZN(n15549) );
  NAND2_X1 U14823 ( .A1(n11675), .A2(n10490), .ZN(n11676) );
  AND2_X1 U14824 ( .A1(n11674), .A2(n11676), .ZN(n16076) );
  AOI21_X1 U14825 ( .B1(n15549), .B2(n11664), .A(n16076), .ZN(n15542) );
  NAND2_X1 U14826 ( .A1(n11674), .A2(n15541), .ZN(n11677) );
  NAND2_X1 U14827 ( .A1(n11679), .A2(n11677), .ZN(n16070) );
  OAI21_X1 U14828 ( .B1(n15542), .B2(n15742), .A(n16070), .ZN(n15527) );
  INV_X1 U14829 ( .A(n11678), .ZN(n11683) );
  NAND2_X1 U14830 ( .A1(n11679), .A2(n16050), .ZN(n11680) );
  AND2_X1 U14831 ( .A1(n11683), .A2(n11680), .ZN(n16052) );
  AOI21_X1 U14832 ( .B1(n15527), .B2(n11664), .A(n16052), .ZN(n15516) );
  INV_X1 U14833 ( .A(n11681), .ZN(n11686) );
  INV_X1 U14834 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U14835 ( .A1(n11683), .A2(n11682), .ZN(n11684) );
  NAND2_X1 U14836 ( .A1(n11686), .A2(n11684), .ZN(n16041) );
  INV_X1 U14837 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16033) );
  NAND2_X1 U14838 ( .A1(n11686), .A2(n16033), .ZN(n11687) );
  AND2_X1 U14839 ( .A1(n11685), .A2(n11687), .ZN(n16035) );
  AOI21_X1 U14840 ( .B1(n15502), .B2(n11664), .A(n16035), .ZN(n12461) );
  XOR2_X1 U14841 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n11685), .Z(
        n12601) );
  OAI21_X1 U14842 ( .B1(n12461), .B2(n15742), .A(n12601), .ZN(n12463) );
  INV_X1 U14843 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20227) );
  AND2_X1 U14844 ( .A1(n20227), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11823) );
  NAND2_X1 U14845 ( .A1(n11823), .A2(n11688), .ZN(n19364) );
  INV_X1 U14846 ( .A(n19364), .ZN(n19344) );
  INV_X1 U14847 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21386) );
  OR2_X1 U14848 ( .A1(n11703), .A2(n21386), .ZN(n11692) );
  AOI22_X1 U14849 ( .A1(n11716), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11690) );
  NAND2_X1 U14850 ( .A1(n11711), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11689) );
  AND2_X1 U14851 ( .A1(n11690), .A2(n11689), .ZN(n11691) );
  AND2_X1 U14852 ( .A1(n11692), .A2(n11691), .ZN(n15534) );
  INV_X1 U14853 ( .A(n15534), .ZN(n11694) );
  NAND2_X1 U14854 ( .A1(n11694), .A2(n11693), .ZN(n11695) );
  INV_X1 U14855 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16315) );
  OR2_X1 U14856 ( .A1(n11703), .A2(n16315), .ZN(n11701) );
  AOI22_X1 U14857 ( .A1(n11716), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11699) );
  NAND2_X1 U14858 ( .A1(n11711), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11698) );
  AND2_X1 U14859 ( .A1(n11699), .A2(n11698), .ZN(n11700) );
  NAND2_X1 U14860 ( .A1(n11701), .A2(n11700), .ZN(n14532) );
  INV_X1 U14861 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11702) );
  OR2_X1 U14862 ( .A1(n11703), .A2(n11702), .ZN(n11707) );
  AOI22_X1 U14863 ( .A1(n11716), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11705) );
  NAND2_X1 U14864 ( .A1(n11711), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11704) );
  AND2_X1 U14865 ( .A1(n11705), .A2(n11704), .ZN(n11706) );
  NAND2_X1 U14866 ( .A1(n11707), .A2(n11706), .ZN(n15511) );
  AOI22_X1 U14867 ( .A1(n11716), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11709) );
  NAND2_X1 U14868 ( .A1(n11711), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U14869 ( .A1(n11709), .A2(n11708), .ZN(n11710) );
  AOI21_X1 U14870 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11710), .ZN(n15496) );
  AOI22_X1 U14871 ( .A1(n11716), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11713) );
  NAND2_X1 U14872 ( .A1(n11711), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11712) );
  NAND2_X1 U14873 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  AOI21_X1 U14874 ( .B1(n11715), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11714), .ZN(n11795) );
  INV_X1 U14875 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14876 ( .A1(n11715), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11718) );
  AOI22_X1 U14877 ( .A1(n11716), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11717) );
  OAI211_X1 U14878 ( .C1(n11720), .C2(n11719), .A(n11718), .B(n11717), .ZN(
        n11721) );
  NAND2_X1 U14879 ( .A1(n11573), .A2(n13680), .ZN(n12652) );
  AND2_X1 U14880 ( .A1(n20238), .A2(n20227), .ZN(n11756) );
  INV_X1 U14881 ( .A(n11756), .ZN(n11750) );
  OR2_X1 U14882 ( .A1(n11722), .A2(n11750), .ZN(n11723) );
  AOI22_X1 U14883 ( .A1(n11412), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n9742), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11725) );
  NAND2_X1 U14884 ( .A1(n11733), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11724) );
  NAND2_X1 U14885 ( .A1(n11725), .A2(n11724), .ZN(n15532) );
  AOI22_X1 U14886 ( .A1(n11412), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11728) );
  NAND2_X1 U14887 ( .A1(n11733), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11727) );
  AND2_X1 U14888 ( .A1(n11728), .A2(n11727), .ZN(n14525) );
  AOI22_X1 U14889 ( .A1(n11412), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11730) );
  NAND2_X1 U14890 ( .A1(n11733), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11729) );
  AND2_X1 U14891 ( .A1(n11730), .A2(n11729), .ZN(n15507) );
  AOI22_X1 U14892 ( .A1(n11412), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11736), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14893 ( .A1(n11733), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11731) );
  AND2_X1 U14894 ( .A1(n11732), .A2(n11731), .ZN(n15491) );
  AOI22_X1 U14895 ( .A1(n11412), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n9742), .B2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11735) );
  NAND2_X1 U14896 ( .A1(n11733), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11734) );
  NAND2_X1 U14897 ( .A1(n11735), .A2(n11734), .ZN(n11797) );
  INV_X1 U14898 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n11825) );
  NAND2_X1 U14899 ( .A1(n9742), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14900 ( .A1(n11737), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n11738) );
  OAI211_X1 U14901 ( .C1(n11740), .C2(n11825), .A(n11739), .B(n11738), .ZN(
        n11741) );
  INV_X1 U14902 ( .A(n13775), .ZN(n13724) );
  NAND2_X1 U14903 ( .A1(n13680), .A2(n13724), .ZN(n11743) );
  OR2_X1 U14904 ( .A1(n11743), .A2(n11742), .ZN(n13114) );
  NAND2_X1 U14905 ( .A1(n12841), .A2(n20227), .ZN(n11757) );
  INV_X1 U14906 ( .A(n11757), .ZN(n13696) );
  NAND2_X1 U14907 ( .A1(n15910), .A2(n19322), .ZN(n11763) );
  INV_X1 U14908 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15552) );
  INV_X1 U14909 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15839) );
  NAND2_X1 U14910 ( .A1(n19534), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11776) );
  NAND2_X1 U14911 ( .A1(n11771), .A2(n11776), .ZN(n11780) );
  INV_X1 U14912 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11745) );
  NOR2_X1 U14913 ( .A1(n11789), .A2(n11745), .ZN(n11781) );
  NAND2_X1 U14914 ( .A1(n19534), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11785) );
  INV_X1 U14915 ( .A(n11785), .ZN(n11748) );
  NOR2_X1 U14916 ( .A1(n11791), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11749) );
  INV_X1 U14917 ( .A(n11771), .ZN(n15537) );
  MUX2_X1 U14918 ( .A(n11749), .B(n15537), .S(n11789), .Z(n11814) );
  NAND3_X1 U14919 ( .A1(n11751), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n11750), 
        .ZN(n11752) );
  NOR2_X1 U14920 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16769) );
  AND2_X1 U14921 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11753) );
  NAND2_X1 U14922 ( .A1(n16769), .A2(n11753), .ZN(n13769) );
  NAND2_X1 U14923 ( .A1(n19364), .A2(n13769), .ZN(n11754) );
  NOR2_X1 U14924 ( .A1(n11754), .A2(n16281), .ZN(n11755) );
  INV_X1 U14925 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11826) );
  INV_X1 U14926 ( .A(n19355), .ZN(n19315) );
  OAI21_X1 U14927 ( .B1(P2_EBX_REG_31__SCAN_IN), .B2(n11756), .A(n12146), .ZN(
        n11758) );
  NAND2_X1 U14928 ( .A1(n11758), .A2(n11757), .ZN(n11759) );
  OR2_X1 U14929 ( .A1(n13114), .A2(n11759), .ZN(n19354) );
  AOI22_X1 U14930 ( .A1(n19315), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n19360), .ZN(n11760) );
  OAI21_X1 U14931 ( .B1(n19375), .B2(n11826), .A(n11760), .ZN(n11761) );
  AOI21_X1 U14932 ( .B1(n11814), .B2(n16722), .A(n11761), .ZN(n11762) );
  OAI211_X1 U14933 ( .C1(n12574), .C2(n19368), .A(n11763), .B(n11762), .ZN(
        n11764) );
  INV_X1 U14934 ( .A(n11764), .ZN(n11765) );
  NAND2_X1 U14935 ( .A1(n10669), .A2(n11765), .ZN(P2_U2824) );
  AND2_X1 U14936 ( .A1(n16094), .A2(n11766), .ZN(n11767) );
  NAND2_X1 U14937 ( .A1(n16086), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11768) );
  NAND2_X1 U14938 ( .A1(n11772), .A2(n21468), .ZN(n11773) );
  INV_X1 U14939 ( .A(n11776), .ZN(n11777) );
  NAND2_X1 U14940 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  NAND2_X1 U14941 ( .A1(n11780), .A2(n11779), .ZN(n15525) );
  NAND2_X1 U14942 ( .A1(n11780), .A2(n11781), .ZN(n11782) );
  NAND2_X1 U14943 ( .A1(n15515), .A2(n11813), .ZN(n16047) );
  AOI21_X1 U14944 ( .B1(n15501), .B2(n11813), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16029) );
  INV_X1 U14945 ( .A(n15501), .ZN(n11787) );
  INV_X1 U14946 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16303) );
  INV_X1 U14947 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n11788) );
  NOR2_X1 U14948 ( .A1(n11789), .A2(n11788), .ZN(n11790) );
  INV_X1 U14949 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11802) );
  OAI21_X1 U14950 ( .B1(n12467), .B2(n11792), .A(n11802), .ZN(n11811) );
  NOR3_X1 U14951 ( .A1(n12467), .A2(n11802), .A3(n11792), .ZN(n11808) );
  NOR2_X1 U14952 ( .A1(n10278), .A2(n11808), .ZN(n11793) );
  NAND2_X1 U14953 ( .A1(n12597), .A2(n16832), .ZN(n11807) );
  OR2_X1 U14954 ( .A1(n11797), .A2(n15489), .ZN(n11798) );
  AND2_X1 U14955 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16316) );
  NAND2_X1 U14956 ( .A1(n16316), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11801) );
  AND2_X1 U14957 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16344) );
  AOI21_X1 U14958 ( .B1(n11801), .B2(n16556), .A(n16327), .ZN(n12568) );
  NAND2_X1 U14959 ( .A1(n16281), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12600) );
  OAI21_X1 U14960 ( .B1(n12568), .B2(n11802), .A(n12600), .ZN(n11804) );
  NAND2_X1 U14961 ( .A1(n16346), .A2(n16344), .ZN(n16329) );
  NOR2_X1 U14962 ( .A1(n16329), .A2(n11801), .ZN(n12571) );
  AND2_X1 U14963 ( .A1(n12571), .A2(n11802), .ZN(n11803) );
  OAI21_X1 U14964 ( .B1(n12465), .B2(n16590), .A(n10634), .ZN(n11805) );
  INV_X1 U14965 ( .A(n11805), .ZN(n11806) );
  NAND3_X1 U14966 ( .A1(n11807), .A2(n10647), .A3(n10633), .ZN(P2_U3016) );
  INV_X1 U14967 ( .A(n11808), .ZN(n11810) );
  NAND2_X1 U14968 ( .A1(n11814), .A2(n11813), .ZN(n11815) );
  XNOR2_X1 U14969 ( .A(n11815), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11816) );
  AND2_X1 U14970 ( .A1(n13685), .A2(n13724), .ZN(n11817) );
  NAND2_X1 U14971 ( .A1(n11818), .A2(n11817), .ZN(n12653) );
  INV_X1 U14972 ( .A(n12653), .ZN(n11821) );
  NAND2_X1 U14973 ( .A1(n12567), .A2(n19484), .ZN(n11832) );
  NAND2_X1 U14974 ( .A1(n11821), .A2(n19513), .ZN(n19490) );
  OR2_X1 U14975 ( .A1(n20180), .A2(n20179), .ZN(n20210) );
  NAND2_X1 U14976 ( .A1(n20210), .A2(n11619), .ZN(n11822) );
  AND2_X1 U14977 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20197) );
  INV_X1 U14978 ( .A(n11823), .ZN(n11824) );
  NAND2_X1 U14979 ( .A1(n11619), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12163) );
  NAND2_X1 U14980 ( .A1(n11824), .A2(n12163), .ZN(n12853) );
  NOR2_X1 U14981 ( .A1(n19333), .A2(n11825), .ZN(n12569) );
  NOR2_X1 U14982 ( .A1(n16283), .A2(n11826), .ZN(n11827) );
  AOI211_X1 U14983 ( .C1(n11828), .C2(n19487), .A(n12569), .B(n11827), .ZN(
        n11829) );
  OAI21_X1 U14984 ( .B1(n12574), .B2(n16287), .A(n11829), .ZN(n11830) );
  NAND3_X1 U14985 ( .A1(n11832), .A2(n10673), .A3(n11831), .ZN(P2_U2983) );
  NAND2_X1 U14986 ( .A1(n12452), .A2(n16122), .ZN(n11838) );
  INV_X1 U14987 ( .A(n16111), .ZN(n11839) );
  NAND2_X1 U14988 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  XNOR2_X1 U14989 ( .A(n11843), .B(n11842), .ZN(n12438) );
  NAND2_X1 U14990 ( .A1(n12438), .A2(n19484), .ZN(n11853) );
  NAND2_X1 U14991 ( .A1(n16281), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12446) );
  OAI21_X1 U14992 ( .B1(n16283), .B2(n21415), .A(n12446), .ZN(n11851) );
  NAND2_X1 U14993 ( .A1(n10575), .A2(n11848), .ZN(n11849) );
  NAND2_X1 U14994 ( .A1(n11697), .A2(n11849), .ZN(n19311) );
  NOR2_X1 U14995 ( .A1(n19311), .A2(n16287), .ZN(n11850) );
  AOI211_X1 U14996 ( .C1(n19487), .C2(n19306), .A(n11851), .B(n11850), .ZN(
        n11852) );
  INV_X1 U14997 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18441) );
  NAND2_X1 U14998 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18477) );
  INV_X1 U14999 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18154) );
  NOR2_X1 U15000 ( .A1(n18477), .A2(n18154), .ZN(n18480) );
  AOI22_X1 U15001 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U15002 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11858) );
  NOR2_X4 U15003 ( .A1(n11864), .A2(n11863), .ZN(n17597) );
  AOI22_X1 U15004 ( .A1(n16668), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17597), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11857) );
  CLKBUF_X3 U15005 ( .A(n11903), .Z(n17548) );
  CLKBUF_X3 U15006 ( .A(n11893), .Z(n17596) );
  AOI22_X1 U15007 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11856) );
  NAND4_X1 U15008 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(
        n11871) );
  AOI22_X1 U15009 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11869) );
  INV_X2 U15010 ( .A(n9720), .ZN(n17580) );
  AOI22_X1 U15011 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U15012 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17553), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11867) );
  INV_X4 U15013 ( .A(n17333), .ZN(n17616) );
  AOI22_X1 U15014 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U15015 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11870) );
  AOI22_X1 U15016 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15017 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11874) );
  INV_X2 U15018 ( .A(n17566), .ZN(n17618) );
  AOI22_X1 U15019 ( .A1(n16668), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U15020 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U15021 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11881) );
  BUF_X2 U15022 ( .A(n12001), .Z(n17612) );
  AOI22_X1 U15023 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U15024 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15025 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9724), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U15026 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11876) );
  NAND4_X1 U15027 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11880) );
  INV_X1 U15028 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n21458) );
  INV_X2 U15029 ( .A(n9720), .ZN(n17567) );
  AOI22_X1 U15030 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11882) );
  OAI21_X1 U15031 ( .B1(n9784), .B2(n21458), .A(n11882), .ZN(n11887) );
  AOI22_X1 U15032 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U15033 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U15034 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U15035 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9737), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U15036 ( .A1(n11970), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U15037 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11893), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11888) );
  INV_X1 U15038 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17654) );
  AOI22_X1 U15039 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9737), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17618), .ZN(n11897) );
  INV_X2 U15040 ( .A(n12532), .ZN(n17594) );
  AOI22_X1 U15041 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17594), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9729), .ZN(n11896) );
  AOI22_X1 U15042 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17563), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U15043 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11893), .ZN(n11894) );
  AOI22_X1 U15044 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17597), .ZN(n11900) );
  AND2_X1 U15045 ( .A1(n18288), .A2(n17808), .ZN(n11946) );
  OAI21_X1 U15046 ( .B1(n9720), .B2(n21268), .A(n11901), .ZN(n11902) );
  AOI22_X1 U15047 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17553), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U15048 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15049 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9727), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15050 ( .A1(n11970), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17597), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U15051 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U15052 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11893), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U15053 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15054 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U15055 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U15056 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11893), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U15057 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15058 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U15059 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U15060 ( .A1(n16668), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11915) );
  NOR2_X1 U15061 ( .A1(n11944), .A2(n17797), .ZN(n11943) );
  AOI22_X1 U15062 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15063 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11927) );
  INV_X1 U15064 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17645) );
  AOI22_X1 U15065 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11893), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11919) );
  OAI21_X1 U15066 ( .B1(n17333), .B2(n17645), .A(n11919), .ZN(n11925) );
  AOI22_X1 U15067 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U15068 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U15069 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9727), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U15070 ( .A1(n11970), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11920) );
  NAND4_X1 U15071 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(
        n11924) );
  AOI211_X1 U15072 ( .C1(n17615), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n11925), .B(n11924), .ZN(n11926) );
  NAND3_X1 U15073 ( .A1(n11928), .A2(n11927), .A3(n11926), .ZN(n12095) );
  NAND2_X1 U15074 ( .A1(n11943), .A2(n12095), .ZN(n11941) );
  NOR2_X1 U15075 ( .A1(n17790), .A2(n11941), .ZN(n11940) );
  AOI22_X1 U15076 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15077 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15078 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11929) );
  OAI21_X1 U15079 ( .B1(n10640), .B2(n21397), .A(n11929), .ZN(n11935) );
  AOI22_X1 U15080 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15081 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U15082 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U15083 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11930) );
  NAND4_X1 U15084 ( .A1(n11933), .A2(n11932), .A3(n11931), .A4(n11930), .ZN(
        n11934) );
  AOI211_X1 U15085 ( .C1(n9722), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n11935), .B(n11934), .ZN(n11936) );
  NAND3_X1 U15086 ( .A1(n11938), .A2(n11937), .A3(n11936), .ZN(n12096) );
  NAND2_X1 U15087 ( .A1(n11940), .A2(n12096), .ZN(n11939) );
  NOR2_X1 U15088 ( .A1(n17783), .A2(n11939), .ZN(n11960) );
  XNOR2_X1 U15089 ( .A(n11939), .B(n12582), .ZN(n18206) );
  XNOR2_X1 U15090 ( .A(n11940), .B(n17786), .ZN(n11954) );
  XOR2_X1 U15091 ( .A(n11941), .B(n17790), .Z(n11942) );
  NAND2_X1 U15092 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11942), .ZN(
        n11953) );
  XNOR2_X1 U15093 ( .A(n10560), .B(n11942), .ZN(n18231) );
  INV_X1 U15094 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18544) );
  INV_X1 U15095 ( .A(n12095), .ZN(n17793) );
  XNOR2_X1 U15096 ( .A(n11943), .B(n17793), .ZN(n18249) );
  XOR2_X1 U15097 ( .A(n17797), .B(n11944), .Z(n11945) );
  NAND2_X1 U15098 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11945), .ZN(
        n11951) );
  INV_X1 U15099 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18556) );
  XNOR2_X1 U15100 ( .A(n18556), .B(n11945), .ZN(n18554) );
  INV_X1 U15101 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18580) );
  XNOR2_X1 U15102 ( .A(n17800), .B(n11946), .ZN(n11947) );
  OR2_X1 U15103 ( .A1(n18580), .A2(n11947), .ZN(n11950) );
  XNOR2_X1 U15104 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11947), .ZN(
        n18270) );
  AOI21_X1 U15105 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17808), .A(
        n18288), .ZN(n11949) );
  INV_X1 U15106 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19237) );
  NOR2_X1 U15107 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17808), .ZN(
        n11948) );
  AOI221_X1 U15108 ( .B1(n18288), .B2(n17808), .C1(n11949), .C2(n19237), .A(
        n11948), .ZN(n18269) );
  NAND2_X1 U15109 ( .A1(n18270), .A2(n18269), .ZN(n18268) );
  NAND2_X1 U15110 ( .A1(n11950), .A2(n18268), .ZN(n18553) );
  NAND2_X1 U15111 ( .A1(n18554), .A2(n18553), .ZN(n18552) );
  NAND2_X1 U15112 ( .A1(n11951), .A2(n18552), .ZN(n18248) );
  NAND2_X1 U15113 ( .A1(n18249), .A2(n18248), .ZN(n11952) );
  NOR2_X1 U15114 ( .A1(n18249), .A2(n18248), .ZN(n18247) );
  AOI21_X2 U15115 ( .B1(n18544), .B2(n11952), .A(n18247), .ZN(n18230) );
  NAND2_X1 U15116 ( .A1(n18231), .A2(n18230), .ZN(n18229) );
  NAND2_X1 U15117 ( .A1(n11953), .A2(n18229), .ZN(n11955) );
  NAND2_X1 U15118 ( .A1(n11954), .A2(n11955), .ZN(n11956) );
  XOR2_X1 U15119 ( .A(n11955), .B(n11954), .Z(n18224) );
  INV_X1 U15120 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18504) );
  NAND2_X1 U15121 ( .A1(n11960), .A2(n11957), .ZN(n11961) );
  NAND2_X1 U15122 ( .A1(n18206), .A2(n18207), .ZN(n18205) );
  NAND2_X1 U15123 ( .A1(n11960), .A2(n11959), .ZN(n11958) );
  OAI211_X1 U15124 ( .C1(n11960), .C2(n11959), .A(n18205), .B(n11958), .ZN(
        n18191) );
  NAND2_X1 U15125 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18191), .ZN(
        n18190) );
  NAND2_X2 U15126 ( .A1(n11961), .A2(n18190), .ZN(n16901) );
  INV_X1 U15127 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18135) );
  INV_X1 U15128 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18338) );
  NAND2_X1 U15129 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18067) );
  INV_X1 U15130 ( .A(n18067), .ZN(n18390) );
  NAND2_X1 U15131 ( .A1(n18390), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18368) );
  INV_X1 U15132 ( .A(n18368), .ZN(n18366) );
  INV_X1 U15133 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18357) );
  NAND2_X1 U15134 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18031) );
  NOR2_X1 U15135 ( .A1(n18357), .A2(n18031), .ZN(n18359) );
  NAND2_X1 U15136 ( .A1(n18366), .A2(n18359), .ZN(n18354) );
  INV_X1 U15137 ( .A(n18354), .ZN(n16903) );
  NAND2_X1 U15138 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16903), .ZN(
        n18344) );
  NOR2_X1 U15139 ( .A1(n18338), .A2(n18344), .ZN(n17982) );
  INV_X1 U15140 ( .A(n17982), .ZN(n17984) );
  INV_X1 U15141 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18296) );
  NOR2_X1 U15142 ( .A1(n17984), .A2(n18296), .ZN(n18321) );
  INV_X1 U15143 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18322) );
  INV_X1 U15144 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18317) );
  NOR2_X1 U15145 ( .A1(n18322), .A2(n18317), .ZN(n18301) );
  INV_X1 U15146 ( .A(n18301), .ZN(n11962) );
  INV_X1 U15147 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18307) );
  INV_X1 U15148 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17921) );
  NOR2_X1 U15149 ( .A1(n18307), .A2(n17921), .ZN(n12128) );
  NAND2_X1 U15150 ( .A1(n18303), .A2(n12128), .ZN(n16867) );
  INV_X1 U15151 ( .A(n16867), .ZN(n16894) );
  AOI22_X1 U15152 ( .A1(n17597), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15153 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15154 ( .A1(n17594), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15155 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U15156 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U15157 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15158 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15159 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U15160 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16668), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15161 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11971) );
  NAND4_X1 U15162 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(
        n11980) );
  AOI22_X1 U15163 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15164 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9728), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15165 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15166 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U15167 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  AOI22_X1 U15168 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17597), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15169 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U15170 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11981) );
  OAI21_X1 U15171 ( .B1(n17505), .B2(n21397), .A(n11981), .ZN(n11984) );
  AOI22_X1 U15172 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15173 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17553), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15174 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15175 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15176 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15177 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11987) );
  NAND4_X1 U15178 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11996) );
  AOI22_X1 U15179 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15180 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15181 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15182 ( .A1(n16668), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11991) );
  NAND4_X1 U15183 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n11995) );
  AOI22_X1 U15184 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15185 ( .A1(n16668), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15186 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15187 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11997) );
  NAND4_X1 U15188 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12007) );
  AOI22_X1 U15189 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U15190 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15191 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15192 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12002) );
  NAND4_X1 U15193 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12006) );
  NOR2_X2 U15194 ( .A1(n12007), .A2(n12006), .ZN(n18645) );
  AOI22_X1 U15195 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15196 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15197 ( .A1(n16668), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U15198 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15199 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15200 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9725), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15201 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15202 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15203 ( .A1(n16668), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15204 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15205 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12015) );
  NAND4_X1 U15206 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12024) );
  AOI22_X1 U15207 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15208 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15209 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15210 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12019) );
  NAND4_X1 U15211 ( .A1(n12022), .A2(n12021), .A3(n12020), .A4(n12019), .ZN(
        n12023) );
  NOR2_X1 U15212 ( .A1(n12024), .A2(n12023), .ZN(n18629) );
  AOI22_X1 U15213 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15214 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15215 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12025) );
  OAI21_X1 U15216 ( .B1(n9784), .B2(n21268), .A(n12025), .ZN(n12031) );
  AOI22_X1 U15217 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15218 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15219 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15220 ( .A1(n17596), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U15221 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12030) );
  AOI211_X1 U15222 ( .C1(n16668), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n12031), .B(n12030), .ZN(n12032) );
  NAND3_X1 U15223 ( .A1(n12034), .A2(n12033), .A3(n12032), .ZN(n12077) );
  INV_X1 U15224 ( .A(n12086), .ZN(n12080) );
  NAND3_X1 U15225 ( .A1(n18625), .A2(n18640), .A3(n18632), .ZN(n12044) );
  INV_X1 U15226 ( .A(n18645), .ZN(n17749) );
  INV_X1 U15227 ( .A(n16778), .ZN(n19063) );
  NAND2_X1 U15228 ( .A1(n18621), .A2(n17815), .ZN(n12083) );
  AOI21_X1 U15229 ( .B1(n17749), .B2(n19063), .A(n12083), .ZN(n12072) );
  AOI21_X1 U15230 ( .B1(n12080), .B2(n12044), .A(n12072), .ZN(n12043) );
  NAND2_X1 U15231 ( .A1(n12086), .A2(n12085), .ZN(n12068) );
  AOI21_X1 U15232 ( .B1(n12044), .B2(n12068), .A(n17815), .ZN(n12042) );
  INV_X1 U15233 ( .A(n12035), .ZN(n12048) );
  AOI22_X1 U15234 ( .A1(n12048), .A2(n18629), .B1(n18632), .B2(n16778), .ZN(
        n12036) );
  INV_X1 U15235 ( .A(n12036), .ZN(n12041) );
  NAND2_X1 U15236 ( .A1(n12084), .A2(n18625), .ZN(n12071) );
  INV_X1 U15237 ( .A(n12071), .ZN(n12037) );
  OAI22_X1 U15238 ( .A1(n18632), .A2(n12039), .B1(n12038), .B2(n12037), .ZN(
        n12040) );
  NOR2_X2 U15239 ( .A1(n12046), .A2(n12089), .ZN(n16687) );
  NAND2_X1 U15240 ( .A1(n18629), .A2(n18625), .ZN(n12087) );
  NAND2_X1 U15241 ( .A1(n18636), .A2(n12085), .ZN(n12069) );
  NAND2_X1 U15242 ( .A1(n18621), .A2(n12478), .ZN(n12047) );
  INV_X1 U15243 ( .A(n12044), .ZN(n12045) );
  NAND2_X1 U15244 ( .A1(n18625), .A2(n19260), .ZN(n12078) );
  NOR2_X1 U15245 ( .A1(n18640), .A2(n12078), .ZN(n12094) );
  OAI22_X1 U15246 ( .A1(n19226), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18613), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12054) );
  INV_X1 U15247 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18611) );
  OAI22_X1 U15248 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18611), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12051), .ZN(n12057) );
  NOR2_X1 U15249 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18611), .ZN(
        n12052) );
  NAND2_X1 U15250 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12051), .ZN(
        n12058) );
  AOI22_X1 U15251 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12057), .B1(
        n12052), .B2(n12058), .ZN(n12062) );
  NAND2_X1 U15252 ( .A1(n12055), .A2(n12054), .ZN(n12053) );
  OAI211_X1 U15253 ( .C1(n12055), .C2(n12054), .A(n12062), .B(n12053), .ZN(
        n12064) );
  OAI21_X1 U15254 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19066), .A(
        n12056), .ZN(n12067) );
  XNOR2_X1 U15255 ( .A(n12056), .B(n12061), .ZN(n12060) );
  AOI21_X1 U15256 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12058), .A(
        n12057), .ZN(n12059) );
  OAI21_X1 U15257 ( .B1(n12064), .B2(n12067), .A(n19054), .ZN(n12581) );
  INV_X1 U15258 ( .A(n12581), .ZN(n19056) );
  INV_X1 U15259 ( .A(n12061), .ZN(n12063) );
  NAND2_X1 U15260 ( .A1(n12063), .A2(n12062), .ZN(n12066) );
  AOI21_X1 U15261 ( .B1(n18632), .B2(n12068), .A(n19059), .ZN(n12076) );
  OAI211_X1 U15262 ( .C1(n18632), .C2(n16778), .A(n12090), .B(n12069), .ZN(
        n12070) );
  NOR2_X1 U15263 ( .A1(n12071), .A2(n12070), .ZN(n12093) );
  INV_X1 U15264 ( .A(n12072), .ZN(n12073) );
  OAI211_X1 U15265 ( .C1(n12075), .C2(n12093), .A(n12074), .B(n12073), .ZN(
        n16693) );
  NAND2_X1 U15266 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19134), .ZN(n19270) );
  INV_X2 U15267 ( .A(n19270), .ZN(n19272) );
  NOR2_X1 U15268 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17000) );
  INV_X1 U15269 ( .A(n17000), .ZN(n19124) );
  AOI21_X1 U15270 ( .B1(n18621), .B2(n12077), .A(n19259), .ZN(n12079) );
  NAND2_X1 U15271 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19254) );
  INV_X1 U15272 ( .A(n19254), .ZN(n19261) );
  AOI21_X1 U15273 ( .B1(n12079), .B2(n12078), .A(n19261), .ZN(n17003) );
  NAND3_X1 U15274 ( .A1(n19054), .A2(n17003), .A3(n12080), .ZN(n12081) );
  NAND2_X1 U15275 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19221), .ZN(n19105) );
  NAND2_X1 U15276 ( .A1(n12084), .A2(n12083), .ZN(n19275) );
  NOR2_X1 U15277 ( .A1(n18632), .A2(n12085), .ZN(n19074) );
  NAND3_X1 U15278 ( .A1(n19074), .A2(n12086), .A3(n12090), .ZN(n12476) );
  INV_X1 U15279 ( .A(n12087), .ZN(n19073) );
  INV_X1 U15280 ( .A(n12089), .ZN(n12092) );
  NAND3_X1 U15281 ( .A1(n10317), .A2(n19260), .A3(n12623), .ZN(n12091) );
  INV_X1 U15282 ( .A(n19064), .ZN(n18462) );
  NAND3_X1 U15283 ( .A1(n9780), .A2(n18595), .A3(n18587), .ZN(n18545) );
  NAND2_X1 U15284 ( .A1(n12094), .A2(n12093), .ZN(n19055) );
  NOR2_X1 U15285 ( .A1(n19055), .A2(n12582), .ZN(n18452) );
  INV_X1 U15286 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18423) );
  NAND2_X1 U15287 ( .A1(n12103), .A2(n12095), .ZN(n12108) );
  INV_X1 U15288 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21317) );
  NOR2_X1 U15289 ( .A1(n17808), .A2(n21317), .ZN(n12097) );
  NOR2_X1 U15290 ( .A1(n18280), .A2(n18287), .ZN(n18279) );
  NOR2_X1 U15291 ( .A1(n12097), .A2(n18279), .ZN(n18267) );
  NOR2_X1 U15292 ( .A1(n18580), .A2(n12099), .ZN(n12100) );
  NAND2_X1 U15293 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  XNOR2_X1 U15294 ( .A(n12114), .B(n12113), .ZN(n18214) );
  INV_X1 U15295 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12116) );
  NOR2_X1 U15296 ( .A1(n18199), .A2(n18509), .ZN(n18198) );
  NOR2_X4 U15297 ( .A1(n18198), .A2(n12116), .ZN(n18475) );
  NAND2_X1 U15298 ( .A1(n18436), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18438) );
  NOR2_X1 U15299 ( .A1(n18441), .A2(n18438), .ZN(n18415) );
  INV_X1 U15300 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21331) );
  NAND3_X1 U15301 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n18301), .ZN(n18295) );
  NOR2_X1 U15302 ( .A1(n21331), .A2(n18295), .ZN(n16900) );
  AND3_X1 U15303 ( .A1(n16903), .A2(n12128), .A3(n16900), .ZN(n12586) );
  INV_X1 U15304 ( .A(n19060), .ZN(n19088) );
  NAND2_X1 U15305 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18415), .ZN(
        n18400) );
  AOI21_X1 U15306 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18500) );
  NOR3_X1 U15307 ( .A1(n10560), .A2(n18556), .A3(n18544), .ZN(n18503) );
  NOR3_X1 U15308 ( .A1(n18504), .A2(n10171), .A3(n12116), .ZN(n18397) );
  NAND2_X1 U15309 ( .A1(n18503), .A2(n18397), .ZN(n12117) );
  OR2_X1 U15310 ( .A1(n18500), .A2(n12117), .ZN(n18412) );
  NOR2_X1 U15311 ( .A1(n18400), .A2(n18412), .ZN(n18391) );
  INV_X1 U15312 ( .A(n18391), .ZN(n12132) );
  INV_X1 U15313 ( .A(n9780), .ZN(n19080) );
  OAI21_X1 U15314 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19080), .A(
        n18502), .ZN(n18564) );
  INV_X1 U15315 ( .A(n18400), .ZN(n16902) );
  NAND2_X1 U15316 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18501) );
  NOR2_X1 U15317 ( .A1(n18501), .A2(n12117), .ZN(n12134) );
  NAND2_X1 U15318 ( .A1(n16902), .A2(n12134), .ZN(n18389) );
  OAI22_X1 U15319 ( .A1(n19088), .A2(n12132), .B1(n18564), .B2(n18389), .ZN(
        n18320) );
  NAND2_X1 U15320 ( .A1(n12586), .A2(n18320), .ZN(n16882) );
  OAI21_X1 U15321 ( .B1(n18508), .B2(n16896), .A(n16882), .ZN(n12118) );
  AOI22_X1 U15322 ( .A1(n16894), .A2(n18598), .B1(n18595), .B2(n12118), .ZN(
        n16708) );
  INV_X1 U15323 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16861) );
  NAND2_X1 U15324 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16861), .ZN(
        n12589) );
  NOR4_X1 U15325 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12121) );
  INV_X1 U15326 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12120) );
  INV_X1 U15327 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12119) );
  INV_X1 U15328 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18417) );
  NAND2_X1 U15329 ( .A1(n18199), .A2(n18417), .ZN(n12122) );
  AND3_X2 U15330 ( .A1(n10243), .A2(n12123), .A3(n12122), .ZN(n18076) );
  INV_X1 U15331 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18396) );
  NOR2_X2 U15332 ( .A1(n18012), .A2(n21331), .ZN(n17988) );
  INV_X1 U15333 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18071) );
  NAND2_X1 U15334 ( .A1(n18071), .A2(n18117), .ZN(n18065) );
  INV_X1 U15335 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18040) );
  NAND2_X1 U15336 ( .A1(n18037), .A2(n18040), .ZN(n18029) );
  NAND3_X1 U15337 ( .A1(n18010), .A2(n18338), .A3(n21331), .ZN(n12124) );
  NAND3_X1 U15338 ( .A1(n17988), .A2(n17975), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12127) );
  NAND2_X1 U15339 ( .A1(n12128), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12137) );
  INV_X1 U15340 ( .A(n12137), .ZN(n12131) );
  AOI21_X1 U15341 ( .B1(n12129), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16850), .ZN(n12584) );
  NOR2_X1 U15342 ( .A1(n17783), .A2(n19055), .ZN(n18514) );
  NAND2_X1 U15343 ( .A1(n18595), .A2(n18514), .ZN(n18485) );
  OAI22_X1 U15344 ( .A1(n16708), .A2(n12589), .B1(n12584), .B2(n18485), .ZN(
        n12130) );
  INV_X1 U15345 ( .A(n12130), .ZN(n12140) );
  NOR2_X1 U15346 ( .A1(n18586), .A2(n18508), .ZN(n18318) );
  NAND2_X1 U15347 ( .A1(n18303), .A2(n12131), .ZN(n16859) );
  INV_X1 U15348 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19212) );
  NAND2_X1 U15349 ( .A1(n19221), .A2(n19212), .ZN(n19216) );
  INV_X1 U15350 ( .A(n19216), .ZN(n19274) );
  INV_X1 U15351 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19263) );
  OR2_X1 U15352 ( .A1(n18344), .A2(n18389), .ZN(n18298) );
  NOR2_X1 U15353 ( .A1(n18295), .A2(n18298), .ZN(n12136) );
  AOI21_X1 U15354 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16900), .A(
        n19064), .ZN(n12133) );
  OAI21_X1 U15355 ( .B1(n18344), .B2(n12132), .A(n19060), .ZN(n18299) );
  INV_X1 U15356 ( .A(n18299), .ZN(n18339) );
  AOI211_X1 U15357 ( .C1(n19060), .C2(n18295), .A(n12133), .B(n18339), .ZN(
        n12135) );
  INV_X1 U15358 ( .A(n12134), .ZN(n18411) );
  NOR2_X1 U15359 ( .A1(n19237), .A2(n18411), .ZN(n18471) );
  NAND2_X1 U15360 ( .A1(n16902), .A2(n18471), .ZN(n18413) );
  OAI21_X1 U15361 ( .B1(n18354), .B2(n18413), .A(n18462), .ZN(n18297) );
  OAI211_X1 U15362 ( .C1(n9780), .C2(n12136), .A(n12135), .B(n18297), .ZN(
        n16700) );
  INV_X1 U15363 ( .A(n9743), .ZN(n18505) );
  OAI211_X1 U15364 ( .C1(n16700), .C2(n12137), .A(n18505), .B(n18595), .ZN(
        n16884) );
  NAND2_X1 U15365 ( .A1(n9732), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n12593) );
  NAND2_X1 U15366 ( .A1(n12140), .A2(n10667), .ZN(P3_U2832) );
  OAI21_X1 U15367 ( .B1(n19541), .B2(n11619), .A(n19977), .ZN(n12161) );
  NOR2_X1 U15368 ( .A1(n20196), .A2(n20205), .ZN(n19975) );
  NAND2_X1 U15369 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19975), .ZN(
        n12158) );
  INV_X1 U15370 ( .A(n12158), .ZN(n12142) );
  NAND2_X1 U15371 ( .A1(n12142), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20030) );
  OAI211_X1 U15372 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n12142), .A(
        n20030), .B(n20180), .ZN(n12143) );
  INV_X1 U15373 ( .A(n12143), .ZN(n12144) );
  AOI21_X1 U15374 ( .B1(n12161), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12144), .ZN(n12145) );
  OAI21_X2 U15375 ( .B1(n13436), .B2(n12163), .A(n12145), .ZN(n12172) );
  INV_X1 U15376 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12147) );
  INV_X1 U15378 ( .A(n12163), .ZN(n12152) );
  NAND2_X1 U15379 ( .A1(n12161), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12150) );
  NAND2_X1 U15380 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n12154), .ZN(
        n19848) );
  NAND2_X1 U15381 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20205), .ZN(
        n19805) );
  NAND2_X1 U15382 ( .A1(n19848), .A2(n19805), .ZN(n19651) );
  NAND2_X1 U15383 ( .A1(n20180), .A2(n19651), .ZN(n19850) );
  NAND2_X1 U15384 ( .A1(n12150), .A2(n19850), .ZN(n12151) );
  AOI22_X1 U15385 ( .A1(n12161), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20180), .B2(n12154), .ZN(n12155) );
  NAND2_X1 U15386 ( .A1(n13490), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12156) );
  NAND2_X1 U15387 ( .A1(n13290), .A2(n13291), .ZN(n13289) );
  NAND2_X1 U15388 ( .A1(n13066), .A2(n12156), .ZN(n12157) );
  INV_X1 U15389 ( .A(n20180), .ZN(n20176) );
  NAND2_X1 U15390 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19743) );
  NAND2_X1 U15391 ( .A1(n19743), .A2(n20196), .ZN(n12159) );
  NAND2_X1 U15392 ( .A1(n12159), .A2(n12158), .ZN(n19652) );
  NOR2_X1 U15393 ( .A1(n20176), .A2(n19652), .ZN(n12160) );
  AOI21_X1 U15394 ( .B1(n12161), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12160), .ZN(n12162) );
  NAND2_X1 U15395 ( .A1(n13490), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12165) );
  NAND2_X1 U15396 ( .A1(n13312), .A2(n13313), .ZN(n13311) );
  INV_X1 U15397 ( .A(n12165), .ZN(n12166) );
  NAND2_X1 U15398 ( .A1(n12167), .A2(n12166), .ZN(n12168) );
  NAND2_X1 U15399 ( .A1(n13311), .A2(n12168), .ZN(n13435) );
  NAND2_X1 U15400 ( .A1(n21501), .A2(n13435), .ZN(n12171) );
  NAND2_X1 U15401 ( .A1(n12169), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12170) );
  NAND2_X1 U15402 ( .A1(n12171), .A2(n12170), .ZN(n13495) );
  NAND2_X1 U15403 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13600) );
  NAND2_X1 U15404 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12174) );
  NOR2_X1 U15405 ( .A1(n13600), .A2(n12174), .ZN(n12175) );
  NAND4_X1 U15406 ( .A1(n13759), .A2(n13755), .A3(n13782), .A4(n12175), .ZN(
        n12176) );
  NOR2_X1 U15407 ( .A1(n14515), .A2(n12176), .ZN(n12177) );
  INV_X1 U15408 ( .A(n13792), .ZN(n12178) );
  NOR2_X2 U15409 ( .A1(n13743), .A2(n12178), .ZN(n13790) );
  AND2_X2 U15410 ( .A1(n13790), .A2(n13803), .ZN(n13801) );
  AOI22_X1 U15411 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n10936), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15412 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12257), .B1(
        n12256), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15413 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12180) );
  NAND4_X1 U15414 ( .A1(n12183), .A2(n12182), .A3(n12181), .A4(n12180), .ZN(
        n12189) );
  AOI22_X1 U15415 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15416 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15417 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15418 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12184) );
  NAND4_X1 U15419 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n12188) );
  OR2_X1 U15420 ( .A1(n12189), .A2(n12188), .ZN(n15900) );
  AOI22_X1 U15421 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10937), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15422 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12257), .B1(
        n12256), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15423 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12190) );
  NAND4_X1 U15424 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12199) );
  AOI22_X1 U15425 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15426 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15427 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15428 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12194) );
  NAND4_X1 U15429 ( .A1(n12197), .A2(n12196), .A3(n12195), .A4(n12194), .ZN(
        n12198) );
  OR2_X1 U15430 ( .A1(n12199), .A2(n12198), .ZN(n15891) );
  AOI22_X1 U15431 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10884), .B1(
        n10089), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15432 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10937), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15433 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12257), .B1(
        n12256), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15434 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U15435 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12209) );
  AOI22_X1 U15436 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15437 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15438 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15439 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U15440 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12208) );
  OR2_X1 U15441 ( .A1(n12209), .A2(n12208), .ZN(n15885) );
  INV_X1 U15442 ( .A(n15885), .ZN(n12210) );
  NOR2_X2 U15443 ( .A1(n15883), .A2(n12210), .ZN(n15878) );
  AOI22_X1 U15444 ( .A1(n10936), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15445 ( .A1(n12256), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15446 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12211) );
  NAND4_X1 U15447 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12220) );
  AOI22_X1 U15448 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15449 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15450 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15451 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12215) );
  NAND4_X1 U15452 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12219) );
  OR2_X1 U15453 ( .A1(n12220), .A2(n12219), .ZN(n15880) );
  NAND2_X1 U15454 ( .A1(n15878), .A2(n15880), .ZN(n15873) );
  AOI22_X1 U15455 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10884), .B1(
        n10089), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15456 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10937), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15457 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12257), .B1(
        n12256), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15458 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12221) );
  NAND4_X1 U15459 ( .A1(n12224), .A2(n12223), .A3(n12222), .A4(n12221), .ZN(
        n12230) );
  AOI22_X1 U15460 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15461 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15462 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15463 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U15464 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12229) );
  NOR2_X1 U15465 ( .A1(n12230), .A2(n12229), .ZN(n15874) );
  AOI22_X1 U15466 ( .A1(n10936), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15467 ( .A1(n12256), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12257), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15468 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12231) );
  NAND4_X1 U15469 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n12240) );
  AOI22_X1 U15470 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15471 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15472 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15473 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12235) );
  NAND4_X1 U15474 ( .A1(n12238), .A2(n12237), .A3(n12236), .A4(n12235), .ZN(
        n12239) );
  OR2_X1 U15475 ( .A1(n12240), .A2(n12239), .ZN(n15870) );
  AOI22_X1 U15476 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10884), .B1(
        n10089), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15477 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10936), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15478 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12257), .B1(
        n12256), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15479 ( .A1(n10882), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12241) );
  NAND4_X1 U15480 ( .A1(n12244), .A2(n12243), .A3(n12242), .A4(n12241), .ZN(
        n12250) );
  AOI22_X1 U15481 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10885), .B1(
        n10862), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15482 ( .A1(n10912), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15483 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15484 ( .A1(n11246), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12245) );
  NAND4_X1 U15485 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(
        n12249) );
  OR2_X1 U15486 ( .A1(n12250), .A2(n12249), .ZN(n15861) );
  AOI22_X1 U15487 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11246), .B1(
        n10912), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15488 ( .A1(n10862), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15489 ( .A1(n10885), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10864), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12252) );
  NAND4_X1 U15490 ( .A1(n12255), .A2(n12254), .A3(n12253), .A4(n12252), .ZN(
        n12263) );
  AOI22_X1 U15491 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10872), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15492 ( .A1(n10883), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10911), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15493 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12256), .B1(
        n10936), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15494 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12257), .B1(
        n10937), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15495 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12262) );
  NOR2_X1 U15496 ( .A1(n12263), .A2(n12262), .ZN(n12295) );
  AOI22_X1 U15497 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12395), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15498 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12368), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12271) );
  XNOR2_X1 U15499 ( .A(n10789), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12403) );
  INV_X1 U15500 ( .A(n12265), .ZN(n13641) );
  INV_X1 U15501 ( .A(n13641), .ZN(n13631) );
  NAND2_X1 U15502 ( .A1(n13631), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U15503 ( .A1(n12398), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12268) );
  NAND2_X1 U15504 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12266) );
  AND4_X1 U15505 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12266), .ZN(
        n12270) );
  NAND4_X1 U15506 ( .A1(n12272), .A2(n12271), .A3(n12403), .A4(n12270), .ZN(
        n12281) );
  AOI22_X1 U15507 ( .A1(n12393), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12395), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12279) );
  NAND2_X1 U15508 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12276) );
  NAND2_X1 U15509 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12274) );
  NAND2_X1 U15510 ( .A1(n13631), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12273) );
  AND4_X1 U15511 ( .A1(n12276), .A2(n12275), .A3(n12274), .A4(n12273), .ZN(
        n12278) );
  AOI22_X1 U15512 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12277) );
  INV_X1 U15513 ( .A(n12403), .ZN(n12390) );
  NAND4_X1 U15514 ( .A1(n12279), .A2(n12278), .A3(n12277), .A4(n12390), .ZN(
        n12280) );
  NAND2_X1 U15515 ( .A1(n12281), .A2(n12280), .ZN(n15846) );
  NOR2_X1 U15516 ( .A1(n19513), .A2(n15846), .ZN(n12282) );
  XOR2_X1 U15517 ( .A(n12295), .B(n12282), .Z(n15847) );
  AOI22_X1 U15518 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15519 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12283) );
  AND2_X1 U15520 ( .A1(n12284), .A2(n12283), .ZN(n12287) );
  AOI22_X1 U15521 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15522 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12285) );
  NAND4_X1 U15523 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12390), .ZN(
        n12294) );
  AOI22_X1 U15524 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15525 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12288) );
  AND2_X1 U15526 ( .A1(n12289), .A2(n12288), .ZN(n12292) );
  AOI22_X1 U15527 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15528 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12290) );
  NAND4_X1 U15529 ( .A1(n12292), .A2(n12403), .A3(n12291), .A4(n12290), .ZN(
        n12293) );
  AND2_X1 U15530 ( .A1(n12294), .A2(n12293), .ZN(n12299) );
  INV_X1 U15531 ( .A(n12299), .ZN(n12301) );
  INV_X1 U15532 ( .A(n12295), .ZN(n12297) );
  INV_X1 U15533 ( .A(n15846), .ZN(n12296) );
  NAND2_X1 U15534 ( .A1(n12297), .A2(n12296), .ZN(n12302) );
  XOR2_X1 U15535 ( .A(n12301), .B(n12302), .Z(n12298) );
  NAND2_X1 U15536 ( .A1(n12298), .A2(n13490), .ZN(n15848) );
  NOR2_X1 U15537 ( .A1(n15847), .A2(n15848), .ZN(n12300) );
  NAND2_X1 U15538 ( .A1(n19513), .A2(n12299), .ZN(n15849) );
  NOR2_X1 U15539 ( .A1(n12302), .A2(n12301), .ZN(n12315) );
  AOI22_X1 U15540 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12304) );
  AND2_X1 U15541 ( .A1(n12304), .A2(n12303), .ZN(n12307) );
  AOI22_X1 U15542 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15543 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12305) );
  NAND4_X1 U15544 ( .A1(n12307), .A2(n12306), .A3(n12305), .A4(n12390), .ZN(
        n12314) );
  AOI22_X1 U15545 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12309) );
  AND2_X1 U15546 ( .A1(n12309), .A2(n12308), .ZN(n12312) );
  AOI22_X1 U15547 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15548 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12310) );
  NAND4_X1 U15549 ( .A1(n12312), .A2(n12403), .A3(n12311), .A4(n12310), .ZN(
        n12313) );
  AND2_X1 U15550 ( .A1(n12314), .A2(n12313), .ZN(n12316) );
  NAND2_X1 U15551 ( .A1(n12315), .A2(n12316), .ZN(n12381) );
  OAI211_X1 U15552 ( .C1(n12315), .C2(n12316), .A(n12381), .B(n13490), .ZN(
        n12335) );
  XNOR2_X2 U15553 ( .A(n12336), .B(n12335), .ZN(n15832) );
  INV_X1 U15554 ( .A(n15832), .ZN(n12339) );
  NAND2_X1 U15555 ( .A1(n19513), .A2(n12316), .ZN(n15842) );
  INV_X1 U15556 ( .A(n15842), .ZN(n12334) );
  AOI22_X1 U15557 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12323) );
  NAND2_X1 U15558 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12320) );
  NAND2_X1 U15559 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12318) );
  NAND2_X1 U15560 ( .A1(n13631), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12317) );
  AND4_X1 U15561 ( .A1(n12320), .A2(n12319), .A3(n12318), .A4(n12317), .ZN(
        n12322) );
  AOI22_X1 U15562 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12321) );
  NAND4_X1 U15563 ( .A1(n12323), .A2(n12322), .A3(n12321), .A4(n12390), .ZN(
        n12332) );
  AOI22_X1 U15564 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U15565 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12327) );
  NAND2_X1 U15566 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12325) );
  NAND2_X1 U15567 ( .A1(n13631), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12324) );
  AND4_X1 U15568 ( .A1(n12327), .A2(n12326), .A3(n12325), .A4(n12324), .ZN(
        n12329) );
  AOI22_X1 U15569 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12328) );
  NAND4_X1 U15570 ( .A1(n12330), .A2(n12329), .A3(n12403), .A4(n12328), .ZN(
        n12331) );
  NAND2_X1 U15571 ( .A1(n12332), .A2(n12331), .ZN(n15834) );
  XNOR2_X1 U15572 ( .A(n12381), .B(n15834), .ZN(n12337) );
  NOR2_X1 U15573 ( .A1(n12337), .A2(n14515), .ZN(n15836) );
  AOI21_X2 U15574 ( .B1(n12339), .B2(n10641), .A(n12338), .ZN(n14514) );
  AOI22_X1 U15575 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12341) );
  AND2_X1 U15576 ( .A1(n12341), .A2(n12340), .ZN(n12344) );
  AOI22_X1 U15577 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15578 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12342) );
  NAND4_X1 U15579 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12390), .ZN(
        n12351) );
  AOI22_X1 U15580 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12346) );
  AND2_X1 U15581 ( .A1(n12346), .A2(n12345), .ZN(n12349) );
  AOI22_X1 U15582 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15583 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12347) );
  NAND4_X1 U15584 ( .A1(n12349), .A2(n12403), .A3(n12348), .A4(n12347), .ZN(
        n12350) );
  NAND2_X1 U15585 ( .A1(n12351), .A2(n12350), .ZN(n12382) );
  AOI22_X1 U15586 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12358) );
  NAND2_X1 U15587 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12355) );
  NAND2_X1 U15588 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12353) );
  NAND2_X1 U15589 ( .A1(n13631), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12352) );
  AND4_X1 U15590 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12357) );
  AOI22_X1 U15591 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12356) );
  NAND4_X1 U15592 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12390), .ZN(
        n12367) );
  AOI22_X1 U15593 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12365) );
  NAND2_X1 U15594 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12362) );
  NAND2_X1 U15595 ( .A1(n12400), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12361) );
  NAND2_X1 U15596 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12360) );
  NAND2_X1 U15597 ( .A1(n13631), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12359) );
  AND4_X1 U15598 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12364) );
  AOI22_X1 U15599 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12363) );
  NAND4_X1 U15600 ( .A1(n12365), .A2(n12364), .A3(n12403), .A4(n12363), .ZN(
        n12366) );
  NAND2_X1 U15601 ( .A1(n12367), .A2(n12366), .ZN(n14519) );
  AOI22_X1 U15602 ( .A1(n12368), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12370) );
  AND2_X1 U15603 ( .A1(n12370), .A2(n12369), .ZN(n12373) );
  AOI22_X1 U15604 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15605 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12371) );
  NAND4_X1 U15606 ( .A1(n12373), .A2(n12372), .A3(n12371), .A4(n12390), .ZN(
        n12380) );
  AOI22_X1 U15607 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15608 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12374) );
  AND2_X1 U15609 ( .A1(n12375), .A2(n12374), .ZN(n12378) );
  AOI22_X1 U15610 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15611 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12376) );
  NAND4_X1 U15612 ( .A1(n12378), .A2(n12403), .A3(n12377), .A4(n12376), .ZN(
        n12379) );
  NAND2_X1 U15613 ( .A1(n12380), .A2(n12379), .ZN(n12385) );
  OR2_X1 U15614 ( .A1(n12381), .A2(n15834), .ZN(n14516) );
  NOR2_X1 U15615 ( .A1(n14516), .A2(n14519), .ZN(n15825) );
  INV_X1 U15616 ( .A(n12382), .ZN(n15828) );
  AND2_X1 U15617 ( .A1(n13063), .A2(n15828), .ZN(n12383) );
  NAND2_X1 U15618 ( .A1(n15825), .A2(n12383), .ZN(n12384) );
  NOR2_X1 U15619 ( .A1(n12384), .A2(n12385), .ZN(n12386) );
  AOI21_X1 U15620 ( .B1(n12385), .B2(n12384), .A(n12386), .ZN(n15820) );
  INV_X1 U15621 ( .A(n12386), .ZN(n12387) );
  AOI22_X1 U15622 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15623 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12388) );
  NAND2_X1 U15624 ( .A1(n12389), .A2(n12388), .ZN(n12408) );
  AOI22_X1 U15625 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U15626 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12391) );
  NAND3_X1 U15627 ( .A1(n12392), .A2(n12391), .A3(n12390), .ZN(n12407) );
  AOI22_X1 U15628 ( .A1(n12394), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12393), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15629 ( .A1(n12395), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13631), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12396) );
  NAND2_X1 U15630 ( .A1(n12397), .A2(n12396), .ZN(n12406) );
  AOI22_X1 U15631 ( .A1(n12399), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12398), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15632 ( .A1(n12401), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12400), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12402) );
  NAND3_X1 U15633 ( .A1(n12404), .A2(n12403), .A3(n12402), .ZN(n12405) );
  OAI22_X1 U15634 ( .A1(n12408), .A2(n12407), .B1(n12406), .B2(n12405), .ZN(
        n12409) );
  NOR2_X1 U15635 ( .A1(n14550), .A2(n20103), .ZN(n12651) );
  INV_X1 U15636 ( .A(n12652), .ZN(n12410) );
  INV_X1 U15637 ( .A(n12411), .ZN(n12413) );
  NAND2_X1 U15638 ( .A1(n12413), .A2(n12412), .ZN(n12414) );
  NAND2_X1 U15639 ( .A1(n16017), .A2(n12415), .ZN(n16023) );
  INV_X1 U15640 ( .A(n13069), .ZN(n19548) );
  NAND2_X1 U15641 ( .A1(n16017), .A2(n19548), .ZN(n16014) );
  NOR2_X1 U15642 ( .A1(n12465), .A2(n16014), .ZN(n12436) );
  NOR2_X1 U15643 ( .A1(n19548), .A2(n19541), .ZN(n12416) );
  NOR4_X1 U15644 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12420) );
  NOR4_X1 U15645 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12419) );
  NOR4_X1 U15646 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12418) );
  NOR4_X1 U15647 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12417) );
  AND4_X1 U15648 ( .A1(n12420), .A2(n12419), .A3(n12418), .A4(n12417), .ZN(
        n12425) );
  NOR4_X1 U15649 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12423) );
  NOR4_X1 U15650 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12422) );
  NOR4_X1 U15651 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12421) );
  INV_X1 U15652 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20113) );
  AND4_X1 U15653 ( .A1(n12423), .A2(n12422), .A3(n12421), .A4(n20113), .ZN(
        n12424) );
  NAND2_X1 U15654 ( .A1(n12425), .A2(n12424), .ZN(n12426) );
  AND2_X2 U15655 ( .A1(n12426), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19499)
         );
  NAND2_X1 U15656 ( .A1(n12941), .A2(n19497), .ZN(n16007) );
  INV_X1 U15657 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n12431) );
  AND2_X1 U15658 ( .A1(n19534), .A2(n13069), .ZN(n12427) );
  INV_X1 U15659 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n12429) );
  NAND2_X1 U15660 ( .A1(n19499), .A2(BUF1_REG_14__SCAN_IN), .ZN(n12428) );
  OAI21_X1 U15661 ( .B1(n19499), .B2(n12429), .A(n12428), .ZN(n13624) );
  AOI22_X1 U15662 ( .A1(n15985), .A2(n13624), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19396), .ZN(n12430) );
  OAI21_X1 U15663 ( .B1(n16007), .B2(n12431), .A(n12430), .ZN(n12432) );
  INV_X1 U15664 ( .A(n12432), .ZN(n12434) );
  NAND2_X1 U15665 ( .A1(n16011), .A2(BUF1_REG_30__SCAN_IN), .ZN(n12433) );
  NAND2_X1 U15666 ( .A1(n12434), .A2(n12433), .ZN(n12435) );
  OAI21_X1 U15667 ( .B1(n10670), .B2(n16023), .A(n12437), .ZN(P2_U2889) );
  NAND2_X1 U15668 ( .A1(n12438), .A2(n16832), .ZN(n12449) );
  XOR2_X1 U15669 ( .A(n12441), .B(n12440), .Z(n19305) );
  INV_X1 U15670 ( .A(n12442), .ZN(n12444) );
  INV_X1 U15671 ( .A(n16381), .ZN(n12443) );
  OAI21_X1 U15672 ( .B1(n12444), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12443), .ZN(n12445) );
  OAI211_X1 U15673 ( .C1(n19311), .C2(n16836), .A(n12446), .B(n12445), .ZN(
        n12447) );
  AOI21_X1 U15674 ( .B1(n16838), .B2(n19305), .A(n12447), .ZN(n12448) );
  OR2_X1 U15675 ( .A1(n12454), .A2(n12455), .ZN(n12456) );
  AND2_X1 U15676 ( .A1(n12453), .A2(n12456), .ZN(n16411) );
  NAND2_X1 U15677 ( .A1(n19359), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16407) );
  NAND2_X1 U15678 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12457) );
  OAI211_X1 U15679 ( .C1(n15605), .C2(n19476), .A(n16407), .B(n12457), .ZN(
        n12458) );
  OAI21_X1 U15680 ( .B1(n16416), .B2(n16299), .A(n12459), .ZN(n12460) );
  INV_X1 U15681 ( .A(n12461), .ZN(n15503) );
  INV_X1 U15682 ( .A(n12601), .ZN(n12462) );
  AOI21_X1 U15683 ( .B1(n15503), .B2(n12462), .A(n19364), .ZN(n12464) );
  OAI21_X1 U15684 ( .B1(n12464), .B2(n19320), .A(n12463), .ZN(n12475) );
  INV_X1 U15685 ( .A(n12465), .ZN(n12466) );
  INV_X1 U15686 ( .A(n12467), .ZN(n12472) );
  INV_X1 U15687 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15688 ( .A1(n19315), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n19360), .ZN(n12468) );
  OAI21_X1 U15689 ( .B1(n19375), .B2(n12469), .A(n12468), .ZN(n12471) );
  NOR2_X1 U15690 ( .A1(n14544), .A2(n19368), .ZN(n12470) );
  AND2_X1 U15691 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17386) );
  AND2_X1 U15692 ( .A1(n18645), .A2(n18632), .ZN(n12477) );
  INV_X1 U15693 ( .A(n17655), .ZN(n17657) );
  NOR2_X1 U15694 ( .A1(n17749), .A2(n17657), .ZN(n16681) );
  AND2_X1 U15695 ( .A1(n17655), .A2(n17749), .ZN(n17658) );
  INV_X1 U15696 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17383) );
  NAND4_X1 U15697 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(P3_EBX_REG_2__SCAN_IN), .ZN(n17611) );
  INV_X1 U15698 ( .A(n17611), .ZN(n12479) );
  INV_X1 U15699 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n21399) );
  INV_X1 U15700 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17315) );
  NAND3_X1 U15701 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n17635), .ZN(n17593) );
  INV_X1 U15702 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17270) );
  INV_X1 U15703 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17243) );
  INV_X1 U15704 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17216) );
  INV_X1 U15705 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17194) );
  INV_X1 U15706 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17171) );
  INV_X1 U15707 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17149) );
  INV_X1 U15708 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17124) );
  INV_X1 U15709 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17382) );
  NAND2_X1 U15710 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17420), .ZN(n17412) );
  INV_X1 U15711 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17384) );
  NAND4_X1 U15712 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17420), .A3(n17386), 
        .A4(n17384), .ZN(n12564) );
  AOI22_X1 U15713 ( .A1(n17594), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15714 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17597), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15715 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15716 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12480) );
  NAND4_X1 U15717 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12489) );
  AOI22_X1 U15718 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15719 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15720 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U15721 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9725), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12484) );
  NAND4_X1 U15722 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12488) );
  NOR2_X1 U15723 ( .A1(n12489), .A2(n12488), .ZN(n17413) );
  AOI22_X1 U15724 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15725 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15726 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17616), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15727 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17594), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12490) );
  NAND4_X1 U15728 ( .A1(n12493), .A2(n12492), .A3(n12491), .A4(n12490), .ZN(
        n12499) );
  AOI22_X1 U15729 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17597), .ZN(n12497) );
  AOI22_X1 U15730 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9722), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15731 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9728), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n16674), .ZN(n12495) );
  AOI22_X1 U15732 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9724), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12494) );
  NAND4_X1 U15733 ( .A1(n12497), .A2(n12496), .A3(n12495), .A4(n12494), .ZN(
        n12498) );
  NOR2_X1 U15734 ( .A1(n12499), .A2(n12498), .ZN(n17421) );
  AOI22_X1 U15735 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U15736 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12509) );
  AOI22_X1 U15737 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12501) );
  OAI21_X1 U15738 ( .B1(n10640), .B2(n21458), .A(n12501), .ZN(n12507) );
  AOI22_X1 U15739 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17597), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15740 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15741 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U15742 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17602), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12502) );
  NAND4_X1 U15743 ( .A1(n12505), .A2(n12504), .A3(n12503), .A4(n12502), .ZN(
        n12506) );
  AOI211_X1 U15744 ( .C1(n9722), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n12507), .B(n12506), .ZN(n12508) );
  NAND3_X1 U15745 ( .A1(n12510), .A2(n12509), .A3(n12508), .ZN(n17425) );
  AOI22_X1 U15746 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17597), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U15747 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12519) );
  INV_X1 U15748 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U15749 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9724), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12511) );
  OAI21_X1 U15750 ( .B1(n10640), .B2(n17393), .A(n12511), .ZN(n12517) );
  AOI22_X1 U15751 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15752 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U15753 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15754 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12512) );
  NAND4_X1 U15755 ( .A1(n12515), .A2(n12514), .A3(n12513), .A4(n12512), .ZN(
        n12516) );
  AOI211_X1 U15756 ( .C1(n17602), .C2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n12517), .B(n12516), .ZN(n12518) );
  NAND3_X1 U15757 ( .A1(n12520), .A2(n12519), .A3(n12518), .ZN(n17426) );
  NAND2_X1 U15758 ( .A1(n17425), .A2(n17426), .ZN(n17424) );
  NOR2_X1 U15759 ( .A1(n17421), .A2(n17424), .ZN(n17418) );
  AOI22_X1 U15760 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15761 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15762 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12521) );
  OAI21_X1 U15763 ( .B1(n17533), .B2(n21268), .A(n12521), .ZN(n12527) );
  AOI22_X1 U15764 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15765 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15766 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15767 ( .A1(n17596), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12522) );
  NAND4_X1 U15768 ( .A1(n12525), .A2(n12524), .A3(n12523), .A4(n12522), .ZN(
        n12526) );
  AOI211_X1 U15769 ( .C1(n17553), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n12527), .B(n12526), .ZN(n12528) );
  NAND3_X1 U15770 ( .A1(n12530), .A2(n12529), .A3(n12528), .ZN(n17417) );
  NAND2_X1 U15771 ( .A1(n17418), .A2(n17417), .ZN(n17416) );
  NOR2_X1 U15772 ( .A1(n17413), .A2(n17416), .ZN(n17683) );
  AOI22_X1 U15773 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12541) );
  AOI22_X1 U15774 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U15775 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12531) );
  OAI21_X1 U15776 ( .B1(n12532), .B2(n17645), .A(n12531), .ZN(n12538) );
  AOI22_X1 U15777 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15778 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12535) );
  AOI22_X1 U15779 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U15780 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12533) );
  NAND4_X1 U15781 ( .A1(n12536), .A2(n12535), .A3(n12534), .A4(n12533), .ZN(
        n12537) );
  AOI211_X1 U15782 ( .C1(n17615), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n12538), .B(n12537), .ZN(n12539) );
  NAND3_X1 U15783 ( .A1(n12541), .A2(n12540), .A3(n12539), .ZN(n17682) );
  NAND2_X1 U15784 ( .A1(n17683), .A2(n17682), .ZN(n17681) );
  AOI22_X1 U15785 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9737), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15786 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15787 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15788 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12542) );
  NAND4_X1 U15789 ( .A1(n12545), .A2(n12544), .A3(n12543), .A4(n12542), .ZN(
        n12551) );
  AOI22_X1 U15790 ( .A1(n17597), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15791 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15792 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15793 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12546) );
  NAND4_X1 U15794 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12550) );
  NOR2_X1 U15795 ( .A1(n12551), .A2(n12550), .ZN(n17403) );
  NOR2_X1 U15796 ( .A1(n17681), .A2(n17403), .ZN(n12562) );
  AOI22_X1 U15797 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15798 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15799 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15800 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12552) );
  NAND4_X1 U15801 ( .A1(n12555), .A2(n12554), .A3(n12553), .A4(n12552), .ZN(
        n12561) );
  AOI22_X1 U15802 ( .A1(n9737), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15803 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9728), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15804 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15805 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12556) );
  NAND4_X1 U15806 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        n12560) );
  NOR2_X1 U15807 ( .A1(n12561), .A2(n12560), .ZN(n17404) );
  XNOR2_X1 U15808 ( .A(n12562), .B(n17404), .ZN(n17672) );
  NAND2_X1 U15809 ( .A1(n17658), .A2(n17672), .ZN(n12563) );
  AOI21_X1 U15810 ( .B1(n13817), .B2(P3_EBX_REG_29__SCAN_IN), .A(n12565), .ZN(
        n12566) );
  INV_X1 U15811 ( .A(n12566), .ZN(P3_U2674) );
  NAND2_X1 U15812 ( .A1(n12567), .A2(n16832), .ZN(n12580) );
  OAI21_X1 U15813 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16846), .A(
        n12568), .ZN(n12570) );
  AOI21_X1 U15814 ( .B1(n12570), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12569), .ZN(n12573) );
  NAND3_X1 U15815 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11819), .ZN(n12572) );
  OAI211_X1 U15816 ( .C1(n12574), .C2(n16836), .A(n12573), .B(n12572), .ZN(
        n12575) );
  AOI21_X1 U15817 ( .B1(n16838), .B2(n15910), .A(n12575), .ZN(n12579) );
  INV_X1 U15818 ( .A(n12576), .ZN(n12577) );
  NAND2_X1 U15819 ( .A1(n12577), .A2(n16640), .ZN(n12578) );
  NAND3_X1 U15820 ( .A1(n12580), .A2(n12579), .A3(n12578), .ZN(P2_U3015) );
  AOI22_X1 U15821 ( .A1(n18261), .A2(n16859), .B1(n18202), .B2(n16865), .ZN(
        n12583) );
  OAI22_X1 U15822 ( .A1(n12584), .A2(n18164), .B1(n12583), .B2(n16861), .ZN(
        n12585) );
  INV_X1 U15823 ( .A(n12585), .ZN(n12596) );
  AOI22_X2 U15824 ( .A1(n18202), .A2(n18475), .B1(n16901), .B2(n18261), .ZN(
        n18167) );
  NOR2_X4 U15825 ( .A1(n18167), .A2(n18400), .ZN(n18068) );
  NAND2_X1 U15826 ( .A1(n12586), .A2(n18068), .ZN(n12590) );
  NAND2_X1 U15827 ( .A1(n19273), .A2(n19212), .ZN(n16998) );
  NAND2_X1 U15828 ( .A1(n19216), .A2(n16998), .ZN(n18604) );
  INV_X1 U15829 ( .A(n18604), .ZN(n19257) );
  NAND2_X1 U15830 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18251) );
  INV_X1 U15832 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21384) );
  NOR2_X1 U15833 ( .A1(n18130), .A2(n18129), .ZN(n18128) );
  INV_X1 U15834 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18112) );
  INV_X1 U15835 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18072) );
  INV_X1 U15836 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17993) );
  INV_X1 U15837 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17952) );
  NAND2_X1 U15838 ( .A1(n12629), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17929) );
  INV_X1 U15839 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17922) );
  INV_X1 U15840 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18285) );
  XOR2_X1 U15841 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n9894), .Z(n17041) );
  OAI21_X1 U15842 ( .B1(n12590), .B2(n12589), .A(n12588), .ZN(n12595) );
  NOR2_X1 U15843 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19273), .ZN(n18051) );
  INV_X1 U15844 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17317) );
  NAND2_X1 U15845 ( .A1(n17317), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19214) );
  INV_X1 U15846 ( .A(n19214), .ZN(n19235) );
  NOR2_X1 U15847 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19266) );
  AOI21_X1 U15848 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19266), .ZN(n19119) );
  INV_X1 U15849 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n17001) );
  NOR3_X1 U15850 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n17001), .ZN(n18964) );
  OAI21_X2 U15851 ( .B1(n18285), .B2(n18008), .A(n18639), .ZN(n18127) );
  INV_X1 U15852 ( .A(n18127), .ZN(n18018) );
  OR2_X1 U15853 ( .A1(n12591), .A2(n18018), .ZN(n16857) );
  NOR2_X1 U15854 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18008), .ZN(
        n16870) );
  INV_X1 U15855 ( .A(n12592), .ZN(n16873) );
  NOR2_X1 U15856 ( .A1(n18285), .A2(n16873), .ZN(n17022) );
  INV_X1 U15857 ( .A(n18051), .ZN(n19123) );
  NAND2_X1 U15858 ( .A1(n18998), .A2(n12591), .ZN(n16874) );
  OAI211_X1 U15859 ( .C1(n17022), .C2(n19123), .A(n18289), .B(n16874), .ZN(
        n16868) );
  NOR2_X1 U15860 ( .A1(n16870), .A2(n16868), .ZN(n16855) );
  OAI221_X1 U15861 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16857), .C1(
        n10483), .C2(n16855), .A(n12593), .ZN(n12594) );
  NAND2_X1 U15862 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12599) );
  OAI211_X1 U15863 ( .C1(n12601), .C2(n19476), .A(n12600), .B(n12599), .ZN(
        n12602) );
  INV_X1 U15864 ( .A(n12602), .ZN(n12603) );
  NAND2_X1 U15865 ( .A1(n12607), .A2(n12606), .ZN(P2_U2984) );
  NOR4_X1 U15866 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12611) );
  NOR4_X1 U15867 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12610) );
  NOR4_X1 U15868 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12609) );
  NOR4_X1 U15869 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12608) );
  AND4_X1 U15870 ( .A1(n12611), .A2(n12610), .A3(n12609), .A4(n12608), .ZN(
        n12616) );
  NOR4_X1 U15871 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_23__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12614) );
  NOR4_X1 U15872 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12613) );
  NOR4_X1 U15873 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12612) );
  INV_X1 U15874 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21114) );
  AND4_X1 U15875 ( .A1(n12614), .A2(n12613), .A3(n12612), .A4(n21114), .ZN(
        n12615) );
  NAND2_X1 U15876 ( .A1(n12616), .A2(n12615), .ZN(n12617) );
  INV_X1 U15877 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21369) );
  NOR3_X1 U15878 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21369), .ZN(n12619) );
  NOR4_X1 U15879 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12618) );
  NAND4_X1 U15880 ( .A1(n20488), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n12619), .A4(
        n12618), .ZN(U214) );
  NOR2_X1 U15881 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12621) );
  NOR4_X1 U15882 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12620) );
  NAND4_X1 U15883 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12621), .A4(n12620), .ZN(n12622) );
  NOR2_X1 U15884 ( .A1(n19497), .A2(n12622), .ZN(n16913) );
  NAND2_X1 U15885 ( .A1(n16913), .A2(U214), .ZN(U212) );
  NOR2_X1 U15886 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12622), .ZN(n16989)
         );
  INV_X1 U15887 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17340) );
  NAND2_X1 U15888 ( .A1(n17349), .A2(n17340), .ZN(n17339) );
  NAND2_X1 U15889 ( .A1(n17323), .A2(n17315), .ZN(n17312) );
  INV_X1 U15890 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17631) );
  NAND2_X1 U15891 ( .A1(n17252), .A2(n17243), .ZN(n17242) );
  NAND2_X1 U15892 ( .A1(n17223), .A2(n17216), .ZN(n17215) );
  NAND2_X1 U15893 ( .A1(n17152), .A2(n17149), .ZN(n17148) );
  INV_X1 U15894 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17104) );
  NOR2_X1 U15895 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17103), .ZN(n17090) );
  INV_X1 U15896 ( .A(n12623), .ZN(n12624) );
  NOR2_X1 U15897 ( .A1(n16687), .A2(n12624), .ZN(n19053) );
  NAND2_X1 U15898 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19260), .ZN(n12625) );
  AOI211_X4 U15899 ( .C1(n17001), .C2(n19254), .A(n12641), .B(n12625), .ZN(
        n17376) );
  AOI211_X1 U15900 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17084), .A(n17074), .B(
        n17365), .ZN(n12646) );
  INV_X1 U15901 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19184) );
  OAI211_X1 U15902 ( .C1(n19259), .C2(n19260), .A(n19254), .B(n17001), .ZN(
        n12640) );
  INV_X1 U15903 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19182) );
  INV_X1 U15904 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19178) );
  INV_X1 U15905 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19175) );
  INV_X1 U15906 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19158) );
  INV_X1 U15907 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19152) );
  INV_X1 U15908 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19143) );
  NAND3_X1 U15909 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17316) );
  NOR2_X1 U15910 ( .A1(n19143), .A2(n17316), .ZN(n17307) );
  NAND2_X1 U15911 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17307), .ZN(n17273) );
  NAND2_X1 U15912 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n17275) );
  NOR3_X1 U15913 ( .A1(n19152), .A2(n17273), .A3(n17275), .ZN(n17235) );
  NAND4_X1 U15914 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17235), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n17230) );
  NOR2_X1 U15915 ( .A1(n19158), .A2(n17230), .ZN(n17214) );
  NAND3_X1 U15916 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17214), .ZN(n17203) );
  NAND2_X1 U15917 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17183) );
  NOR2_X1 U15918 ( .A1(n17203), .A2(n17183), .ZN(n17163) );
  NAND2_X1 U15919 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17163), .ZN(n17143) );
  NAND2_X1 U15920 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n17144) );
  NOR2_X1 U15921 ( .A1(n17143), .A2(n17144), .ZN(n17135) );
  NAND2_X1 U15922 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17135), .ZN(n17127) );
  NOR2_X1 U15923 ( .A1(n19175), .A2(n17127), .ZN(n17108) );
  NAND2_X1 U15924 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17108), .ZN(n17097) );
  NOR2_X1 U15925 ( .A1(n19178), .A2(n17097), .ZN(n17089) );
  NAND2_X1 U15926 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17089), .ZN(n17080) );
  NOR2_X1 U15927 ( .A1(n19182), .A2(n17080), .ZN(n12627) );
  NAND2_X1 U15928 ( .A1(n17353), .A2(n12627), .ZN(n17020) );
  INV_X1 U15929 ( .A(n19105), .ZN(n19115) );
  NAND2_X1 U15930 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19273), .ZN(n19113) );
  INV_X1 U15931 ( .A(n19113), .ZN(n18932) );
  NOR4_X4 U15932 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n19221), .ZN(n17338) );
  NOR2_X1 U15933 ( .A1(n9732), .A2(n17338), .ZN(n17264) );
  INV_X1 U15934 ( .A(n17264), .ZN(n12626) );
  OAI221_X1 U15935 ( .B1(n17366), .B2(P3_REIP_REG_26__SCAN_IN), .C1(n17366), 
        .C2(n12627), .A(n17372), .ZN(n17072) );
  INV_X1 U15936 ( .A(n17072), .ZN(n17057) );
  AOI21_X1 U15937 ( .B1(n19184), .B2(n17020), .A(n17057), .ZN(n12645) );
  NAND2_X1 U15938 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n12628), .ZN(
        n12632) );
  NAND3_X1 U15939 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n12633), .ZN(n17925) );
  INV_X1 U15940 ( .A(n12629), .ZN(n17923) );
  NOR2_X1 U15941 ( .A1(n18285), .A2(n17923), .ZN(n17024) );
  AOI21_X1 U15942 ( .B1(n17952), .B2(n17925), .A(n17024), .ZN(n17954) );
  INV_X1 U15943 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17965) );
  NAND2_X1 U15944 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12633), .ZN(
        n12631) );
  INV_X1 U15945 ( .A(n17925), .ZN(n12630) );
  AOI21_X1 U15946 ( .B1(n17965), .B2(n12631), .A(n12630), .ZN(n17968) );
  INV_X1 U15947 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17978) );
  AOI22_X1 U15948 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12633), .B1(
        n12632), .B2(n17978), .ZN(n17981) );
  NOR2_X1 U15949 ( .A1(n18285), .A2(n18017), .ZN(n12637) );
  NAND3_X1 U15950 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(n12637), .ZN(n17999) );
  AOI21_X1 U15951 ( .B1(n17993), .B2(n17999), .A(n12633), .ZN(n17997) );
  INV_X1 U15952 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17117) );
  NAND2_X1 U15953 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12637), .ZN(
        n12634) );
  INV_X1 U15954 ( .A(n17999), .ZN(n17963) );
  AOI21_X1 U15955 ( .B1(n17117), .B2(n12634), .A(n17963), .ZN(n18009) );
  NOR2_X1 U15956 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18285), .ZN(
        n17199) );
  AND2_X1 U15957 ( .A1(n12635), .A2(n17199), .ZN(n12636) );
  NOR2_X1 U15958 ( .A1(n12639), .A2(n12636), .ZN(n17130) );
  INV_X1 U15959 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17138) );
  NAND2_X1 U15960 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n12635), .ZN(
        n18007) );
  AOI21_X1 U15961 ( .B1(n17138), .B2(n18007), .A(n12637), .ZN(n18035) );
  NOR2_X1 U15962 ( .A1(n17130), .A2(n18035), .ZN(n17129) );
  NOR2_X1 U15963 ( .A1(n17129), .A2(n12639), .ZN(n17120) );
  INV_X1 U15964 ( .A(n12637), .ZN(n12638) );
  XNOR2_X1 U15965 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12638), .ZN(
        n18022) );
  NOR2_X1 U15966 ( .A1(n17120), .A2(n18022), .ZN(n17119) );
  NOR2_X1 U15967 ( .A1(n17981), .A2(n17092), .ZN(n17091) );
  INV_X1 U15968 ( .A(n17338), .ZN(n19118) );
  AOI211_X1 U15969 ( .C1(n17954), .C2(n9879), .A(n17026), .B(n19118), .ZN(
        n12644) );
  INV_X1 U15970 ( .A(n12640), .ZN(n19103) );
  AOI211_X4 U15971 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19260), .A(n19103), .B(
        n12641), .ZN(n17377) );
  INV_X1 U15972 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n12642) );
  OAI22_X1 U15973 ( .A1(n17952), .A2(n17363), .B1(n17334), .B2(n12642), .ZN(
        n12643) );
  OR4_X1 U15974 ( .A1(n12646), .A2(n12645), .A3(n12644), .A4(n12643), .ZN(
        P3_U2645) );
  NAND2_X1 U15975 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19410) );
  INV_X1 U15976 ( .A(n19410), .ZN(n16768) );
  AND2_X1 U15977 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16768), .ZN(n13772) );
  INV_X1 U15978 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20207) );
  NAND2_X1 U15979 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20207), .ZN(n13726) );
  NOR2_X1 U15980 ( .A1(n20238), .A2(n13726), .ZN(n13771) );
  NOR3_X1 U15981 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n12647) );
  NOR4_X1 U15982 ( .A1(n16769), .A2(n13772), .A3(n13771), .A4(n12647), .ZN(
        P2_U3178) );
  NOR2_X1 U15983 ( .A1(n11220), .A2(n13775), .ZN(n19406) );
  NAND2_X1 U15984 ( .A1(n19406), .A2(n13680), .ZN(n15810) );
  INV_X1 U15985 ( .A(n15810), .ZN(n12649) );
  INV_X1 U15986 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20243) );
  INV_X1 U15987 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16648) );
  AND2_X1 U15988 ( .A1(n20180), .A2(n16648), .ZN(n14547) );
  INV_X1 U15989 ( .A(n14547), .ZN(n12648) );
  OAI211_X1 U15990 ( .C1(n12649), .C2(n20243), .A(n13114), .B(n12648), .ZN(
        P2_U2814) );
  INV_X1 U15991 ( .A(n14549), .ZN(n20235) );
  INV_X1 U15992 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n12650) );
  INV_X1 U15993 ( .A(n20179), .ZN(n16664) );
  OAI22_X1 U15994 ( .A1(n20235), .A2(n12650), .B1(n13726), .B2(n16664), .ZN(
        P2_U2816) );
  NOR3_X1 U15995 ( .A1(n12652), .A2(n12651), .A3(n12841), .ZN(n13688) );
  NOR2_X1 U15996 ( .A1(n13688), .A2(n13775), .ZN(n20224) );
  OAI21_X1 U15997 ( .B1(n20224), .B2(n12654), .A(n12653), .ZN(P2_U2819) );
  AND2_X2 U15998 ( .A1(n13438), .A2(n12958), .ZN(n12780) );
  AOI22_X1 U15999 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U16000 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U16001 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12658) );
  AND2_X2 U16002 ( .A1(n12662), .A2(n12958), .ZN(n14486) );
  AND2_X2 U16003 ( .A1(n12656), .A2(n12962), .ZN(n14482) );
  AOI22_X1 U16004 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12657) );
  AND2_X2 U16005 ( .A1(n12963), .A2(n12661), .ZN(n12768) );
  AOI22_X1 U16006 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12994), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12666) );
  AND2_X2 U16007 ( .A1(n12664), .A2(n13438), .ZN(n14488) );
  AND2_X2 U16008 ( .A1(n13438), .A2(n13451), .ZN(n14449) );
  AOI22_X1 U16009 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U16010 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U16011 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U16012 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U16013 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U16014 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U16015 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12677) );
  AOI22_X1 U16016 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U16017 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12994), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12675) );
  INV_X2 U16018 ( .A(n12888), .ZN(n12797) );
  XNOR2_X1 U16019 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12716) );
  NAND2_X1 U16020 ( .A1(n12708), .A2(n12716), .ZN(n12680) );
  NAND2_X1 U16021 ( .A1(n20905), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12679) );
  NAND2_X1 U16022 ( .A1(n12680), .A2(n12679), .ZN(n12704) );
  XNOR2_X1 U16023 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12703) );
  XNOR2_X1 U16024 ( .A(n12704), .B(n12703), .ZN(n12801) );
  INV_X1 U16025 ( .A(n12801), .ZN(n12734) );
  NAND2_X1 U16026 ( .A1(n13833), .A2(n12734), .ZN(n12707) );
  AOI22_X1 U16027 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U16028 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U16029 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12682) );
  NAND4_X1 U16030 ( .A1(n12684), .A2(n12683), .A3(n12682), .A4(n12681), .ZN(
        n12690) );
  AOI22_X1 U16031 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12780), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U16032 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14488), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U16033 ( .A1(n14449), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12994), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U16034 ( .A1(n14474), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12685) );
  NAND4_X1 U16035 ( .A1(n12688), .A2(n12687), .A3(n12686), .A4(n12685), .ZN(
        n12689) );
  AND2_X2 U16036 ( .A1(n12691), .A2(n12797), .ZN(n12900) );
  INV_X2 U16037 ( .A(n12900), .ZN(n14853) );
  AOI22_X1 U16038 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U16039 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14235), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U16040 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U16041 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12692) );
  NAND4_X1 U16042 ( .A1(n12695), .A2(n12694), .A3(n12693), .A4(n12692), .ZN(
        n12701) );
  AOI22_X1 U16043 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U16044 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12696) );
  NAND4_X1 U16045 ( .A1(n12699), .A2(n12698), .A3(n12697), .A4(n12696), .ZN(
        n12700) );
  NAND2_X1 U16046 ( .A1(n12691), .A2(n12813), .ZN(n12702) );
  NAND2_X1 U16047 ( .A1(n12704), .A2(n12703), .ZN(n12706) );
  NAND2_X1 U16048 ( .A1(n20830), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12705) );
  NAND2_X1 U16049 ( .A1(n12706), .A2(n12705), .ZN(n12729) );
  XNOR2_X1 U16050 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12728) );
  XNOR2_X1 U16051 ( .A(n12729), .B(n12728), .ZN(n12800) );
  NOR2_X1 U16052 ( .A1(n13835), .A2(n12734), .ZN(n12725) );
  AND2_X2 U16053 ( .A1(n12813), .A2(n12814), .ZN(n14376) );
  INV_X1 U16054 ( .A(n12708), .ZN(n12715) );
  NAND2_X1 U16055 ( .A1(n16728), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12709) );
  AND2_X1 U16056 ( .A1(n12715), .A2(n12709), .ZN(n12712) );
  NAND2_X1 U16057 ( .A1(n13833), .A2(n12712), .ZN(n12710) );
  NAND2_X1 U16058 ( .A1(n12730), .A2(n12710), .ZN(n12714) );
  INV_X1 U16059 ( .A(n12711), .ZN(n13013) );
  OAI211_X1 U16060 ( .C1(n13013), .C2(n12823), .A(n12732), .B(n12712), .ZN(
        n12713) );
  XNOR2_X1 U16061 ( .A(n12716), .B(n12715), .ZN(n12804) );
  NAND2_X1 U16062 ( .A1(n13833), .A2(n20506), .ZN(n12717) );
  NAND2_X1 U16063 ( .A1(n12898), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12718) );
  OAI211_X1 U16064 ( .C1(n13835), .C2(n12804), .A(n12717), .B(n12718), .ZN(
        n12720) );
  NAND2_X1 U16065 ( .A1(n12718), .A2(n20506), .ZN(n12719) );
  OAI22_X1 U16066 ( .A1(n12721), .A2(n12720), .B1(n12731), .B2(n12804), .ZN(
        n12723) );
  NAND2_X1 U16067 ( .A1(n12721), .A2(n12720), .ZN(n12722) );
  NAND2_X1 U16068 ( .A1(n12723), .A2(n12722), .ZN(n12724) );
  OAI21_X1 U16069 ( .B1(n12735), .B2(n12725), .A(n12724), .ZN(n12738) );
  NOR2_X1 U16070 ( .A1(n12726), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12727) );
  AOI21_X1 U16071 ( .B1(n12729), .B2(n12728), .A(n12727), .ZN(n12743) );
  INV_X1 U16072 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20484) );
  NOR2_X1 U16073 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20484), .ZN(
        n12746) );
  AND2_X1 U16074 ( .A1(n12743), .A2(n12746), .ZN(n12802) );
  AOI22_X1 U16075 ( .A1(n12731), .A2(n12802), .B1(n12749), .B2(n12800), .ZN(
        n12737) );
  INV_X1 U16076 ( .A(n12732), .ZN(n12733) );
  NAND4_X1 U16077 ( .A1(n12735), .A2(n12734), .A3(n13833), .A4(n12733), .ZN(
        n12736) );
  NAND3_X1 U16078 ( .A1(n12738), .A2(n12737), .A3(n12736), .ZN(n12740) );
  NAND2_X1 U16079 ( .A1(n13835), .A2(n12802), .ZN(n12739) );
  NAND2_X1 U16080 ( .A1(n12740), .A2(n12739), .ZN(n12742) );
  NAND2_X1 U16081 ( .A1(n21091), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12741) );
  NAND2_X1 U16082 ( .A1(n12742), .A2(n12741), .ZN(n12751) );
  INV_X1 U16083 ( .A(n12743), .ZN(n12745) );
  INV_X1 U16084 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13580) );
  NOR2_X1 U16085 ( .A1(n13580), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12744) );
  INV_X1 U16086 ( .A(n12746), .ZN(n12747) );
  NAND2_X1 U16087 ( .A1(n12749), .A2(n12806), .ZN(n12750) );
  AOI22_X1 U16088 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U16089 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U16090 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12761) );
  AOI22_X1 U16091 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U16092 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U16093 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U16094 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U16095 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U16096 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14484), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U16097 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U16098 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12994), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12766) );
  NAND2_X1 U16099 ( .A1(n12767), .A2(n12766), .ZN(n12772) );
  AOI22_X1 U16100 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U16101 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12769) );
  NAND2_X1 U16102 ( .A1(n12770), .A2(n12769), .ZN(n12771) );
  NAND2_X2 U16103 ( .A1(n12774), .A2(n12773), .ZN(n12892) );
  AOI22_X1 U16104 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12779) );
  AOI22_X1 U16105 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U16106 ( .A1(n14449), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12994), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U16107 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U16108 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U16109 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14488), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12782) );
  AOI22_X1 U16110 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12781) );
  NAND2_X2 U16111 ( .A1(n12785), .A2(n9786), .ZN(n12819) );
  AOI22_X1 U16112 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U16113 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U16114 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U16115 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12786) );
  NAND4_X1 U16116 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12795) );
  AOI22_X1 U16117 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U16118 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U16119 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12994), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12790) );
  NAND4_X1 U16120 ( .A1(n12793), .A2(n12792), .A3(n12791), .A4(n12790), .ZN(
        n12794) );
  NAND2_X1 U16121 ( .A1(n21090), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16750) );
  OR2_X1 U16122 ( .A1(n16750), .A2(n21091), .ZN(n20246) );
  INV_X1 U16123 ( .A(n12892), .ZN(n12815) );
  NAND2_X1 U16124 ( .A1(n12815), .A2(n12813), .ZN(n12796) );
  NOR2_X1 U16125 ( .A1(n12796), .A2(n13208), .ZN(n12799) );
  NOR3_X1 U16126 ( .A1(n12802), .A2(n12801), .A3(n12800), .ZN(n12803) );
  AND2_X1 U16127 ( .A1(n12804), .A2(n12803), .ZN(n12805) );
  NOR2_X1 U16128 ( .A1(n12806), .A2(n12805), .ZN(n13319) );
  NAND2_X1 U16129 ( .A1(n12902), .A2(n13319), .ZN(n12868) );
  NOR2_X2 U16130 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20908) );
  NAND2_X1 U16131 ( .A1(n20908), .A2(n21090), .ZN(n20249) );
  INV_X1 U16132 ( .A(n20249), .ZN(n14717) );
  AOI21_X1 U16133 ( .B1(n12832), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14717), 
        .ZN(n12807) );
  NAND2_X1 U16134 ( .A1(n13073), .A2(n12807), .ZN(P1_U2801) );
  NAND2_X1 U16135 ( .A1(n13328), .A2(n14853), .ZN(n12809) );
  NAND2_X1 U16136 ( .A1(n12897), .A2(n12868), .ZN(n12808) );
  NAND2_X1 U16137 ( .A1(n12809), .A2(n12808), .ZN(n20247) );
  NAND2_X1 U16138 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21102) );
  INV_X1 U16139 ( .A(n21102), .ZN(n21094) );
  NAND2_X1 U16140 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21108) );
  OAI21_X1 U16141 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n21108), .ZN(n12896) );
  OR2_X1 U16142 ( .A1(n12896), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n16765) );
  NAND2_X1 U16143 ( .A1(n14416), .A2(n16765), .ZN(n12810) );
  NAND2_X1 U16144 ( .A1(n12810), .A2(n21102), .ZN(n12865) );
  OAI21_X1 U16145 ( .B1(n14853), .B2(n21094), .A(n12865), .ZN(n12811) );
  NOR2_X1 U16146 ( .A1(n20247), .A2(n12811), .ZN(n16741) );
  OR2_X1 U16147 ( .A1(n16741), .A2(n20246), .ZN(n12829) );
  INV_X1 U16148 ( .A(n12829), .ZN(n20255) );
  INV_X1 U16149 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12831) );
  NAND2_X1 U16150 ( .A1(n12880), .A2(n12871), .ZN(n12882) );
  NOR2_X1 U16151 ( .A1(n15472), .A2(n12691), .ZN(n13327) );
  INV_X1 U16152 ( .A(n14866), .ZN(n12817) );
  NAND2_X1 U16153 ( .A1(n12817), .A2(n12823), .ZN(n12954) );
  AND2_X1 U16154 ( .A1(n12889), .A2(n12954), .ZN(n13340) );
  INV_X1 U16155 ( .A(n13339), .ZN(n12961) );
  AOI21_X1 U16156 ( .B1(n15472), .B2(n12797), .A(n12862), .ZN(n12824) );
  NAND2_X1 U16157 ( .A1(n12871), .A2(n13333), .ZN(n12822) );
  NAND2_X1 U16158 ( .A1(n12898), .A2(n12819), .ZN(n12820) );
  NAND2_X1 U16159 ( .A1(n12820), .A2(n20532), .ZN(n12870) );
  INV_X1 U16160 ( .A(n12870), .ZN(n12821) );
  AND2_X1 U16161 ( .A1(n12822), .A2(n12821), .ZN(n12950) );
  AND2_X1 U16162 ( .A1(n12824), .A2(n12950), .ZN(n12869) );
  NAND2_X1 U16163 ( .A1(n12824), .A2(n12900), .ZN(n12960) );
  NAND2_X1 U16164 ( .A1(n16744), .A2(n12960), .ZN(n13334) );
  NOR2_X1 U16165 ( .A1(n13334), .A2(n12825), .ZN(n12826) );
  MUX2_X1 U16166 ( .A(n12961), .B(n12826), .S(n13328), .Z(n12827) );
  OAI21_X1 U16167 ( .B1(n13319), .B2(n10413), .A(n12827), .ZN(n12828) );
  NAND2_X1 U16168 ( .A1(n12828), .A2(n20532), .ZN(n16743) );
  OR2_X1 U16169 ( .A1(n12829), .A2(n16743), .ZN(n12830) );
  OAI21_X1 U16170 ( .B1(n20255), .B2(n12831), .A(n12830), .ZN(P1_U3484) );
  INV_X1 U16171 ( .A(n20908), .ZN(n21030) );
  NAND2_X1 U16172 ( .A1(n14540), .A2(n21091), .ZN(n13243) );
  NOR2_X1 U16173 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21090), .ZN(n14327) );
  NAND3_X1 U16174 ( .A1(n21102), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n14327), 
        .ZN(n12833) );
  NAND3_X1 U16175 ( .A1(n21030), .A2(n13243), .A3(n12833), .ZN(n12834) );
  NOR2_X1 U16176 ( .A1(n14557), .A2(n12834), .ZN(n12838) );
  NOR2_X1 U16177 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16753) );
  NOR2_X1 U16178 ( .A1(n12838), .A2(n16753), .ZN(n12840) );
  INV_X1 U16179 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20832) );
  OAI21_X1 U16180 ( .B1(n16765), .B2(n20832), .A(n14381), .ZN(n12835) );
  NAND3_X1 U16181 ( .A1(n12835), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n21102), 
        .ZN(n12837) );
  INV_X1 U16182 ( .A(n13382), .ZN(n13090) );
  NAND2_X1 U16183 ( .A1(n20506), .A2(n16765), .ZN(n13318) );
  INV_X1 U16184 ( .A(n13318), .ZN(n12836) );
  AOI22_X1 U16185 ( .A1(n12837), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13090), 
        .B2(n12836), .ZN(n12839) );
  INV_X1 U16186 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21105) );
  AOI22_X1 U16187 ( .A1(n12840), .A2(n12839), .B1(n12838), .B2(n21105), .ZN(
        P1_U3485) );
  INV_X1 U16188 ( .A(n12841), .ZN(n12842) );
  OR2_X1 U16189 ( .A1(n11220), .A2(n12842), .ZN(n12847) );
  NOR2_X1 U16190 ( .A1(n13765), .A2(n13630), .ZN(n13068) );
  INV_X1 U16191 ( .A(n12843), .ZN(n12844) );
  NOR2_X1 U16192 ( .A1(n13068), .A2(n12844), .ZN(n12845) );
  OAI211_X1 U16193 ( .C1(n12847), .C2(n19405), .A(n12846), .B(n12845), .ZN(
        n13691) );
  NAND2_X1 U16194 ( .A1(n13691), .A2(n13724), .ZN(n12849) );
  NAND2_X1 U16195 ( .A1(n13772), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n16772) );
  NAND2_X1 U16196 ( .A1(n11619), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13701) );
  AND2_X1 U16197 ( .A1(n16772), .A2(n13701), .ZN(n12848) );
  NAND2_X1 U16198 ( .A1(n12849), .A2(n12848), .ZN(n16666) );
  NOR2_X1 U16199 ( .A1(n11220), .A2(n12850), .ZN(n13687) );
  NAND4_X1 U16200 ( .A1(n16666), .A2(n20179), .A3(n19513), .A4(n13687), .ZN(
        n12851) );
  OAI21_X1 U16201 ( .B1(n11199), .B2(n16666), .A(n12851), .ZN(P2_U3595) );
  AOI21_X1 U16202 ( .B1(n13181), .B2(n15809), .A(n12852), .ZN(n16831) );
  INV_X1 U16203 ( .A(n12853), .ZN(n12855) );
  INV_X1 U16204 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12854) );
  AOI21_X1 U16205 ( .B1(n16283), .B2(n12855), .A(n12854), .ZN(n12860) );
  NAND2_X1 U16206 ( .A1(n12856), .A2(n13181), .ZN(n12857) );
  NAND2_X1 U16207 ( .A1(n12858), .A2(n12857), .ZN(n16841) );
  NAND2_X1 U16208 ( .A1(n19359), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16834) );
  OAI21_X1 U16209 ( .B1(n19490), .B2(n16841), .A(n16834), .ZN(n12859) );
  AOI211_X1 U16210 ( .C1(n16831), .C2(n19484), .A(n12860), .B(n12859), .ZN(
        n12861) );
  OAI21_X1 U16211 ( .B1(n16835), .B2(n16287), .A(n12861), .ZN(P2_U3014) );
  AND2_X1 U16212 ( .A1(n12902), .A2(n20506), .ZN(n14537) );
  INV_X1 U16213 ( .A(n16765), .ZN(n13320) );
  NAND2_X1 U16214 ( .A1(n14537), .A2(n13320), .ZN(n13029) );
  NAND3_X1 U16215 ( .A1(n12864), .A2(n12863), .A3(n20532), .ZN(n12901) );
  AOI21_X1 U16216 ( .B1(n13029), .B2(n12901), .A(n12865), .ZN(n12866) );
  MUX2_X1 U16217 ( .A(n12866), .B(n13339), .S(n13328), .Z(n12876) );
  NAND2_X1 U16218 ( .A1(n12691), .A2(n21102), .ZN(n12867) );
  OAI22_X1 U16219 ( .A1(n13328), .A2(n12960), .B1(n12868), .B2(n12867), .ZN(
        n13202) );
  OR2_X1 U16220 ( .A1(n12869), .A2(n12902), .ZN(n12873) );
  NOR2_X2 U16221 ( .A1(n12870), .A2(n12812), .ZN(n12911) );
  NAND2_X1 U16222 ( .A1(n12911), .A2(n13205), .ZN(n12893) );
  AOI21_X1 U16223 ( .B1(n14376), .B2(n13018), .A(n12797), .ZN(n12872) );
  NAND2_X1 U16224 ( .A1(n12893), .A2(n12872), .ZN(n12886) );
  NAND2_X1 U16225 ( .A1(n12873), .A2(n12886), .ZN(n13326) );
  INV_X1 U16226 ( .A(n13326), .ZN(n12874) );
  INV_X1 U16227 ( .A(n20246), .ZN(n13203) );
  NAND2_X1 U16228 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16824) );
  INV_X1 U16229 ( .A(n16824), .ZN(n13457) );
  NAND2_X1 U16230 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13457), .ZN(n16829) );
  INV_X1 U16231 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20254) );
  NOR2_X1 U16232 ( .A1(n16829), .A2(n20254), .ZN(n12877) );
  AOI21_X1 U16233 ( .B1(n16730), .B2(n13203), .A(n12877), .ZN(n12936) );
  NAND2_X1 U16234 ( .A1(n21091), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n12878) );
  NAND2_X1 U16235 ( .A1(n12936), .A2(n12878), .ZN(n15487) );
  NAND2_X1 U16236 ( .A1(n12813), .A2(n12819), .ZN(n12879) );
  INV_X1 U16237 ( .A(n12880), .ZN(n12881) );
  NAND2_X1 U16238 ( .A1(n12884), .A2(n12883), .ZN(n12885) );
  NAND2_X1 U16239 ( .A1(n12885), .A2(n12797), .ZN(n12918) );
  NAND2_X1 U16240 ( .A1(n12918), .A2(n12886), .ZN(n12952) );
  INV_X4 U16241 ( .A(n12887), .ZN(n14318) );
  NOR2_X1 U16242 ( .A1(n12892), .A2(n12891), .ZN(n12899) );
  NAND2_X1 U16243 ( .A1(n12893), .A2(n15472), .ZN(n12910) );
  NAND3_X1 U16244 ( .A1(n12956), .A2(n12894), .A3(n12910), .ZN(n12895) );
  OAI21_X1 U16245 ( .B1(n12952), .B2(n12895), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12904) );
  NAND2_X1 U16246 ( .A1(n12904), .A2(n10402), .ZN(n12924) );
  NAND2_X1 U16247 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12927) );
  OAI21_X1 U16248 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n12927), .ZN(n20835) );
  NAND2_X1 U16249 ( .A1(n16750), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12921) );
  OAI21_X1 U16250 ( .B1(n13243), .B2(n20835), .A(n12921), .ZN(n12905) );
  INV_X1 U16251 ( .A(n12905), .ZN(n12906) );
  NAND2_X1 U16252 ( .A1(n12924), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12909) );
  INV_X1 U16253 ( .A(n16750), .ZN(n12907) );
  MUX2_X1 U16254 ( .A(n12907), .B(n13243), .S(n20953), .Z(n12908) );
  NAND2_X1 U16255 ( .A1(n12909), .A2(n12908), .ZN(n12988) );
  OR2_X1 U16256 ( .A1(n12910), .A2(n12691), .ZN(n12919) );
  INV_X1 U16257 ( .A(n12911), .ZN(n12912) );
  NAND2_X1 U16258 ( .A1(n12912), .A2(n14381), .ZN(n12917) );
  NAND3_X1 U16259 ( .A1(n14866), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14540), 
        .ZN(n12915) );
  NAND2_X1 U16260 ( .A1(n13205), .A2(n12892), .ZN(n12916) );
  INV_X1 U16261 ( .A(n12987), .ZN(n12920) );
  INV_X1 U16262 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15469) );
  NAND2_X1 U16263 ( .A1(n12921), .A2(n15469), .ZN(n12922) );
  NAND2_X1 U16264 ( .A1(n12923), .A2(n12922), .ZN(n12946) );
  NAND2_X1 U16265 ( .A1(n16750), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12925) );
  INV_X1 U16266 ( .A(n13243), .ZN(n12931) );
  INV_X1 U16267 ( .A(n12927), .ZN(n12926) );
  NAND2_X1 U16268 ( .A1(n12926), .A2(n20830), .ZN(n20606) );
  NAND2_X1 U16269 ( .A1(n12927), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U16270 ( .A1(n20606), .A2(n12928), .ZN(n20501) );
  NAND2_X1 U16271 ( .A1(n12929), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12933) );
  INV_X1 U16272 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20834) );
  NOR3_X1 U16273 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20830), .A3(
        n20905), .ZN(n20751) );
  NAND2_X1 U16274 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20751), .ZN(
        n20745) );
  NAND2_X1 U16275 ( .A1(n20834), .A2(n20745), .ZN(n12930) );
  NAND3_X1 U16276 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21028) );
  INV_X1 U16277 ( .A(n21028), .ZN(n21036) );
  NAND2_X1 U16278 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21036), .ZN(
        n21029) );
  AOI22_X1 U16279 ( .A1(n12931), .A2(n20776), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16750), .ZN(n12932) );
  INV_X1 U16280 ( .A(n20648), .ZN(n20911) );
  XNOR2_X1 U16281 ( .A(n12934), .B(n13580), .ZN(n20319) );
  INV_X1 U16282 ( .A(n14540), .ZN(n15485) );
  OR4_X1 U16283 ( .A1(n20319), .A2(n12936), .A3(n15485), .A4(n12935), .ZN(
        n12937) );
  OAI21_X1 U16284 ( .B1(n15487), .B2(n13580), .A(n12937), .ZN(P1_U3468) );
  INV_X1 U16285 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n21457) );
  INV_X1 U16286 ( .A(n12939), .ZN(n12940) );
  XNOR2_X1 U16287 ( .A(n12938), .B(n12940), .ZN(n16580) );
  INV_X1 U16288 ( .A(n16580), .ZN(n19367) );
  INV_X1 U16289 ( .A(n12941), .ZN(n12942) );
  INV_X1 U16290 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U16291 ( .A1(n19499), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12943) );
  OAI21_X1 U16292 ( .B1(n19499), .B2(n12944), .A(n12943), .ZN(n19543) );
  INV_X1 U16293 ( .A(n19543), .ZN(n12945) );
  OAI222_X1 U16294 ( .A1(n21457), .A2(n16017), .B1(n19367), .B2(n16015), .C1(
        n19403), .C2(n12945), .ZN(P2_U2913) );
  NOR2_X1 U16295 ( .A1(n12950), .A2(n14414), .ZN(n12951) );
  NOR2_X1 U16296 ( .A1(n12952), .A2(n12951), .ZN(n13342) );
  INV_X1 U16297 ( .A(n12953), .ZN(n13199) );
  AND2_X1 U16298 ( .A1(n12901), .A2(n12954), .ZN(n12955) );
  AND4_X1 U16299 ( .A1(n13199), .A2(n12956), .A3(n12955), .A4(n12935), .ZN(
        n12957) );
  NAND2_X1 U16300 ( .A1(n13342), .A2(n12957), .ZN(n15474) );
  INV_X1 U16301 ( .A(n15474), .ZN(n14538) );
  OR2_X1 U16302 ( .A1(n12949), .A2(n14538), .ZN(n12970) );
  XNOR2_X1 U16303 ( .A(n12958), .B(n10007), .ZN(n12973) );
  INV_X1 U16304 ( .A(n12973), .ZN(n12959) );
  NOR2_X1 U16305 ( .A1(n13442), .A2(n12959), .ZN(n12968) );
  AND2_X1 U16306 ( .A1(n12961), .A2(n12960), .ZN(n13440) );
  INV_X1 U16307 ( .A(n14537), .ZN(n16727) );
  INV_X1 U16308 ( .A(n12962), .ZN(n12965) );
  INV_X1 U16309 ( .A(n12963), .ZN(n12964) );
  NAND2_X1 U16310 ( .A1(n12965), .A2(n12964), .ZN(n12966) );
  OAI22_X1 U16311 ( .A1(n13440), .A2(n12973), .B1(n16727), .B2(n12966), .ZN(
        n12967) );
  AOI21_X1 U16312 ( .B1(n14538), .B2(n12968), .A(n12967), .ZN(n12969) );
  NAND2_X1 U16313 ( .A1(n12970), .A2(n12969), .ZN(n13448) );
  NOR2_X1 U16314 ( .A1(n21090), .A2(n13344), .ZN(n15478) );
  INV_X1 U16315 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20481) );
  INV_X1 U16316 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16317 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20481), .B2(n12971), .ZN(
        n15476) );
  INV_X1 U16318 ( .A(n16754), .ZN(n15480) );
  AOI222_X1 U16319 ( .A1(n13448), .A2(n14540), .B1(n15478), .B2(n15476), .C1(
        n12973), .C2(n15480), .ZN(n12975) );
  INV_X1 U16320 ( .A(n15487), .ZN(n14542) );
  NAND2_X1 U16321 ( .A1(n14542), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12974) );
  OAI21_X1 U16322 ( .B1(n12975), .B2(n14542), .A(n12974), .ZN(P1_U3472) );
  INV_X1 U16323 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14882) );
  OR2_X1 U16324 ( .A1(n14314), .A2(n14882), .ZN(n12978) );
  NAND2_X1 U16325 ( .A1(n14318), .A2(n14882), .ZN(n12977) );
  NAND2_X1 U16326 ( .A1(n12978), .A2(n12977), .ZN(n13079) );
  INV_X1 U16327 ( .A(n13079), .ZN(n12981) );
  OR2_X1 U16328 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12980) );
  AND2_X1 U16329 ( .A1(n12981), .A2(n12980), .ZN(n14885) );
  INV_X1 U16330 ( .A(n14885), .ZN(n13028) );
  NAND2_X1 U16331 ( .A1(n13328), .A2(n13339), .ZN(n12985) );
  NAND3_X1 U16332 ( .A1(n13333), .A2(n14551), .A3(n12819), .ZN(n13198) );
  INV_X1 U16333 ( .A(n13198), .ZN(n12983) );
  NAND3_X1 U16334 ( .A1(n12982), .A2(n14409), .A3(n12983), .ZN(n12984) );
  NAND2_X1 U16335 ( .A1(n12985), .A2(n12984), .ZN(n12986) );
  AOI22_X1 U16336 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16337 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16338 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16339 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12989) );
  NAND4_X1 U16340 ( .A1(n12992), .A2(n12991), .A3(n12990), .A4(n12989), .ZN(
        n13000) );
  AOI22_X1 U16341 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14476), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16342 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16343 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U16344 ( .A1(n14487), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12995) );
  NAND4_X1 U16345 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n12999) );
  INV_X1 U16346 ( .A(n13381), .ZN(n13098) );
  INV_X1 U16347 ( .A(n14380), .ZN(n14388) );
  NAND2_X1 U16348 ( .A1(n13098), .A2(n14388), .ZN(n13092) );
  AOI22_X1 U16349 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16350 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U16351 ( .A1(n14450), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U16352 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13001) );
  NAND4_X1 U16353 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13010) );
  AOI22_X1 U16354 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U16355 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U16356 ( .A1(n12775), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16357 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13005) );
  NAND4_X1 U16358 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  MUX2_X1 U16359 ( .A(n14357), .B(n13092), .S(n13402), .Z(n13011) );
  NAND2_X1 U16360 ( .A1(n13830), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13017) );
  INV_X1 U16361 ( .A(n13012), .ZN(n13015) );
  OAI21_X1 U16362 ( .B1(n13402), .B2(n21091), .A(n13013), .ZN(n13014) );
  NAND2_X1 U16363 ( .A1(n20567), .A2(n13018), .ZN(n13019) );
  NAND2_X1 U16364 ( .A1(n13019), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13026) );
  AND2_X1 U16365 ( .A1(n13021), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13389) );
  INV_X1 U16366 ( .A(n13389), .ZN(n13581) );
  NAND2_X1 U16367 ( .A1(n13022), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13024) );
  INV_X2 U16368 ( .A(n9862), .ZN(n14504) );
  NAND2_X1 U16369 ( .A1(n14504), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13023) );
  OAI211_X1 U16370 ( .C1(n13581), .C2(n16728), .A(n13024), .B(n13023), .ZN(
        n13025) );
  AOI21_X1 U16371 ( .B1(n13020), .B2(n13984), .A(n13025), .ZN(n13107) );
  OR2_X1 U16372 ( .A1(n13026), .A2(n13107), .ZN(n13110) );
  NAND2_X1 U16373 ( .A1(n13026), .A2(n13107), .ZN(n13027) );
  NAND2_X1 U16374 ( .A1(n13110), .A2(n13027), .ZN(n14888) );
  NAND2_X2 U16375 ( .A1(n20355), .A2(n20532), .ZN(n14932) );
  OAI222_X1 U16376 ( .A1(n13028), .A2(n14930), .B1(n14882), .B2(n20355), .C1(
        n14888), .C2(n14932), .ZN(P1_U2872) );
  INV_X1 U16377 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13035) );
  INV_X1 U16378 ( .A(n13029), .ZN(n13031) );
  NAND2_X1 U16379 ( .A1(n12691), .A2(n13320), .ZN(n13030) );
  NOR2_X1 U16380 ( .A1(n12897), .A2(n13030), .ZN(n16752) );
  NOR2_X1 U16381 ( .A1(n13031), .A2(n16752), .ZN(n13032) );
  NAND2_X1 U16382 ( .A1(n13033), .A2(n12816), .ZN(n13368) );
  NOR2_X1 U16383 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16824), .ZN(n20372) );
  AOI22_X1 U16384 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20372), .B1(n16767), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13034) );
  OAI21_X1 U16385 ( .B1(n13035), .B2(n13368), .A(n13034), .ZN(P1_U2920) );
  INV_X1 U16386 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U16387 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20372), .B1(n16767), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13036) );
  OAI21_X1 U16388 ( .B1(n13037), .B2(n13368), .A(n13036), .ZN(P1_U2919) );
  INV_X1 U16389 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U16390 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20382), .B1(n16767), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13038) );
  OAI21_X1 U16391 ( .B1(n13039), .B2(n13368), .A(n13038), .ZN(P1_U2911) );
  INV_X1 U16392 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U16393 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20382), .B1(n16767), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13040) );
  OAI21_X1 U16394 ( .B1(n13041), .B2(n13368), .A(n13040), .ZN(P1_U2912) );
  INV_X1 U16395 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16396 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20382), .B1(n16767), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13042) );
  OAI21_X1 U16397 ( .B1(n13043), .B2(n13368), .A(n13042), .ZN(P1_U2907) );
  INV_X1 U16398 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16399 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20382), .B1(n16767), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13044) );
  OAI21_X1 U16400 ( .B1(n13045), .B2(n13368), .A(n13044), .ZN(P1_U2908) );
  INV_X1 U16401 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U16402 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20382), .B1(n16767), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13046) );
  OAI21_X1 U16403 ( .B1(n13047), .B2(n13368), .A(n13046), .ZN(P1_U2909) );
  INV_X1 U16404 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U16405 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20382), .B1(n16767), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13048) );
  OAI21_X1 U16406 ( .B1(n14963), .B2(n13368), .A(n13048), .ZN(P1_U2913) );
  INV_X1 U16407 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16408 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20372), .B1(n16767), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13049) );
  OAI21_X1 U16409 ( .B1(n13050), .B2(n13368), .A(n13049), .ZN(P1_U2917) );
  INV_X1 U16410 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U16411 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20372), .B1(n16767), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13051) );
  OAI21_X1 U16412 ( .B1(n13052), .B2(n13368), .A(n13051), .ZN(P1_U2918) );
  INV_X1 U16413 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19455) );
  XNOR2_X1 U16414 ( .A(n13054), .B(n13053), .ZN(n16572) );
  INV_X1 U16415 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n13056) );
  NAND2_X1 U16416 ( .A1(n19499), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13055) );
  OAI21_X1 U16417 ( .B1(n19499), .B2(n13056), .A(n13055), .ZN(n19552) );
  INV_X1 U16418 ( .A(n19552), .ZN(n13057) );
  OAI222_X1 U16419 ( .A1(n19455), .A2(n16017), .B1(n16572), .B2(n16015), .C1(
        n19403), .C2(n13057), .ZN(P2_U2912) );
  NAND2_X1 U16420 ( .A1(n13059), .A2(n13058), .ZN(n13060) );
  NAND2_X1 U16421 ( .A1(n9867), .A2(n13060), .ZN(n16559) );
  INV_X1 U16422 ( .A(n19403), .ZN(n13625) );
  INV_X1 U16423 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17778) );
  NAND2_X1 U16424 ( .A1(n19499), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13061) );
  OAI21_X1 U16425 ( .B1(n19499), .B2(n17778), .A(n13061), .ZN(n15945) );
  AOI22_X1 U16426 ( .A1(n13625), .A2(n15945), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19396), .ZN(n13062) );
  OAI21_X1 U16427 ( .B1(n16559), .B2(n16015), .A(n13062), .ZN(P2_U2911) );
  NAND2_X1 U16428 ( .A1(n13063), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13064) );
  NAND4_X1 U16429 ( .A1(n13064), .A2(n19541), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19977), .ZN(n13065) );
  OAI21_X1 U16430 ( .B1(n13068), .B2(n13067), .A(n13724), .ZN(n15824) );
  NAND2_X1 U16431 ( .A1(n15887), .A2(n13069), .ZN(n15897) );
  MUX2_X1 U16432 ( .A(n16835), .B(n13070), .S(n9733), .Z(n13071) );
  OAI21_X1 U16433 ( .B1(n19501), .B2(n15897), .A(n13071), .ZN(P2_U2887) );
  NOR2_X1 U16434 ( .A1(n14381), .A2(n21102), .ZN(n13072) );
  OR2_X1 U16435 ( .A1(n20392), .A2(n20506), .ZN(n13278) );
  INV_X1 U16436 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n21259) );
  NOR2_X2 U16437 ( .A1(n20392), .A2(n12691), .ZN(n20405) );
  INV_X1 U16438 ( .A(n20405), .ZN(n13076) );
  INV_X1 U16439 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13117) );
  NOR2_X1 U16440 ( .A1(n20485), .A2(n13117), .ZN(n13074) );
  AOI21_X1 U16441 ( .B1(DATAI_15_), .B2(n20485), .A(n13074), .ZN(n14992) );
  INV_X1 U16442 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13075) );
  OAI222_X1 U16443 ( .A1(n13278), .A2(n21259), .B1(n13076), .B2(n14992), .C1(
        n13075), .C2(n13269), .ZN(P1_U2967) );
  MUX2_X1 U16444 ( .A(n13427), .B(n14414), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n13078) );
  OR2_X1 U16445 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13077) );
  XNOR2_X1 U16446 ( .A(n14873), .B(n14416), .ZN(n20470) );
  INV_X1 U16447 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14874) );
  INV_X1 U16448 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16449 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16450 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13082) );
  AOI22_X1 U16451 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13081) );
  AOI22_X1 U16452 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13080) );
  NAND4_X1 U16453 ( .A1(n13083), .A2(n13082), .A3(n13081), .A4(n13080), .ZN(
        n13089) );
  AOI22_X1 U16454 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16455 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U16456 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16457 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13084) );
  NAND4_X1 U16458 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13088) );
  NAND2_X1 U16459 ( .A1(n13090), .A2(n13401), .ZN(n13091) );
  OAI211_X1 U16460 ( .C1(n13835), .C2(n13093), .A(n13092), .B(n13091), .ZN(
        n13094) );
  INV_X1 U16461 ( .A(n13094), .ZN(n13095) );
  NAND2_X1 U16462 ( .A1(n13098), .A2(n13401), .ZN(n13099) );
  NAND2_X1 U16463 ( .A1(n13100), .A2(n13400), .ZN(n13101) );
  NAND2_X1 U16464 ( .A1(n20568), .A2(n13984), .ZN(n13106) );
  AOI22_X1 U16465 ( .A1(n14504), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n13022), .ZN(n13104) );
  NAND2_X1 U16466 ( .A1(n13389), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13103) );
  AND2_X1 U16467 ( .A1(n13104), .A2(n13103), .ZN(n13105) );
  NAND2_X1 U16468 ( .A1(n13106), .A2(n13105), .ZN(n13112) );
  INV_X1 U16469 ( .A(n13107), .ZN(n13108) );
  NOR2_X1 U16470 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14328) );
  OR2_X1 U16471 ( .A1(n13108), .A2(n14468), .ZN(n13109) );
  NAND2_X1 U16472 ( .A1(n13110), .A2(n13109), .ZN(n13111) );
  NAND2_X1 U16473 ( .A1(n13112), .A2(n13111), .ZN(n13393) );
  OR2_X1 U16474 ( .A1(n13112), .A2(n13111), .ZN(n13113) );
  NAND2_X1 U16475 ( .A1(n13393), .A2(n13113), .ZN(n14880) );
  OAI222_X1 U16476 ( .A1(n20470), .A2(n14930), .B1(n14874), .B2(n20355), .C1(
        n14880), .C2(n14932), .ZN(P1_U2871) );
  INV_X1 U16477 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13121) );
  NOR2_X1 U16478 ( .A1(n13114), .A2(n20103), .ZN(n13115) );
  INV_X1 U16479 ( .A(n13115), .ZN(n13116) );
  NOR2_X2 U16480 ( .A1(n13116), .A2(n19513), .ZN(n13222) );
  INV_X1 U16481 ( .A(n13222), .ZN(n13120) );
  INV_X1 U16482 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n13118) );
  MUX2_X1 U16483 ( .A(n13118), .B(n13117), .S(n19499), .Z(n13740) );
  INV_X1 U16484 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13119) );
  OAI222_X1 U16485 ( .A1(n13121), .A2(n13154), .B1(n13120), .B2(n13740), .C1(
        n13119), .C2(n19408), .ZN(P2_U2982) );
  AOI22_X1 U16486 ( .A1(n9734), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n13177), .ZN(n13124) );
  INV_X1 U16487 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U16488 ( .A1(n19499), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13122) );
  OAI21_X1 U16489 ( .B1(n19499), .B2(n13123), .A(n13122), .ZN(n15915) );
  NAND2_X1 U16490 ( .A1(n13222), .A2(n15915), .ZN(n13155) );
  NAND2_X1 U16491 ( .A1(n13124), .A2(n13155), .ZN(P2_U2980) );
  AOI22_X1 U16492 ( .A1(n9734), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n13136), .ZN(n13127) );
  INV_X1 U16493 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n13126) );
  NAND2_X1 U16494 ( .A1(n19499), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13125) );
  OAI21_X1 U16495 ( .B1(n19499), .B2(n13126), .A(n13125), .ZN(n15923) );
  NAND2_X1 U16496 ( .A1(n13222), .A2(n15923), .ZN(n13157) );
  NAND2_X1 U16497 ( .A1(n13127), .A2(n13157), .ZN(P2_U2979) );
  AOI22_X1 U16498 ( .A1(n9734), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n13136), .ZN(n13130) );
  INV_X1 U16499 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U16500 ( .A1(n19499), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13128) );
  OAI21_X1 U16501 ( .B1(n19499), .B2(n13129), .A(n13128), .ZN(n14521) );
  NAND2_X1 U16502 ( .A1(n13222), .A2(n14521), .ZN(n13159) );
  NAND2_X1 U16503 ( .A1(n13130), .A2(n13159), .ZN(P2_U2978) );
  AOI22_X1 U16504 ( .A1(n9734), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n13136), .ZN(n13133) );
  INV_X1 U16505 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n13132) );
  NAND2_X1 U16506 ( .A1(n19499), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13131) );
  OAI21_X1 U16507 ( .B1(n19499), .B2(n13132), .A(n13131), .ZN(n15938) );
  NAND2_X1 U16508 ( .A1(n13222), .A2(n15938), .ZN(n13161) );
  NAND2_X1 U16509 ( .A1(n13133), .A2(n13161), .ZN(P2_U2976) );
  AOI22_X1 U16510 ( .A1(n9734), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_7__SCAN_IN), .B2(n13136), .ZN(n13134) );
  NAND2_X1 U16511 ( .A1(n13222), .A2(n19552), .ZN(n13163) );
  NAND2_X1 U16512 ( .A1(n13134), .A2(n13163), .ZN(P2_U2974) );
  AOI22_X1 U16513 ( .A1(n9734), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_6__SCAN_IN), .B2(n13136), .ZN(n13135) );
  NAND2_X1 U16514 ( .A1(n13222), .A2(n19543), .ZN(n13169) );
  NAND2_X1 U16515 ( .A1(n13135), .A2(n13169), .ZN(P2_U2973) );
  AOI22_X1 U16516 ( .A1(n9734), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n13136), .ZN(n13139) );
  INV_X1 U16517 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n13138) );
  NAND2_X1 U16518 ( .A1(n19499), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13137) );
  OAI21_X1 U16519 ( .B1(n19499), .B2(n13138), .A(n13137), .ZN(n19535) );
  NAND2_X1 U16520 ( .A1(n13222), .A2(n19535), .ZN(n13173) );
  NAND2_X1 U16521 ( .A1(n13139), .A2(n13173), .ZN(P2_U2972) );
  AOI22_X1 U16522 ( .A1(n9734), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n13177), .ZN(n13142) );
  NAND2_X1 U16523 ( .A1(n19497), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13141) );
  NAND2_X1 U16524 ( .A1(n19499), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13140) );
  AND2_X1 U16525 ( .A1(n13141), .A2(n13140), .ZN(n19382) );
  INV_X1 U16526 ( .A(n19382), .ZN(n19530) );
  NAND2_X1 U16527 ( .A1(n13222), .A2(n19530), .ZN(n13171) );
  NAND2_X1 U16528 ( .A1(n13142), .A2(n13171), .ZN(P2_U2971) );
  AOI22_X1 U16529 ( .A1(n9734), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n13177), .ZN(n13145) );
  NAND2_X1 U16530 ( .A1(n19497), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13144) );
  NAND2_X1 U16531 ( .A1(n19499), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13143) );
  AND2_X1 U16532 ( .A1(n13144), .A2(n13143), .ZN(n19389) );
  INV_X1 U16533 ( .A(n19389), .ZN(n19525) );
  NAND2_X1 U16534 ( .A1(n13222), .A2(n19525), .ZN(n13165) );
  NAND2_X1 U16535 ( .A1(n13145), .A2(n13165), .ZN(P2_U2970) );
  AOI22_X1 U16536 ( .A1(n9734), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n13177), .ZN(n13147) );
  INV_X1 U16537 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18624) );
  NAND2_X1 U16538 ( .A1(n19499), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13146) );
  OAI21_X1 U16539 ( .B1(n19499), .B2(n18624), .A(n13146), .ZN(n19520) );
  NAND2_X1 U16540 ( .A1(n13222), .A2(n19520), .ZN(n13175) );
  NAND2_X1 U16541 ( .A1(n13147), .A2(n13175), .ZN(P2_U2969) );
  AOI22_X1 U16542 ( .A1(n9734), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_1__SCAN_IN), .B2(n13177), .ZN(n13150) );
  NAND2_X1 U16543 ( .A1(n19497), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U16544 ( .A1(n19499), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13148) );
  AND2_X1 U16545 ( .A1(n13149), .A2(n13148), .ZN(n19395) );
  INV_X1 U16546 ( .A(n19395), .ZN(n19515) );
  NAND2_X1 U16547 ( .A1(n13222), .A2(n19515), .ZN(n13167) );
  NAND2_X1 U16548 ( .A1(n13150), .A2(n13167), .ZN(P2_U2968) );
  AOI22_X1 U16549 ( .A1(n9734), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n13177), .ZN(n13153) );
  NAND2_X1 U16550 ( .A1(n19497), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U16551 ( .A1(n19499), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13151) );
  AND2_X1 U16552 ( .A1(n13152), .A2(n13151), .ZN(n19404) );
  INV_X1 U16553 ( .A(n19404), .ZN(n19506) );
  NAND2_X1 U16554 ( .A1(n13222), .A2(n19506), .ZN(n13178) );
  NAND2_X1 U16555 ( .A1(n13153), .A2(n13178), .ZN(P2_U2967) );
  AOI22_X1 U16556 ( .A1(n9734), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13177), .ZN(n13156) );
  NAND2_X1 U16557 ( .A1(n13156), .A2(n13155), .ZN(P2_U2965) );
  AOI22_X1 U16558 ( .A1(n9734), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n13177), .ZN(n13158) );
  NAND2_X1 U16559 ( .A1(n13158), .A2(n13157), .ZN(P2_U2964) );
  AOI22_X1 U16560 ( .A1(n9734), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13177), .ZN(n13160) );
  NAND2_X1 U16561 ( .A1(n13160), .A2(n13159), .ZN(P2_U2963) );
  AOI22_X1 U16562 ( .A1(n9734), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n13177), .ZN(n13162) );
  NAND2_X1 U16563 ( .A1(n13162), .A2(n13161), .ZN(P2_U2961) );
  AOI22_X1 U16564 ( .A1(n9734), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(
        P2_EAX_REG_23__SCAN_IN), .B2(n13177), .ZN(n13164) );
  NAND2_X1 U16565 ( .A1(n13164), .A2(n13163), .ZN(P2_U2959) );
  AOI22_X1 U16566 ( .A1(n9734), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n13177), .ZN(n13166) );
  NAND2_X1 U16567 ( .A1(n13166), .A2(n13165), .ZN(P2_U2955) );
  AOI22_X1 U16568 ( .A1(n9734), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n13177), .ZN(n13168) );
  NAND2_X1 U16569 ( .A1(n13168), .A2(n13167), .ZN(P2_U2953) );
  AOI22_X1 U16570 ( .A1(n9734), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n13177), .ZN(n13170) );
  NAND2_X1 U16571 ( .A1(n13170), .A2(n13169), .ZN(P2_U2958) );
  AOI22_X1 U16572 ( .A1(n9734), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13177), .ZN(n13172) );
  NAND2_X1 U16573 ( .A1(n13172), .A2(n13171), .ZN(P2_U2956) );
  AOI22_X1 U16574 ( .A1(n9734), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n13177), .ZN(n13174) );
  NAND2_X1 U16575 ( .A1(n13174), .A2(n13173), .ZN(P2_U2957) );
  AOI22_X1 U16576 ( .A1(n9734), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n13177), .ZN(n13176) );
  NAND2_X1 U16577 ( .A1(n13176), .A2(n13175), .ZN(P2_U2954) );
  AOI22_X1 U16578 ( .A1(n9734), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n13177), .ZN(n13179) );
  NAND2_X1 U16579 ( .A1(n13179), .A2(n13178), .ZN(P2_U2952) );
  AOI211_X1 U16580 ( .C1(n13181), .C2(n16654), .A(n13180), .B(n16846), .ZN(
        n13195) );
  NAND2_X1 U16581 ( .A1(n13183), .A2(n13182), .ZN(n13184) );
  XNOR2_X1 U16582 ( .A(n13184), .B(n16654), .ZN(n19482) );
  INV_X1 U16583 ( .A(n13185), .ZN(n13186) );
  OAI21_X1 U16584 ( .B1(n13187), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13186), .ZN(n19491) );
  OAI22_X1 U16585 ( .A1(n16625), .A2(n19482), .B1(n16842), .B2(n19491), .ZN(
        n13194) );
  OR2_X1 U16586 ( .A1(n13189), .A2(n13188), .ZN(n13190) );
  NAND2_X1 U16587 ( .A1(n13191), .A2(n13190), .ZN(n20203) );
  AOI22_X1 U16588 ( .A1(n16633), .A2(n19494), .B1(n16838), .B2(n20203), .ZN(
        n13192) );
  INV_X1 U16589 ( .A(n19333), .ZN(n19359) );
  NAND2_X1 U16590 ( .A1(n19359), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19488) );
  OAI211_X1 U16591 ( .C1(n16627), .C2(n16654), .A(n13192), .B(n19488), .ZN(
        n13193) );
  OR3_X1 U16592 ( .A1(n13195), .A2(n13194), .A3(n13193), .ZN(P2_U3045) );
  INV_X1 U16593 ( .A(n13196), .ZN(n13197) );
  NAND2_X1 U16594 ( .A1(n13197), .A2(n21102), .ZN(n13200) );
  OAI22_X1 U16595 ( .A1(n13328), .A2(n13200), .B1(n13199), .B2(n13198), .ZN(
        n13201) );
  INV_X2 U16596 ( .A(n14552), .ZN(n15007) );
  NAND2_X1 U16597 ( .A1(n13205), .A2(n20532), .ZN(n13206) );
  NAND2_X2 U16598 ( .A1(n15007), .A2(n13206), .ZN(n15009) );
  NOR2_X1 U16599 ( .A1(n14551), .A2(n12813), .ZN(n13207) );
  OR2_X1 U16600 ( .A1(n14552), .A2(n13208), .ZN(n14250) );
  INV_X1 U16601 ( .A(n14250), .ZN(n13209) );
  NAND2_X1 U16602 ( .A1(n20485), .A2(DATAI_1_), .ZN(n13212) );
  NAND2_X1 U16603 ( .A1(n20488), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13211) );
  AND2_X1 U16604 ( .A1(n13212), .A2(n13211), .ZN(n20508) );
  INV_X1 U16605 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20380) );
  OAI222_X1 U16606 ( .A1(n15009), .A2(n14880), .B1(n15006), .B2(n20508), .C1(
        n15007), .C2(n20380), .ZN(P1_U2903) );
  NAND2_X1 U16607 ( .A1(n20485), .A2(DATAI_0_), .ZN(n13214) );
  NAND2_X1 U16608 ( .A1(n20488), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13213) );
  AND2_X1 U16609 ( .A1(n13214), .A2(n13213), .ZN(n20499) );
  INV_X1 U16610 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20385) );
  OAI222_X1 U16611 ( .A1(n15009), .A2(n14888), .B1(n15006), .B2(n20499), .C1(
        n15007), .C2(n20385), .ZN(P1_U2904) );
  INV_X1 U16612 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19450) );
  NAND2_X1 U16613 ( .A1(n9734), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13216) );
  INV_X1 U16614 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17768) );
  NAND2_X1 U16615 ( .A1(n19499), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13215) );
  OAI21_X1 U16616 ( .B1(n19499), .B2(n17768), .A(n13215), .ZN(n15930) );
  NAND2_X1 U16617 ( .A1(n13222), .A2(n15930), .ZN(n13220) );
  OAI211_X1 U16618 ( .C1(n19450), .C2(n19408), .A(n13216), .B(n13220), .ZN(
        P2_U2977) );
  INV_X1 U16619 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n21340) );
  NAND2_X1 U16620 ( .A1(n9734), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13217) );
  NAND2_X1 U16621 ( .A1(n13222), .A2(n15945), .ZN(n13218) );
  OAI211_X1 U16622 ( .C1(n21340), .C2(n19408), .A(n13217), .B(n13218), .ZN(
        P2_U2960) );
  INV_X1 U16623 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19453) );
  NAND2_X1 U16624 ( .A1(n9734), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13219) );
  OAI211_X1 U16625 ( .C1(n19453), .C2(n19408), .A(n13219), .B(n13218), .ZN(
        P2_U2975) );
  INV_X1 U16626 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19419) );
  NAND2_X1 U16627 ( .A1(n9734), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13221) );
  OAI211_X1 U16628 ( .C1(n19419), .C2(n19408), .A(n13221), .B(n13220), .ZN(
        P2_U2962) );
  INV_X1 U16629 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19442) );
  NAND2_X1 U16630 ( .A1(n9734), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13223) );
  NAND2_X1 U16631 ( .A1(n13222), .A2(n13624), .ZN(n13224) );
  OAI211_X1 U16632 ( .C1(n19442), .C2(n19408), .A(n13223), .B(n13224), .ZN(
        P2_U2981) );
  INV_X1 U16633 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n21272) );
  NAND2_X1 U16634 ( .A1(n9734), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13225) );
  OAI211_X1 U16635 ( .C1(n21272), .C2(n19408), .A(n13225), .B(n13224), .ZN(
        P2_U2966) );
  NAND2_X1 U16636 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n14327), .ZN(n16822) );
  INV_X1 U16637 ( .A(n16822), .ZN(n13226) );
  NAND2_X1 U16638 ( .A1(n20908), .A2(n13226), .ZN(n20487) );
  INV_X1 U16639 ( .A(n13402), .ZN(n13227) );
  NAND2_X1 U16640 ( .A1(n14381), .A2(n13227), .ZN(n13231) );
  AND2_X1 U16641 ( .A1(n12797), .A2(n12892), .ZN(n13395) );
  INV_X1 U16642 ( .A(n13395), .ZN(n13230) );
  INV_X1 U16643 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13344) );
  NAND3_X1 U16644 ( .A1(n13231), .A2(n13230), .A3(n13344), .ZN(n13228) );
  AOI21_X1 U16645 ( .B1(n20490), .B2(n14376), .A(n13228), .ZN(n13240) );
  NAND2_X1 U16646 ( .A1(n13231), .A2(n13230), .ZN(n13236) );
  NOR2_X1 U16647 ( .A1(n13232), .A2(n13236), .ZN(n13234) );
  OAI21_X1 U16648 ( .B1(n13236), .B2(n14376), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13233) );
  AOI21_X1 U16649 ( .B1(n13235), .B2(n13234), .A(n13233), .ZN(n13239) );
  OR2_X1 U16650 ( .A1(n13237), .A2(n13236), .ZN(n13238) );
  NOR2_X1 U16651 ( .A1(n13240), .A2(n10052), .ZN(n13337) );
  OR2_X2 U16652 ( .A1(n13243), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20457) );
  INV_X1 U16653 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13242) );
  NOR2_X1 U16654 ( .A1(n20457), .A2(n13242), .ZN(n13352) );
  NAND2_X1 U16655 ( .A1(n21030), .A2(n13243), .ZN(n13244) );
  NAND2_X1 U16656 ( .A1(n13244), .A2(n21091), .ZN(n13245) );
  NAND2_X1 U16657 ( .A1(n21091), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13247) );
  NAND2_X1 U16658 ( .A1(n20832), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13246) );
  AND2_X1 U16659 ( .A1(n13247), .A2(n13246), .ZN(n13413) );
  INV_X1 U16660 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13248) );
  AOI21_X1 U16661 ( .B1(n15138), .B2(n13413), .A(n13248), .ZN(n13249) );
  AOI211_X1 U16662 ( .C1(n13337), .C2(n20429), .A(n13352), .B(n13249), .ZN(
        n13250) );
  OAI21_X1 U16663 ( .B1(n20487), .B2(n14888), .A(n13250), .ZN(P1_U2999) );
  INV_X1 U16664 ( .A(n13278), .ZN(n20393) );
  AOI22_X1 U16665 ( .A1(n20393), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20417), .ZN(n13254) );
  NAND2_X1 U16666 ( .A1(n20485), .A2(DATAI_4_), .ZN(n13252) );
  NAND2_X1 U16667 ( .A1(n20488), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13251) );
  AND2_X1 U16668 ( .A1(n13252), .A2(n13251), .ZN(n20520) );
  INV_X1 U16669 ( .A(n20520), .ZN(n13253) );
  NAND2_X1 U16670 ( .A1(n20405), .A2(n13253), .ZN(n13299) );
  NAND2_X1 U16671 ( .A1(n13254), .A2(n13299), .ZN(P1_U2956) );
  AOI22_X1 U16672 ( .A1(n20393), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20417), .ZN(n13258) );
  NAND2_X1 U16673 ( .A1(n20485), .A2(DATAI_5_), .ZN(n13256) );
  NAND2_X1 U16674 ( .A1(n20488), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13255) );
  AND2_X1 U16675 ( .A1(n13256), .A2(n13255), .ZN(n20524) );
  INV_X1 U16676 ( .A(n20524), .ZN(n13257) );
  NAND2_X1 U16677 ( .A1(n20405), .A2(n13257), .ZN(n13297) );
  NAND2_X1 U16678 ( .A1(n13258), .A2(n13297), .ZN(P1_U2957) );
  AOI22_X1 U16679 ( .A1(n20393), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20417), .ZN(n13260) );
  INV_X1 U16680 ( .A(DATAI_6_), .ZN(n21322) );
  INV_X1 U16681 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16949) );
  MUX2_X1 U16682 ( .A(n21322), .B(n16949), .S(n20488), .Z(n20528) );
  INV_X1 U16683 ( .A(n20528), .ZN(n13259) );
  NAND2_X1 U16684 ( .A1(n20405), .A2(n13259), .ZN(n13309) );
  NAND2_X1 U16685 ( .A1(n13260), .A2(n13309), .ZN(P1_U2958) );
  AOI22_X1 U16686 ( .A1(n20393), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20417), .ZN(n13264) );
  NAND2_X1 U16687 ( .A1(n20485), .A2(DATAI_3_), .ZN(n13262) );
  NAND2_X1 U16688 ( .A1(n20488), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13261) );
  AND2_X1 U16689 ( .A1(n13262), .A2(n13261), .ZN(n20516) );
  INV_X1 U16690 ( .A(n20516), .ZN(n13263) );
  NAND2_X1 U16691 ( .A1(n20405), .A2(n13263), .ZN(n13301) );
  NAND2_X1 U16692 ( .A1(n13264), .A2(n13301), .ZN(P1_U2955) );
  AOI22_X1 U16693 ( .A1(n20393), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20417), .ZN(n13268) );
  NAND2_X1 U16694 ( .A1(n20485), .A2(DATAI_7_), .ZN(n13266) );
  NAND2_X1 U16695 ( .A1(n20488), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13265) );
  AND2_X1 U16696 ( .A1(n13266), .A2(n13265), .ZN(n20536) );
  INV_X1 U16697 ( .A(n20536), .ZN(n13267) );
  NAND2_X1 U16698 ( .A1(n20405), .A2(n13267), .ZN(n13307) );
  NAND2_X1 U16699 ( .A1(n13268), .A2(n13307), .ZN(P1_U2959) );
  INV_X1 U16700 ( .A(n13269), .ZN(n20417) );
  AOI22_X1 U16701 ( .A1(n20393), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20417), .ZN(n13273) );
  INV_X1 U16702 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13270) );
  NOR2_X1 U16703 ( .A1(n20485), .A2(n13270), .ZN(n13271) );
  AOI21_X1 U16704 ( .B1(DATAI_14_), .B2(n20485), .A(n13271), .ZN(n14993) );
  INV_X1 U16705 ( .A(n14993), .ZN(n13272) );
  NAND2_X1 U16706 ( .A1(n20405), .A2(n13272), .ZN(n13287) );
  NAND2_X1 U16707 ( .A1(n13273), .A2(n13287), .ZN(P1_U2966) );
  NAND2_X1 U16708 ( .A1(n9867), .A2(n13275), .ZN(n13276) );
  NAND2_X1 U16709 ( .A1(n13274), .A2(n13276), .ZN(n16540) );
  INV_X1 U16710 ( .A(n15938), .ZN(n13277) );
  INV_X1 U16711 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n21406) );
  OAI222_X1 U16712 ( .A1(n16540), .A2(n16015), .B1(n13277), .B2(n19403), .C1(
        n21406), .C2(n16017), .ZN(P2_U2910) );
  AOI22_X1 U16713 ( .A1(n20418), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20417), .ZN(n13280) );
  INV_X1 U16714 ( .A(n20499), .ZN(n13279) );
  NAND2_X1 U16715 ( .A1(n20405), .A2(n13279), .ZN(n13295) );
  NAND2_X1 U16716 ( .A1(n13280), .A2(n13295), .ZN(P1_U2952) );
  AOI22_X1 U16717 ( .A1(n20418), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20417), .ZN(n13284) );
  NAND2_X1 U16718 ( .A1(n20485), .A2(DATAI_2_), .ZN(n13282) );
  NAND2_X1 U16719 ( .A1(n20488), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13281) );
  AND2_X1 U16720 ( .A1(n13282), .A2(n13281), .ZN(n20512) );
  INV_X1 U16721 ( .A(n20512), .ZN(n13283) );
  NAND2_X1 U16722 ( .A1(n20405), .A2(n13283), .ZN(n13303) );
  NAND2_X1 U16723 ( .A1(n13284), .A2(n13303), .ZN(P1_U2954) );
  AOI22_X1 U16724 ( .A1(n20418), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20417), .ZN(n13286) );
  INV_X1 U16725 ( .A(n20508), .ZN(n13285) );
  NAND2_X1 U16726 ( .A1(n20405), .A2(n13285), .ZN(n13305) );
  NAND2_X1 U16727 ( .A1(n13286), .A2(n13305), .ZN(P1_U2953) );
  AOI22_X1 U16728 ( .A1(n20418), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20417), .ZN(n13288) );
  NAND2_X1 U16729 ( .A1(n13288), .A2(n13287), .ZN(P1_U2951) );
  INV_X1 U16730 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13293) );
  MUX2_X1 U16731 ( .A(n13293), .B(n10830), .S(n15887), .Z(n13294) );
  OAI21_X1 U16732 ( .B1(n19502), .B2(n15897), .A(n13294), .ZN(P2_U2886) );
  AOI22_X1 U16733 ( .A1(n20418), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20417), .ZN(n13296) );
  NAND2_X1 U16734 ( .A1(n13296), .A2(n13295), .ZN(P1_U2937) );
  AOI22_X1 U16735 ( .A1(n20418), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20417), .ZN(n13298) );
  NAND2_X1 U16736 ( .A1(n13298), .A2(n13297), .ZN(P1_U2942) );
  AOI22_X1 U16737 ( .A1(n20418), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20417), .ZN(n13300) );
  NAND2_X1 U16738 ( .A1(n13300), .A2(n13299), .ZN(P1_U2941) );
  AOI22_X1 U16739 ( .A1(n20418), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20417), .ZN(n13302) );
  NAND2_X1 U16740 ( .A1(n13302), .A2(n13301), .ZN(P1_U2940) );
  AOI22_X1 U16741 ( .A1(n20418), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20417), .ZN(n13304) );
  NAND2_X1 U16742 ( .A1(n13304), .A2(n13303), .ZN(P1_U2939) );
  AOI22_X1 U16743 ( .A1(n20418), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20417), .ZN(n13306) );
  NAND2_X1 U16744 ( .A1(n13306), .A2(n13305), .ZN(P1_U2938) );
  AOI22_X1 U16745 ( .A1(n20418), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20417), .ZN(n13308) );
  NAND2_X1 U16746 ( .A1(n13308), .A2(n13307), .ZN(P1_U2944) );
  AOI22_X1 U16747 ( .A1(n20418), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20417), .ZN(n13310) );
  NAND2_X1 U16748 ( .A1(n13310), .A2(n13309), .ZN(P1_U2943) );
  NOR2_X1 U16749 ( .A1(n13315), .A2(n9733), .ZN(n13316) );
  AOI21_X1 U16750 ( .B1(P2_EBX_REG_2__SCAN_IN), .B2(n9733), .A(n13316), .ZN(
        n13317) );
  OAI21_X1 U16751 ( .B1(n20190), .B2(n15897), .A(n13317), .ZN(P2_U2885) );
  NAND3_X1 U16752 ( .A1(n13319), .A2(n21102), .A3(n13318), .ZN(n13325) );
  OAI21_X1 U16753 ( .B1(n20506), .B2(n13320), .A(n21102), .ZN(n14336) );
  OAI211_X1 U16754 ( .C1(n12901), .C2(n14336), .A(n12816), .B(n13208), .ZN(
        n13321) );
  INV_X1 U16755 ( .A(n13321), .ZN(n13322) );
  MUX2_X1 U16756 ( .A(n13325), .B(n13324), .S(n13323), .Z(n13330) );
  AOI21_X1 U16757 ( .B1(n13328), .B2(n13327), .A(n13326), .ZN(n13329) );
  AOI21_X2 U16758 ( .B1(n13330), .B2(n13329), .A(n20246), .ZN(n13345) );
  OAI21_X1 U16759 ( .B1(n13331), .B2(n13333), .A(n13332), .ZN(n13335) );
  OR2_X1 U16760 ( .A1(n13335), .A2(n13334), .ZN(n13336) );
  NAND2_X2 U16761 ( .A1(n13345), .A2(n13336), .ZN(n15456) );
  INV_X1 U16762 ( .A(n13337), .ZN(n13354) );
  OAI22_X1 U16763 ( .A1(n13331), .A2(n12812), .B1(n12897), .B2(n20506), .ZN(
        n13338) );
  INV_X1 U16764 ( .A(n15339), .ZN(n13350) );
  NAND2_X1 U16765 ( .A1(n13345), .A2(n13339), .ZN(n20452) );
  INV_X1 U16766 ( .A(n20452), .ZN(n15398) );
  NAND3_X1 U16767 ( .A1(n13342), .A2(n13341), .A3(n13340), .ZN(n13343) );
  AND2_X1 U16768 ( .A1(n13345), .A2(n13343), .ZN(n15341) );
  NAND2_X1 U16769 ( .A1(n15341), .A2(n13344), .ZN(n13348) );
  INV_X1 U16770 ( .A(n13345), .ZN(n13346) );
  NAND2_X1 U16771 ( .A1(n13346), .A2(n20457), .ZN(n13347) );
  NAND2_X1 U16772 ( .A1(n13348), .A2(n13347), .ZN(n14423) );
  AOI21_X1 U16773 ( .B1(n15398), .B2(n13344), .A(n14423), .ZN(n20482) );
  NOR3_X1 U16774 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15398), .A3(
        n15341), .ZN(n13349) );
  AOI21_X1 U16775 ( .B1(n13350), .B2(n20482), .A(n13349), .ZN(n13351) );
  AOI211_X1 U16776 ( .C1(n14885), .C2(n20454), .A(n13352), .B(n13351), .ZN(
        n13353) );
  OAI21_X1 U16777 ( .B1(n15456), .B2(n13354), .A(n13353), .ZN(P1_U3031) );
  INV_X1 U16778 ( .A(n13355), .ZN(n13358) );
  NAND2_X1 U16779 ( .A1(n13274), .A2(n13356), .ZN(n13357) );
  NAND2_X1 U16780 ( .A1(n13358), .A2(n13357), .ZN(n16520) );
  AOI22_X1 U16781 ( .A1(n13625), .A2(n15930), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19396), .ZN(n13359) );
  OAI21_X1 U16782 ( .B1(n16520), .B2(n16015), .A(n13359), .ZN(P2_U2909) );
  INV_X1 U16783 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13361) );
  AOI22_X1 U16784 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13360) );
  OAI21_X1 U16785 ( .B1(n13361), .B2(n13368), .A(n13360), .ZN(P1_U2916) );
  INV_X1 U16786 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13363) );
  AOI22_X1 U16787 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13362) );
  OAI21_X1 U16788 ( .B1(n13363), .B2(n13368), .A(n13362), .ZN(P1_U2914) );
  AOI22_X1 U16789 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13364) );
  OAI21_X1 U16790 ( .B1(n14948), .B2(n13368), .A(n13364), .ZN(P1_U2910) );
  INV_X1 U16791 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13366) );
  AOI22_X1 U16792 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13365) );
  OAI21_X1 U16793 ( .B1(n13366), .B2(n13368), .A(n13365), .ZN(P1_U2915) );
  INV_X1 U16794 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21235) );
  AOI22_X1 U16795 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20382), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20381), .ZN(n13367) );
  OAI21_X1 U16796 ( .B1(n21235), .B2(n13368), .A(n13367), .ZN(P1_U2906) );
  AOI22_X1 U16797 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U16798 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U16799 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U16800 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13371) );
  NAND4_X1 U16801 ( .A1(n13374), .A2(n13373), .A3(n13372), .A4(n13371), .ZN(
        n13380) );
  AOI22_X1 U16802 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U16803 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13377) );
  AOI22_X1 U16804 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U16805 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13375) );
  NAND4_X1 U16806 ( .A1(n13378), .A2(n13377), .A3(n13376), .A4(n13375), .ZN(
        n13379) );
  INV_X1 U16807 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13383) );
  INV_X1 U16808 ( .A(n13984), .ZN(n13874) );
  INV_X1 U16809 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13387) );
  XNOR2_X1 U16810 ( .A(n13387), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20345) );
  NAND2_X1 U16811 ( .A1(n13022), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13899) );
  OAI21_X1 U16812 ( .B1(n20345), .B2(n14468), .A(n13899), .ZN(n13388) );
  AOI21_X1 U16813 ( .B1(n14504), .B2(P1_EAX_REG_2__SCAN_IN), .A(n13388), .ZN(
        n13391) );
  NAND2_X1 U16814 ( .A1(n13389), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13390) );
  NAND2_X1 U16815 ( .A1(n14503), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13461) );
  OAI21_X1 U16816 ( .B1(n9808), .B2(n13394), .A(n13462), .ZN(n20342) );
  INV_X1 U16817 ( .A(n14376), .ZN(n14356) );
  NAND2_X1 U16818 ( .A1(n13402), .A2(n13401), .ZN(n13530) );
  XNOR2_X1 U16819 ( .A(n13530), .B(n13529), .ZN(n13396) );
  AOI21_X1 U16820 ( .B1(n13396), .B2(n14381), .A(n13395), .ZN(n13397) );
  INV_X1 U16821 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20463) );
  NAND2_X1 U16822 ( .A1(n20463), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13399) );
  NAND2_X1 U16823 ( .A1(n20481), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13398) );
  MUX2_X1 U16824 ( .A(n13399), .B(n13398), .S(n13545), .Z(n13409) );
  XNOR2_X1 U16825 ( .A(n13402), .B(n13401), .ZN(n13403) );
  INV_X1 U16826 ( .A(n14381), .ZN(n14387) );
  OAI211_X1 U16827 ( .C1(n13403), .C2(n14387), .A(n12863), .B(n12813), .ZN(
        n13404) );
  INV_X1 U16828 ( .A(n13404), .ZN(n13405) );
  NAND2_X1 U16829 ( .A1(n13545), .A2(n20481), .ZN(n13406) );
  NAND3_X1 U16830 ( .A1(n10159), .A2(n13406), .A3(n20463), .ZN(n13408) );
  OAI211_X1 U16831 ( .C1(n13545), .C2(n20481), .A(n13546), .B(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13407) );
  NAND3_X1 U16832 ( .A1(n13409), .A2(n13408), .A3(n13407), .ZN(n13410) );
  NAND2_X1 U16833 ( .A1(n13411), .A2(n13410), .ZN(n13548) );
  OAI21_X1 U16834 ( .B1(n13411), .B2(n13410), .A(n13548), .ZN(n13412) );
  INV_X1 U16835 ( .A(n13412), .ZN(n20462) );
  INV_X1 U16836 ( .A(n20345), .ZN(n13415) );
  INV_X1 U16837 ( .A(n20457), .ZN(n20436) );
  AOI22_X1 U16838 ( .A1(n20421), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20436), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13414) );
  OAI21_X1 U16839 ( .B1(n20433), .B2(n13415), .A(n13414), .ZN(n13416) );
  AOI21_X1 U16840 ( .B1(n20462), .B2(n20429), .A(n13416), .ZN(n13417) );
  OAI21_X1 U16841 ( .B1(n20342), .B2(n20487), .A(n13417), .ZN(P1_U2997) );
  OAI21_X1 U16842 ( .B1(n13418), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13544), .ZN(n20473) );
  MUX2_X1 U16843 ( .A(n20433), .B(n15138), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13420) );
  INV_X1 U16844 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13419) );
  OR2_X1 U16845 ( .A1(n20457), .A2(n13419), .ZN(n20469) );
  OAI211_X1 U16846 ( .C1(n20473), .C2(n20253), .A(n13420), .B(n20469), .ZN(
        n13421) );
  INV_X1 U16847 ( .A(n13421), .ZN(n13422) );
  OAI21_X1 U16848 ( .B1(n20487), .B2(n14880), .A(n13422), .ZN(P1_U2998) );
  OAI21_X1 U16849 ( .B1(n13355), .B2(n13424), .A(n13423), .ZN(n16513) );
  INV_X1 U16850 ( .A(n14521), .ZN(n13425) );
  INV_X1 U16851 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19448) );
  OAI222_X1 U16852 ( .A1(n16513), .A2(n16015), .B1(n13425), .B2(n19403), .C1(
        n19448), .C2(n16017), .ZN(P2_U2908) );
  INV_X1 U16853 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20378) );
  OAI222_X1 U16854 ( .A1(n15009), .A2(n20342), .B1(n15006), .B2(n20512), .C1(
        n15007), .C2(n20378), .ZN(P1_U2902) );
  NOR2_X1 U16855 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13428) );
  NOR2_X1 U16856 ( .A1(n13429), .A2(n13428), .ZN(n13430) );
  NAND2_X1 U16857 ( .A1(n13431), .A2(n13430), .ZN(n13589) );
  OR2_X1 U16858 ( .A1(n13431), .A2(n13430), .ZN(n13432) );
  NAND2_X1 U16859 ( .A1(n13589), .A2(n13432), .ZN(n20332) );
  INV_X1 U16860 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13433) );
  OAI222_X1 U16861 ( .A1(n20332), .A2(n14930), .B1(n13433), .B2(n20355), .C1(
        n20342), .C2(n14932), .ZN(P1_U2870) );
  XNOR2_X2 U16862 ( .A(n21501), .B(n13435), .ZN(n19807) );
  MUX2_X1 U16863 ( .A(n13436), .B(n11032), .S(n9733), .Z(n13437) );
  OAI21_X1 U16864 ( .B1(n19807), .B2(n15897), .A(n13437), .ZN(P2_U2884) );
  INV_X1 U16865 ( .A(n20775), .ZN(n13447) );
  XNOR2_X1 U16866 ( .A(n12963), .B(n12726), .ZN(n13445) );
  MUX2_X1 U16867 ( .A(n13438), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n12958), .Z(n13439) );
  INV_X1 U16868 ( .A(n12958), .ZN(n15470) );
  AOI211_X1 U16869 ( .C1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n15470), .A(
        n13441), .B(n14230), .ZN(n15484) );
  NOR3_X1 U16870 ( .A1(n15474), .A2(n15484), .A3(n13442), .ZN(n13443) );
  AOI211_X1 U16871 ( .C1(n14537), .C2(n13445), .A(n13444), .B(n13443), .ZN(
        n13446) );
  OAI21_X1 U16872 ( .B1(n13447), .B2(n14538), .A(n13446), .ZN(n15483) );
  MUX2_X1 U16873 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15483), .S(
        n16730), .Z(n16737) );
  NOR2_X1 U16874 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21090), .ZN(n13453) );
  AOI22_X1 U16875 ( .A1(n16737), .A2(n21090), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13453), .ZN(n13450) );
  MUX2_X1 U16876 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13448), .S(
        n16730), .Z(n16735) );
  AOI22_X1 U16877 ( .A1(n13453), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16735), .B2(n21090), .ZN(n13449) );
  NOR2_X1 U16878 ( .A1(n13450), .A2(n13449), .ZN(n16747) );
  INV_X1 U16879 ( .A(n13451), .ZN(n15471) );
  NAND2_X1 U16880 ( .A1(n16747), .A2(n15471), .ZN(n13458) );
  OAI21_X1 U16881 ( .B1(n20319), .B2(n12935), .A(n16730), .ZN(n13455) );
  INV_X1 U16882 ( .A(n16730), .ZN(n13452) );
  AOI21_X1 U16883 ( .B1(n13452), .B2(n13580), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13454) );
  AOI22_X1 U16884 ( .A1(n13455), .A2(n13454), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13453), .ZN(n16745) );
  AND3_X1 U16885 ( .A1(n13458), .A2(n16745), .A3(n20254), .ZN(n13456) );
  AND3_X1 U16886 ( .A1(n13458), .A2(n16745), .A3(n13457), .ZN(n16758) );
  INV_X1 U16887 ( .A(n13020), .ZN(n14881) );
  INV_X1 U16888 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20913) );
  NAND2_X1 U16889 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20913), .ZN(n15465) );
  INV_X1 U16890 ( .A(n15465), .ZN(n15460) );
  OAI22_X1 U16891 ( .A1(n20567), .A2(n21030), .B1(n14881), .B2(n15460), .ZN(
        n13459) );
  OAI21_X1 U16892 ( .B1(n16758), .B2(n13459), .A(n20483), .ZN(n13460) );
  OAI21_X1 U16893 ( .B1(n20483), .B2(n20953), .A(n13460), .ZN(P1_U3478) );
  AOI22_X1 U16894 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13467) );
  INV_X1 U16895 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n21319) );
  AOI22_X1 U16896 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U16897 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U16898 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13464) );
  NAND4_X1 U16899 ( .A1(n13467), .A2(n13466), .A3(n13465), .A4(n13464), .ZN(
        n13473) );
  AOI22_X1 U16900 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U16901 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U16902 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U16903 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13468) );
  NAND4_X1 U16904 ( .A1(n13471), .A2(n13470), .A3(n13469), .A4(n13468), .ZN(
        n13472) );
  AOI22_X1 U16905 ( .A1(n13833), .A2(n13537), .B1(n13830), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U16906 ( .A1(n15462), .A2(n13984), .ZN(n13483) );
  INV_X1 U16908 ( .A(n13476), .ZN(n13478) );
  INV_X1 U16909 ( .A(n13577), .ZN(n13477) );
  OAI21_X1 U16910 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13478), .A(
        n13477), .ZN(n14857) );
  AOI22_X1 U16911 ( .A1(n14502), .A2(n14857), .B1(n14503), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13480) );
  NAND2_X1 U16912 ( .A1(n14504), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n13479) );
  OAI211_X1 U16913 ( .C1(n13581), .C2(n10219), .A(n13480), .B(n13479), .ZN(
        n13481) );
  INV_X1 U16914 ( .A(n13481), .ZN(n13482) );
  NAND2_X1 U16915 ( .A1(n13892), .A2(n13904), .ZN(n13610) );
  OAI21_X1 U16916 ( .B1(n13892), .B2(n13904), .A(n13610), .ZN(n14870) );
  INV_X1 U16917 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14860) );
  NAND2_X1 U16918 ( .A1(n14413), .A2(n14860), .ZN(n13486) );
  NAND2_X1 U16919 ( .A1(n14314), .A2(n9973), .ZN(n13484) );
  OAI211_X1 U16920 ( .C1(n14416), .C2(P1_EBX_REG_3__SCAN_IN), .A(n13484), .B(
        n14414), .ZN(n13485) );
  NAND2_X1 U16921 ( .A1(n13486), .A2(n13485), .ZN(n13585) );
  XOR2_X1 U16922 ( .A(n13589), .B(n13585), .Z(n14862) );
  INV_X1 U16923 ( .A(n14862), .ZN(n20444) );
  AOI22_X1 U16924 ( .A1(n20350), .A2(n20444), .B1(n14922), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13487) );
  OAI21_X1 U16925 ( .B1(n14870), .B2(n14932), .A(n13487), .ZN(P1_U2869) );
  INV_X1 U16926 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19446) );
  INV_X1 U16927 ( .A(n15923), .ZN(n13489) );
  XNOR2_X1 U16928 ( .A(n13423), .B(n13488), .ZN(n16497) );
  OAI222_X1 U16929 ( .A1(n16017), .A2(n19446), .B1(n13489), .B2(n19403), .C1(
        n16497), .C2(n16015), .ZN(P2_U2907) );
  INV_X1 U16930 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20376) );
  OAI222_X1 U16931 ( .A1(n15009), .A2(n14870), .B1(n15006), .B2(n20516), .C1(
        n15007), .C2(n20376), .ZN(P1_U2901) );
  AND2_X1 U16932 ( .A1(n13490), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13493) );
  NAND2_X1 U16933 ( .A1(n13491), .A2(n13493), .ZN(n13601) );
  INV_X1 U16934 ( .A(n13492), .ZN(n13494) );
  OR3_X1 U16935 ( .A1(n13495), .A2(n13494), .A3(n13493), .ZN(n13496) );
  NAND2_X1 U16936 ( .A1(n13601), .A2(n13496), .ZN(n19378) );
  NOR2_X1 U16937 ( .A1(n13499), .A2(n13498), .ZN(n13500) );
  OR2_X1 U16938 ( .A1(n13497), .A2(n13500), .ZN(n16607) );
  NOR2_X1 U16939 ( .A1(n16607), .A2(n9733), .ZN(n13501) );
  AOI21_X1 U16940 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n9733), .A(n13501), .ZN(
        n13502) );
  OAI21_X1 U16941 ( .B1(n19378), .B2(n15897), .A(n13502), .ZN(P2_U2883) );
  AOI22_X1 U16942 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U16943 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14476), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13505) );
  AOI22_X1 U16944 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13504) );
  AOI22_X1 U16945 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13503) );
  NAND4_X1 U16946 ( .A1(n13506), .A2(n13505), .A3(n13504), .A4(n13503), .ZN(
        n13512) );
  AOI22_X1 U16947 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n14477), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13510) );
  AOI22_X1 U16948 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14171), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13509) );
  AOI22_X1 U16949 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13508) );
  AOI22_X1 U16950 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13507) );
  NAND4_X1 U16951 ( .A1(n13510), .A2(n13509), .A3(n13508), .A4(n13507), .ZN(
        n13511) );
  NAND2_X1 U16952 ( .A1(n13833), .A2(n13539), .ZN(n13514) );
  NAND2_X1 U16953 ( .A1(n13830), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13513) );
  NAND2_X1 U16954 ( .A1(n13514), .A2(n13513), .ZN(n13536) );
  AOI22_X1 U16955 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14475), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13519) );
  AOI22_X1 U16956 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U16957 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U16958 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13516) );
  NAND4_X1 U16959 ( .A1(n13519), .A2(n13518), .A3(n13517), .A4(n13516), .ZN(
        n13525) );
  INV_X1 U16960 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n21323) );
  AOI22_X1 U16961 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U16962 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U16963 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U16964 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13520) );
  NAND4_X1 U16965 ( .A1(n13523), .A2(n13522), .A3(n13521), .A4(n13520), .ZN(
        n13524) );
  OR2_X1 U16966 ( .A1(n13525), .A2(n13524), .ZN(n14368) );
  NAND2_X1 U16967 ( .A1(n13833), .A2(n14368), .ZN(n13527) );
  NAND2_X1 U16968 ( .A1(n13830), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13526) );
  NAND2_X1 U16969 ( .A1(n13527), .A2(n13526), .ZN(n13528) );
  NAND2_X1 U16970 ( .A1(n13530), .A2(n13529), .ZN(n13538) );
  AND2_X1 U16971 ( .A1(n13537), .A2(n13539), .ZN(n13531) );
  NAND2_X1 U16972 ( .A1(n13538), .A2(n13531), .ZN(n14367) );
  XNOR2_X1 U16973 ( .A(n14367), .B(n14368), .ZN(n13532) );
  NAND2_X1 U16974 ( .A1(n13532), .A2(n14381), .ZN(n13533) );
  INV_X1 U16975 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13555) );
  INV_X1 U16976 ( .A(n13537), .ZN(n13534) );
  XNOR2_X1 U16977 ( .A(n13538), .B(n13534), .ZN(n13535) );
  NAND2_X1 U16978 ( .A1(n13538), .A2(n13537), .ZN(n13540) );
  XNOR2_X1 U16979 ( .A(n13540), .B(n13539), .ZN(n13541) );
  NAND2_X1 U16980 ( .A1(n13541), .A2(n14381), .ZN(n13542) );
  NAND3_X1 U16981 ( .A1(n13543), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13549) );
  OAI21_X1 U16982 ( .B1(n13551), .B2(n13550), .A(n14364), .ZN(n16802) );
  NOR2_X1 U16983 ( .A1(n20463), .A2(n20481), .ZN(n20450) );
  INV_X2 U16984 ( .A(n15426), .ZN(n20460) );
  INV_X1 U16985 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13561) );
  NOR2_X1 U16986 ( .A1(n13561), .A2(n9973), .ZN(n20434) );
  OAI21_X1 U16987 ( .B1(n13344), .B2(n20481), .A(n20463), .ZN(n20438) );
  AND3_X1 U16988 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20434), .A3(
        n20438), .ZN(n15406) );
  NOR2_X1 U16989 ( .A1(n20452), .A2(n15406), .ZN(n13552) );
  NOR2_X1 U16990 ( .A1(n14423), .A2(n13552), .ZN(n15432) );
  OAI221_X1 U16991 ( .B1(n20450), .B2(n20460), .C1(n20434), .C2(n20460), .A(
        n15432), .ZN(n13553) );
  INV_X1 U16992 ( .A(n13553), .ZN(n15442) );
  NAND2_X1 U16993 ( .A1(n20434), .A2(n13555), .ZN(n15443) );
  NAND2_X1 U16994 ( .A1(n20464), .A2(n20450), .ZN(n15444) );
  NAND2_X1 U16995 ( .A1(n15444), .A2(n20452), .ZN(n15407) );
  NAND2_X1 U16996 ( .A1(n20438), .A2(n15407), .ZN(n20449) );
  OAI22_X1 U16997 ( .A1(n15442), .A2(n13555), .B1(n15443), .B2(n20449), .ZN(
        n13554) );
  INV_X1 U16998 ( .A(n13554), .ZN(n13567) );
  NAND2_X1 U16999 ( .A1(n14413), .A2(n20304), .ZN(n13558) );
  OAI21_X1 U17000 ( .B1(n14318), .B2(n13555), .A(n14314), .ZN(n13556) );
  OAI21_X1 U17001 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n14416), .A(n13556), .ZN(
        n13557) );
  INV_X1 U17002 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13559) );
  NAND2_X1 U17003 ( .A1(n14319), .A2(n13559), .ZN(n13563) );
  NAND2_X1 U17004 ( .A1(n14409), .A2(n13559), .ZN(n13560) );
  OAI211_X1 U17005 ( .C1(n14318), .C2(n13561), .A(n13560), .B(n14314), .ZN(
        n13562) );
  AOI21_X1 U17006 ( .B1(n13565), .B2(n13590), .A(n14256), .ZN(n20307) );
  AOI22_X1 U17007 ( .A1(n20454), .A2(n20307), .B1(n20436), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n13566) );
  OAI211_X1 U17008 ( .C1(n16802), .C2(n15456), .A(n13567), .B(n13566), .ZN(
        P1_U3026) );
  XOR2_X1 U17009 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13601), .Z(n13573)
         );
  OR2_X1 U17010 ( .A1(n13497), .A2(n13569), .ZN(n13570) );
  NAND2_X1 U17011 ( .A1(n13568), .A2(n13570), .ZN(n16597) );
  MUX2_X1 U17012 ( .A(n16597), .B(n13571), .S(n9733), .Z(n13572) );
  OAI21_X1 U17013 ( .B1(n13573), .B2(n15897), .A(n13572), .ZN(P2_U2882) );
  AND2_X1 U17014 ( .A1(n13984), .A2(n13574), .ZN(n13575) );
  NAND2_X1 U17015 ( .A1(n13576), .A2(n13575), .ZN(n13584) );
  OAI21_X1 U17016 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13577), .A(
        n13611), .ZN(n20432) );
  OAI21_X1 U17017 ( .B1(n20832), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13022), .ZN(n13579) );
  NAND2_X1 U17018 ( .A1(n14504), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13578) );
  OAI211_X1 U17019 ( .C1(n13581), .C2(n13580), .A(n13579), .B(n13578), .ZN(
        n13582) );
  OAI21_X1 U17020 ( .B1(n14468), .B2(n20432), .A(n13582), .ZN(n13583) );
  XNOR2_X1 U17021 ( .A(n13610), .B(n13891), .ZN(n20427) );
  INV_X1 U17022 ( .A(n20427), .ZN(n13598) );
  INV_X1 U17023 ( .A(n13585), .ZN(n13588) );
  INV_X1 U17024 ( .A(n13586), .ZN(n13587) );
  OAI21_X1 U17025 ( .B1(n13589), .B2(n13588), .A(n13587), .ZN(n13591) );
  AND2_X1 U17026 ( .A1(n13591), .A2(n13590), .ZN(n20437) );
  AOI22_X1 U17027 ( .A1(n20350), .A2(n20437), .B1(n14922), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13592) );
  OAI21_X1 U17028 ( .B1(n13598), .B2(n14932), .A(n13592), .ZN(P1_U2868) );
  XNOR2_X1 U17029 ( .A(n20423), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13594) );
  NOR2_X1 U17030 ( .A1(n13594), .A2(n13593), .ZN(n20422) );
  AOI21_X1 U17031 ( .B1(n13594), .B2(n13593), .A(n20422), .ZN(n20446) );
  NAND2_X1 U17032 ( .A1(n20446), .A2(n20429), .ZN(n13597) );
  AND2_X1 U17033 ( .A1(n20436), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20443) );
  NOR2_X1 U17034 ( .A1(n20433), .A2(n14857), .ZN(n13595) );
  AOI211_X1 U17035 ( .C1(n20421), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20443), .B(n13595), .ZN(n13596) );
  OAI211_X1 U17036 ( .C1(n20487), .C2(n14870), .A(n13597), .B(n13596), .ZN(
        P1_U2996) );
  INV_X1 U17037 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20374) );
  OAI222_X1 U17038 ( .A1(n15009), .A2(n13598), .B1(n20374), .B2(n15007), .C1(
        n15006), .C2(n20520), .ZN(P1_U2900) );
  INV_X1 U17039 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13608) );
  INV_X1 U17040 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13599) );
  NOR2_X1 U17041 ( .A1(n13601), .A2(n13599), .ZN(n13602) );
  OAI211_X1 U17042 ( .C1(n13602), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15904), .B(n13754), .ZN(n13607) );
  NAND2_X1 U17043 ( .A1(n13568), .A2(n13603), .ZN(n13604) );
  NAND2_X1 U17044 ( .A1(n13732), .A2(n13604), .ZN(n19369) );
  INV_X1 U17045 ( .A(n19369), .ZN(n13605) );
  NAND2_X1 U17046 ( .A1(n13605), .A2(n15887), .ZN(n13606) );
  OAI211_X1 U17047 ( .C1(n15887), .C2(n13608), .A(n13607), .B(n13606), .ZN(
        P2_U2881) );
  INV_X1 U17048 ( .A(n13891), .ZN(n13609) );
  INV_X1 U17049 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13614) );
  OAI21_X1 U17050 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13612), .A(
        n13838), .ZN(n20313) );
  NAND2_X1 U17051 ( .A1(n20313), .A2(n14502), .ZN(n13613) );
  OAI21_X1 U17052 ( .B1(n13614), .B2(n13899), .A(n13613), .ZN(n13615) );
  AOI21_X1 U17053 ( .B1(n14504), .B2(P1_EAX_REG_5__SCAN_IN), .A(n13615), .ZN(
        n13616) );
  NOR2_X1 U17054 ( .A1(n13618), .A2(n13905), .ZN(n13619) );
  INV_X1 U17055 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20371) );
  OAI222_X1 U17056 ( .A1(n15009), .A2(n16803), .B1(n20524), .B2(n15006), .C1(
        n15007), .C2(n20371), .ZN(P1_U2899) );
  NOR2_X1 U17057 ( .A1(n13621), .A2(n13622), .ZN(n13623) );
  OR2_X1 U17058 ( .A1(n13620), .A2(n13623), .ZN(n16475) );
  AOI22_X1 U17059 ( .A1(n13625), .A2(n13624), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19396), .ZN(n13626) );
  OAI21_X1 U17060 ( .B1(n16475), .B2(n16015), .A(n13626), .ZN(P2_U2905) );
  INV_X1 U17061 ( .A(n13661), .ZN(n13653) );
  NAND2_X1 U17062 ( .A1(n13663), .A2(n13627), .ZN(n13658) );
  NAND2_X1 U17063 ( .A1(n13663), .A2(n10789), .ZN(n13628) );
  AND2_X1 U17064 ( .A1(n13658), .A2(n13628), .ZN(n13646) );
  NOR2_X1 U17065 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13635) );
  NOR2_X1 U17066 ( .A1(n13629), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13643) );
  INV_X1 U17067 ( .A(n13630), .ZN(n13681) );
  OR2_X1 U17068 ( .A1(n13682), .A2(n13681), .ZN(n13639) );
  OAI21_X1 U17069 ( .B1(n13631), .B2(n13643), .A(n13639), .ZN(n13634) );
  AOI21_X1 U17070 ( .B1(n13632), .B2(n11363), .A(n13631), .ZN(n13644) );
  INV_X1 U17071 ( .A(n13643), .ZN(n13638) );
  NAND2_X1 U17072 ( .A1(n13644), .A2(n13638), .ZN(n13633) );
  OAI211_X1 U17073 ( .C1(n13646), .C2(n13635), .A(n13634), .B(n13633), .ZN(
        n13636) );
  AOI21_X1 U17074 ( .B1(n19479), .B2(n13653), .A(n13636), .ZN(n16660) );
  NOR2_X1 U17075 ( .A1(n13691), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13637) );
  AOI21_X1 U17076 ( .B1(n16660), .B2(n13691), .A(n13637), .ZN(n13675) );
  OR2_X1 U17077 ( .A1(n13436), .A2(n13661), .ZN(n13651) );
  NAND2_X1 U17078 ( .A1(n13639), .A2(n13638), .ZN(n13642) );
  NAND3_X1 U17079 ( .A1(n13663), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13640) );
  NAND3_X1 U17080 ( .A1(n13642), .A2(n13641), .A3(n13640), .ZN(n13648) );
  INV_X1 U17081 ( .A(n13644), .ZN(n13645) );
  NAND3_X1 U17082 ( .A1(n13638), .A2(n13646), .A3(n13645), .ZN(n13647) );
  MUX2_X1 U17083 ( .A(n13648), .B(n13647), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13649) );
  INV_X1 U17084 ( .A(n13649), .ZN(n13650) );
  AND2_X1 U17085 ( .A1(n13651), .A2(n13650), .ZN(n16665) );
  NOR2_X1 U17086 ( .A1(n13691), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13652) );
  AOI21_X1 U17087 ( .B1(n16665), .B2(n13691), .A(n13652), .ZN(n13676) );
  AOI21_X1 U17088 ( .B1(n13675), .B2(n20196), .A(n13676), .ZN(n13673) );
  NAND2_X1 U17089 ( .A1(n19494), .A2(n13653), .ZN(n13660) );
  OAI21_X1 U17090 ( .B1(n13656), .B2(n13655), .A(n13662), .ZN(n13657) );
  AND2_X1 U17091 ( .A1(n13658), .A2(n13657), .ZN(n13659) );
  NAND2_X1 U17092 ( .A1(n13660), .A2(n13659), .ZN(n16655) );
  OR2_X1 U17093 ( .A1(n16835), .A2(n13661), .ZN(n13667) );
  INV_X1 U17094 ( .A(n13662), .ZN(n13665) );
  INV_X1 U17095 ( .A(n13663), .ZN(n13664) );
  MUX2_X1 U17096 ( .A(n13665), .B(n13664), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13666) );
  AND2_X1 U17097 ( .A1(n13667), .A2(n13666), .ZN(n16649) );
  INV_X1 U17098 ( .A(n16649), .ZN(n13668) );
  OAI22_X1 U17099 ( .A1(n16655), .A2(n20205), .B1(n13668), .B2(n12154), .ZN(
        n13671) );
  NAND2_X1 U17100 ( .A1(n16655), .A2(n20205), .ZN(n13670) );
  INV_X1 U17101 ( .A(n13691), .ZN(n13669) );
  AOI21_X1 U17102 ( .B1(n13671), .B2(n13670), .A(n13669), .ZN(n13674) );
  OAI21_X1 U17103 ( .B1(n13675), .B2(n20196), .A(n13674), .ZN(n13672) );
  AOI211_X1 U17104 ( .C1(n13673), .C2(n13672), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n13695) );
  INV_X1 U17105 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21284) );
  NAND3_X1 U17106 ( .A1(n13674), .A2(n20196), .A3(n21284), .ZN(n13679) );
  INV_X1 U17107 ( .A(n13675), .ZN(n13678) );
  INV_X1 U17108 ( .A(n13676), .ZN(n13677) );
  AOI21_X1 U17109 ( .B1(n13679), .B2(n13678), .A(n13677), .ZN(n13694) );
  INV_X1 U17110 ( .A(n13680), .ZN(n13684) );
  MUX2_X1 U17111 ( .A(n13682), .B(n13681), .S(n13765), .Z(n13683) );
  AOI21_X1 U17112 ( .B1(n11573), .B2(n13684), .A(n13683), .ZN(n20223) );
  INV_X1 U17113 ( .A(n20223), .ZN(n13693) );
  AOI22_X1 U17114 ( .A1(n13687), .A2(n19513), .B1(n13686), .B2(n13685), .ZN(
        n13690) );
  OAI21_X1 U17115 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n13688), .ZN(n13689) );
  OAI211_X1 U17116 ( .C1(n13691), .C2(n11199), .A(n13690), .B(n13689), .ZN(
        n13692) );
  NOR4_X1 U17117 ( .A1(n13695), .A2(n13694), .A3(n13693), .A4(n13692), .ZN(
        n13776) );
  AOI21_X1 U17118 ( .B1(n13776), .B2(n16648), .A(n11619), .ZN(n13700) );
  NAND3_X1 U17119 ( .A1(n13697), .A2(n20226), .A3(n13696), .ZN(n13699) );
  NOR2_X1 U17120 ( .A1(n13698), .A2(n20207), .ZN(n20234) );
  NAND2_X1 U17121 ( .A1(n13699), .A2(n20234), .ZN(n13766) );
  INV_X1 U17122 ( .A(n13730), .ZN(n13767) );
  INV_X1 U17123 ( .A(n13772), .ZN(n16773) );
  OAI211_X1 U17124 ( .C1(n13767), .C2(n19977), .A(n16773), .B(n13701), .ZN(
        P2_U3593) );
  INV_X1 U17125 ( .A(n19520), .ZN(n13717) );
  OR2_X1 U17126 ( .A1(n13703), .A2(n13702), .ZN(n13704) );
  NAND2_X1 U17127 ( .A1(n13705), .A2(n13704), .ZN(n20194) );
  XNOR2_X1 U17128 ( .A(n20190), .B(n20194), .ZN(n13713) );
  NOR2_X1 U17129 ( .A1(n20199), .A2(n20203), .ZN(n13710) );
  AOI21_X1 U17130 ( .B1(n20199), .B2(n20203), .A(n13710), .ZN(n19391) );
  OR2_X1 U17131 ( .A1(n13707), .A2(n13706), .ZN(n13709) );
  AND2_X1 U17132 ( .A1(n13709), .A2(n13708), .ZN(n19400) );
  NAND2_X1 U17133 ( .A1(n20211), .A2(n19400), .ZN(n19399) );
  NAND2_X1 U17134 ( .A1(n19391), .A2(n19399), .ZN(n19390) );
  INV_X1 U17135 ( .A(n13710), .ZN(n13711) );
  NAND2_X1 U17136 ( .A1(n19390), .A2(n13711), .ZN(n13712) );
  NAND2_X1 U17137 ( .A1(n13712), .A2(n13713), .ZN(n16019) );
  OAI21_X1 U17138 ( .B1(n13713), .B2(n13712), .A(n16019), .ZN(n13714) );
  NAND2_X1 U17139 ( .A1(n13714), .A2(n19398), .ZN(n13716) );
  AOI22_X1 U17140 ( .A1(n19397), .A2(n20194), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19396), .ZN(n13715) );
  OAI211_X1 U17141 ( .C1(n13717), .C2(n19403), .A(n13716), .B(n13715), .ZN(
        P2_U2917) );
  AND2_X1 U17142 ( .A1(n13719), .A2(n13718), .ZN(n13720) );
  NOR2_X1 U17143 ( .A1(n13621), .A2(n13720), .ZN(n16488) );
  INV_X1 U17144 ( .A(n16488), .ZN(n13722) );
  INV_X1 U17145 ( .A(n15915), .ZN(n13721) );
  INV_X1 U17146 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19444) );
  OAI222_X1 U17147 ( .A1(n13722), .A2(n16015), .B1(n13721), .B2(n19403), .C1(
        n19444), .C2(n16017), .ZN(P2_U2906) );
  INV_X1 U17148 ( .A(n20307), .ZN(n13723) );
  INV_X1 U17149 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20304) );
  OAI222_X1 U17150 ( .A1(n13723), .A2(n14930), .B1(n20355), .B2(n20304), .C1(
        n16803), .C2(n14932), .ZN(P1_U2867) );
  NOR3_X1 U17151 ( .A1(n20103), .A2(n16664), .A3(n11619), .ZN(n13725) );
  NOR2_X1 U17152 ( .A1(n13725), .A2(n13724), .ZN(n13729) );
  INV_X1 U17153 ( .A(n13726), .ZN(n13727) );
  OAI211_X1 U17154 ( .C1(n13730), .C2(n13727), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n20103), .ZN(n13728) );
  OAI211_X1 U17155 ( .C1(n13730), .C2(n13729), .A(n13728), .B(n19364), .ZN(
        P2_U3177) );
  XOR2_X1 U17156 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13754), .Z(n13736)
         );
  AND2_X1 U17157 ( .A1(n13732), .A2(n13731), .ZN(n13733) );
  OR2_X1 U17158 ( .A1(n13733), .A2(n13751), .ZN(n16566) );
  MUX2_X1 U17159 ( .A(n16566), .B(n13734), .S(n9733), .Z(n13735) );
  OAI21_X1 U17160 ( .B1(n13736), .B2(n15897), .A(n13735), .ZN(P2_U2880) );
  OR2_X1 U17161 ( .A1(n13620), .A2(n13738), .ZN(n13739) );
  NAND2_X1 U17162 ( .A1(n13737), .A2(n13739), .ZN(n16457) );
  OAI222_X1 U17163 ( .A1(n16457), .A2(n16015), .B1(n16017), .B2(n13119), .C1(
        n13740), .C2(n19403), .ZN(P2_U2904) );
  AOI21_X1 U17164 ( .B1(n13741), .B2(n9865), .A(n13787), .ZN(n16509) );
  NAND2_X1 U17165 ( .A1(n16509), .A2(n15887), .ZN(n13747) );
  INV_X1 U17166 ( .A(n13742), .ZN(n13745) );
  OAI211_X1 U17167 ( .C1(n13745), .C2(n13744), .A(n15904), .B(n13789), .ZN(
        n13746) );
  OAI211_X1 U17168 ( .C1(n15887), .C2(n13748), .A(n13747), .B(n13746), .ZN(
        P2_U2876) );
  OR2_X1 U17169 ( .A1(n13751), .A2(n13750), .ZN(n13752) );
  NAND2_X1 U17170 ( .A1(n13749), .A2(n13752), .ZN(n16551) );
  INV_X1 U17171 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13753) );
  NOR2_X1 U17172 ( .A1(n13754), .A2(n13753), .ZN(n13756) );
  NAND2_X1 U17173 ( .A1(n13756), .A2(n13755), .ZN(n13781) );
  OAI211_X1 U17174 ( .C1(n13756), .C2(n13755), .A(n13781), .B(n15904), .ZN(
        n13758) );
  NAND2_X1 U17175 ( .A1(n9733), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13757) );
  OAI211_X1 U17176 ( .C1(n16551), .C2(n9733), .A(n13758), .B(n13757), .ZN(
        P2_U2879) );
  INV_X1 U17177 ( .A(n13759), .ZN(n13780) );
  XNOR2_X1 U17178 ( .A(n13781), .B(n13780), .ZN(n13764) );
  INV_X1 U17179 ( .A(n13760), .ZN(n13778) );
  NAND2_X1 U17180 ( .A1(n13749), .A2(n13761), .ZN(n13762) );
  NAND2_X1 U17181 ( .A1(n13778), .A2(n13762), .ZN(n16531) );
  MUX2_X1 U17182 ( .A(n11092), .B(n16531), .S(n15887), .Z(n13763) );
  OAI21_X1 U17183 ( .B1(n13764), .B2(n15897), .A(n13763), .ZN(P2_U2878) );
  INV_X1 U17184 ( .A(n16769), .ZN(n20232) );
  OAI22_X1 U17185 ( .A1(n16771), .A2(n20232), .B1(n20238), .B2(n13766), .ZN(
        n13768) );
  MUX2_X1 U17186 ( .A(n13768), .B(n13767), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n13774) );
  INV_X1 U17187 ( .A(n13769), .ZN(n13770) );
  AOI211_X1 U17188 ( .C1(n20216), .C2(n13772), .A(n13771), .B(n13770), .ZN(
        n13773) );
  OAI211_X1 U17189 ( .C1(n13776), .C2(n13775), .A(n13774), .B(n13773), .ZN(
        P2_U3176) );
  NAND2_X1 U17190 ( .A1(n13778), .A2(n13777), .ZN(n13779) );
  NAND2_X1 U17191 ( .A1(n9865), .A2(n13779), .ZN(n16524) );
  NOR2_X1 U17192 ( .A1(n13781), .A2(n13780), .ZN(n13783) );
  OAI211_X1 U17193 ( .C1(n13783), .C2(n13782), .A(n15904), .B(n13742), .ZN(
        n13785) );
  NAND2_X1 U17194 ( .A1(n9733), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13784) );
  OAI211_X1 U17195 ( .C1(n16524), .C2(n9733), .A(n13785), .B(n13784), .ZN(
        P2_U2877) );
  OR2_X1 U17196 ( .A1(n13787), .A2(n13786), .ZN(n13788) );
  AND2_X1 U17197 ( .A1(n13799), .A2(n13788), .ZN(n16500) );
  INV_X1 U17198 ( .A(n16500), .ZN(n13796) );
  INV_X1 U17199 ( .A(n13789), .ZN(n13793) );
  INV_X1 U17200 ( .A(n13790), .ZN(n13791) );
  OAI211_X1 U17201 ( .C1(n13793), .C2(n13792), .A(n13791), .B(n15904), .ZN(
        n13795) );
  NAND2_X1 U17202 ( .A1(n9733), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13794) );
  OAI211_X1 U17203 ( .C1(n13796), .C2(n15824), .A(n13795), .B(n13794), .ZN(
        P2_U2875) );
  INV_X1 U17204 ( .A(n13797), .ZN(n13807) );
  NAND2_X1 U17205 ( .A1(n13799), .A2(n13798), .ZN(n13800) );
  NAND2_X1 U17206 ( .A1(n13807), .A2(n13800), .ZN(n16485) );
  OAI211_X1 U17207 ( .C1(n13790), .C2(n13803), .A(n13802), .B(n15904), .ZN(
        n13805) );
  NAND2_X1 U17208 ( .A1(n9733), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13804) );
  OAI211_X1 U17209 ( .C1(n16485), .C2(n9733), .A(n13805), .B(n13804), .ZN(
        P2_U2874) );
  AND2_X1 U17210 ( .A1(n13807), .A2(n13806), .ZN(n13809) );
  OR2_X1 U17211 ( .A1(n13809), .A2(n13808), .ZN(n16470) );
  OAI211_X1 U17212 ( .C1(n13801), .C2(n12179), .A(n15904), .B(n13811), .ZN(
        n13813) );
  NAND2_X1 U17213 ( .A1(n9733), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13812) );
  OAI211_X1 U17214 ( .C1(n16470), .C2(n9733), .A(n13813), .B(n13812), .ZN(
        P2_U2873) );
  NAND3_X1 U17215 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19210)
         );
  NAND2_X1 U17216 ( .A1(n16698), .A2(n17317), .ZN(n13814) );
  NOR2_X1 U17217 ( .A1(n17602), .A2(n13814), .ZN(n18603) );
  INV_X1 U17218 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17006) );
  OAI221_X1 U17219 ( .B1(n19210), .B2(n18603), .C1(n19210), .C2(n17006), .A(
        n18690), .ZN(n18610) );
  INV_X1 U17220 ( .A(n18610), .ZN(n18606) );
  INV_X1 U17221 ( .A(n18251), .ZN(n18124) );
  NOR2_X1 U17222 ( .A1(n19257), .A2(n18124), .ZN(n16684) );
  AOI21_X1 U17223 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n16684), .ZN(n16685) );
  NOR2_X1 U17224 ( .A1(n18606), .A2(n16685), .ZN(n13816) );
  NAND2_X1 U17225 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19066), .ZN(n18649) );
  NAND2_X1 U17226 ( .A1(n18649), .A2(n18610), .ZN(n16683) );
  OR2_X1 U17227 ( .A1(n18964), .A2(n16683), .ZN(n13815) );
  MUX2_X1 U17228 ( .A(n13816), .B(n13815), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  XOR2_X1 U17229 ( .A(n17403), .B(n17681), .Z(n17676) );
  INV_X1 U17230 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n13818) );
  INV_X1 U17231 ( .A(n17412), .ZN(n17415) );
  NAND3_X1 U17232 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n13818), .A3(n17415), 
        .ZN(n13819) );
  AOI22_X1 U17233 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13823) );
  AOI22_X1 U17234 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13822) );
  AOI22_X1 U17235 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13821) );
  AOI22_X1 U17236 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13820) );
  NAND4_X1 U17237 ( .A1(n13823), .A2(n13822), .A3(n13821), .A4(n13820), .ZN(
        n13829) );
  AOI22_X1 U17238 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U17239 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13826) );
  AOI22_X1 U17240 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13825) );
  AOI22_X1 U17241 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13824) );
  NAND4_X1 U17242 ( .A1(n13827), .A2(n13826), .A3(n13825), .A4(n13824), .ZN(
        n13828) );
  OR2_X1 U17243 ( .A1(n13829), .A2(n13828), .ZN(n14378) );
  NAND2_X1 U17244 ( .A1(n13833), .A2(n14378), .ZN(n13832) );
  NAND2_X1 U17245 ( .A1(n13830), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13831) );
  INV_X1 U17246 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13836) );
  NAND2_X1 U17247 ( .A1(n13833), .A2(n14380), .ZN(n13834) );
  OAI21_X1 U17248 ( .B1(n13836), .B2(n13835), .A(n13834), .ZN(n13837) );
  NAND2_X1 U17249 ( .A1(n14375), .A2(n13984), .ZN(n13844) );
  INV_X1 U17250 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13841) );
  OAI21_X1 U17251 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13839), .A(
        n13885), .ZN(n20290) );
  NAND2_X1 U17252 ( .A1(n20290), .A2(n14502), .ZN(n13840) );
  OAI21_X1 U17253 ( .B1(n13841), .B2(n13899), .A(n13840), .ZN(n13842) );
  AOI21_X1 U17254 ( .B1(n14504), .B2(P1_EAX_REG_7__SCAN_IN), .A(n13842), .ZN(
        n13843) );
  NAND2_X1 U17255 ( .A1(n13844), .A2(n13843), .ZN(n14839) );
  INV_X1 U17256 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n15002) );
  AOI22_X1 U17257 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13848) );
  AOI22_X1 U17258 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13847) );
  AOI22_X1 U17259 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17260 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13845) );
  NAND4_X1 U17261 ( .A1(n13848), .A2(n13847), .A3(n13846), .A4(n13845), .ZN(
        n13854) );
  AOI22_X1 U17262 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14473), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13852) );
  AOI22_X1 U17263 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14476), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13851) );
  AOI22_X1 U17264 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U17265 ( .A1(n14487), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13849) );
  NAND4_X1 U17266 ( .A1(n13852), .A2(n13851), .A3(n13850), .A4(n13849), .ZN(
        n13853) );
  OAI21_X1 U17267 ( .B1(n13854), .B2(n13853), .A(n13984), .ZN(n13857) );
  INV_X1 U17268 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13855) );
  XNOR2_X1 U17269 ( .A(n13885), .B(n13855), .ZN(n15223) );
  AOI22_X1 U17270 ( .A1(n15223), .A2(n14502), .B1(n14503), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13856) );
  OAI211_X1 U17271 ( .C1(n9862), .C2(n15002), .A(n13857), .B(n13856), .ZN(
        n14840) );
  AOI22_X1 U17272 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13861) );
  AOI22_X1 U17273 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13860) );
  AOI22_X1 U17274 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13859) );
  AOI22_X1 U17275 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13858) );
  NAND4_X1 U17276 ( .A1(n13861), .A2(n13860), .A3(n13859), .A4(n13858), .ZN(
        n13867) );
  AOI22_X1 U17277 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U17278 ( .A1(n14228), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13864) );
  AOI22_X1 U17279 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13863) );
  AOI22_X1 U17280 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13862) );
  NAND4_X1 U17281 ( .A1(n13865), .A2(n13864), .A3(n13863), .A4(n13862), .ZN(
        n13866) );
  NOR2_X1 U17282 ( .A1(n13867), .A2(n13866), .ZN(n13873) );
  NAND2_X1 U17283 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13868) );
  INV_X1 U17284 ( .A(n13869), .ZN(n13887) );
  INV_X1 U17285 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21477) );
  NAND2_X1 U17286 ( .A1(n13887), .A2(n21477), .ZN(n13870) );
  NAND2_X1 U17287 ( .A1(n13968), .A2(n13870), .ZN(n16784) );
  AOI22_X1 U17288 ( .A1(n16784), .A2(n14502), .B1(n14503), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13872) );
  NAND2_X1 U17289 ( .A1(n14504), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13871) );
  OAI211_X1 U17290 ( .C1(n13874), .C2(n13873), .A(n13872), .B(n13871), .ZN(
        n14910) );
  AND2_X1 U17291 ( .A1(n14840), .A2(n14910), .ZN(n13890) );
  INV_X1 U17292 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15001) );
  AOI22_X1 U17293 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U17294 ( .A1(n14228), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U17295 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U17296 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13875) );
  NAND4_X1 U17297 ( .A1(n13878), .A2(n13877), .A3(n13876), .A4(n13875), .ZN(
        n13884) );
  AOI22_X1 U17298 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14171), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U17299 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13881) );
  AOI22_X1 U17300 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U17301 ( .A1(n12775), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13879) );
  NAND4_X1 U17302 ( .A1(n13882), .A2(n13881), .A3(n13880), .A4(n13879), .ZN(
        n13883) );
  OAI21_X1 U17303 ( .B1(n13884), .B2(n13883), .A(n13984), .ZN(n13889) );
  INV_X1 U17304 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21256) );
  OAI21_X1 U17305 ( .B1(n13885), .B2(n13855), .A(n21256), .ZN(n13886) );
  NAND2_X1 U17306 ( .A1(n13887), .A2(n13886), .ZN(n20274) );
  AOI22_X1 U17307 ( .A1(n20274), .A2(n14502), .B1(n14503), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13888) );
  OAI211_X1 U17308 ( .C1(n9862), .C2(n15001), .A(n13889), .B(n13888), .ZN(
        n14915) );
  INV_X1 U17309 ( .A(n13893), .ZN(n13894) );
  INV_X1 U17310 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13900) );
  OAI21_X1 U17311 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13897), .A(
        n13896), .ZN(n20301) );
  NAND2_X1 U17312 ( .A1(n20301), .A2(n14502), .ZN(n13898) );
  OAI21_X1 U17313 ( .B1(n13900), .B2(n13899), .A(n13898), .ZN(n13901) );
  AOI21_X1 U17314 ( .B1(n14504), .B2(P1_EAX_REG_6__SCAN_IN), .A(n13901), .ZN(
        n13902) );
  AOI22_X1 U17315 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14476), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17316 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U17317 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U17318 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n14230), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13906) );
  NAND4_X1 U17319 ( .A1(n13909), .A2(n13908), .A3(n13907), .A4(n13906), .ZN(
        n13915) );
  AOI22_X1 U17320 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14171), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17321 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U17322 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U17323 ( .A1(n12775), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13910) );
  NAND4_X1 U17324 ( .A1(n13913), .A2(n13912), .A3(n13911), .A4(n13910), .ZN(
        n13914) );
  OAI21_X1 U17325 ( .B1(n13915), .B2(n13914), .A(n13984), .ZN(n13920) );
  NAND2_X1 U17326 ( .A1(n14504), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n13919) );
  INV_X1 U17327 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13967) );
  INV_X1 U17328 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13916) );
  XNOR2_X1 U17329 ( .A(n13970), .B(n13916), .ZN(n15184) );
  NAND2_X1 U17330 ( .A1(n15184), .A2(n14502), .ZN(n13918) );
  NAND2_X1 U17331 ( .A1(n14503), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13917) );
  NAND4_X1 U17332 ( .A1(n13920), .A2(n13919), .A3(n13918), .A4(n13917), .ZN(
        n14814) );
  AOI22_X1 U17333 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13924) );
  AOI22_X1 U17334 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13923) );
  AOI22_X1 U17335 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13922) );
  AOI22_X1 U17336 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13921) );
  NAND4_X1 U17337 ( .A1(n13924), .A2(n13923), .A3(n13922), .A4(n13921), .ZN(
        n13930) );
  AOI22_X1 U17338 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14171), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U17339 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U17340 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U17341 ( .A1(n14472), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13925) );
  NAND4_X1 U17342 ( .A1(n13928), .A2(n13927), .A3(n13926), .A4(n13925), .ZN(
        n13929) );
  OAI21_X1 U17343 ( .B1(n13930), .B2(n13929), .A(n13984), .ZN(n13936) );
  NAND2_X1 U17344 ( .A1(n14504), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13935) );
  INV_X1 U17345 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13932) );
  XNOR2_X1 U17346 ( .A(n13948), .B(n13932), .ZN(n15177) );
  NAND2_X1 U17347 ( .A1(n15177), .A2(n14502), .ZN(n13934) );
  NAND2_X1 U17348 ( .A1(n14503), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13933) );
  NAND4_X1 U17349 ( .A1(n13936), .A2(n13935), .A3(n13934), .A4(n13933), .ZN(
        n14802) );
  AND2_X1 U17350 ( .A1(n14814), .A2(n14802), .ZN(n14766) );
  AOI22_X1 U17351 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U17352 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17353 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13938) );
  AOI22_X1 U17354 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13937) );
  NAND4_X1 U17355 ( .A1(n13940), .A2(n13939), .A3(n13938), .A4(n13937), .ZN(
        n13946) );
  AOI22_X1 U17356 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U17357 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13943) );
  AOI22_X1 U17358 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13942) );
  AOI22_X1 U17359 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13941) );
  NAND4_X1 U17360 ( .A1(n13944), .A2(n13943), .A3(n13942), .A4(n13941), .ZN(
        n13945) );
  OR2_X1 U17361 ( .A1(n13946), .A2(n13945), .ZN(n13947) );
  AOI22_X1 U17362 ( .A1(n13984), .A2(n13947), .B1(n14503), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13951) );
  INV_X1 U17363 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14792) );
  OR2_X2 U17364 ( .A1(n13962), .A2(n14792), .ZN(n14001) );
  INV_X1 U17365 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14775) );
  XNOR2_X1 U17366 ( .A(n14001), .B(n14775), .ZN(n15155) );
  NAND2_X1 U17367 ( .A1(n15155), .A2(n14502), .ZN(n13950) );
  OAI211_X1 U17368 ( .C1(n9862), .C2(n21259), .A(n13951), .B(n13950), .ZN(
        n14769) );
  AOI22_X1 U17369 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U17370 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U17371 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U17372 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13952) );
  NAND4_X1 U17373 ( .A1(n13955), .A2(n13954), .A3(n13953), .A4(n13952), .ZN(
        n13961) );
  AOI22_X1 U17374 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14476), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13959) );
  AOI22_X1 U17375 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13958) );
  AOI22_X1 U17376 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U17377 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13956) );
  NAND4_X1 U17378 ( .A1(n13959), .A2(n13958), .A3(n13957), .A4(n13956), .ZN(
        n13960) );
  OAI21_X1 U17379 ( .B1(n13961), .B2(n13960), .A(n13984), .ZN(n13966) );
  NAND2_X1 U17380 ( .A1(n14504), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13965) );
  XNOR2_X1 U17381 ( .A(n13962), .B(n14792), .ZN(n15166) );
  NAND2_X1 U17382 ( .A1(n15166), .A2(n14502), .ZN(n13964) );
  NAND2_X1 U17383 ( .A1(n14503), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13963) );
  NAND4_X1 U17384 ( .A1(n13966), .A2(n13965), .A3(n13964), .A4(n13963), .ZN(
        n14781) );
  NAND2_X1 U17385 ( .A1(n14504), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n13972) );
  NAND2_X1 U17386 ( .A1(n13968), .A2(n13967), .ZN(n13969) );
  NAND2_X1 U17387 ( .A1(n13970), .A2(n13969), .ZN(n15193) );
  AOI22_X1 U17388 ( .A1(n15193), .A2(n14502), .B1(n14503), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13971) );
  NAND2_X1 U17389 ( .A1(n13972), .A2(n13971), .ZN(n14799) );
  AOI22_X1 U17390 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13976) );
  AOI22_X1 U17391 ( .A1(n14450), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U17392 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17393 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13973) );
  NAND4_X1 U17394 ( .A1(n13976), .A2(n13975), .A3(n13974), .A4(n13973), .ZN(
        n13982) );
  AOI22_X1 U17395 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13980) );
  AOI22_X1 U17396 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13979) );
  AOI22_X1 U17397 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13978) );
  AOI22_X1 U17398 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13977) );
  NAND4_X1 U17399 ( .A1(n13980), .A2(n13979), .A3(n13978), .A4(n13977), .ZN(
        n13981) );
  OR2_X1 U17400 ( .A1(n13982), .A2(n13981), .ZN(n13983) );
  AND2_X1 U17401 ( .A1(n13984), .A2(n13983), .ZN(n14829) );
  OR2_X1 U17402 ( .A1(n14799), .A2(n14829), .ZN(n13985) );
  NAND2_X1 U17403 ( .A1(n13986), .A2(n9874), .ZN(n14750) );
  AOI22_X1 U17404 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14229), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U17405 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13989) );
  AOI22_X1 U17406 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13988) );
  AOI22_X1 U17407 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13987) );
  NAND4_X1 U17408 ( .A1(n13990), .A2(n13989), .A3(n13988), .A4(n13987), .ZN(
        n13998) );
  AOI22_X1 U17409 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13996) );
  AOI21_X1 U17410 ( .B1(n14450), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n14502), .ZN(n13992) );
  NAND2_X1 U17411 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13991) );
  AND2_X1 U17412 ( .A1(n13992), .A2(n13991), .ZN(n13995) );
  AOI22_X1 U17413 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13994) );
  AOI22_X1 U17414 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13993) );
  NAND4_X1 U17415 ( .A1(n13996), .A2(n13995), .A3(n13994), .A4(n13993), .ZN(
        n13997) );
  NAND2_X1 U17416 ( .A1(n14465), .A2(n14468), .ZN(n14107) );
  OAI21_X1 U17417 ( .B1(n13998), .B2(n13997), .A(n14107), .ZN(n14000) );
  AOI22_X1 U17418 ( .A1(n14504), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13022), .ZN(n13999) );
  NAND2_X1 U17419 ( .A1(n14000), .A2(n13999), .ZN(n14003) );
  OR2_X2 U17420 ( .A1(n14001), .A2(n14775), .ZN(n14014) );
  XNOR2_X1 U17421 ( .A(n14014), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15140) );
  NAND2_X1 U17422 ( .A1(n15140), .A2(n14328), .ZN(n14002) );
  NAND2_X1 U17423 ( .A1(n14003), .A2(n14002), .ZN(n14751) );
  AOI22_X1 U17424 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14171), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14007) );
  AOI22_X1 U17425 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14229), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17426 ( .A1(n14450), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14005) );
  AOI22_X1 U17427 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14004) );
  NAND4_X1 U17428 ( .A1(n14007), .A2(n14006), .A3(n14005), .A4(n14004), .ZN(
        n14013) );
  AOI22_X1 U17429 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14011) );
  AOI22_X1 U17430 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14010) );
  AOI22_X1 U17431 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14009) );
  AOI22_X1 U17432 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14008) );
  NAND4_X1 U17433 ( .A1(n14011), .A2(n14010), .A3(n14009), .A4(n14008), .ZN(
        n14012) );
  NOR2_X1 U17434 ( .A1(n14013), .A2(n14012), .ZN(n14019) );
  INV_X1 U17435 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14016) );
  XNOR2_X1 U17436 ( .A(n14020), .B(n14016), .ZN(n15131) );
  NAND2_X1 U17437 ( .A1(n15131), .A2(n14328), .ZN(n14018) );
  AOI22_X1 U17438 ( .A1(n14504), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n14503), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14017) );
  OAI211_X1 U17439 ( .C1(n14019), .C2(n14465), .A(n14018), .B(n14017), .ZN(
        n14739) );
  XNOR2_X1 U17440 ( .A(n14039), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15120) );
  NAND2_X1 U17441 ( .A1(n15120), .A2(n14328), .ZN(n14038) );
  AOI22_X1 U17442 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14025) );
  AOI22_X1 U17443 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14024) );
  AOI22_X1 U17444 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14023) );
  AOI22_X1 U17445 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14022) );
  NAND4_X1 U17446 ( .A1(n14025), .A2(n14024), .A3(n14023), .A4(n14022), .ZN(
        n14034) );
  NAND2_X1 U17447 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14027) );
  NAND2_X1 U17448 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14026) );
  AND3_X1 U17449 ( .A1(n14027), .A2(n14468), .A3(n14026), .ZN(n14032) );
  AOI22_X1 U17450 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14031) );
  AOI22_X1 U17451 ( .A1(n14472), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U17452 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14029) );
  NAND4_X1 U17453 ( .A1(n14032), .A2(n14031), .A3(n14030), .A4(n14029), .ZN(
        n14033) );
  OAI21_X1 U17454 ( .B1(n14034), .B2(n14033), .A(n14107), .ZN(n14036) );
  AOI22_X1 U17455 ( .A1(n14504), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13022), .ZN(n14035) );
  NAND2_X1 U17456 ( .A1(n14036), .A2(n14035), .ZN(n14037) );
  INV_X1 U17457 ( .A(n14041), .ZN(n14043) );
  INV_X1 U17458 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14042) );
  NAND2_X1 U17459 ( .A1(n14043), .A2(n14042), .ZN(n14044) );
  NAND2_X1 U17460 ( .A1(n14076), .A2(n14044), .ZN(n15112) );
  AOI22_X1 U17461 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14048) );
  AOI22_X1 U17462 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14047) );
  AOI22_X1 U17463 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14046) );
  AOI22_X1 U17464 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14045) );
  NAND4_X1 U17465 ( .A1(n14048), .A2(n14047), .A3(n14046), .A4(n14045), .ZN(
        n14054) );
  AOI22_X1 U17466 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U17467 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U17468 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14050) );
  AOI22_X1 U17469 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14049) );
  NAND4_X1 U17470 ( .A1(n14052), .A2(n14051), .A3(n14050), .A4(n14049), .ZN(
        n14053) );
  NOR2_X1 U17471 ( .A1(n14054), .A2(n14053), .ZN(n14058) );
  NAND2_X1 U17472 ( .A1(n13022), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14055) );
  NAND2_X1 U17473 ( .A1(n14468), .A2(n14055), .ZN(n14056) );
  AOI21_X1 U17474 ( .B1(n14504), .B2(P1_EAX_REG_19__SCAN_IN), .A(n14056), .ZN(
        n14057) );
  OAI21_X1 U17475 ( .B1(n14465), .B2(n14058), .A(n14057), .ZN(n14059) );
  NAND2_X1 U17476 ( .A1(n14060), .A2(n14059), .ZN(n14706) );
  XNOR2_X1 U17477 ( .A(n14076), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15104) );
  AOI22_X1 U17478 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U17479 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14171), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U17480 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14229), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14062) );
  AOI22_X1 U17481 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14061) );
  NAND4_X1 U17482 ( .A1(n14064), .A2(n14063), .A3(n14062), .A4(n14061), .ZN(
        n14070) );
  AOI22_X1 U17483 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U17484 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14067) );
  AOI22_X1 U17485 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14476), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14066) );
  AOI22_X1 U17486 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14065) );
  NAND4_X1 U17487 ( .A1(n14068), .A2(n14067), .A3(n14066), .A4(n14065), .ZN(
        n14069) );
  NOR2_X1 U17488 ( .A1(n14070), .A2(n14069), .ZN(n14073) );
  INV_X1 U17489 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15100) );
  AOI21_X1 U17490 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15100), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14071) );
  AOI21_X1 U17491 ( .B1(n14504), .B2(P1_EAX_REG_20__SCAN_IN), .A(n14071), .ZN(
        n14072) );
  OAI21_X1 U17492 ( .B1(n14465), .B2(n14073), .A(n14072), .ZN(n14074) );
  INV_X1 U17493 ( .A(n14074), .ZN(n14075) );
  AOI21_X1 U17494 ( .B1(n15104), .B2(n14502), .A(n14075), .ZN(n14692) );
  AND2_X2 U17495 ( .A1(n14691), .A2(n14692), .ZN(n14681) );
  INV_X1 U17496 ( .A(n14078), .ZN(n14079) );
  INV_X1 U17497 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15092) );
  NAND2_X1 U17498 ( .A1(n14079), .A2(n15092), .ZN(n14080) );
  AND2_X1 U17499 ( .A1(n14114), .A2(n14080), .ZN(n15094) );
  INV_X1 U17500 ( .A(n14465), .ZN(n14499) );
  AOI22_X1 U17501 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U17502 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14171), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17503 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17504 ( .A1(n14228), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14081) );
  NAND4_X1 U17505 ( .A1(n14084), .A2(n14083), .A3(n14082), .A4(n14081), .ZN(
        n14090) );
  AOI22_X1 U17506 ( .A1(n14472), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14229), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14088) );
  AOI22_X1 U17507 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14087) );
  AOI22_X1 U17508 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U17509 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14085) );
  NAND4_X1 U17510 ( .A1(n14088), .A2(n14087), .A3(n14086), .A4(n14085), .ZN(
        n14089) );
  OR2_X1 U17511 ( .A1(n14090), .A2(n14089), .ZN(n14093) );
  NAND2_X1 U17512 ( .A1(n13022), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14091) );
  OAI211_X1 U17513 ( .C1(n9862), .C2(n13366), .A(n14468), .B(n14091), .ZN(
        n14092) );
  AOI21_X1 U17514 ( .B1(n14499), .B2(n14093), .A(n14092), .ZN(n14094) );
  AOI21_X1 U17515 ( .B1(n15094), .B2(n14502), .A(n14094), .ZN(n14682) );
  XNOR2_X1 U17516 ( .A(n14114), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15081) );
  NAND2_X1 U17517 ( .A1(n15081), .A2(n14328), .ZN(n14113) );
  AOI22_X1 U17518 ( .A1(n13515), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U17519 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14476), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14097) );
  AOI22_X1 U17520 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U17521 ( .A1(n14450), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14095) );
  NAND4_X1 U17522 ( .A1(n14098), .A2(n14097), .A3(n14096), .A4(n14095), .ZN(
        n14109) );
  NAND2_X1 U17523 ( .A1(n14099), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14101) );
  NAND2_X1 U17524 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14100) );
  AND3_X1 U17525 ( .A1(n14101), .A2(n14100), .A3(n14468), .ZN(n14106) );
  AOI22_X1 U17526 ( .A1(n14102), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14105) );
  AOI22_X1 U17527 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12768), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17528 ( .A1(n14472), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14103) );
  NAND4_X1 U17529 ( .A1(n14106), .A2(n14105), .A3(n14104), .A4(n14103), .ZN(
        n14108) );
  OAI21_X1 U17530 ( .B1(n14109), .B2(n14108), .A(n14107), .ZN(n14111) );
  AOI22_X1 U17531 ( .A1(n14504), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13022), .ZN(n14110) );
  NAND2_X1 U17532 ( .A1(n14111), .A2(n14110), .ZN(n14112) );
  NAND2_X1 U17533 ( .A1(n14113), .A2(n14112), .ZN(n14666) );
  INV_X1 U17534 ( .A(n14116), .ZN(n14117) );
  INV_X1 U17535 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14140) );
  NAND2_X1 U17536 ( .A1(n14117), .A2(n14140), .ZN(n14118) );
  NAND2_X1 U17537 ( .A1(n14165), .A2(n14118), .ZN(n15074) );
  AOI22_X1 U17538 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U17539 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17540 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14229), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17541 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14120) );
  NAND4_X1 U17542 ( .A1(n14123), .A2(n14122), .A3(n14121), .A4(n14120), .ZN(
        n14129) );
  AOI22_X1 U17543 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U17544 ( .A1(n14450), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17545 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17546 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14124) );
  NAND4_X1 U17547 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14124), .ZN(
        n14128) );
  NOR2_X1 U17548 ( .A1(n14129), .A2(n14128), .ZN(n14147) );
  AOI22_X1 U17549 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14133) );
  AOI22_X1 U17550 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U17551 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U17552 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14130) );
  NAND4_X1 U17553 ( .A1(n14133), .A2(n14132), .A3(n14131), .A4(n14130), .ZN(
        n14139) );
  AOI22_X1 U17554 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U17555 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14136) );
  AOI22_X1 U17556 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14135) );
  AOI22_X1 U17557 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14134) );
  NAND4_X1 U17558 ( .A1(n14137), .A2(n14136), .A3(n14135), .A4(n14134), .ZN(
        n14138) );
  NOR2_X1 U17559 ( .A1(n14139), .A2(n14138), .ZN(n14146) );
  XNOR2_X1 U17560 ( .A(n14147), .B(n14146), .ZN(n14143) );
  AOI21_X1 U17561 ( .B1(n14140), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14141) );
  AOI21_X1 U17562 ( .B1(n14504), .B2(P1_EAX_REG_23__SCAN_IN), .A(n14141), .ZN(
        n14142) );
  OAI21_X1 U17563 ( .B1(n14143), .B2(n14465), .A(n14142), .ZN(n14144) );
  NAND2_X1 U17564 ( .A1(n14145), .A2(n14144), .ZN(n14654) );
  XNOR2_X1 U17565 ( .A(n14165), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15065) );
  NOR2_X1 U17566 ( .A1(n14147), .A2(n14146), .ZN(n14179) );
  INV_X1 U17567 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n21304) );
  AOI22_X1 U17568 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14151) );
  AOI22_X1 U17569 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14150) );
  AOI22_X1 U17570 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U17571 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14148) );
  NAND4_X1 U17572 ( .A1(n14151), .A2(n14150), .A3(n14149), .A4(n14148), .ZN(
        n14157) );
  AOI22_X1 U17573 ( .A1(n14171), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14155) );
  AOI22_X1 U17574 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U17575 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17576 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14152) );
  NAND4_X1 U17577 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14156) );
  OR2_X1 U17578 ( .A1(n14157), .A2(n14156), .ZN(n14178) );
  INV_X1 U17579 ( .A(n14178), .ZN(n14158) );
  XNOR2_X1 U17580 ( .A(n14179), .B(n14158), .ZN(n14161) );
  NAND2_X1 U17581 ( .A1(n13022), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14159) );
  OAI211_X1 U17582 ( .C1(n9862), .C2(n13041), .A(n14468), .B(n14159), .ZN(
        n14160) );
  AOI21_X1 U17583 ( .B1(n14161), .B2(n14499), .A(n14160), .ZN(n14162) );
  AOI21_X1 U17584 ( .B1(n15065), .B2(n14328), .A(n14162), .ZN(n14643) );
  INV_X1 U17585 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15063) );
  INV_X1 U17586 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14163) );
  OAI21_X1 U17587 ( .B1(n14165), .B2(n15063), .A(n14163), .ZN(n14166) );
  NAND2_X1 U17588 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14164) );
  OR2_X2 U17589 ( .A1(n14165), .A2(n14164), .ZN(n14185) );
  NAND2_X1 U17590 ( .A1(n14166), .A2(n14185), .ZN(n15056) );
  AOI22_X1 U17591 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14476), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U17592 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14169) );
  AOI22_X1 U17593 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U17594 ( .A1(n14472), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14167) );
  NAND4_X1 U17595 ( .A1(n14170), .A2(n14169), .A3(n14168), .A4(n14167), .ZN(
        n14177) );
  AOI22_X1 U17596 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14175) );
  AOI22_X1 U17597 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14171), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14174) );
  AOI22_X1 U17598 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14173) );
  AOI22_X1 U17599 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14172) );
  NAND4_X1 U17600 ( .A1(n14175), .A2(n14174), .A3(n14173), .A4(n14172), .ZN(
        n14176) );
  NOR2_X1 U17601 ( .A1(n14177), .A2(n14176), .ZN(n14188) );
  NAND2_X1 U17602 ( .A1(n14179), .A2(n14178), .ZN(n14187) );
  XNOR2_X1 U17603 ( .A(n14188), .B(n14187), .ZN(n14180) );
  NOR2_X1 U17604 ( .A1(n14180), .A2(n14465), .ZN(n14183) );
  NAND2_X1 U17605 ( .A1(n13022), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14181) );
  OAI211_X1 U17606 ( .C1(n9862), .C2(n13039), .A(n14468), .B(n14181), .ZN(
        n14182) );
  OAI22_X1 U17607 ( .A1(n15056), .A2(n14468), .B1(n14183), .B2(n14182), .ZN(
        n14630) );
  INV_X1 U17608 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n21412) );
  NAND2_X1 U17609 ( .A1(n14185), .A2(n21412), .ZN(n14186) );
  NAND2_X1 U17610 ( .A1(n14206), .A2(n14186), .ZN(n15047) );
  NOR2_X1 U17611 ( .A1(n14188), .A2(n14187), .ZN(n14219) );
  AOI22_X1 U17612 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U17613 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14191) );
  AOI22_X1 U17614 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U17615 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14189) );
  NAND4_X1 U17616 ( .A1(n14192), .A2(n14191), .A3(n14190), .A4(n14189), .ZN(
        n14198) );
  AOI22_X1 U17617 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U17618 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14195) );
  INV_X1 U17619 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n21335) );
  AOI22_X1 U17620 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U17621 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14193) );
  NAND4_X1 U17622 ( .A1(n14196), .A2(n14195), .A3(n14194), .A4(n14193), .ZN(
        n14197) );
  OR2_X1 U17623 ( .A1(n14198), .A2(n14197), .ZN(n14218) );
  XNOR2_X1 U17624 ( .A(n14219), .B(n14218), .ZN(n14201) );
  OAI21_X1 U17625 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21412), .A(n14468), 
        .ZN(n14199) );
  AOI21_X1 U17626 ( .B1(n14504), .B2(P1_EAX_REG_26__SCAN_IN), .A(n14199), .ZN(
        n14200) );
  OAI21_X1 U17627 ( .B1(n14201), .B2(n14465), .A(n14200), .ZN(n14202) );
  NAND2_X1 U17628 ( .A1(n14203), .A2(n14202), .ZN(n14616) );
  INV_X1 U17629 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14205) );
  NAND2_X1 U17631 ( .A1(n14206), .A2(n14205), .ZN(n14207) );
  NAND2_X1 U17632 ( .A1(n14324), .A2(n14207), .ZN(n15038) );
  AOI22_X1 U17633 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n14477), .B1(
        n14230), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14211) );
  AOI22_X1 U17634 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14210) );
  AOI22_X1 U17635 ( .A1(n14229), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14209) );
  AOI22_X1 U17636 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14208) );
  NAND4_X1 U17637 ( .A1(n14211), .A2(n14210), .A3(n14209), .A4(n14208), .ZN(
        n14217) );
  AOI22_X1 U17638 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14171), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14215) );
  AOI22_X1 U17639 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n14475), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14214) );
  AOI22_X1 U17640 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14450), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14213) );
  AOI22_X1 U17641 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14212) );
  NAND4_X1 U17642 ( .A1(n14215), .A2(n14214), .A3(n14213), .A4(n14212), .ZN(
        n14216) );
  NOR2_X1 U17643 ( .A1(n14217), .A2(n14216), .ZN(n14227) );
  NAND2_X1 U17644 ( .A1(n14219), .A2(n14218), .ZN(n14226) );
  XNOR2_X1 U17645 ( .A(n14227), .B(n14226), .ZN(n14223) );
  NAND2_X1 U17646 ( .A1(n13022), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14220) );
  NAND2_X1 U17647 ( .A1(n14468), .A2(n14220), .ZN(n14221) );
  AOI21_X1 U17648 ( .B1(n14504), .B2(P1_EAX_REG_27__SCAN_IN), .A(n14221), .ZN(
        n14222) );
  OAI21_X1 U17649 ( .B1(n14223), .B2(n14465), .A(n14222), .ZN(n14224) );
  NAND2_X1 U17650 ( .A1(n14225), .A2(n14224), .ZN(n14598) );
  XNOR2_X1 U17651 ( .A(n14324), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15031) );
  INV_X1 U17652 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15027) );
  OAI21_X1 U17653 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15027), .A(n14468), 
        .ZN(n14244) );
  NOR2_X1 U17654 ( .A1(n14227), .A2(n14226), .ZN(n14462) );
  AOI22_X1 U17655 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14228), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14234) );
  AOI22_X1 U17656 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14233) );
  AOI22_X1 U17657 ( .A1(n12780), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14229), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14232) );
  AOI22_X1 U17658 ( .A1(n14230), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14231) );
  NAND4_X1 U17659 ( .A1(n14234), .A2(n14233), .A3(n14232), .A4(n14231), .ZN(
        n14241) );
  AOI22_X1 U17660 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U17661 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14238) );
  AOI22_X1 U17662 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U17663 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14236) );
  NAND4_X1 U17664 ( .A1(n14239), .A2(n14238), .A3(n14237), .A4(n14236), .ZN(
        n14240) );
  OR2_X1 U17665 ( .A1(n14241), .A2(n14240), .ZN(n14461) );
  XNOR2_X1 U17666 ( .A(n14462), .B(n14461), .ZN(n14242) );
  NOR2_X1 U17667 ( .A1(n14242), .A2(n14465), .ZN(n14243) );
  AOI211_X1 U17668 ( .C1(n14504), .C2(P1_EAX_REG_28__SCAN_IN), .A(n14244), .B(
        n14243), .ZN(n14245) );
  AOI21_X1 U17669 ( .B1(n14328), .B2(n15031), .A(n14245), .ZN(n14246) );
  OR2_X1 U17670 ( .A1(n14250), .A2(n20485), .ZN(n14556) );
  INV_X1 U17671 ( .A(DATAI_12_), .ZN(n14248) );
  INV_X1 U17672 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14247) );
  MUX2_X1 U17673 ( .A(n14248), .B(n14247), .S(n20488), .Z(n20400) );
  OAI22_X1 U17674 ( .A1(n14986), .A2(n20400), .B1(n15007), .B2(n13045), .ZN(
        n14249) );
  AOI21_X1 U17675 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14988), .A(n14249), .ZN(
        n14252) );
  NOR2_X2 U17676 ( .A1(n14250), .A2(n20488), .ZN(n14989) );
  NAND2_X1 U17677 ( .A1(n14989), .A2(DATAI_28_), .ZN(n14251) );
  OAI211_X1 U17678 ( .C1(n15028), .C2(n15009), .A(n14252), .B(n14251), .ZN(
        P1_U2876) );
  INV_X1 U17679 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14323) );
  INV_X1 U17680 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20354) );
  NAND2_X1 U17681 ( .A1(n14319), .A2(n20354), .ZN(n14255) );
  INV_X1 U17682 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15445) );
  NAND2_X1 U17683 ( .A1(n14409), .A2(n20354), .ZN(n14253) );
  OAI211_X1 U17684 ( .C1(n14318), .C2(n15445), .A(n14253), .B(n14314), .ZN(
        n14254) );
  INV_X1 U17685 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16811) );
  OAI21_X1 U17686 ( .B1(n14318), .B2(n16811), .A(n14314), .ZN(n14257) );
  OAI21_X1 U17687 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n14416), .A(n14257), .ZN(
        n14258) );
  OAI21_X1 U17688 ( .B1(n14317), .B2(P1_EBX_REG_7__SCAN_IN), .A(n14258), .ZN(
        n14929) );
  INV_X1 U17689 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14259) );
  NAND2_X1 U17690 ( .A1(n14319), .A2(n14259), .ZN(n14262) );
  INV_X1 U17691 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15450) );
  NAND2_X1 U17692 ( .A1(n14409), .A2(n14259), .ZN(n14260) );
  OAI211_X1 U17693 ( .C1(n14318), .C2(n15450), .A(n14260), .B(n14314), .ZN(
        n14261) );
  NAND2_X1 U17694 ( .A1(n14262), .A2(n14261), .ZN(n14844) );
  INV_X1 U17695 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U17696 ( .A1(n14413), .A2(n14921), .ZN(n14265) );
  INV_X1 U17697 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15422) );
  OAI21_X1 U17698 ( .B1(n14318), .B2(n15422), .A(n14314), .ZN(n14263) );
  OAI21_X1 U17699 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n14416), .A(n14263), .ZN(
        n14264) );
  MUX2_X1 U17700 ( .A(n14319), .B(n14318), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n14267) );
  NOR2_X1 U17701 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14266) );
  NOR2_X1 U17702 ( .A1(n14267), .A2(n14266), .ZN(n14913) );
  INV_X1 U17703 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14268) );
  NAND2_X1 U17704 ( .A1(n14319), .A2(n14268), .ZN(n14272) );
  INV_X1 U17705 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14270) );
  NAND2_X1 U17706 ( .A1(n14409), .A2(n14268), .ZN(n14269) );
  OAI211_X1 U17707 ( .C1(n14318), .C2(n14270), .A(n14269), .B(n14314), .ZN(
        n14271) );
  NAND2_X1 U17708 ( .A1(n14272), .A2(n14271), .ZN(n14817) );
  INV_X1 U17709 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21449) );
  NAND2_X1 U17710 ( .A1(n14413), .A2(n21449), .ZN(n14275) );
  INV_X1 U17711 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15416) );
  OAI21_X1 U17712 ( .B1(n14318), .B2(n15416), .A(n14314), .ZN(n14273) );
  OAI21_X1 U17713 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(n14416), .A(n14273), .ZN(
        n14274) );
  MUX2_X1 U17714 ( .A(n14319), .B(n14318), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n14279) );
  NOR2_X1 U17715 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14278) );
  NOR2_X1 U17716 ( .A1(n14279), .A2(n14278), .ZN(n14785) );
  INV_X1 U17717 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15344) );
  NAND2_X1 U17718 ( .A1(n14314), .A2(n15344), .ZN(n14280) );
  OAI211_X1 U17719 ( .C1(P1_EBX_REG_13__SCAN_IN), .C2(n14416), .A(n14280), .B(
        n14414), .ZN(n14281) );
  OAI21_X1 U17720 ( .B1(n14317), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14281), .ZN(
        n14805) );
  NAND2_X1 U17721 ( .A1(n14785), .A2(n14805), .ZN(n14282) );
  INV_X1 U17722 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21351) );
  OAI21_X1 U17723 ( .B1(n14318), .B2(n21351), .A(n14314), .ZN(n14283) );
  OAI21_X1 U17724 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(n14416), .A(n14283), .ZN(
        n14284) );
  OAI21_X1 U17725 ( .B1(n14317), .B2(P1_EBX_REG_15__SCAN_IN), .A(n14284), .ZN(
        n14770) );
  MUX2_X1 U17726 ( .A(n13427), .B(n14414), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n14285) );
  OAI21_X1 U17727 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n14418), .A(
        n14285), .ZN(n14754) );
  MUX2_X1 U17728 ( .A(n14319), .B(n14318), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n14287) );
  NOR2_X1 U17729 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14286) );
  NOR2_X1 U17730 ( .A1(n14287), .A2(n14286), .ZN(n14732) );
  INV_X1 U17731 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15355) );
  NAND2_X1 U17732 ( .A1(n14314), .A2(n15355), .ZN(n14288) );
  OAI211_X1 U17733 ( .C1(P1_EBX_REG_17__SCAN_IN), .C2(n14416), .A(n14288), .B(
        n14414), .ZN(n14289) );
  OAI21_X1 U17734 ( .B1(n14317), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14289), .ZN(
        n14740) );
  NAND2_X1 U17735 ( .A1(n14732), .A2(n14740), .ZN(n14290) );
  INV_X1 U17736 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21383) );
  NAND2_X1 U17737 ( .A1(n14319), .A2(n21383), .ZN(n14293) );
  INV_X1 U17738 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15318) );
  NAND2_X1 U17739 ( .A1(n14409), .A2(n21383), .ZN(n14291) );
  OAI211_X1 U17740 ( .C1(n14318), .C2(n15318), .A(n14291), .B(n14314), .ZN(
        n14292) );
  AND2_X1 U17741 ( .A1(n14293), .A2(n14292), .ZN(n14694) );
  INV_X1 U17742 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U17743 ( .A1(n14314), .A2(n15312), .ZN(n14294) );
  OAI211_X1 U17744 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n14416), .A(n14294), .B(
        n14414), .ZN(n14295) );
  OAI21_X1 U17745 ( .B1(n14317), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14295), .ZN(
        n14708) );
  AND2_X1 U17746 ( .A1(n14694), .A2(n14708), .ZN(n14296) );
  MUX2_X1 U17747 ( .A(n13427), .B(n14414), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14298) );
  OR2_X1 U17748 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14297) );
  NAND2_X1 U17749 ( .A1(n14298), .A2(n14297), .ZN(n14678) );
  INV_X1 U17750 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14900) );
  NAND2_X1 U17751 ( .A1(n14413), .A2(n14900), .ZN(n14301) );
  INV_X1 U17752 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U17753 ( .A1(n14314), .A2(n14403), .ZN(n14299) );
  OAI211_X1 U17754 ( .C1(P1_EBX_REG_21__SCAN_IN), .C2(n14416), .A(n14299), .B(
        n14414), .ZN(n14300) );
  AND2_X1 U17755 ( .A1(n14301), .A2(n14300), .ZN(n14683) );
  NOR2_X1 U17756 ( .A1(n14678), .A2(n14683), .ZN(n14302) );
  INV_X1 U17757 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14303) );
  NAND2_X1 U17758 ( .A1(n14413), .A2(n14303), .ZN(n14306) );
  INV_X1 U17759 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21417) );
  NAND2_X1 U17760 ( .A1(n14314), .A2(n21417), .ZN(n14304) );
  OAI211_X1 U17761 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n14416), .A(n14304), .B(
        n14414), .ZN(n14305) );
  AND2_X1 U17762 ( .A1(n14306), .A2(n14305), .ZN(n14658) );
  MUX2_X1 U17763 ( .A(n13427), .B(n14414), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14307) );
  OAI21_X1 U17764 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14418), .A(
        n14307), .ZN(n14647) );
  INV_X1 U17765 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14308) );
  NAND2_X1 U17766 ( .A1(n14413), .A2(n14308), .ZN(n14311) );
  INV_X1 U17767 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U17768 ( .A1(n14314), .A2(n15269), .ZN(n14309) );
  OAI211_X1 U17769 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n14416), .A(n14309), .B(
        n14414), .ZN(n14310) );
  AND2_X1 U17770 ( .A1(n14311), .A2(n14310), .ZN(n14632) );
  MUX2_X1 U17771 ( .A(n14319), .B(n14318), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14313) );
  NOR2_X1 U17772 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14312) );
  NOR2_X1 U17773 ( .A1(n14313), .A2(n14312), .ZN(n14617) );
  INV_X1 U17774 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15035) );
  NAND2_X1 U17775 ( .A1(n14314), .A2(n15035), .ZN(n14315) );
  OAI211_X1 U17776 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n14416), .A(n14315), .B(
        n14414), .ZN(n14316) );
  OAI21_X1 U17777 ( .B1(n14317), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14316), .ZN(
        n14601) );
  MUX2_X1 U17778 ( .A(n14319), .B(n14318), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14321) );
  NOR2_X1 U17779 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14320) );
  NOR2_X1 U17780 ( .A1(n14321), .A2(n14320), .ZN(n14322) );
  OAI21_X1 U17781 ( .B1(n14603), .B2(n14322), .A(n14587), .ZN(n14331) );
  OAI222_X1 U17782 ( .A1(n14932), .A2(n15028), .B1(n14323), .B2(n20355), .C1(
        n14331), .C2(n14930), .ZN(P1_U2844) );
  INV_X1 U17783 ( .A(n14469), .ZN(n14325) );
  NAND2_X1 U17784 ( .A1(n14325), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14326) );
  INV_X1 U17785 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14562) );
  NAND2_X1 U17786 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16753), .ZN(n16756) );
  NAND2_X1 U17787 ( .A1(n14328), .A2(n14327), .ZN(n14329) );
  OAI211_X1 U17788 ( .C1(n16756), .C2(n21091), .A(n20457), .B(n14329), .ZN(
        n14330) );
  NAND2_X1 U17789 ( .A1(n14872), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14334) );
  INV_X1 U17790 ( .A(n14331), .ZN(n15248) );
  AND2_X1 U17791 ( .A1(n12888), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14332) );
  NAND2_X1 U17792 ( .A1(n20506), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14346) );
  AND2_X1 U17793 ( .A1(n21102), .A2(n20832), .ZN(n16751) );
  NOR2_X1 U17794 ( .A1(n14346), .A2(n16751), .ZN(n14333) );
  AND2_X2 U17795 ( .A1(n14350), .A2(n14333), .ZN(n20333) );
  INV_X1 U17796 ( .A(n14334), .ZN(n14335) );
  INV_X1 U17797 ( .A(n15031), .ZN(n14353) );
  NOR2_X1 U17798 ( .A1(n14336), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14348) );
  AND2_X1 U17799 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14756) );
  NAND3_X1 U17800 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14789) );
  INV_X1 U17801 ( .A(n14789), .ZN(n14337) );
  AND2_X1 U17802 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n14337), .ZN(n14755) );
  AND3_X1 U17803 ( .A1(n14756), .A2(n14755), .A3(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n14716) );
  NAND4_X1 U17804 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14709)
         );
  NAND2_X1 U17805 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14713) );
  INV_X1 U17806 ( .A(n14713), .ZN(n14698) );
  NAND4_X1 U17807 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14698), .A3(
        P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n14338) );
  NAND4_X1 U17808 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14711)
         );
  NOR3_X1 U17809 ( .A1(n14709), .A2(n14338), .A3(n14711), .ZN(n14339) );
  AND2_X1 U17810 ( .A1(n14716), .A2(n14339), .ZN(n14667) );
  AND3_X1 U17811 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n14340) );
  NAND2_X1 U17812 ( .A1(n14667), .A2(n14340), .ZN(n14342) );
  INV_X1 U17813 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21148) );
  NOR2_X1 U17814 ( .A1(n14342), .A2(n21148), .ZN(n14341) );
  AND2_X1 U17815 ( .A1(n20337), .A2(n14341), .ZN(n14634) );
  NAND2_X1 U17816 ( .A1(n14634), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14608) );
  INV_X1 U17817 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21155) );
  INV_X1 U17818 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21152) );
  NOR3_X1 U17819 ( .A1(n14608), .A2(n21155), .A3(n21152), .ZN(n14563) );
  NAND2_X1 U17820 ( .A1(n20322), .A2(n14872), .ZN(n14714) );
  INV_X1 U17821 ( .A(n14342), .ZN(n14644) );
  NAND2_X1 U17822 ( .A1(n14872), .A2(n14644), .ZN(n14633) );
  NAND3_X1 U17823 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_26__SCAN_IN), .ZN(n14343) );
  NOR2_X1 U17824 ( .A1(n14633), .A2(n14343), .ZN(n14606) );
  NAND3_X1 U17825 ( .A1(n14606), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14344) );
  NAND2_X1 U17826 ( .A1(n14714), .A2(n14344), .ZN(n14590) );
  INV_X1 U17827 ( .A(n14590), .ZN(n14345) );
  OAI21_X1 U17828 ( .B1(n14563), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14345), 
        .ZN(n14352) );
  INV_X1 U17829 ( .A(n14346), .ZN(n14347) );
  NOR2_X1 U17830 ( .A1(n14348), .A2(n14347), .ZN(n14349) );
  NAND2_X1 U17831 ( .A1(n14350), .A2(n14349), .ZN(n20305) );
  AND2_X2 U17832 ( .A1(n14872), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20335) );
  AOI22_X1 U17833 ( .A1(n20334), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20335), .ZN(n14351) );
  OAI211_X1 U17834 ( .C1(n20330), .C2(n14353), .A(n14352), .B(n14351), .ZN(
        n14354) );
  AOI21_X1 U17835 ( .B1(n15248), .B2(n20333), .A(n14354), .ZN(n14355) );
  OAI21_X1 U17836 ( .B1(n15028), .B2(n14856), .A(n14355), .ZN(P1_U2812) );
  NOR2_X1 U17837 ( .A1(n14357), .A2(n14356), .ZN(n14358) );
  NAND2_X1 U17838 ( .A1(n14392), .A2(n14270), .ZN(n15173) );
  NAND2_X1 U17839 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14359) );
  INV_X1 U17840 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15377) );
  NAND3_X1 U17841 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14360) );
  NAND2_X1 U17842 ( .A1(n10120), .A2(n14360), .ZN(n14361) );
  NAND2_X1 U17843 ( .A1(n14362), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14363) );
  NAND3_X1 U17844 ( .A1(n14366), .A2(n14376), .A3(n14365), .ZN(n14372) );
  INV_X1 U17845 ( .A(n14367), .ZN(n14369) );
  NAND2_X1 U17846 ( .A1(n14369), .A2(n14368), .ZN(n14377) );
  XNOR2_X1 U17847 ( .A(n14377), .B(n14378), .ZN(n14370) );
  NAND2_X1 U17848 ( .A1(n14370), .A2(n14381), .ZN(n14371) );
  NAND2_X1 U17849 ( .A1(n14372), .A2(n14371), .ZN(n16797) );
  OR2_X1 U17850 ( .A1(n16797), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14373) );
  NAND2_X1 U17851 ( .A1(n16797), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14374) );
  NAND2_X1 U17852 ( .A1(n14375), .A2(n14376), .ZN(n14384) );
  INV_X1 U17853 ( .A(n14377), .ZN(n14379) );
  NAND2_X1 U17854 ( .A1(n14379), .A2(n14378), .ZN(n14389) );
  XNOR2_X1 U17855 ( .A(n14389), .B(n14380), .ZN(n14382) );
  NAND2_X1 U17856 ( .A1(n14382), .A2(n14381), .ZN(n14383) );
  NAND2_X1 U17857 ( .A1(n14384), .A2(n14383), .ZN(n14386) );
  OR3_X1 U17858 ( .A1(n14389), .A2(n14388), .A3(n14387), .ZN(n14390) );
  NAND2_X1 U17859 ( .A1(n14392), .A2(n14390), .ZN(n15219) );
  OR2_X1 U17860 ( .A1(n15219), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14391) );
  NAND2_X1 U17861 ( .A1(n15219), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15208) );
  NOR2_X1 U17862 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14396) );
  NAND2_X1 U17863 ( .A1(n14392), .A2(n15355), .ZN(n14398) );
  NOR2_X1 U17864 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14399) );
  INV_X1 U17865 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15198) );
  NAND2_X1 U17866 ( .A1(n15198), .A2(n15416), .ZN(n15170) );
  NAND2_X1 U17867 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U17868 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14401) );
  NOR2_X1 U17869 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14402) );
  AND2_X1 U17870 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14434) );
  NAND2_X1 U17871 ( .A1(n14434), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15259) );
  INV_X1 U17872 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15277) );
  NAND3_X1 U17873 ( .A1(n21417), .A2(n15269), .A3(n15277), .ZN(n15024) );
  NOR2_X1 U17874 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14405) );
  AND2_X1 U17875 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14422) );
  INV_X1 U17876 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15227) );
  MUX2_X1 U17877 ( .A(n14406), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .S(
        n15210), .Z(n14407) );
  XNOR2_X1 U17878 ( .A(n14408), .B(n12971), .ZN(n14513) );
  OR2_X1 U17879 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14411) );
  INV_X1 U17880 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14412) );
  NAND2_X1 U17881 ( .A1(n14409), .A2(n14412), .ZN(n14410) );
  AND2_X1 U17882 ( .A1(n14411), .A2(n14410), .ZN(n14571) );
  AOI22_X1 U17883 ( .A1(n14571), .A2(n14414), .B1(n14413), .B2(n14412), .ZN(
        n14588) );
  AND2_X1 U17884 ( .A1(n14416), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14415) );
  AOI21_X1 U17885 ( .B1(n14418), .B2(P1_EBX_REG_31__SCAN_IN), .A(n14415), .ZN(
        n14419) );
  AND2_X1 U17886 ( .A1(n14416), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14417) );
  AOI21_X1 U17887 ( .B1(n14418), .B2(P1_EBX_REG_30__SCAN_IN), .A(n14417), .ZN(
        n14573) );
  XNOR2_X1 U17888 ( .A(n14419), .B(n14573), .ZN(n14420) );
  MUX2_X1 U17889 ( .A(n14420), .B(n14419), .S(n10452), .Z(n14421) );
  INV_X1 U17890 ( .A(n20475), .ZN(n15345) );
  INV_X1 U17891 ( .A(n14422), .ZN(n14442) );
  NAND2_X1 U17892 ( .A1(n15345), .A2(n20459), .ZN(n14437) );
  NAND2_X1 U17893 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14424) );
  AND2_X1 U17894 ( .A1(n20475), .A2(n14424), .ZN(n14433) );
  NAND3_X1 U17895 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15427) );
  NAND2_X1 U17896 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14425) );
  NOR2_X1 U17897 ( .A1(n15427), .A2(n14425), .ZN(n15417) );
  AND2_X1 U17898 ( .A1(n15417), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15408) );
  AND4_X1 U17899 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n20434), .A4(n20438), .ZN(
        n14426) );
  NAND2_X1 U17900 ( .A1(n15408), .A2(n14426), .ZN(n15336) );
  NAND3_X1 U17901 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20450), .A3(
        n20434), .ZN(n15425) );
  INV_X1 U17902 ( .A(n15425), .ZN(n15396) );
  AND2_X1 U17903 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15396), .ZN(
        n14427) );
  NAND2_X1 U17904 ( .A1(n15408), .A2(n14427), .ZN(n15340) );
  OAI21_X1 U17905 ( .B1(n15426), .B2(n15336), .A(n15340), .ZN(n14430) );
  AND3_X1 U17906 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15335) );
  AND3_X1 U17907 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U17908 ( .A1(n15335), .A2(n14428), .ZN(n15313) );
  NOR2_X1 U17909 ( .A1(n15313), .A2(n15088), .ZN(n14429) );
  NAND2_X1 U17910 ( .A1(n14430), .A2(n14429), .ZN(n14431) );
  NAND2_X1 U17911 ( .A1(n14431), .A2(n20475), .ZN(n14432) );
  NAND2_X1 U17912 ( .A1(n14432), .A2(n20459), .ZN(n15304) );
  OR2_X1 U17913 ( .A1(n14433), .A2(n15304), .ZN(n15287) );
  INV_X1 U17914 ( .A(n14434), .ZN(n15258) );
  AND2_X1 U17915 ( .A1(n20475), .A2(n15258), .ZN(n14435) );
  NOR2_X1 U17916 ( .A1(n15287), .A2(n14435), .ZN(n15270) );
  NAND2_X1 U17917 ( .A1(n15270), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15261) );
  OR2_X1 U17918 ( .A1(n15261), .A2(n15269), .ZN(n14436) );
  AND2_X1 U17919 ( .A1(n14436), .A2(n14437), .ZN(n15253) );
  AOI21_X1 U17920 ( .B1(n14442), .B2(n14437), .A(n15253), .ZN(n15239) );
  OAI211_X1 U17921 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15345), .A(
        n15239), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15231) );
  NAND3_X1 U17922 ( .A1(n15231), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14437), .ZN(n14445) );
  INV_X1 U17923 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21160) );
  NOR2_X1 U17924 ( .A1(n20457), .A2(n21160), .ZN(n14508) );
  INV_X1 U17925 ( .A(n14508), .ZN(n14444) );
  INV_X1 U17926 ( .A(n15340), .ZN(n15337) );
  NAND2_X1 U17927 ( .A1(n20464), .A2(n15337), .ZN(n14438) );
  OR2_X1 U17928 ( .A1(n20452), .A2(n15336), .ZN(n15311) );
  NAND2_X1 U17929 ( .A1(n14438), .A2(n15311), .ZN(n15386) );
  NOR2_X1 U17930 ( .A1(n15313), .A2(n15312), .ZN(n14439) );
  NAND2_X1 U17931 ( .A1(n15386), .A2(n14439), .ZN(n15309) );
  NAND2_X1 U17932 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14440) );
  NOR2_X1 U17933 ( .A1(n15309), .A2(n14440), .ZN(n15294) );
  NAND2_X1 U17934 ( .A1(n15294), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15289) );
  INV_X1 U17935 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14441) );
  OR3_X2 U17936 ( .A1(n15289), .A2(n15259), .A3(n14441), .ZN(n15250) );
  NOR2_X1 U17937 ( .A1(n15250), .A2(n14442), .ZN(n15237) );
  NAND4_X1 U17938 ( .A1(n15237), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n12971), .ZN(n14443) );
  NAND3_X1 U17939 ( .A1(n14445), .A2(n14444), .A3(n14443), .ZN(n14446) );
  AOI21_X1 U17940 ( .B1(n14889), .B2(n20454), .A(n14446), .ZN(n14447) );
  OAI21_X1 U17941 ( .B1(n14513), .B2(n15456), .A(n14447), .ZN(P1_U3000) );
  OAI21_X1 U17942 ( .B1(n14448), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14469), .ZN(n15019) );
  AOI22_X1 U17943 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14449), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U17944 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14453) );
  AOI22_X1 U17945 ( .A1(n14450), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14452) );
  AOI22_X1 U17946 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14451) );
  NAND4_X1 U17947 ( .A1(n14454), .A2(n14453), .A3(n14452), .A4(n14451), .ZN(
        n14460) );
  AOI22_X1 U17948 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14458) );
  AOI22_X1 U17949 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14457) );
  AOI22_X1 U17950 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U17951 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14455) );
  NAND4_X1 U17952 ( .A1(n14458), .A2(n14457), .A3(n14456), .A4(n14455), .ZN(
        n14459) );
  NOR2_X1 U17953 ( .A1(n14460), .A2(n14459), .ZN(n14471) );
  NAND2_X1 U17954 ( .A1(n14462), .A2(n14461), .ZN(n14470) );
  XNOR2_X1 U17955 ( .A(n14471), .B(n14470), .ZN(n14466) );
  AOI21_X1 U17956 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n13022), .A(
        n14502), .ZN(n14464) );
  NAND2_X1 U17957 ( .A1(n14504), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n14463) );
  OAI211_X1 U17958 ( .C1(n14466), .C2(n14465), .A(n14464), .B(n14463), .ZN(
        n14467) );
  OAI21_X1 U17959 ( .B1(n15019), .B2(n14468), .A(n14467), .ZN(n14585) );
  XNOR2_X1 U17960 ( .A(n14469), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14576) );
  NOR2_X1 U17961 ( .A1(n14471), .A2(n14470), .ZN(n14496) );
  AOI22_X1 U17962 ( .A1(n14473), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14472), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U17963 ( .A1(n14475), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14474), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14480) );
  AOI22_X1 U17964 ( .A1(n14476), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12775), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U17965 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14028), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14478) );
  NAND4_X1 U17966 ( .A1(n14481), .A2(n14480), .A3(n14479), .A4(n14478), .ZN(
        n14494) );
  AOI22_X1 U17967 ( .A1(n14483), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14482), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U17968 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14102), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U17969 ( .A1(n14486), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14485), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14490) );
  AOI22_X1 U17970 ( .A1(n14488), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14487), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14489) );
  NAND4_X1 U17971 ( .A1(n14492), .A2(n14491), .A3(n14490), .A4(n14489), .ZN(
        n14493) );
  NOR2_X1 U17972 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  XNOR2_X1 U17973 ( .A(n14496), .B(n14495), .ZN(n14500) );
  OAI21_X1 U17974 ( .B1(n20832), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n13022), .ZN(n14497) );
  OAI21_X1 U17975 ( .B1(n9862), .B2(n21235), .A(n14497), .ZN(n14498) );
  AOI21_X1 U17976 ( .B1(n14500), .B2(n14499), .A(n14498), .ZN(n14501) );
  NAND2_X1 U17977 ( .A1(n14583), .A2(n14569), .ZN(n14507) );
  AOI22_X1 U17978 ( .A1(n14504), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n14503), .ZN(n14505) );
  INV_X1 U17979 ( .A(n14505), .ZN(n14506) );
  XNOR2_X2 U17980 ( .A(n14507), .B(n14506), .ZN(n14559) );
  AOI21_X1 U17981 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14508), .ZN(n14509) );
  OAI21_X1 U17982 ( .B1(n14510), .B2(n20433), .A(n14509), .ZN(n14511) );
  AOI21_X1 U17983 ( .B1(n14559), .B2(n20428), .A(n14511), .ZN(n14512) );
  OAI21_X1 U17984 ( .B1(n14513), .B2(n20253), .A(n14512), .ZN(P1_U2968) );
  INV_X1 U17985 ( .A(n14514), .ZN(n14518) );
  AOI211_X1 U17986 ( .C1(n14519), .C2(n14516), .A(n14515), .B(n15825), .ZN(
        n14517) );
  NAND2_X1 U17987 ( .A1(n14518), .A2(n14517), .ZN(n15827) );
  OAI21_X1 U17988 ( .B1(n14518), .B2(n14517), .A(n15827), .ZN(n14520) );
  INV_X1 U17989 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n14523) );
  AOI22_X1 U17990 ( .A1(n15985), .A2(n14521), .B1(n19396), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n14522) );
  OAI21_X1 U17991 ( .B1(n16007), .B2(n14523), .A(n14522), .ZN(n14528) );
  NAND2_X1 U17992 ( .A1(n14524), .A2(n14525), .ZN(n14526) );
  NAND2_X1 U17993 ( .A1(n9828), .A2(n14526), .ZN(n16325) );
  NOR2_X1 U17994 ( .A1(n16325), .A2(n16014), .ZN(n14527) );
  AOI211_X1 U17995 ( .C1(n16011), .C2(BUF1_REG_27__SCAN_IN), .A(n14528), .B(
        n14527), .ZN(n14529) );
  OAI21_X1 U17996 ( .B1(n14536), .B2(n16023), .A(n14529), .ZN(P2_U2892) );
  NOR2_X1 U17997 ( .A1(n14531), .A2(n14532), .ZN(n14533) );
  OR2_X1 U17998 ( .A1(n14530), .A2(n14533), .ZN(n15521) );
  NOR2_X1 U17999 ( .A1(n15521), .A2(n9733), .ZN(n14534) );
  AOI21_X1 U18000 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n9733), .A(n14534), .ZN(
        n14535) );
  OAI21_X1 U18001 ( .B1(n14536), .B2(n15897), .A(n14535), .ZN(P2_U2860) );
  AOI21_X1 U18002 ( .B1(n14537), .B2(n14540), .A(n14542), .ZN(n14543) );
  OAI22_X1 U18003 ( .A1(n14881), .A2(n14538), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15472), .ZN(n16725) );
  OAI22_X1 U18004 ( .A1(n16754), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21090), .ZN(n14539) );
  AOI21_X1 U18005 ( .B1(n16725), .B2(n14540), .A(n14539), .ZN(n14541) );
  OAI22_X1 U18006 ( .A1(n14543), .A2(n16728), .B1(n14542), .B2(n14541), .ZN(
        P1_U3474) );
  NOR2_X1 U18007 ( .A1(n14544), .A2(n9733), .ZN(n14545) );
  AOI21_X1 U18008 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n9733), .A(n14545), .ZN(
        n14546) );
  OAI21_X1 U18009 ( .B1(n10670), .B2(n15897), .A(n14546), .ZN(P2_U2857) );
  OAI21_X1 U18010 ( .B1(n14547), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n14549), 
        .ZN(n14548) );
  OAI21_X1 U18011 ( .B1(n14550), .B2(n14549), .A(n14548), .ZN(P2_U3612) );
  INV_X1 U18012 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n14555) );
  NAND3_X1 U18013 ( .A1(n14559), .A2(n14551), .A3(n15007), .ZN(n14554) );
  AOI22_X1 U18014 ( .A1(n14989), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14552), .ZN(n14553) );
  OAI211_X1 U18015 ( .C1(n14556), .C2(n14555), .A(n14554), .B(n14553), .ZN(
        P1_U2873) );
  OR2_X1 U18016 ( .A1(n14717), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14558) );
  MUX2_X1 U18017 ( .A(n14558), .B(n10602), .S(n14557), .Z(P1_U3487) );
  INV_X1 U18018 ( .A(n14559), .ZN(n14568) );
  INV_X1 U18019 ( .A(n14714), .ZN(n20286) );
  INV_X1 U18020 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21158) );
  INV_X1 U18021 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21162) );
  NOR2_X1 U18022 ( .A1(n21158), .A2(n21162), .ZN(n14560) );
  OAI21_X1 U18023 ( .B1(n20286), .B2(n14560), .A(n14590), .ZN(n14577) );
  INV_X1 U18024 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14561) );
  OAI22_X1 U18025 ( .A1(n14562), .A2(n16781), .B1(n20305), .B2(n14561), .ZN(
        n14565) );
  NAND2_X1 U18026 ( .A1(n14563), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14594) );
  NOR4_X1 U18027 ( .A1(n14594), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21162), 
        .A4(n21158), .ZN(n14564) );
  AOI211_X1 U18028 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14577), .A(n14565), 
        .B(n14564), .ZN(n14567) );
  NAND2_X1 U18029 ( .A1(n14889), .A2(n20333), .ZN(n14566) );
  OAI211_X1 U18030 ( .C1(n14568), .C2(n14856), .A(n14567), .B(n14566), .ZN(
        P1_U2809) );
  XOR2_X1 U18031 ( .A(n14569), .B(n14583), .Z(n15014) );
  INV_X1 U18032 ( .A(n15014), .ZN(n14936) );
  INV_X1 U18033 ( .A(n14587), .ZN(n14572) );
  INV_X1 U18034 ( .A(n14576), .ZN(n15012) );
  NOR2_X1 U18035 ( .A1(n14594), .A2(n21158), .ZN(n14578) );
  OAI21_X1 U18036 ( .B1(n14578), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14577), 
        .ZN(n14580) );
  AOI22_X1 U18037 ( .A1(n20334), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20335), .ZN(n14579) );
  OAI211_X1 U18038 ( .C1(n15012), .C2(n20330), .A(n14580), .B(n14579), .ZN(
        n14581) );
  AOI21_X1 U18039 ( .B1(n15232), .B2(n20333), .A(n14581), .ZN(n14582) );
  OAI21_X1 U18040 ( .B1(n14936), .B2(n14856), .A(n14582), .ZN(P1_U2810) );
  AOI21_X1 U18041 ( .B1(n14585), .B2(n14584), .A(n14583), .ZN(n15021) );
  INV_X1 U18042 ( .A(n15021), .ZN(n14942) );
  AOI21_X1 U18043 ( .B1(n14588), .B2(n14587), .A(n14586), .ZN(n15241) );
  INV_X1 U18044 ( .A(n15019), .ZN(n14592) );
  AOI22_X1 U18045 ( .A1(n20334), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20335), .ZN(n14589) );
  OAI21_X1 U18046 ( .B1(n14590), .B2(n21158), .A(n14589), .ZN(n14591) );
  AOI21_X1 U18047 ( .B1(n20344), .B2(n14592), .A(n14591), .ZN(n14593) );
  OAI21_X1 U18048 ( .B1(n14594), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14593), 
        .ZN(n14595) );
  AOI21_X1 U18049 ( .B1(n15241), .B2(n20333), .A(n14595), .ZN(n14596) );
  OAI21_X1 U18050 ( .B1(n14942), .B2(n14856), .A(n14596), .ZN(P1_U2811) );
  AND2_X1 U18051 ( .A1(n14597), .A2(n14598), .ZN(n14600) );
  OR2_X1 U18052 ( .A1(n14600), .A2(n14599), .ZN(n15036) );
  INV_X1 U18053 ( .A(n14601), .ZN(n14605) );
  INV_X1 U18054 ( .A(n14602), .ZN(n14604) );
  AOI21_X1 U18055 ( .B1(n14605), .B2(n14604), .A(n14603), .ZN(n15254) );
  NOR2_X1 U18056 ( .A1(n20330), .A2(n15038), .ZN(n14612) );
  INV_X1 U18057 ( .A(n14606), .ZN(n14607) );
  NAND2_X1 U18058 ( .A1(n14714), .A2(n14607), .ZN(n14619) );
  INV_X1 U18059 ( .A(n14608), .ZN(n14621) );
  NAND3_X1 U18060 ( .A1(n14621), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n21155), 
        .ZN(n14610) );
  AOI22_X1 U18061 ( .A1(n20334), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20335), .ZN(n14609) );
  OAI211_X1 U18062 ( .C1(n14619), .C2(n21155), .A(n14610), .B(n14609), .ZN(
        n14611) );
  AOI211_X1 U18063 ( .C1(n15254), .C2(n20333), .A(n14612), .B(n14611), .ZN(
        n14613) );
  OAI21_X1 U18064 ( .B1(n15036), .B2(n14856), .A(n14613), .ZN(P1_U2813) );
  INV_X1 U18065 ( .A(n14597), .ZN(n14615) );
  AOI21_X1 U18066 ( .B1(n14616), .B2(n14629), .A(n14615), .ZN(n15049) );
  INV_X1 U18067 ( .A(n15049), .ZN(n14952) );
  NOR2_X1 U18068 ( .A1(n14631), .A2(n14617), .ZN(n14618) );
  OR2_X1 U18069 ( .A1(n14602), .A2(n14618), .ZN(n15264) );
  INV_X1 U18070 ( .A(n15264), .ZN(n14625) );
  AOI22_X1 U18071 ( .A1(n20334), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20335), .ZN(n14623) );
  INV_X1 U18072 ( .A(n14619), .ZN(n14620) );
  OAI21_X1 U18073 ( .B1(n14621), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14620), 
        .ZN(n14622) );
  OAI211_X1 U18074 ( .C1(n20330), .C2(n15047), .A(n14623), .B(n14622), .ZN(
        n14624) );
  AOI21_X1 U18075 ( .B1(n14625), .B2(n20333), .A(n14624), .ZN(n14626) );
  OAI21_X1 U18076 ( .B1(n14952), .B2(n14856), .A(n14626), .ZN(P1_U2814) );
  AOI21_X1 U18077 ( .B1(n14630), .B2(n14628), .A(n14614), .ZN(n15058) );
  INV_X1 U18078 ( .A(n15058), .ZN(n14958) );
  AOI21_X1 U18079 ( .B1(n14632), .B2(n14649), .A(n14631), .ZN(n15273) );
  NAND2_X1 U18080 ( .A1(n14714), .A2(n14633), .ZN(n14660) );
  OAI21_X1 U18081 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n20322), .A(n14660), 
        .ZN(n14638) );
  INV_X1 U18082 ( .A(n14634), .ZN(n14636) );
  AOI22_X1 U18083 ( .A1(n20334), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20335), .ZN(n14635) );
  OAI21_X1 U18084 ( .B1(n14636), .B2(P1_REIP_REG_25__SCAN_IN), .A(n14635), 
        .ZN(n14637) );
  AOI21_X1 U18085 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n14638), .A(n14637), 
        .ZN(n14639) );
  OAI21_X1 U18086 ( .B1(n20330), .B2(n15056), .A(n14639), .ZN(n14640) );
  AOI21_X1 U18087 ( .B1(n15273), .B2(n20333), .A(n14640), .ZN(n14641) );
  OAI21_X1 U18088 ( .B1(n14958), .B2(n14856), .A(n14641), .ZN(P1_U2815) );
  OAI21_X1 U18089 ( .B1(n14642), .B2(n14643), .A(n14628), .ZN(n15066) );
  AOI22_X1 U18090 ( .A1(n20334), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20335), .ZN(n14646) );
  NAND3_X1 U18091 ( .A1(n20337), .A2(n14644), .A3(n21148), .ZN(n14645) );
  OAI211_X1 U18092 ( .C1(n14660), .C2(n21148), .A(n14646), .B(n14645), .ZN(
        n14651) );
  NAND2_X1 U18093 ( .A1(n14656), .A2(n14647), .ZN(n14648) );
  NAND2_X1 U18094 ( .A1(n14649), .A2(n14648), .ZN(n15276) );
  NOR2_X1 U18095 ( .A1(n15276), .A2(n20294), .ZN(n14650) );
  AOI211_X1 U18096 ( .C1(n20344), .C2(n15065), .A(n14651), .B(n14650), .ZN(
        n14652) );
  OAI21_X1 U18097 ( .B1(n15066), .B2(n14856), .A(n14652), .ZN(P1_U2816) );
  AND2_X1 U18098 ( .A1(n10624), .A2(n14654), .ZN(n14655) );
  OR2_X1 U18099 ( .A1(n14642), .A2(n14655), .ZN(n15071) );
  INV_X1 U18100 ( .A(n14656), .ZN(n14657) );
  AOI21_X1 U18101 ( .B1(n14658), .B2(n14675), .A(n14657), .ZN(n15291) );
  NOR2_X1 U18102 ( .A1(n20330), .A2(n15074), .ZN(n14663) );
  INV_X1 U18103 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15091) );
  INV_X1 U18104 ( .A(n14667), .ZN(n14684) );
  NOR3_X1 U18105 ( .A1(n20322), .A2(n15091), .A3(n14684), .ZN(n14669) );
  AOI21_X1 U18106 ( .B1(n14669), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14661) );
  AOI22_X1 U18107 ( .A1(n20334), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20335), .ZN(n14659) );
  OAI21_X1 U18108 ( .B1(n14661), .B2(n14660), .A(n14659), .ZN(n14662) );
  AOI211_X1 U18109 ( .C1(n15291), .C2(n20333), .A(n14663), .B(n14662), .ZN(
        n14664) );
  OAI21_X1 U18110 ( .B1(n15071), .B2(n14856), .A(n14664), .ZN(P1_U2817) );
  AOI21_X1 U18111 ( .B1(n14666), .B2(n14665), .A(n14653), .ZN(n15085) );
  INV_X1 U18112 ( .A(n15085), .ZN(n14970) );
  NAND2_X1 U18113 ( .A1(n14872), .A2(n14667), .ZN(n14668) );
  AND2_X1 U18114 ( .A1(n14714), .A2(n14668), .ZN(n14699) );
  AOI21_X1 U18115 ( .B1(n20337), .B2(n15091), .A(n14699), .ZN(n14672) );
  INV_X1 U18116 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21146) );
  AOI22_X1 U18117 ( .A1(n20334), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20335), .ZN(n14671) );
  NAND2_X1 U18118 ( .A1(n14669), .A2(n21146), .ZN(n14670) );
  OAI211_X1 U18119 ( .C1(n14672), .C2(n21146), .A(n14671), .B(n14670), .ZN(
        n14673) );
  AOI21_X1 U18120 ( .B1(n15081), .B2(n20344), .A(n14673), .ZN(n14680) );
  INV_X1 U18121 ( .A(n14683), .ZN(n14674) );
  NAND2_X1 U18122 ( .A1(n14695), .A2(n14674), .ZN(n14677) );
  INV_X1 U18123 ( .A(n14675), .ZN(n14676) );
  AOI21_X1 U18124 ( .B1(n14678), .B2(n14677), .A(n14676), .ZN(n15299) );
  NAND2_X1 U18125 ( .A1(n15299), .A2(n20333), .ZN(n14679) );
  OAI211_X1 U18126 ( .C1(n14970), .C2(n14856), .A(n14680), .B(n14679), .ZN(
        P1_U2818) );
  OAI21_X1 U18127 ( .B1(n14681), .B2(n14682), .A(n14665), .ZN(n15095) );
  XNOR2_X1 U18128 ( .A(n14695), .B(n14683), .ZN(n15305) );
  INV_X1 U18129 ( .A(n15094), .ZN(n14688) );
  OAI22_X1 U18130 ( .A1(n15092), .A2(n16781), .B1(n20305), .B2(n14900), .ZN(
        n14686) );
  NOR3_X1 U18131 ( .A1(n20322), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14684), 
        .ZN(n14685) );
  AOI211_X1 U18132 ( .C1(n14699), .C2(P1_REIP_REG_21__SCAN_IN), .A(n14686), 
        .B(n14685), .ZN(n14687) );
  OAI21_X1 U18133 ( .B1(n14688), .B2(n20330), .A(n14687), .ZN(n14689) );
  AOI21_X1 U18134 ( .B1(n15305), .B2(n20333), .A(n14689), .ZN(n14690) );
  OAI21_X1 U18135 ( .B1(n15095), .B2(n14856), .A(n14690), .ZN(P1_U2819) );
  NOR2_X1 U18136 ( .A1(n14691), .A2(n14692), .ZN(n14693) );
  OR2_X1 U18137 ( .A1(n14681), .A2(n14693), .ZN(n15101) );
  AOI21_X1 U18138 ( .B1(n14733), .B2(n14708), .A(n14694), .ZN(n14696) );
  NOR2_X1 U18139 ( .A1(n14696), .A2(n14695), .ZN(n15322) );
  INV_X1 U18140 ( .A(n15104), .ZN(n14703) );
  AOI22_X1 U18141 ( .A1(n20334), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20335), .ZN(n14702) );
  INV_X1 U18142 ( .A(n14709), .ZN(n14697) );
  NAND2_X1 U18143 ( .A1(n20337), .A2(n14697), .ZN(n20309) );
  NOR2_X1 U18144 ( .A1(n14711), .A2(n20309), .ZN(n20272) );
  AND2_X1 U18145 ( .A1(n14698), .A2(n20272), .ZN(n14822) );
  AND2_X1 U18146 ( .A1(n14755), .A2(n14822), .ZN(n14773) );
  NAND3_X1 U18147 ( .A1(n14773), .A2(P1_REIP_REG_17__SCAN_IN), .A3(n14756), 
        .ZN(n14728) );
  INV_X1 U18148 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15110) );
  INV_X1 U18149 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21140) );
  NOR3_X1 U18150 ( .A1(n14728), .A2(n15110), .A3(n21140), .ZN(n14700) );
  OAI21_X1 U18151 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n14700), .A(n14699), 
        .ZN(n14701) );
  OAI211_X1 U18152 ( .C1(n20330), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14704) );
  AOI21_X1 U18153 ( .B1(n15322), .B2(n20333), .A(n14704), .ZN(n14705) );
  OAI21_X1 U18154 ( .B1(n15101), .B2(n14856), .A(n14705), .ZN(P1_U2820) );
  AND2_X1 U18155 ( .A1(n9801), .A2(n14706), .ZN(n14707) );
  OR2_X1 U18156 ( .A1(n14707), .A2(n14691), .ZN(n15109) );
  XOR2_X1 U18157 ( .A(n14708), .B(n14733), .Z(n15329) );
  INV_X1 U18158 ( .A(n14872), .ZN(n20331) );
  OR2_X1 U18159 ( .A1(n20331), .A2(n14709), .ZN(n14710) );
  AND2_X1 U18160 ( .A1(n14714), .A2(n14710), .ZN(n20302) );
  AND2_X1 U18161 ( .A1(n14714), .A2(n14711), .ZN(n14712) );
  OR2_X1 U18162 ( .A1(n20302), .A2(n14712), .ZN(n20273) );
  AND2_X1 U18163 ( .A1(n14714), .A2(n14713), .ZN(n14715) );
  NOR2_X1 U18164 ( .A1(n20273), .A2(n14715), .ZN(n16790) );
  OAI21_X1 U18165 ( .B1(n14716), .B2(n20322), .A(n16790), .ZN(n14744) );
  NAND2_X1 U18166 ( .A1(n14744), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14722) );
  XNOR2_X1 U18167 ( .A(P1_REIP_REG_19__SCAN_IN), .B(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14719) );
  NAND2_X1 U18168 ( .A1(n20335), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14718) );
  NAND2_X1 U18169 ( .A1(n14872), .A2(n14717), .ZN(n20314) );
  OAI211_X1 U18170 ( .C1(n14728), .C2(n14719), .A(n14718), .B(n20314), .ZN(
        n14720) );
  AOI21_X1 U18171 ( .B1(n20334), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14720), .ZN(
        n14721) );
  OAI211_X1 U18172 ( .C1(n20330), .C2(n15112), .A(n14722), .B(n14721), .ZN(
        n14723) );
  AOI21_X1 U18173 ( .B1(n15329), .B2(n20333), .A(n14723), .ZN(n14724) );
  OAI21_X1 U18174 ( .B1(n15109), .B2(n14856), .A(n14724), .ZN(P1_U2821) );
  INV_X1 U18175 ( .A(n14725), .ZN(n14726) );
  OAI21_X1 U18176 ( .B1(n14726), .B2(n9901), .A(n9801), .ZN(n15123) );
  INV_X1 U18177 ( .A(n15120), .ZN(n14731) );
  NAND2_X1 U18178 ( .A1(n20335), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14727) );
  OAI211_X1 U18179 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n14728), .A(n14727), 
        .B(n20314), .ZN(n14729) );
  AOI21_X1 U18180 ( .B1(n20334), .B2(P1_EBX_REG_18__SCAN_IN), .A(n14729), .ZN(
        n14730) );
  OAI21_X1 U18181 ( .B1(n20330), .B2(n14731), .A(n14730), .ZN(n14736) );
  INV_X1 U18182 ( .A(n14741), .ZN(n14753) );
  AOI21_X1 U18183 ( .B1(n14753), .B2(n14740), .A(n14732), .ZN(n14734) );
  OR2_X1 U18184 ( .A1(n14734), .A2(n14733), .ZN(n15352) );
  NOR2_X1 U18185 ( .A1(n15352), .A2(n20294), .ZN(n14735) );
  AOI211_X1 U18186 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n14744), .A(n14736), 
        .B(n14735), .ZN(n14737) );
  OAI21_X1 U18187 ( .B1(n15123), .B2(n14856), .A(n14737), .ZN(P1_U2822) );
  OAI21_X1 U18188 ( .B1(n14738), .B2(n14739), .A(n14725), .ZN(n15128) );
  XNOR2_X1 U18189 ( .A(n14741), .B(n14740), .ZN(n15358) );
  INV_X1 U18190 ( .A(n20314), .ZN(n20296) );
  AOI21_X1 U18191 ( .B1(n20335), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20296), .ZN(n14743) );
  NAND2_X1 U18192 ( .A1(n20334), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14742) );
  OAI211_X1 U18193 ( .C1(n20330), .C2(n15131), .A(n14743), .B(n14742), .ZN(
        n14748) );
  INV_X1 U18194 ( .A(n14744), .ZN(n14746) );
  AOI21_X1 U18195 ( .B1(n14773), .B2(n14756), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n14745) );
  NOR2_X1 U18196 ( .A1(n14746), .A2(n14745), .ZN(n14747) );
  AOI211_X1 U18197 ( .C1(n20333), .C2(n15358), .A(n14748), .B(n14747), .ZN(
        n14749) );
  OAI21_X1 U18198 ( .B1(n15128), .B2(n14856), .A(n14749), .ZN(P1_U2823) );
  AND2_X1 U18199 ( .A1(n14750), .A2(n14751), .ZN(n14752) );
  OR2_X1 U18200 ( .A1(n14752), .A2(n14738), .ZN(n15142) );
  AOI21_X1 U18201 ( .B1(n14754), .B2(n14772), .A(n14753), .ZN(n15365) );
  INV_X1 U18202 ( .A(n15140), .ZN(n14762) );
  OAI21_X1 U18203 ( .B1(n14755), .B2(n20286), .A(n16790), .ZN(n14790) );
  NAND2_X1 U18204 ( .A1(n14790), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n14761) );
  INV_X1 U18205 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15137) );
  INV_X1 U18206 ( .A(n14756), .ZN(n14757) );
  OAI211_X1 U18207 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14773), .B(n14757), .ZN(n14758) );
  OAI211_X1 U18208 ( .C1(n16781), .C2(n15137), .A(n20314), .B(n14758), .ZN(
        n14759) );
  AOI21_X1 U18209 ( .B1(n20334), .B2(P1_EBX_REG_16__SCAN_IN), .A(n14759), .ZN(
        n14760) );
  OAI211_X1 U18210 ( .C1(n20330), .C2(n14762), .A(n14761), .B(n14760), .ZN(
        n14763) );
  AOI21_X1 U18211 ( .B1(n15365), .B2(n20333), .A(n14763), .ZN(n14764) );
  OAI21_X1 U18212 ( .B1(n15142), .B2(n14856), .A(n14764), .ZN(P1_U2824) );
  NAND2_X1 U18213 ( .A1(n14911), .A2(n14829), .ZN(n14768) );
  INV_X1 U18214 ( .A(n14766), .ZN(n14767) );
  AND2_X1 U18215 ( .A1(n14803), .A2(n14781), .ZN(n14782) );
  OAI21_X1 U18216 ( .B1(n14782), .B2(n14769), .A(n14750), .ZN(n15153) );
  OR2_X1 U18217 ( .A1(n14787), .A2(n14770), .ZN(n14771) );
  AND2_X1 U18218 ( .A1(n14772), .A2(n14771), .ZN(n15371) );
  NAND2_X1 U18219 ( .A1(n14790), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14778) );
  INV_X1 U18220 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21135) );
  AOI21_X1 U18221 ( .B1(n14773), .B2(n21135), .A(n20296), .ZN(n14774) );
  OAI21_X1 U18222 ( .B1(n14775), .B2(n16781), .A(n14774), .ZN(n14776) );
  AOI21_X1 U18223 ( .B1(n20334), .B2(P1_EBX_REG_15__SCAN_IN), .A(n14776), .ZN(
        n14777) );
  OAI211_X1 U18224 ( .C1(n20330), .C2(n15155), .A(n14778), .B(n14777), .ZN(
        n14779) );
  AOI21_X1 U18225 ( .B1(n20333), .B2(n15371), .A(n14779), .ZN(n14780) );
  OAI21_X1 U18226 ( .B1(n15153), .B2(n14856), .A(n14780), .ZN(P1_U2825) );
  INV_X1 U18227 ( .A(n14781), .ZN(n14784) );
  INV_X1 U18228 ( .A(n14803), .ZN(n14783) );
  AOI21_X1 U18229 ( .B1(n14784), .B2(n14783), .A(n14782), .ZN(n15168) );
  INV_X1 U18230 ( .A(n15168), .ZN(n14994) );
  INV_X1 U18231 ( .A(n14818), .ZN(n14786) );
  AOI21_X1 U18232 ( .B1(n14786), .B2(n14805), .A(n14785), .ZN(n14788) );
  OR2_X1 U18233 ( .A1(n14788), .A2(n14787), .ZN(n15380) );
  INV_X1 U18234 ( .A(n15380), .ZN(n14797) );
  INV_X1 U18235 ( .A(n14822), .ZN(n14832) );
  NOR2_X1 U18236 ( .A1(n14832), .A2(n14789), .ZN(n14791) );
  OAI21_X1 U18237 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14791), .A(n14790), 
        .ZN(n14795) );
  OAI21_X1 U18238 ( .B1(n16781), .B2(n14792), .A(n20314), .ZN(n14793) );
  AOI21_X1 U18239 ( .B1(n20334), .B2(P1_EBX_REG_14__SCAN_IN), .A(n14793), .ZN(
        n14794) );
  OAI211_X1 U18240 ( .C1(n20330), .C2(n15166), .A(n14795), .B(n14794), .ZN(
        n14796) );
  AOI21_X1 U18241 ( .B1(n20333), .B2(n14797), .A(n14796), .ZN(n14798) );
  OAI21_X1 U18242 ( .B1(n14994), .B2(n14856), .A(n14798), .ZN(P1_U2826) );
  OAI21_X1 U18243 ( .B1(n14911), .B2(n14799), .A(n14800), .ZN(n14830) );
  INV_X1 U18244 ( .A(n14829), .ZN(n14801) );
  OAI21_X1 U18245 ( .B1(n14830), .B2(n14801), .A(n14800), .ZN(n14815) );
  NAND2_X1 U18246 ( .A1(n14815), .A2(n14814), .ZN(n14813) );
  INV_X1 U18247 ( .A(n14802), .ZN(n14804) );
  AOI21_X1 U18248 ( .B1(n14813), .B2(n14804), .A(n14803), .ZN(n15179) );
  INV_X1 U18249 ( .A(n15179), .ZN(n14996) );
  XNOR2_X1 U18250 ( .A(n14818), .B(n14805), .ZN(n15391) );
  INV_X1 U18251 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21127) );
  INV_X1 U18252 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21129) );
  NOR4_X1 U18253 ( .A1(n21127), .A2(n21129), .A3(P1_REIP_REG_13__SCAN_IN), 
        .A4(n14832), .ZN(n14806) );
  AOI211_X1 U18254 ( .C1(n20335), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n14806), .B(n20296), .ZN(n14808) );
  NAND2_X1 U18255 ( .A1(n20334), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n14807) );
  OAI211_X1 U18256 ( .C1(n20330), .C2(n15177), .A(n14808), .B(n14807), .ZN(
        n14811) );
  NAND2_X1 U18257 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14809) );
  INV_X1 U18258 ( .A(n16790), .ZN(n14836) );
  AOI21_X1 U18259 ( .B1(n20337), .B2(n14809), .A(n14836), .ZN(n14824) );
  INV_X1 U18260 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21131) );
  NOR2_X1 U18261 ( .A1(n14824), .A2(n21131), .ZN(n14810) );
  AOI211_X1 U18262 ( .C1(n20333), .C2(n15391), .A(n14811), .B(n14810), .ZN(
        n14812) );
  OAI21_X1 U18263 ( .B1(n14996), .B2(n14856), .A(n14812), .ZN(P1_U2827) );
  OAI21_X1 U18264 ( .B1(n14815), .B2(n14814), .A(n14813), .ZN(n15188) );
  OAI21_X1 U18265 ( .B1(n14816), .B2(n14828), .A(n14817), .ZN(n14819) );
  AND2_X1 U18266 ( .A1(n14819), .A2(n14818), .ZN(n15405) );
  AOI21_X1 U18267 ( .B1(n20335), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20296), .ZN(n14821) );
  NAND2_X1 U18268 ( .A1(n20334), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n14820) );
  OAI211_X1 U18269 ( .C1(n20330), .C2(n15184), .A(n14821), .B(n14820), .ZN(
        n14826) );
  AOI21_X1 U18270 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n14822), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14823) );
  NOR2_X1 U18271 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  AOI211_X1 U18272 ( .C1(n15405), .C2(n20333), .A(n14826), .B(n14825), .ZN(
        n14827) );
  OAI21_X1 U18273 ( .B1(n15188), .B2(n14856), .A(n14827), .ZN(P1_U2828) );
  XNOR2_X1 U18274 ( .A(n14816), .B(n14828), .ZN(n15412) );
  XNOR2_X1 U18275 ( .A(n14830), .B(n14829), .ZN(n15195) );
  NAND2_X1 U18276 ( .A1(n15195), .A2(n20298), .ZN(n14838) );
  NAND2_X1 U18277 ( .A1(n20335), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14831) );
  OAI211_X1 U18278 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n14832), .A(n14831), 
        .B(n20314), .ZN(n14833) );
  AOI21_X1 U18279 ( .B1(n20334), .B2(P1_EBX_REG_11__SCAN_IN), .A(n14833), .ZN(
        n14834) );
  OAI21_X1 U18280 ( .B1(n20330), .B2(n15193), .A(n14834), .ZN(n14835) );
  AOI21_X1 U18281 ( .B1(n14836), .B2(P1_REIP_REG_11__SCAN_IN), .A(n14835), 
        .ZN(n14837) );
  OAI211_X1 U18282 ( .C1(n15412), .C2(n20294), .A(n14838), .B(n14837), .ZN(
        P1_U2829) );
  NAND2_X1 U18283 ( .A1(n15004), .A2(n15005), .ZN(n14926) );
  INV_X1 U18284 ( .A(n14839), .ZN(n14927) );
  INV_X1 U18285 ( .A(n14840), .ZN(n14841) );
  AND2_X1 U18286 ( .A1(n14924), .A2(n14841), .ZN(n14842) );
  INV_X1 U18287 ( .A(n15223), .ZN(n14849) );
  INV_X1 U18288 ( .A(n14918), .ZN(n14843) );
  AOI21_X1 U18289 ( .B1(n14844), .B2(n14928), .A(n14843), .ZN(n15446) );
  AOI22_X1 U18290 ( .A1(n20333), .A2(n15446), .B1(P1_REIP_REG_8__SCAN_IN), 
        .B2(n20273), .ZN(n14845) );
  AND2_X1 U18291 ( .A1(n20314), .A2(n14845), .ZN(n14847) );
  NAND2_X1 U18292 ( .A1(n20335), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14846) );
  OAI211_X1 U18293 ( .C1(n20305), .C2(n14259), .A(n14847), .B(n14846), .ZN(
        n14848) );
  AOI21_X1 U18294 ( .B1(n20344), .B2(n14849), .A(n14848), .ZN(n14852) );
  NAND3_X1 U18295 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14850) );
  OR3_X1 U18296 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14850), .A3(n20309), .ZN(
        n14851) );
  OAI211_X1 U18297 ( .C1(n15221), .C2(n14856), .A(n14852), .B(n14851), .ZN(
        P1_U2832) );
  NOR2_X1 U18298 ( .A1(n14853), .A2(n13022), .ZN(n14854) );
  NAND2_X1 U18299 ( .A1(n14872), .A2(n14854), .ZN(n14855) );
  NAND2_X1 U18300 ( .A1(n14856), .A2(n14855), .ZN(n20327) );
  INV_X1 U18301 ( .A(n14857), .ZN(n14865) );
  OAI221_X1 U18302 ( .B1(n20322), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20322), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n14872), .ZN(n14858) );
  AOI22_X1 U18303 ( .A1(n20335), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n14858), .ZN(n14859) );
  OAI21_X1 U18304 ( .B1(n14860), .B2(n20305), .A(n14859), .ZN(n14864) );
  INV_X1 U18305 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21115) );
  NAND4_X1 U18306 ( .A1(n20337), .A2(P1_REIP_REG_2__SCAN_IN), .A3(n21115), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n14861) );
  OAI21_X1 U18307 ( .B1(n20294), .B2(n14862), .A(n14861), .ZN(n14863) );
  AOI211_X1 U18308 ( .C1(n20344), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        n14869) );
  NOR2_X1 U18309 ( .A1(n14866), .A2(n13022), .ZN(n14867) );
  AND2_X1 U18310 ( .A1(n14872), .A2(n14867), .ZN(n20338) );
  NAND2_X1 U18311 ( .A1(n20775), .A2(n20338), .ZN(n14868) );
  OAI211_X1 U18312 ( .C1(n14870), .C2(n20341), .A(n14869), .B(n14868), .ZN(
        P1_U2837) );
  MUX2_X1 U18313 ( .A(n20330), .B(n16781), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14879) );
  INV_X1 U18314 ( .A(n20338), .ZN(n20318) );
  OAI22_X1 U18315 ( .A1(n20318), .A2(n14871), .B1(n13419), .B2(n14872), .ZN(
        n14877) );
  INV_X1 U18316 ( .A(n14873), .ZN(n14875) );
  OAI22_X1 U18317 ( .A1(n20294), .A2(n14875), .B1(n14874), .B2(n20305), .ZN(
        n14876) );
  AOI211_X1 U18318 ( .C1(n20337), .C2(n13419), .A(n14877), .B(n14876), .ZN(
        n14878) );
  OAI211_X1 U18319 ( .C1(n20341), .C2(n14880), .A(n14879), .B(n14878), .ZN(
        P1_U2839) );
  OAI22_X1 U18320 ( .A1(n14882), .A2(n20305), .B1(n20318), .B2(n14881), .ZN(
        n14884) );
  NOR2_X1 U18321 ( .A1(n20286), .A2(n13242), .ZN(n14883) );
  AOI211_X1 U18322 ( .C1(n14885), .C2(n20333), .A(n14884), .B(n14883), .ZN(
        n14887) );
  OAI21_X1 U18323 ( .B1(n20344), .B2(n20335), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14886) );
  OAI211_X1 U18324 ( .C1(n20341), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        P1_U2840) );
  INV_X1 U18325 ( .A(n14889), .ZN(n14890) );
  OAI22_X1 U18326 ( .A1(n14890), .A2(n14930), .B1(n20355), .B2(n14561), .ZN(
        P1_U2841) );
  OAI21_X1 U18327 ( .B1(n14936), .B2(n14932), .A(n14891), .ZN(P1_U2842) );
  AOI22_X1 U18328 ( .A1(n15241), .A2(n20350), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14922), .ZN(n14892) );
  OAI21_X1 U18329 ( .B1(n14942), .B2(n14932), .A(n14892), .ZN(P1_U2843) );
  AOI22_X1 U18330 ( .A1(n15254), .A2(n20350), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14922), .ZN(n14893) );
  OAI21_X1 U18331 ( .B1(n15036), .B2(n14932), .A(n14893), .ZN(P1_U2845) );
  INV_X1 U18332 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14894) );
  OAI222_X1 U18333 ( .A1(n14932), .A2(n14952), .B1(n14894), .B2(n20355), .C1(
        n15264), .C2(n14930), .ZN(P1_U2846) );
  AOI22_X1 U18334 ( .A1(n15273), .A2(n20350), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14922), .ZN(n14895) );
  OAI21_X1 U18335 ( .B1(n14958), .B2(n14932), .A(n14895), .ZN(P1_U2847) );
  INV_X1 U18336 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14896) );
  OAI222_X1 U18337 ( .A1(n14932), .A2(n15066), .B1(n14896), .B2(n20355), .C1(
        n15276), .C2(n14930), .ZN(P1_U2848) );
  AOI22_X1 U18338 ( .A1(n15291), .A2(n20350), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14922), .ZN(n14897) );
  OAI21_X1 U18339 ( .B1(n15071), .B2(n14932), .A(n14897), .ZN(P1_U2849) );
  AOI22_X1 U18340 ( .A1(n15299), .A2(n20350), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14922), .ZN(n14898) );
  OAI21_X1 U18341 ( .B1(n14970), .B2(n14932), .A(n14898), .ZN(P1_U2850) );
  INV_X1 U18342 ( .A(n15305), .ZN(n14899) );
  OAI222_X1 U18343 ( .A1(n15095), .A2(n14932), .B1(n14900), .B2(n20355), .C1(
        n14930), .C2(n14899), .ZN(P1_U2851) );
  INV_X1 U18344 ( .A(n15322), .ZN(n14901) );
  OAI222_X1 U18345 ( .A1(n15101), .A2(n14932), .B1(n21383), .B2(n20355), .C1(
        n14901), .C2(n14930), .ZN(P1_U2852) );
  AOI22_X1 U18346 ( .A1(n15329), .A2(n20350), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14922), .ZN(n14902) );
  OAI21_X1 U18347 ( .B1(n15109), .B2(n14932), .A(n14902), .ZN(P1_U2853) );
  INV_X1 U18348 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14903) );
  OAI222_X1 U18349 ( .A1(n15123), .A2(n14932), .B1(n14903), .B2(n20355), .C1(
        n15352), .C2(n14930), .ZN(P1_U2854) );
  AOI22_X1 U18350 ( .A1(n15358), .A2(n20350), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14922), .ZN(n14904) );
  OAI21_X1 U18351 ( .B1(n15128), .B2(n14932), .A(n14904), .ZN(P1_U2855) );
  AOI22_X1 U18352 ( .A1(n15365), .A2(n20350), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14922), .ZN(n14905) );
  OAI21_X1 U18353 ( .B1(n15142), .B2(n14932), .A(n14905), .ZN(P1_U2856) );
  AOI22_X1 U18354 ( .A1(n15371), .A2(n20350), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14922), .ZN(n14906) );
  OAI21_X1 U18355 ( .B1(n15153), .B2(n14932), .A(n14906), .ZN(P1_U2857) );
  INV_X1 U18356 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14907) );
  OAI222_X1 U18357 ( .A1(n14994), .A2(n14932), .B1(n14907), .B2(n20355), .C1(
        n15380), .C2(n14930), .ZN(P1_U2858) );
  AOI22_X1 U18358 ( .A1(n15391), .A2(n20350), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14922), .ZN(n14908) );
  OAI21_X1 U18359 ( .B1(n14996), .B2(n14932), .A(n14908), .ZN(P1_U2859) );
  AOI22_X1 U18360 ( .A1(n15405), .A2(n20350), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14922), .ZN(n14909) );
  OAI21_X1 U18361 ( .B1(n15188), .B2(n14932), .A(n14909), .ZN(P1_U2860) );
  INV_X1 U18362 ( .A(n15195), .ZN(n14998) );
  OAI222_X1 U18363 ( .A1(n14998), .A2(n14932), .B1(n21449), .B2(n20355), .C1(
        n14930), .C2(n15412), .ZN(P1_U2861) );
  NAND2_X1 U18364 ( .A1(n14916), .A2(n14915), .ZN(n14914) );
  INV_X1 U18365 ( .A(n14910), .ZN(n14912) );
  AOI21_X1 U18366 ( .B1(n14914), .B2(n14912), .A(n14911), .ZN(n16786) );
  INV_X1 U18367 ( .A(n16786), .ZN(n15000) );
  INV_X1 U18368 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21465) );
  OAI21_X1 U18369 ( .B1(n14919), .B2(n14913), .A(n14816), .ZN(n15421) );
  OAI222_X1 U18370 ( .A1(n15000), .A2(n14932), .B1(n20355), .B2(n21465), .C1(
        n15421), .C2(n14930), .ZN(P1_U2862) );
  OAI21_X1 U18371 ( .B1(n14916), .B2(n14915), .A(n14914), .ZN(n15213) );
  AND2_X1 U18372 ( .A1(n14918), .A2(n14917), .ZN(n14920) );
  OR2_X1 U18373 ( .A1(n14920), .A2(n14919), .ZN(n20270) );
  OAI222_X1 U18374 ( .A1(n15213), .A2(n14932), .B1(n14921), .B2(n20355), .C1(
        n20270), .C2(n14930), .ZN(P1_U2863) );
  AOI22_X1 U18375 ( .A1(n15446), .A2(n20350), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14922), .ZN(n14923) );
  OAI21_X1 U18376 ( .B1(n15221), .B2(n14932), .A(n14923), .ZN(P1_U2864) );
  INV_X1 U18377 ( .A(n14924), .ZN(n14925) );
  AOI21_X1 U18378 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n20287) );
  INV_X1 U18379 ( .A(n20287), .ZN(n15003) );
  INV_X1 U18380 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14931) );
  OAI21_X1 U18381 ( .B1(n9896), .B2(n14929), .A(n14928), .ZN(n20280) );
  OAI222_X1 U18382 ( .A1(n15003), .A2(n14932), .B1(n14931), .B2(n20355), .C1(
        n20280), .C2(n14930), .ZN(P1_U2865) );
  OAI22_X1 U18383 ( .A1(n14986), .A2(n14993), .B1(n15007), .B2(n21235), .ZN(
        n14933) );
  AOI21_X1 U18384 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14988), .A(n14933), .ZN(
        n14935) );
  NAND2_X1 U18385 ( .A1(n14989), .A2(DATAI_30_), .ZN(n14934) );
  OAI211_X1 U18386 ( .C1(n14936), .C2(n15009), .A(n14935), .B(n14934), .ZN(
        P1_U2874) );
  INV_X1 U18387 ( .A(DATAI_13_), .ZN(n14938) );
  INV_X1 U18388 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14937) );
  MUX2_X1 U18389 ( .A(n14938), .B(n14937), .S(n20488), .Z(n20403) );
  OAI22_X1 U18390 ( .A1(n14986), .A2(n20403), .B1(n15007), .B2(n13043), .ZN(
        n14939) );
  AOI21_X1 U18391 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14988), .A(n14939), .ZN(
        n14941) );
  NAND2_X1 U18392 ( .A1(n14989), .A2(DATAI_29_), .ZN(n14940) );
  OAI211_X1 U18393 ( .C1(n14942), .C2(n15009), .A(n14941), .B(n14940), .ZN(
        P1_U2875) );
  INV_X1 U18394 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16940) );
  NOR2_X1 U18395 ( .A1(n20485), .A2(n16940), .ZN(n14943) );
  AOI21_X1 U18396 ( .B1(DATAI_11_), .B2(n20485), .A(n14943), .ZN(n20397) );
  OAI22_X1 U18397 ( .A1(n14986), .A2(n20397), .B1(n15007), .B2(n13047), .ZN(
        n14944) );
  AOI21_X1 U18398 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14988), .A(n14944), .ZN(
        n14946) );
  NAND2_X1 U18399 ( .A1(n14989), .A2(DATAI_27_), .ZN(n14945) );
  OAI211_X1 U18400 ( .C1(n15036), .C2(n15009), .A(n14946), .B(n14945), .ZN(
        P1_U2877) );
  INV_X1 U18401 ( .A(DATAI_10_), .ZN(n14947) );
  INV_X1 U18402 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16942) );
  MUX2_X1 U18403 ( .A(n14947), .B(n16942), .S(n20488), .Z(n20394) );
  INV_X1 U18404 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14948) );
  OAI22_X1 U18405 ( .A1(n14986), .A2(n20394), .B1(n15007), .B2(n14948), .ZN(
        n14949) );
  AOI21_X1 U18406 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14988), .A(n14949), .ZN(
        n14951) );
  NAND2_X1 U18407 ( .A1(n14989), .A2(DATAI_26_), .ZN(n14950) );
  OAI211_X1 U18408 ( .C1(n14952), .C2(n15009), .A(n14951), .B(n14950), .ZN(
        P1_U2878) );
  INV_X1 U18409 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14953) );
  NOR2_X1 U18410 ( .A1(n20485), .A2(n14953), .ZN(n14954) );
  AOI21_X1 U18411 ( .B1(DATAI_9_), .B2(n20485), .A(n14954), .ZN(n20389) );
  OAI22_X1 U18412 ( .A1(n14986), .A2(n20389), .B1(n15007), .B2(n13039), .ZN(
        n14955) );
  AOI21_X1 U18413 ( .B1(n14988), .B2(BUF1_REG_25__SCAN_IN), .A(n14955), .ZN(
        n14957) );
  NAND2_X1 U18414 ( .A1(n14989), .A2(DATAI_25_), .ZN(n14956) );
  OAI211_X1 U18415 ( .C1(n14958), .C2(n15009), .A(n14957), .B(n14956), .ZN(
        P1_U2879) );
  INV_X1 U18416 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16945) );
  NOR2_X1 U18417 ( .A1(n20485), .A2(n16945), .ZN(n14959) );
  AOI21_X1 U18418 ( .B1(DATAI_8_), .B2(n20485), .A(n14959), .ZN(n20386) );
  OAI22_X1 U18419 ( .A1(n14986), .A2(n20386), .B1(n15007), .B2(n13041), .ZN(
        n14960) );
  AOI21_X1 U18420 ( .B1(BUF1_REG_24__SCAN_IN), .B2(n14988), .A(n14960), .ZN(
        n14962) );
  NAND2_X1 U18421 ( .A1(n14989), .A2(DATAI_24_), .ZN(n14961) );
  OAI211_X1 U18422 ( .C1(n15066), .C2(n15009), .A(n14962), .B(n14961), .ZN(
        P1_U2880) );
  OAI22_X1 U18423 ( .A1(n14986), .A2(n20536), .B1(n15007), .B2(n14963), .ZN(
        n14964) );
  AOI21_X1 U18424 ( .B1(n14988), .B2(BUF1_REG_23__SCAN_IN), .A(n14964), .ZN(
        n14966) );
  NAND2_X1 U18425 ( .A1(n14989), .A2(DATAI_23_), .ZN(n14965) );
  OAI211_X1 U18426 ( .C1(n15071), .C2(n15009), .A(n14966), .B(n14965), .ZN(
        P1_U2881) );
  OAI22_X1 U18427 ( .A1(n14986), .A2(n20528), .B1(n15007), .B2(n13363), .ZN(
        n14967) );
  AOI21_X1 U18428 ( .B1(n14988), .B2(BUF1_REG_22__SCAN_IN), .A(n14967), .ZN(
        n14969) );
  NAND2_X1 U18429 ( .A1(n14989), .A2(DATAI_22_), .ZN(n14968) );
  OAI211_X1 U18430 ( .C1(n14970), .C2(n15009), .A(n14969), .B(n14968), .ZN(
        P1_U2882) );
  OAI22_X1 U18431 ( .A1(n14986), .A2(n20524), .B1(n15007), .B2(n13366), .ZN(
        n14971) );
  AOI21_X1 U18432 ( .B1(n14988), .B2(BUF1_REG_21__SCAN_IN), .A(n14971), .ZN(
        n14973) );
  NAND2_X1 U18433 ( .A1(n14989), .A2(DATAI_21_), .ZN(n14972) );
  OAI211_X1 U18434 ( .C1(n15095), .C2(n15009), .A(n14973), .B(n14972), .ZN(
        P1_U2883) );
  OAI22_X1 U18435 ( .A1(n14986), .A2(n20520), .B1(n15007), .B2(n13361), .ZN(
        n14974) );
  AOI21_X1 U18436 ( .B1(n14988), .B2(BUF1_REG_20__SCAN_IN), .A(n14974), .ZN(
        n14976) );
  NAND2_X1 U18437 ( .A1(n14989), .A2(DATAI_20_), .ZN(n14975) );
  OAI211_X1 U18438 ( .C1(n15101), .C2(n15009), .A(n14976), .B(n14975), .ZN(
        P1_U2884) );
  OAI22_X1 U18439 ( .A1(n14986), .A2(n20516), .B1(n15007), .B2(n13050), .ZN(
        n14977) );
  AOI21_X1 U18440 ( .B1(n14988), .B2(BUF1_REG_19__SCAN_IN), .A(n14977), .ZN(
        n14979) );
  NAND2_X1 U18441 ( .A1(n14989), .A2(DATAI_19_), .ZN(n14978) );
  OAI211_X1 U18442 ( .C1(n15109), .C2(n15009), .A(n14979), .B(n14978), .ZN(
        P1_U2885) );
  OAI22_X1 U18443 ( .A1(n14986), .A2(n20512), .B1(n15007), .B2(n13052), .ZN(
        n14980) );
  AOI21_X1 U18444 ( .B1(n14988), .B2(BUF1_REG_18__SCAN_IN), .A(n14980), .ZN(
        n14982) );
  NAND2_X1 U18445 ( .A1(n14989), .A2(DATAI_18_), .ZN(n14981) );
  OAI211_X1 U18446 ( .C1(n15123), .C2(n15009), .A(n14982), .B(n14981), .ZN(
        P1_U2886) );
  OAI22_X1 U18447 ( .A1(n14986), .A2(n20508), .B1(n15007), .B2(n13037), .ZN(
        n14983) );
  AOI21_X1 U18448 ( .B1(n14988), .B2(BUF1_REG_17__SCAN_IN), .A(n14983), .ZN(
        n14985) );
  NAND2_X1 U18449 ( .A1(n14989), .A2(DATAI_17_), .ZN(n14984) );
  OAI211_X1 U18450 ( .C1(n15128), .C2(n15009), .A(n14985), .B(n14984), .ZN(
        P1_U2887) );
  OAI22_X1 U18451 ( .A1(n14986), .A2(n20499), .B1(n15007), .B2(n13035), .ZN(
        n14987) );
  AOI21_X1 U18452 ( .B1(n14988), .B2(BUF1_REG_16__SCAN_IN), .A(n14987), .ZN(
        n14991) );
  NAND2_X1 U18453 ( .A1(n14989), .A2(DATAI_16_), .ZN(n14990) );
  OAI211_X1 U18454 ( .C1(n15142), .C2(n15009), .A(n14991), .B(n14990), .ZN(
        P1_U2888) );
  OAI222_X1 U18455 ( .A1(n15009), .A2(n15153), .B1(n15006), .B2(n14992), .C1(
        n21259), .C2(n15007), .ZN(P1_U2889) );
  INV_X1 U18456 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20358) );
  OAI222_X1 U18457 ( .A1(n14994), .A2(n15009), .B1(n14993), .B2(n15006), .C1(
        n20358), .C2(n15007), .ZN(P1_U2890) );
  INV_X1 U18458 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14995) );
  OAI222_X1 U18459 ( .A1(n14996), .A2(n15009), .B1(n20403), .B2(n15006), .C1(
        n14995), .C2(n15007), .ZN(P1_U2891) );
  INV_X1 U18460 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14997) );
  OAI222_X1 U18461 ( .A1(n15188), .A2(n15009), .B1(n20400), .B2(n15006), .C1(
        n14997), .C2(n15007), .ZN(P1_U2892) );
  OAI222_X1 U18462 ( .A1(n14998), .A2(n15009), .B1(n20397), .B2(n15006), .C1(
        n20362), .C2(n15007), .ZN(P1_U2893) );
  INV_X1 U18463 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14999) );
  OAI222_X1 U18464 ( .A1(n15009), .A2(n15000), .B1(n20394), .B2(n15006), .C1(
        n14999), .C2(n15007), .ZN(P1_U2894) );
  OAI222_X1 U18465 ( .A1(n15213), .A2(n15009), .B1(n20389), .B2(n15006), .C1(
        n15001), .C2(n15007), .ZN(P1_U2895) );
  OAI222_X1 U18466 ( .A1(n15221), .A2(n15009), .B1(n20386), .B2(n15006), .C1(
        n15002), .C2(n15007), .ZN(P1_U2896) );
  INV_X1 U18467 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20367) );
  OAI222_X1 U18468 ( .A1(n15009), .A2(n15003), .B1(n20536), .B2(n15006), .C1(
        n15007), .C2(n20367), .ZN(P1_U2897) );
  XOR2_X1 U18469 ( .A(n15005), .B(n15004), .Z(n20352) );
  INV_X1 U18470 ( .A(n20352), .ZN(n15008) );
  INV_X1 U18471 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20369) );
  OAI222_X1 U18472 ( .A1(n15009), .A2(n15008), .B1(n15007), .B2(n20369), .C1(
        n15006), .C2(n20528), .ZN(P1_U2898) );
  XNOR2_X1 U18473 ( .A(n15010), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15235) );
  NOR2_X1 U18474 ( .A1(n20457), .A2(n21162), .ZN(n15229) );
  AOI21_X1 U18475 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15229), .ZN(n15011) );
  OAI21_X1 U18476 ( .B1(n15012), .B2(n20433), .A(n15011), .ZN(n15013) );
  AOI21_X1 U18477 ( .B1(n15014), .B2(n20428), .A(n15013), .ZN(n15015) );
  OAI21_X1 U18478 ( .B1(n20253), .B2(n15235), .A(n15015), .ZN(P1_U2969) );
  XNOR2_X1 U18479 ( .A(n10120), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15016) );
  XNOR2_X1 U18480 ( .A(n15017), .B(n15016), .ZN(n15243) );
  NOR2_X1 U18481 ( .A1(n20457), .A2(n21158), .ZN(n15236) );
  AOI21_X1 U18482 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15236), .ZN(n15018) );
  OAI21_X1 U18483 ( .B1(n15019), .B2(n20433), .A(n15018), .ZN(n15020) );
  AOI21_X1 U18484 ( .B1(n15021), .B2(n20428), .A(n15020), .ZN(n15022) );
  OAI21_X1 U18485 ( .B1(n15243), .B2(n20253), .A(n15022), .ZN(P1_U2970) );
  NAND2_X1 U18486 ( .A1(n15210), .A2(n15259), .ZN(n15042) );
  NAND2_X1 U18487 ( .A1(n15023), .A2(n15042), .ZN(n15026) );
  MUX2_X1 U18488 ( .A(n15035), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15210), .Z(n15025) );
  INV_X1 U18489 ( .A(n20433), .ZN(n15141) );
  NAND2_X1 U18490 ( .A1(n20436), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15244) );
  OAI21_X1 U18491 ( .B1(n15138), .B2(n15027), .A(n15244), .ZN(n15030) );
  NOR2_X1 U18492 ( .A1(n15028), .A2(n20487), .ZN(n15029) );
  AOI211_X2 U18493 ( .C1(n15141), .C2(n15031), .A(n15030), .B(n15029), .ZN(
        n15032) );
  INV_X1 U18494 ( .A(n15036), .ZN(n15040) );
  NOR2_X1 U18495 ( .A1(n20457), .A2(n21155), .ZN(n15252) );
  AOI21_X1 U18496 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15252), .ZN(n15037) );
  OAI21_X1 U18497 ( .B1(n20433), .B2(n15038), .A(n15037), .ZN(n15039) );
  AOI21_X1 U18498 ( .B1(n15040), .B2(n20428), .A(n15039), .ZN(n15041) );
  OAI211_X1 U18499 ( .C1(n10420), .C2(n15023), .A(n15043), .B(n15042), .ZN(
        n15044) );
  XOR2_X1 U18500 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15044), .Z(
        n15267) );
  OR2_X1 U18501 ( .A1(n20457), .A2(n21152), .ZN(n15263) );
  INV_X1 U18502 ( .A(n15263), .ZN(n15045) );
  AOI21_X1 U18503 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15045), .ZN(n15046) );
  OAI21_X1 U18504 ( .B1(n20433), .B2(n15047), .A(n15046), .ZN(n15048) );
  AOI21_X1 U18505 ( .B1(n15049), .B2(n20428), .A(n15048), .ZN(n15050) );
  OAI21_X1 U18506 ( .B1(n20253), .B2(n15267), .A(n15050), .ZN(P1_U2973) );
  INV_X1 U18507 ( .A(n15023), .ZN(n15051) );
  NAND3_X1 U18508 ( .A1(n15051), .A2(n21417), .A3(n15277), .ZN(n15053) );
  NAND2_X1 U18509 ( .A1(n15061), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15052) );
  MUX2_X1 U18510 ( .A(n15053), .B(n15052), .S(n15210), .Z(n15054) );
  XNOR2_X1 U18511 ( .A(n15054), .B(n15269), .ZN(n15275) );
  INV_X1 U18512 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21150) );
  OR2_X1 U18513 ( .A1(n20457), .A2(n21150), .ZN(n15268) );
  NAND2_X1 U18514 ( .A1(n20421), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15055) );
  OAI211_X1 U18515 ( .C1(n20433), .C2(n15056), .A(n15268), .B(n15055), .ZN(
        n15057) );
  AOI21_X1 U18516 ( .B1(n15058), .B2(n20428), .A(n15057), .ZN(n15059) );
  OAI21_X1 U18517 ( .B1(n20253), .B2(n15275), .A(n15059), .ZN(P1_U2974) );
  NOR2_X1 U18518 ( .A1(n15061), .A2(n15023), .ZN(n15060) );
  MUX2_X1 U18519 ( .A(n15061), .B(n15060), .S(n15189), .Z(n15062) );
  XNOR2_X1 U18520 ( .A(n15062), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15285) );
  NOR2_X1 U18521 ( .A1(n20457), .A2(n21148), .ZN(n15281) );
  NOR2_X1 U18522 ( .A1(n15138), .A2(n15063), .ZN(n15064) );
  AOI211_X1 U18523 ( .C1(n15141), .C2(n15065), .A(n15281), .B(n15064), .ZN(
        n15069) );
  INV_X1 U18524 ( .A(n15066), .ZN(n15067) );
  NAND2_X1 U18525 ( .A1(n15067), .A2(n20428), .ZN(n15068) );
  OAI211_X1 U18526 ( .C1(n15285), .C2(n20253), .A(n15069), .B(n15068), .ZN(
        P1_U2975) );
  XNOR2_X1 U18527 ( .A(n10120), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15070) );
  XNOR2_X1 U18528 ( .A(n15023), .B(n15070), .ZN(n15293) );
  INV_X1 U18529 ( .A(n15071), .ZN(n15076) );
  INV_X1 U18530 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15072) );
  NOR2_X1 U18531 ( .A1(n20457), .A2(n15072), .ZN(n15286) );
  AOI21_X1 U18532 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15286), .ZN(n15073) );
  OAI21_X1 U18533 ( .B1(n20433), .B2(n15074), .A(n15073), .ZN(n15075) );
  AOI21_X1 U18534 ( .B1(n15076), .B2(n20428), .A(n15075), .ZN(n15077) );
  OAI21_X1 U18535 ( .B1(n15293), .B2(n20253), .A(n15077), .ZN(P1_U2976) );
  NAND2_X1 U18536 ( .A1(n15078), .A2(n15079), .ZN(n15080) );
  XOR2_X1 U18537 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15080), .Z(
        n15301) );
  INV_X1 U18538 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15083) );
  NAND2_X1 U18539 ( .A1(n15141), .A2(n15081), .ZN(n15082) );
  OR2_X1 U18540 ( .A1(n20457), .A2(n21146), .ZN(n15295) );
  OAI211_X1 U18541 ( .C1(n15138), .C2(n15083), .A(n15082), .B(n15295), .ZN(
        n15084) );
  AOI21_X1 U18542 ( .B1(n15085), .B2(n20428), .A(n15084), .ZN(n15086) );
  OAI21_X1 U18543 ( .B1(n15301), .B2(n20253), .A(n15086), .ZN(P1_U2977) );
  XNOR2_X1 U18544 ( .A(n15189), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15116) );
  INV_X1 U18545 ( .A(n15106), .ZN(n15334) );
  NOR2_X1 U18546 ( .A1(n15334), .A2(n15088), .ZN(n15090) );
  NOR2_X1 U18547 ( .A1(n20457), .A2(n15091), .ZN(n15303) );
  NOR2_X1 U18548 ( .A1(n15138), .A2(n15092), .ZN(n15093) );
  AOI211_X1 U18549 ( .C1(n15141), .C2(n15094), .A(n15303), .B(n15093), .ZN(
        n15098) );
  INV_X1 U18550 ( .A(n15095), .ZN(n15096) );
  NAND2_X1 U18551 ( .A1(n15096), .A2(n20428), .ZN(n15097) );
  OAI211_X1 U18552 ( .C1(n15308), .C2(n20253), .A(n15098), .B(n15097), .ZN(
        P1_U2978) );
  XNOR2_X1 U18553 ( .A(n15099), .B(n15318), .ZN(n15324) );
  INV_X1 U18554 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21143) );
  OR2_X1 U18555 ( .A1(n20457), .A2(n21143), .ZN(n15317) );
  OAI21_X1 U18556 ( .B1(n15138), .B2(n15100), .A(n15317), .ZN(n15103) );
  NOR2_X1 U18557 ( .A1(n15101), .A2(n20487), .ZN(n15102) );
  AOI211_X1 U18558 ( .C1(n15141), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        n15105) );
  OAI21_X1 U18559 ( .B1(n15324), .B2(n20253), .A(n15105), .ZN(P1_U2979) );
  NOR2_X1 U18560 ( .A1(n15210), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15107) );
  MUX2_X1 U18561 ( .A(n15107), .B(n15210), .S(n15106), .Z(n15108) );
  XNOR2_X1 U18562 ( .A(n15108), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15332) );
  INV_X1 U18563 ( .A(n15109), .ZN(n15114) );
  NOR2_X1 U18564 ( .A1(n20457), .A2(n15110), .ZN(n15327) );
  AOI21_X1 U18565 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15327), .ZN(n15111) );
  OAI21_X1 U18566 ( .B1(n20433), .B2(n15112), .A(n15111), .ZN(n15113) );
  AOI21_X1 U18567 ( .B1(n15114), .B2(n20428), .A(n15113), .ZN(n15115) );
  OAI21_X1 U18568 ( .B1(n15332), .B2(n20253), .A(n15115), .ZN(P1_U2980) );
  NAND2_X1 U18569 ( .A1(n15117), .A2(n15116), .ZN(n15333) );
  NAND3_X1 U18570 ( .A1(n15334), .A2(n20429), .A3(n15333), .ZN(n15122) );
  NOR2_X1 U18571 ( .A1(n20457), .A2(n21140), .ZN(n15348) );
  INV_X1 U18572 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15118) );
  NOR2_X1 U18573 ( .A1(n15138), .A2(n15118), .ZN(n15119) );
  AOI211_X1 U18574 ( .C1(n15141), .C2(n15120), .A(n15348), .B(n15119), .ZN(
        n15121) );
  OAI211_X1 U18575 ( .C1(n20487), .C2(n15123), .A(n15122), .B(n15121), .ZN(
        P1_U2981) );
  INV_X1 U18576 ( .A(n15125), .ZN(n15126) );
  NAND2_X1 U18577 ( .A1(n15210), .A2(n21351), .ZN(n15149) );
  OAI21_X1 U18578 ( .B1(n15148), .B2(n15127), .A(n15149), .ZN(n15136) );
  XNOR2_X1 U18579 ( .A(n15189), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15135) );
  INV_X1 U18580 ( .A(n15128), .ZN(n15133) );
  INV_X1 U18581 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15129) );
  NOR2_X1 U18582 ( .A1(n20457), .A2(n15129), .ZN(n15357) );
  AOI21_X1 U18583 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15357), .ZN(n15130) );
  OAI21_X1 U18584 ( .B1(n20433), .B2(n15131), .A(n15130), .ZN(n15132) );
  AOI21_X1 U18585 ( .B1(n15133), .B2(n20428), .A(n15132), .ZN(n15134) );
  OAI21_X1 U18586 ( .B1(n15360), .B2(n20253), .A(n15134), .ZN(P1_U2982) );
  XNOR2_X1 U18587 ( .A(n15136), .B(n15135), .ZN(n15368) );
  INV_X1 U18588 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21137) );
  NOR2_X1 U18589 ( .A1(n20457), .A2(n21137), .ZN(n15364) );
  NOR2_X1 U18590 ( .A1(n15138), .A2(n15137), .ZN(n15139) );
  AOI211_X1 U18591 ( .C1(n15141), .C2(n15140), .A(n15364), .B(n15139), .ZN(
        n15145) );
  INV_X1 U18592 ( .A(n15142), .ZN(n15143) );
  NAND2_X1 U18593 ( .A1(n15143), .A2(n20428), .ZN(n15144) );
  OAI211_X1 U18594 ( .C1(n15368), .C2(n20253), .A(n15145), .B(n15144), .ZN(
        P1_U2983) );
  INV_X1 U18595 ( .A(n15146), .ZN(n15147) );
  NOR2_X1 U18596 ( .A1(n15148), .A2(n15147), .ZN(n15152) );
  NAND2_X1 U18597 ( .A1(n15150), .A2(n15149), .ZN(n15151) );
  XNOR2_X1 U18598 ( .A(n15152), .B(n15151), .ZN(n15375) );
  INV_X1 U18599 ( .A(n15153), .ZN(n15157) );
  NOR2_X1 U18600 ( .A1(n20457), .A2(n21135), .ZN(n15369) );
  AOI21_X1 U18601 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15369), .ZN(n15154) );
  OAI21_X1 U18602 ( .B1(n20433), .B2(n15155), .A(n15154), .ZN(n15156) );
  AOI21_X1 U18603 ( .B1(n15157), .B2(n20428), .A(n15156), .ZN(n15158) );
  OAI21_X1 U18604 ( .B1(n15375), .B2(n20253), .A(n15158), .ZN(P1_U2984) );
  INV_X1 U18605 ( .A(n15159), .ZN(n15162) );
  INV_X1 U18606 ( .A(n15160), .ZN(n15161) );
  AOI22_X1 U18607 ( .A1(n15162), .A2(n15161), .B1(n15189), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15164) );
  XNOR2_X1 U18608 ( .A(n10120), .B(n15377), .ZN(n15163) );
  XNOR2_X1 U18609 ( .A(n15164), .B(n15163), .ZN(n15385) );
  INV_X1 U18610 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21132) );
  NOR2_X1 U18611 ( .A1(n20457), .A2(n21132), .ZN(n15382) );
  AOI21_X1 U18612 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15382), .ZN(n15165) );
  OAI21_X1 U18613 ( .B1(n20433), .B2(n15166), .A(n15165), .ZN(n15167) );
  AOI21_X1 U18614 ( .B1(n15168), .B2(n20428), .A(n15167), .ZN(n15169) );
  OAI21_X1 U18615 ( .B1(n15385), .B2(n20253), .A(n15169), .ZN(P1_U2985) );
  AOI22_X1 U18616 ( .A1(n15199), .A2(n15171), .B1(n15189), .B2(n15170), .ZN(
        n15183) );
  INV_X1 U18617 ( .A(n15173), .ZN(n15172) );
  AOI21_X1 U18618 ( .B1(n15189), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15172), .ZN(n15182) );
  NAND2_X1 U18619 ( .A1(n15183), .A2(n15182), .ZN(n15181) );
  NAND2_X1 U18620 ( .A1(n15181), .A2(n15173), .ZN(n15174) );
  XOR2_X1 U18621 ( .A(n15175), .B(n15174), .Z(n15394) );
  NOR2_X1 U18622 ( .A1(n20457), .A2(n21131), .ZN(n15389) );
  AOI21_X1 U18623 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15389), .ZN(n15176) );
  OAI21_X1 U18624 ( .B1(n20433), .B2(n15177), .A(n15176), .ZN(n15178) );
  AOI21_X1 U18625 ( .B1(n15179), .B2(n20428), .A(n15178), .ZN(n15180) );
  OAI21_X1 U18626 ( .B1(n15394), .B2(n20253), .A(n15180), .ZN(P1_U2986) );
  OAI21_X1 U18627 ( .B1(n15183), .B2(n15182), .A(n15181), .ZN(n15395) );
  NAND2_X1 U18628 ( .A1(n15395), .A2(n20429), .ZN(n15187) );
  NOR2_X1 U18629 ( .A1(n20457), .A2(n21129), .ZN(n15404) );
  NOR2_X1 U18630 ( .A1(n20433), .A2(n15184), .ZN(n15185) );
  AOI211_X1 U18631 ( .C1(n20421), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15404), .B(n15185), .ZN(n15186) );
  OAI211_X1 U18632 ( .C1(n20487), .C2(n15188), .A(n15187), .B(n15186), .ZN(
        P1_U2987) );
  NOR2_X1 U18633 ( .A1(n15189), .A2(n15198), .ZN(n15190) );
  NOR3_X1 U18634 ( .A1(n15124), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15210), .ZN(n15202) );
  AOI21_X1 U18635 ( .B1(n15199), .B2(n15190), .A(n15202), .ZN(n15191) );
  XNOR2_X1 U18636 ( .A(n15191), .B(n15416), .ZN(n15420) );
  NOR2_X1 U18637 ( .A1(n20457), .A2(n21127), .ZN(n15414) );
  AOI21_X1 U18638 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15414), .ZN(n15192) );
  OAI21_X1 U18639 ( .B1(n20433), .B2(n15193), .A(n15192), .ZN(n15194) );
  AOI21_X1 U18640 ( .B1(n15195), .B2(n20428), .A(n15194), .ZN(n15196) );
  OAI21_X1 U18641 ( .B1(n15420), .B2(n20253), .A(n15196), .ZN(P1_U2988) );
  NOR2_X1 U18642 ( .A1(n15197), .A2(n15198), .ZN(n15201) );
  XNOR2_X1 U18643 ( .A(n15199), .B(n15198), .ZN(n15200) );
  MUX2_X1 U18644 ( .A(n15201), .B(n15200), .S(n10120), .Z(n15203) );
  NOR2_X1 U18645 ( .A1(n15203), .A2(n15202), .ZN(n15435) );
  INV_X1 U18646 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15204) );
  NOR2_X1 U18647 ( .A1(n20457), .A2(n15204), .ZN(n15424) );
  AOI21_X1 U18648 ( .B1(n20421), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15424), .ZN(n15205) );
  OAI21_X1 U18649 ( .B1(n20433), .B2(n16784), .A(n15205), .ZN(n15206) );
  AOI21_X1 U18650 ( .B1(n16786), .B2(n20428), .A(n15206), .ZN(n15207) );
  OAI21_X1 U18651 ( .B1(n15435), .B2(n20253), .A(n15207), .ZN(P1_U2989) );
  NAND2_X1 U18652 ( .A1(n15209), .A2(n15208), .ZN(n15212) );
  XNOR2_X1 U18653 ( .A(n10120), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15211) );
  XNOR2_X1 U18654 ( .A(n15212), .B(n15211), .ZN(n15441) );
  INV_X1 U18655 ( .A(n15213), .ZN(n20276) );
  INV_X1 U18656 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15214) );
  OR2_X1 U18657 ( .A1(n20457), .A2(n15214), .ZN(n15436) );
  NAND2_X1 U18658 ( .A1(n20421), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15215) );
  OAI211_X1 U18659 ( .C1(n20433), .C2(n20274), .A(n15436), .B(n15215), .ZN(
        n15216) );
  AOI21_X1 U18660 ( .B1(n20276), .B2(n20428), .A(n15216), .ZN(n15217) );
  OAI21_X1 U18661 ( .B1(n15441), .B2(n20253), .A(n15217), .ZN(P1_U2990) );
  XOR2_X1 U18662 ( .A(n15219), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(
        n15220) );
  XNOR2_X1 U18663 ( .A(n15218), .B(n15220), .ZN(n15455) );
  INV_X1 U18664 ( .A(n15221), .ZN(n15225) );
  NAND2_X1 U18665 ( .A1(n20436), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15447) );
  NAND2_X1 U18666 ( .A1(n20421), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15222) );
  OAI211_X1 U18667 ( .C1(n20433), .C2(n15223), .A(n15447), .B(n15222), .ZN(
        n15224) );
  AOI21_X1 U18668 ( .B1(n15225), .B2(n20428), .A(n15224), .ZN(n15226) );
  OAI21_X1 U18669 ( .B1(n15455), .B2(n20253), .A(n15226), .ZN(P1_U2991) );
  INV_X1 U18670 ( .A(n15237), .ZN(n15228) );
  OAI21_X1 U18671 ( .B1(n15228), .B2(n14406), .A(n15227), .ZN(n15230) );
  AOI21_X1 U18672 ( .B1(n15231), .B2(n15230), .A(n15229), .ZN(n15234) );
  NAND2_X1 U18673 ( .A1(n15232), .A2(n20454), .ZN(n15233) );
  OAI211_X1 U18674 ( .C1(n15235), .C2(n15456), .A(n15234), .B(n15233), .ZN(
        P1_U3001) );
  AOI21_X1 U18675 ( .B1(n15237), .B2(n14406), .A(n15236), .ZN(n15238) );
  OAI21_X1 U18676 ( .B1(n15239), .B2(n14406), .A(n15238), .ZN(n15240) );
  AOI21_X1 U18677 ( .B1(n15241), .B2(n20454), .A(n15240), .ZN(n15242) );
  OAI21_X1 U18678 ( .B1(n15243), .B2(n15456), .A(n15242), .ZN(P1_U3002) );
  XNOR2_X1 U18679 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U18680 ( .A1(n15253), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15245) );
  OAI211_X1 U18681 ( .C1(n15250), .C2(n15246), .A(n15245), .B(n15244), .ZN(
        n15247) );
  AOI21_X1 U18682 ( .B1(n15248), .B2(n20454), .A(n15247), .ZN(n15249) );
  NOR2_X1 U18683 ( .A1(n15250), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15251) );
  AOI211_X1 U18684 ( .C1(n15253), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15252), .B(n15251), .ZN(n15256) );
  NAND2_X1 U18685 ( .A1(n15254), .A2(n20454), .ZN(n15255) );
  OAI211_X1 U18686 ( .C1(n15257), .C2(n15456), .A(n15256), .B(n15255), .ZN(
        P1_U3004) );
  NOR3_X1 U18687 ( .A1(n15289), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15258), .ZN(n15272) );
  NOR2_X1 U18688 ( .A1(n15289), .A2(n15259), .ZN(n15260) );
  OAI22_X1 U18689 ( .A1(n15272), .A2(n15261), .B1(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15260), .ZN(n15262) );
  OAI211_X1 U18690 ( .C1(n15264), .C2(n20471), .A(n15263), .B(n15262), .ZN(
        n15265) );
  INV_X1 U18691 ( .A(n15265), .ZN(n15266) );
  OAI21_X1 U18692 ( .B1(n15267), .B2(n15456), .A(n15266), .ZN(P1_U3005) );
  OAI21_X1 U18693 ( .B1(n15270), .B2(n15269), .A(n15268), .ZN(n15271) );
  AOI211_X1 U18694 ( .C1(n15273), .C2(n20454), .A(n15272), .B(n15271), .ZN(
        n15274) );
  OAI21_X1 U18695 ( .B1(n15275), .B2(n15456), .A(n15274), .ZN(P1_U3006) );
  NOR2_X1 U18696 ( .A1(n15276), .A2(n20471), .ZN(n15283) );
  NOR3_X1 U18697 ( .A1(n15289), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n21417), .ZN(n15282) );
  INV_X1 U18698 ( .A(n15287), .ZN(n15279) );
  OAI21_X1 U18699 ( .B1(n20464), .B2(n15398), .A(n21417), .ZN(n15278) );
  AOI21_X1 U18700 ( .B1(n15279), .B2(n15278), .A(n15277), .ZN(n15280) );
  NOR4_X1 U18701 ( .A1(n15283), .A2(n15282), .A3(n15281), .A4(n15280), .ZN(
        n15284) );
  OAI21_X1 U18702 ( .B1(n15285), .B2(n15456), .A(n15284), .ZN(P1_U3007) );
  AOI21_X1 U18703 ( .B1(n15287), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15286), .ZN(n15288) );
  OAI21_X1 U18704 ( .B1(n15289), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15288), .ZN(n15290) );
  AOI21_X1 U18705 ( .B1(n15291), .B2(n20454), .A(n15290), .ZN(n15292) );
  OAI21_X1 U18706 ( .B1(n15293), .B2(n15456), .A(n15292), .ZN(P1_U3008) );
  INV_X1 U18707 ( .A(n15294), .ZN(n15297) );
  NOR3_X1 U18708 ( .A1(n15309), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15318), .ZN(n15302) );
  OAI21_X1 U18709 ( .B1(n15302), .B2(n15304), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15296) );
  OAI211_X1 U18710 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15297), .A(
        n15296), .B(n15295), .ZN(n15298) );
  AOI21_X1 U18711 ( .B1(n15299), .B2(n20454), .A(n15298), .ZN(n15300) );
  OAI21_X1 U18712 ( .B1(n15301), .B2(n15456), .A(n15300), .ZN(P1_U3009) );
  AOI211_X1 U18713 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15304), .A(
        n15303), .B(n15302), .ZN(n15307) );
  NAND2_X1 U18714 ( .A1(n15305), .A2(n20454), .ZN(n15306) );
  OAI211_X1 U18715 ( .C1(n15308), .C2(n15456), .A(n15307), .B(n15306), .ZN(
        P1_U3010) );
  NOR2_X1 U18716 ( .A1(n15309), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15321) );
  NOR2_X1 U18717 ( .A1(n15313), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15328) );
  INV_X1 U18718 ( .A(n15341), .ZN(n15310) );
  NAND2_X1 U18719 ( .A1(n15311), .A2(n15310), .ZN(n15343) );
  NAND2_X1 U18720 ( .A1(n15339), .A2(n15312), .ZN(n15316) );
  OAI21_X1 U18721 ( .B1(n15340), .B2(n15313), .A(n15426), .ZN(n15315) );
  OAI21_X1 U18722 ( .B1(n15336), .B2(n15313), .A(n15398), .ZN(n15314) );
  NAND4_X1 U18723 ( .A1(n20459), .A2(n15316), .A3(n15315), .A4(n15314), .ZN(
        n15325) );
  AOI21_X1 U18724 ( .B1(n15328), .B2(n15343), .A(n15325), .ZN(n15319) );
  OAI21_X1 U18725 ( .B1(n15319), .B2(n15318), .A(n15317), .ZN(n15320) );
  AOI211_X1 U18726 ( .C1(n15322), .C2(n20454), .A(n15321), .B(n15320), .ZN(
        n15323) );
  OAI21_X1 U18727 ( .B1(n15324), .B2(n15456), .A(n15323), .ZN(P1_U3011) );
  AND2_X1 U18728 ( .A1(n15325), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15326) );
  AOI211_X1 U18729 ( .C1(n15328), .C2(n15386), .A(n15327), .B(n15326), .ZN(
        n15331) );
  NAND2_X1 U18730 ( .A1(n15329), .A2(n20454), .ZN(n15330) );
  OAI211_X1 U18731 ( .C1(n15332), .C2(n15456), .A(n15331), .B(n15330), .ZN(
        P1_U3012) );
  NAND3_X1 U18732 ( .A1(n15334), .A2(n20477), .A3(n15333), .ZN(n15351) );
  INV_X1 U18733 ( .A(n15335), .ZN(n15346) );
  INV_X1 U18734 ( .A(n15336), .ZN(n15378) );
  NAND2_X1 U18735 ( .A1(n15337), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15338) );
  AOI22_X1 U18736 ( .A1(n15341), .A2(n15340), .B1(n15339), .B2(n15338), .ZN(
        n15342) );
  OAI211_X1 U18737 ( .C1(n15378), .C2(n20452), .A(n20459), .B(n15342), .ZN(
        n15390) );
  AOI21_X1 U18738 ( .B1(n15344), .B2(n15343), .A(n15390), .ZN(n15376) );
  OAI21_X1 U18739 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15345), .A(
        n15376), .ZN(n15372) );
  AOI21_X1 U18740 ( .B1(n20475), .B2(n15346), .A(n15372), .ZN(n15353) );
  INV_X1 U18741 ( .A(n15353), .ZN(n15349) );
  AND3_X1 U18742 ( .A1(n15386), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15370) );
  INV_X1 U18743 ( .A(n15370), .ZN(n15362) );
  NOR3_X1 U18744 ( .A1(n15362), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15346), .ZN(n15347) );
  AOI211_X1 U18745 ( .C1(n15349), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15348), .B(n15347), .ZN(n15350) );
  OAI211_X1 U18746 ( .C1(n20471), .C2(n15352), .A(n15351), .B(n15350), .ZN(
        P1_U3013) );
  NAND3_X1 U18747 ( .A1(n15370), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15354) );
  AOI21_X1 U18748 ( .B1(n15355), .B2(n15354), .A(n15353), .ZN(n15356) );
  AOI211_X1 U18749 ( .C1(n20454), .C2(n15358), .A(n15357), .B(n15356), .ZN(
        n15359) );
  OAI21_X1 U18750 ( .B1(n15360), .B2(n15456), .A(n15359), .ZN(P1_U3014) );
  XNOR2_X1 U18751 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15361) );
  NOR2_X1 U18752 ( .A1(n15362), .A2(n15361), .ZN(n15363) );
  AOI211_X1 U18753 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15372), .A(
        n15364), .B(n15363), .ZN(n15367) );
  NAND2_X1 U18754 ( .A1(n15365), .A2(n20454), .ZN(n15366) );
  OAI211_X1 U18755 ( .C1(n15368), .C2(n15456), .A(n15367), .B(n15366), .ZN(
        P1_U3015) );
  AOI21_X1 U18756 ( .B1(n15370), .B2(n21351), .A(n15369), .ZN(n15374) );
  AOI22_X1 U18757 ( .A1(n15372), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20454), .B2(n15371), .ZN(n15373) );
  OAI211_X1 U18758 ( .C1(n15375), .C2(n15456), .A(n15374), .B(n15373), .ZN(
        P1_U3016) );
  INV_X1 U18759 ( .A(n15376), .ZN(n15383) );
  NAND4_X1 U18760 ( .A1(n15407), .A2(n15378), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n15377), .ZN(n15379) );
  OAI21_X1 U18761 ( .B1(n15380), .B2(n20471), .A(n15379), .ZN(n15381) );
  AOI211_X1 U18762 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15383), .A(
        n15382), .B(n15381), .ZN(n15384) );
  OAI21_X1 U18763 ( .B1(n15385), .B2(n15456), .A(n15384), .ZN(P1_U3017) );
  INV_X1 U18764 ( .A(n15386), .ZN(n15387) );
  NOR2_X1 U18765 ( .A1(n15387), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15388) );
  AOI211_X1 U18766 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15390), .A(
        n15389), .B(n15388), .ZN(n15393) );
  NAND2_X1 U18767 ( .A1(n15391), .A2(n20454), .ZN(n15392) );
  OAI211_X1 U18768 ( .C1(n15394), .C2(n15456), .A(n15393), .B(n15392), .ZN(
        P1_U3018) );
  INV_X1 U18769 ( .A(n15395), .ZN(n15411) );
  INV_X1 U18770 ( .A(n15444), .ZN(n15401) );
  NAND2_X1 U18771 ( .A1(n15417), .A2(n15396), .ZN(n15399) );
  INV_X1 U18772 ( .A(n15408), .ZN(n15397) );
  AOI22_X1 U18773 ( .A1(n15426), .A2(n15399), .B1(n15398), .B2(n15397), .ZN(
        n15400) );
  NAND2_X1 U18774 ( .A1(n15432), .A2(n15400), .ZN(n15415) );
  AOI21_X1 U18775 ( .B1(n15401), .B2(n15416), .A(n15415), .ZN(n15402) );
  NOR2_X1 U18776 ( .A1(n15402), .A2(n14270), .ZN(n15403) );
  AOI211_X1 U18777 ( .C1(n20454), .C2(n15405), .A(n15404), .B(n15403), .ZN(
        n15410) );
  NAND3_X1 U18778 ( .A1(n15449), .A2(n15408), .A3(n14270), .ZN(n15409) );
  OAI211_X1 U18779 ( .C1(n15411), .C2(n15456), .A(n15410), .B(n15409), .ZN(
        P1_U3019) );
  NOR2_X1 U18780 ( .A1(n15412), .A2(n20471), .ZN(n15413) );
  AOI211_X1 U18781 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15415), .A(
        n15414), .B(n15413), .ZN(n15419) );
  NAND3_X1 U18782 ( .A1(n15449), .A2(n15417), .A3(n15416), .ZN(n15418) );
  OAI211_X1 U18783 ( .C1(n15420), .C2(n15456), .A(n15419), .B(n15418), .ZN(
        P1_U3020) );
  INV_X1 U18784 ( .A(n15421), .ZN(n16783) );
  INV_X1 U18785 ( .A(n15449), .ZN(n16820) );
  NOR4_X1 U18786 ( .A1(n16820), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15422), .A4(n15427), .ZN(n15423) );
  AOI211_X1 U18787 ( .C1(n20454), .C2(n16783), .A(n15424), .B(n15423), .ZN(
        n15434) );
  NOR3_X1 U18788 ( .A1(n16820), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n15427), .ZN(n15437) );
  NAND2_X1 U18789 ( .A1(n15426), .A2(n15425), .ZN(n15429) );
  INV_X1 U18790 ( .A(n15427), .ZN(n15428) );
  NAND2_X1 U18791 ( .A1(n15429), .A2(n15428), .ZN(n15430) );
  NAND2_X1 U18792 ( .A1(n20475), .A2(n15430), .ZN(n15431) );
  NAND2_X1 U18793 ( .A1(n15432), .A2(n15431), .ZN(n15439) );
  OAI21_X1 U18794 ( .B1(n15437), .B2(n15439), .A(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15433) );
  OAI211_X1 U18795 ( .C1(n15435), .C2(n15456), .A(n15434), .B(n15433), .ZN(
        P1_U3021) );
  OAI21_X1 U18796 ( .B1(n20270), .B2(n20471), .A(n15436), .ZN(n15438) );
  AOI211_X1 U18797 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15439), .A(
        n15438), .B(n15437), .ZN(n15440) );
  OAI21_X1 U18798 ( .B1(n15441), .B2(n15456), .A(n15440), .ZN(P1_U3022) );
  OAI21_X1 U18799 ( .B1(n15444), .B2(n15443), .A(n15442), .ZN(n16816) );
  AOI21_X1 U18800 ( .B1(n15445), .B2(n20475), .A(n16816), .ZN(n16810) );
  INV_X1 U18801 ( .A(n16810), .ZN(n15453) );
  INV_X1 U18802 ( .A(n15446), .ZN(n15448) );
  OAI21_X1 U18803 ( .B1(n15448), .B2(n20471), .A(n15447), .ZN(n15452) );
  NAND2_X1 U18804 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15449), .ZN(
        n16812) );
  AOI221_X1 U18805 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15450), .C2(n16811), .A(
        n16812), .ZN(n15451) );
  AOI211_X1 U18806 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n15453), .A(
        n15452), .B(n15451), .ZN(n15454) );
  OAI21_X1 U18807 ( .B1(n15456), .B2(n15455), .A(n15454), .ZN(P1_U3023) );
  OAI21_X1 U18808 ( .B1(n20568), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20908), 
        .ZN(n15457) );
  OAI22_X1 U18809 ( .A1(n15457), .A2(n20748), .B1(n14871), .B2(n15460), .ZN(
        n15458) );
  MUX2_X1 U18810 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15458), .S(
        n20483), .Z(P1_U3477) );
  INV_X1 U18811 ( .A(n20748), .ZN(n20612) );
  AOI21_X1 U18812 ( .B1(n20612), .B2(n20489), .A(n21030), .ZN(n20877) );
  OAI21_X1 U18813 ( .B1(n20489), .B2(n20612), .A(n20877), .ZN(n15459) );
  OAI21_X1 U18814 ( .B1(n15460), .B2(n12949), .A(n15459), .ZN(n15461) );
  MUX2_X1 U18815 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15461), .S(
        n20483), .Z(P1_U3476) );
  NAND2_X1 U18816 ( .A1(n20873), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15463) );
  AOI22_X1 U18817 ( .A1(n15463), .A2(n15462), .B1(n20748), .B2(n20742), .ZN(
        n15467) );
  OR2_X1 U18818 ( .A1(n20568), .A2(n20832), .ZN(n20804) );
  NOR2_X1 U18819 ( .A1(n20804), .A2(n21030), .ZN(n15464) );
  AND2_X1 U18820 ( .A1(n20987), .A2(n15464), .ZN(n20957) );
  AOI21_X1 U18821 ( .B1(n15465), .B2(n20775), .A(n20957), .ZN(n15466) );
  OAI21_X1 U18822 ( .B1(n15467), .B2(n21030), .A(n15466), .ZN(n15468) );
  MUX2_X1 U18823 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15468), .S(
        n20483), .Z(P1_U3475) );
  NAND2_X1 U18824 ( .A1(n15471), .A2(n15470), .ZN(n15475) );
  OAI22_X1 U18825 ( .A1(n16727), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15475), .B2(n15472), .ZN(n15473) );
  AOI21_X1 U18826 ( .B1(n20988), .B2(n15474), .A(n15473), .ZN(n16729) );
  INV_X1 U18827 ( .A(n15475), .ZN(n15479) );
  INV_X1 U18828 ( .A(n15476), .ZN(n15477) );
  AOI22_X1 U18829 ( .A1(n15480), .A2(n15479), .B1(n15478), .B2(n15477), .ZN(
        n15481) );
  OAI21_X1 U18830 ( .B1(n16729), .B2(n15485), .A(n15481), .ZN(n15482) );
  MUX2_X1 U18831 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15482), .S(
        n15487), .Z(P1_U3473) );
  INV_X1 U18832 ( .A(n15483), .ZN(n15486) );
  OAI22_X1 U18833 ( .A1(n15486), .A2(n15485), .B1(n15484), .B2(n16754), .ZN(
        n15488) );
  MUX2_X1 U18834 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15488), .S(
        n15487), .Z(P1_U3469) );
  INV_X1 U18835 ( .A(n15489), .ZN(n15493) );
  NAND2_X1 U18836 ( .A1(n15490), .A2(n15491), .ZN(n15492) );
  AOI22_X1 U18837 ( .A1(n19315), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19360), .ZN(n15494) );
  OAI21_X1 U18838 ( .B1(n19375), .B2(n16033), .A(n15494), .ZN(n15500) );
  NAND2_X1 U18839 ( .A1(n15495), .A2(n15496), .ZN(n15497) );
  NAND2_X1 U18840 ( .A1(n15498), .A2(n15497), .ZN(n16308) );
  NOR2_X1 U18841 ( .A1(n16308), .A2(n19368), .ZN(n15499) );
  AOI211_X1 U18842 ( .C1(n16722), .C2(n15501), .A(n15500), .B(n15499), .ZN(
        n15506) );
  AOI21_X1 U18843 ( .B1(n15502), .B2(n16035), .A(n19364), .ZN(n15504) );
  OAI21_X1 U18844 ( .B1(n19320), .B2(n15504), .A(n15503), .ZN(n15505) );
  OAI211_X1 U18845 ( .C1(n19366), .C2(n16300), .A(n15506), .B(n15505), .ZN(
        P2_U2826) );
  NAND2_X1 U18846 ( .A1(n9828), .A2(n15507), .ZN(n15508) );
  NAND2_X1 U18847 ( .A1(n15490), .A2(n15508), .ZN(n15922) );
  INV_X1 U18848 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20157) );
  NAND2_X1 U18849 ( .A1(n19337), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15510) );
  NAND2_X1 U18850 ( .A1(n19360), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15509) );
  OAI211_X1 U18851 ( .C1(n19355), .C2(n20157), .A(n15510), .B(n15509), .ZN(
        n15514) );
  OR2_X1 U18852 ( .A1(n14530), .A2(n15511), .ZN(n15512) );
  NAND2_X1 U18853 ( .A1(n15495), .A2(n15512), .ZN(n16321) );
  NOR2_X1 U18854 ( .A1(n16321), .A2(n19368), .ZN(n15513) );
  AOI211_X1 U18855 ( .C1(n16722), .C2(n15515), .A(n15514), .B(n15513), .ZN(
        n15520) );
  INV_X1 U18856 ( .A(n15516), .ZN(n15528) );
  INV_X1 U18857 ( .A(n16041), .ZN(n15517) );
  AOI21_X1 U18858 ( .B1(n15528), .B2(n15517), .A(n19364), .ZN(n15518) );
  OAI21_X1 U18859 ( .B1(n15518), .B2(n19320), .A(n15502), .ZN(n15519) );
  OAI211_X1 U18860 ( .C1(n19366), .C2(n15922), .A(n15520), .B(n15519), .ZN(
        P2_U2827) );
  INV_X1 U18861 ( .A(n15521), .ZN(n16332) );
  INV_X1 U18862 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20156) );
  NAND2_X1 U18863 ( .A1(n19360), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15522) );
  OAI21_X1 U18864 ( .B1(n19355), .B2(n20156), .A(n15522), .ZN(n15523) );
  AOI21_X1 U18865 ( .B1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19337), .A(
        n15523), .ZN(n15524) );
  OAI21_X1 U18866 ( .B1(n15525), .B2(n19356), .A(n15524), .ZN(n15526) );
  AOI21_X1 U18867 ( .B1(n16332), .B2(n19324), .A(n15526), .ZN(n15531) );
  AOI21_X1 U18868 ( .B1(n15527), .B2(n16052), .A(n19364), .ZN(n15529) );
  OAI21_X1 U18869 ( .B1(n19320), .B2(n15529), .A(n15528), .ZN(n15530) );
  OAI211_X1 U18870 ( .C1(n19366), .C2(n16325), .A(n15531), .B(n15530), .ZN(
        P2_U2828) );
  OR2_X1 U18871 ( .A1(n11726), .A2(n15532), .ZN(n15533) );
  NAND2_X1 U18872 ( .A1(n14524), .A2(n15533), .ZN(n16339) );
  AND2_X1 U18873 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  OR2_X1 U18874 ( .A1(n15536), .A2(n14531), .ZN(n16349) );
  INV_X1 U18875 ( .A(n16349), .ZN(n15547) );
  OAI211_X1 U18876 ( .C1(n15538), .C2(n15839), .A(n15537), .B(n16722), .ZN(
        n15540) );
  AOI22_X1 U18877 ( .A1(n19315), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19360), .ZN(n15539) );
  OAI211_X1 U18878 ( .C1(n19375), .C2(n15541), .A(n15540), .B(n15539), .ZN(
        n15546) );
  OAI21_X1 U18879 ( .B1(n15542), .B2(n16070), .A(n19344), .ZN(n15544) );
  INV_X1 U18880 ( .A(n15527), .ZN(n15543) );
  AOI21_X1 U18881 ( .B1(n16718), .B2(n15544), .A(n15543), .ZN(n15545) );
  AOI211_X1 U18882 ( .C1(n19324), .C2(n15547), .A(n15546), .B(n15545), .ZN(
        n15548) );
  OAI21_X1 U18883 ( .B1(n16339), .B2(n19366), .A(n15548), .ZN(P2_U2829) );
  INV_X1 U18884 ( .A(n16078), .ZN(n15558) );
  AOI21_X1 U18885 ( .B1(n15549), .B2(n16076), .A(n19364), .ZN(n15551) );
  INV_X1 U18886 ( .A(n15542), .ZN(n15550) );
  OAI21_X1 U18887 ( .B1(n19320), .B2(n15551), .A(n15550), .ZN(n15555) );
  INV_X1 U18888 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20151) );
  OAI22_X1 U18889 ( .A1(n19354), .A2(n15552), .B1(n19355), .B2(n20151), .ZN(
        n15553) );
  AOI21_X1 U18890 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19337), .A(
        n15553), .ZN(n15554) );
  OAI211_X1 U18891 ( .C1(n19356), .C2(n15556), .A(n15555), .B(n15554), .ZN(
        n15557) );
  AOI21_X1 U18892 ( .B1(n15558), .B2(n19324), .A(n15557), .ZN(n15559) );
  OAI21_X1 U18893 ( .B1(n15944), .B2(n19366), .A(n15559), .ZN(P2_U2830) );
  AND2_X1 U18894 ( .A1(n15862), .A2(n15576), .ZN(n15578) );
  OR2_X1 U18895 ( .A1(n15578), .A2(n15560), .ZN(n15561) );
  NAND2_X1 U18896 ( .A1(n15562), .A2(n15561), .ZN(n16362) );
  XOR2_X1 U18897 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n15563), .Z(n15570) );
  AOI22_X1 U18898 ( .A1(n19315), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19360), .ZN(n15564) );
  OAI21_X1 U18899 ( .B1(n19375), .B2(n15565), .A(n15564), .ZN(n15569) );
  OAI21_X1 U18900 ( .B1(n15582), .B2(n16089), .A(n19344), .ZN(n15567) );
  INV_X1 U18901 ( .A(n15549), .ZN(n15566) );
  AOI21_X1 U18902 ( .B1(n16718), .B2(n15567), .A(n15566), .ZN(n15568) );
  AOI211_X1 U18903 ( .C1(n16722), .C2(n15570), .A(n15569), .B(n15568), .ZN(
        n15575) );
  OR2_X1 U18904 ( .A1(n15571), .A2(n15587), .ZN(n15589) );
  AND2_X1 U18905 ( .A1(n15589), .A2(n15572), .ZN(n15573) );
  NOR2_X1 U18906 ( .A1(n11570), .A2(n15573), .ZN(n16359) );
  NAND2_X1 U18907 ( .A1(n16359), .A2(n19322), .ZN(n15574) );
  OAI211_X1 U18908 ( .C1(n19368), .C2(n16362), .A(n15575), .B(n15574), .ZN(
        P2_U2831) );
  NOR2_X1 U18909 ( .A1(n15862), .A2(n15576), .ZN(n15577) );
  AOI22_X1 U18910 ( .A1(n19315), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19360), .ZN(n15579) );
  OAI21_X1 U18911 ( .B1(n19375), .B2(n16096), .A(n15579), .ZN(n15585) );
  INV_X1 U18912 ( .A(n15580), .ZN(n16716) );
  INV_X1 U18913 ( .A(n16098), .ZN(n15581) );
  OAI21_X1 U18914 ( .B1(n16716), .B2(n15581), .A(n19344), .ZN(n15583) );
  AOI21_X1 U18915 ( .B1(n16718), .B2(n15583), .A(n15582), .ZN(n15584) );
  AOI211_X1 U18916 ( .C1(n16722), .C2(n15586), .A(n15585), .B(n15584), .ZN(
        n15591) );
  NAND2_X1 U18917 ( .A1(n15571), .A2(n15587), .ZN(n15588) );
  NAND2_X1 U18918 ( .A1(n16375), .A2(n19322), .ZN(n15590) );
  OAI211_X1 U18919 ( .C1(n19368), .C2(n16372), .A(n15591), .B(n15590), .ZN(
        P2_U2832) );
  NAND2_X1 U18920 ( .A1(n9853), .A2(n15592), .ZN(n15593) );
  NAND2_X1 U18921 ( .A1(n12440), .A2(n15593), .ZN(n16402) );
  AOI21_X1 U18922 ( .B1(n15594), .B2(n12453), .A(n11847), .ZN(n16400) );
  XNOR2_X1 U18923 ( .A(n15595), .B(n16116), .ZN(n15601) );
  INV_X1 U18924 ( .A(n15596), .ZN(n15599) );
  NOR2_X1 U18925 ( .A1(n19375), .A2(n11661), .ZN(n15598) );
  INV_X1 U18926 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20143) );
  OAI22_X1 U18927 ( .A1(n19354), .A2(n15877), .B1(n19355), .B2(n20143), .ZN(
        n15597) );
  AOI211_X1 U18928 ( .C1(n15599), .C2(n16722), .A(n15598), .B(n15597), .ZN(
        n15600) );
  OAI21_X1 U18929 ( .B1(n15601), .B2(n19364), .A(n15600), .ZN(n15602) );
  AOI21_X1 U18930 ( .B1(n16400), .B2(n19324), .A(n15602), .ZN(n15603) );
  OAI21_X1 U18931 ( .B1(n16402), .B2(n19366), .A(n15603), .ZN(P2_U2835) );
  INV_X1 U18932 ( .A(n16411), .ZN(n15616) );
  NOR2_X1 U18933 ( .A1(n15742), .A2(n15604), .ZN(n15606) );
  XNOR2_X1 U18934 ( .A(n15606), .B(n15605), .ZN(n15612) );
  INV_X1 U18935 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20141) );
  INV_X1 U18936 ( .A(n19354), .ZN(n19360) );
  AOI21_X1 U18937 ( .B1(n19360), .B2(P2_EBX_REG_19__SCAN_IN), .A(n19359), .ZN(
        n15607) );
  OAI21_X1 U18938 ( .B1(n19355), .B2(n20141), .A(n15607), .ZN(n15608) );
  AOI21_X1 U18939 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19337), .A(
        n15608), .ZN(n15609) );
  OAI21_X1 U18940 ( .B1(n15610), .B2(n19356), .A(n15609), .ZN(n15611) );
  AOI21_X1 U18941 ( .B1(n15612), .B2(n19344), .A(n15611), .ZN(n15615) );
  XNOR2_X1 U18942 ( .A(n15613), .B(n9895), .ZN(n16412) );
  NAND2_X1 U18943 ( .A1(n16412), .A2(n19322), .ZN(n15614) );
  OAI211_X1 U18944 ( .C1(n15616), .C2(n19368), .A(n15615), .B(n15614), .ZN(
        P2_U2836) );
  INV_X1 U18945 ( .A(n15613), .ZN(n15620) );
  NAND2_X1 U18946 ( .A1(n15617), .A2(n15618), .ZN(n15619) );
  NAND2_X1 U18947 ( .A1(n15620), .A2(n15619), .ZN(n16422) );
  INV_X1 U18948 ( .A(n15621), .ZN(n15622) );
  AOI21_X1 U18949 ( .B1(n15623), .B2(n15622), .A(n12454), .ZN(n16425) );
  NAND2_X1 U18950 ( .A1(n15624), .A2(n16722), .ZN(n15628) );
  OAI21_X1 U18951 ( .B1(n19354), .B2(n15625), .A(n19333), .ZN(n15626) );
  AOI21_X1 U18952 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n19315), .A(n15626), 
        .ZN(n15627) );
  OAI211_X1 U18953 ( .C1(n19375), .C2(n15629), .A(n15628), .B(n15627), .ZN(
        n15634) );
  INV_X1 U18954 ( .A(n15631), .ZN(n15630) );
  OAI21_X1 U18955 ( .B1(n19364), .B2(n15630), .A(n16718), .ZN(n15632) );
  NOR2_X1 U18956 ( .A1(n15816), .A2(n15631), .ZN(n19326) );
  MUX2_X1 U18957 ( .A(n15632), .B(n19326), .S(n16127), .Z(n15633) );
  AOI211_X1 U18958 ( .C1(n16425), .C2(n19324), .A(n15634), .B(n15633), .ZN(
        n15635) );
  OAI21_X1 U18959 ( .B1(n16422), .B2(n19366), .A(n15635), .ZN(P2_U2837) );
  INV_X1 U18960 ( .A(n19341), .ZN(n15636) );
  AOI21_X1 U18961 ( .B1(n19344), .B2(n15636), .A(n19320), .ZN(n15638) );
  NAND2_X1 U18962 ( .A1(n15787), .A2(n19341), .ZN(n15637) );
  MUX2_X1 U18963 ( .A(n15638), .B(n15637), .S(n19338), .Z(n15648) );
  NOR2_X1 U18964 ( .A1(n13808), .A2(n15640), .ZN(n15641) );
  OR2_X1 U18965 ( .A1(n15639), .A2(n15641), .ZN(n15909) );
  INV_X1 U18966 ( .A(n15909), .ZN(n16465) );
  NAND2_X1 U18967 ( .A1(n19360), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n15642) );
  OAI211_X1 U18968 ( .C1(n19355), .C2(n20134), .A(n19333), .B(n15642), .ZN(
        n15643) );
  AOI21_X1 U18969 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19337), .A(
        n15643), .ZN(n15644) );
  OAI21_X1 U18970 ( .B1(n15645), .B2(n19356), .A(n15644), .ZN(n15646) );
  AOI21_X1 U18971 ( .B1(n16465), .B2(n19324), .A(n15646), .ZN(n15647) );
  OAI211_X1 U18972 ( .C1(n19366), .C2(n16457), .A(n15648), .B(n15647), .ZN(
        P2_U2840) );
  NAND2_X1 U18973 ( .A1(n15787), .A2(n15649), .ZN(n15652) );
  INV_X1 U18974 ( .A(n15649), .ZN(n15650) );
  AOI21_X1 U18975 ( .B1(n19344), .B2(n15650), .A(n19320), .ZN(n15651) );
  MUX2_X1 U18976 ( .A(n15652), .B(n15651), .S(n16162), .Z(n15660) );
  INV_X1 U18977 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20132) );
  NAND2_X1 U18978 ( .A1(n19337), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15654) );
  AOI21_X1 U18979 ( .B1(n19360), .B2(P2_EBX_REG_14__SCAN_IN), .A(n19359), .ZN(
        n15653) );
  OAI211_X1 U18980 ( .C1(n19355), .C2(n20132), .A(n15654), .B(n15653), .ZN(
        n15655) );
  AOI21_X1 U18981 ( .B1(n15656), .B2(n16722), .A(n15655), .ZN(n15657) );
  OAI21_X1 U18982 ( .B1(n16470), .B2(n19368), .A(n15657), .ZN(n15658) );
  INV_X1 U18983 ( .A(n15658), .ZN(n15659) );
  OAI211_X1 U18984 ( .C1(n19366), .C2(n16475), .A(n15660), .B(n15659), .ZN(
        P2_U2841) );
  NOR2_X1 U18985 ( .A1(n15742), .A2(n15661), .ZN(n15662) );
  XOR2_X1 U18986 ( .A(n16175), .B(n15662), .Z(n15671) );
  INV_X1 U18987 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15665) );
  NAND2_X1 U18988 ( .A1(n19337), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15664) );
  AOI21_X1 U18989 ( .B1(n19360), .B2(P2_EBX_REG_13__SCAN_IN), .A(n19359), .ZN(
        n15663) );
  OAI211_X1 U18990 ( .C1(n19355), .C2(n15665), .A(n15664), .B(n15663), .ZN(
        n15666) );
  AOI21_X1 U18991 ( .B1(n15667), .B2(n16722), .A(n15666), .ZN(n15668) );
  OAI21_X1 U18992 ( .B1(n16485), .B2(n19368), .A(n15668), .ZN(n15669) );
  AOI21_X1 U18993 ( .B1(n16488), .B2(n19322), .A(n15669), .ZN(n15670) );
  OAI21_X1 U18994 ( .B1(n15671), .B2(n19364), .A(n15670), .ZN(P2_U2842) );
  INV_X1 U18995 ( .A(n15672), .ZN(n15673) );
  NAND2_X1 U18996 ( .A1(n11664), .A2(n15673), .ZN(n15689) );
  XOR2_X1 U18997 ( .A(n15689), .B(n16185), .Z(n15682) );
  NAND2_X1 U18998 ( .A1(n16500), .A2(n19324), .ZN(n15680) );
  INV_X1 U18999 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20129) );
  OAI22_X1 U19000 ( .A1(n15675), .A2(n19356), .B1(n15674), .B2(n19375), .ZN(
        n15676) );
  INV_X1 U19001 ( .A(n15676), .ZN(n15677) );
  OAI211_X1 U19002 ( .C1(n20129), .C2(n19355), .A(n15677), .B(n19333), .ZN(
        n15678) );
  AOI21_X1 U19003 ( .B1(n19360), .B2(P2_EBX_REG_12__SCAN_IN), .A(n15678), .ZN(
        n15679) );
  OAI211_X1 U19004 ( .C1(n16497), .C2(n19366), .A(n15680), .B(n15679), .ZN(
        n15681) );
  AOI21_X1 U19005 ( .B1(n15682), .B2(n19344), .A(n15681), .ZN(n15683) );
  INV_X1 U19006 ( .A(n15683), .ZN(P2_U2843) );
  INV_X1 U19007 ( .A(n16190), .ZN(n15695) );
  INV_X1 U19008 ( .A(n16513), .ZN(n15693) );
  INV_X1 U19009 ( .A(n16509), .ZN(n15688) );
  AOI22_X1 U19010 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19337), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19360), .ZN(n15684) );
  OAI211_X1 U19011 ( .C1(n19355), .C2(n20127), .A(n15684), .B(n19333), .ZN(
        n15685) );
  AOI21_X1 U19012 ( .B1(n15686), .B2(n16722), .A(n15685), .ZN(n15687) );
  OAI21_X1 U19013 ( .B1(n15688), .B2(n19368), .A(n15687), .ZN(n15692) );
  AOI211_X1 U19014 ( .C1(n16190), .C2(n15690), .A(n19364), .B(n15689), .ZN(
        n15691) );
  AOI211_X1 U19015 ( .C1(n19322), .C2(n15693), .A(n15692), .B(n15691), .ZN(
        n15694) );
  OAI21_X1 U19016 ( .B1(n15695), .B2(n16718), .A(n15694), .ZN(P2_U2844) );
  NAND2_X1 U19017 ( .A1(n15787), .A2(n15696), .ZN(n15699) );
  INV_X1 U19018 ( .A(n15696), .ZN(n15697) );
  AOI21_X1 U19019 ( .B1(n19344), .B2(n15697), .A(n19320), .ZN(n15698) );
  MUX2_X1 U19020 ( .A(n15699), .B(n15698), .S(n16209), .Z(n15707) );
  INV_X1 U19021 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20125) );
  INV_X1 U19022 ( .A(n15700), .ZN(n15701) );
  AOI22_X1 U19023 ( .A1(P2_EBX_REG_10__SCAN_IN), .A2(n19360), .B1(n15701), 
        .B2(n16722), .ZN(n15702) );
  OAI211_X1 U19024 ( .C1(n20125), .C2(n19355), .A(n15702), .B(n19333), .ZN(
        n15703) );
  AOI21_X1 U19025 ( .B1(n19337), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15703), .ZN(n15704) );
  OAI21_X1 U19026 ( .B1(n16524), .B2(n19368), .A(n15704), .ZN(n15705) );
  INV_X1 U19027 ( .A(n15705), .ZN(n15706) );
  OAI211_X1 U19028 ( .C1(n16520), .C2(n19366), .A(n15707), .B(n15706), .ZN(
        P2_U2845) );
  NOR2_X1 U19029 ( .A1(n15742), .A2(n15708), .ZN(n15709) );
  XNOR2_X1 U19030 ( .A(n15709), .B(n16218), .ZN(n15716) );
  NOR2_X1 U19031 ( .A1(n16540), .A2(n19366), .ZN(n15715) );
  AOI22_X1 U19032 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19315), .B1(n16722), 
        .B2(n15710), .ZN(n15711) );
  OAI211_X1 U19033 ( .C1(n11092), .C2(n19354), .A(n15711), .B(n19333), .ZN(
        n15712) );
  AOI21_X1 U19034 ( .B1(n19337), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n15712), .ZN(n15713) );
  OAI21_X1 U19035 ( .B1(n16531), .B2(n19368), .A(n15713), .ZN(n15714) );
  AOI211_X1 U19036 ( .C1(n15716), .C2(n19344), .A(n15715), .B(n15714), .ZN(
        n15717) );
  INV_X1 U19037 ( .A(n15717), .ZN(P2_U2846) );
  NAND2_X1 U19038 ( .A1(n15787), .A2(n15718), .ZN(n15721) );
  INV_X1 U19039 ( .A(n15718), .ZN(n15719) );
  AOI21_X1 U19040 ( .B1(n19344), .B2(n15719), .A(n19320), .ZN(n15720) );
  MUX2_X1 U19041 ( .A(n15721), .B(n15720), .S(n16234), .Z(n15729) );
  INV_X1 U19042 ( .A(n16551), .ZN(n15727) );
  INV_X1 U19043 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20121) );
  NAND2_X1 U19044 ( .A1(n19360), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15722) );
  OAI211_X1 U19045 ( .C1(n19355), .C2(n20121), .A(n19333), .B(n15722), .ZN(
        n15723) );
  AOI21_X1 U19046 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19337), .A(
        n15723), .ZN(n15724) );
  OAI21_X1 U19047 ( .B1(n15725), .B2(n19356), .A(n15724), .ZN(n15726) );
  AOI21_X1 U19048 ( .B1(n15727), .B2(n19324), .A(n15726), .ZN(n15728) );
  OAI211_X1 U19049 ( .C1(n16559), .C2(n19366), .A(n15729), .B(n15728), .ZN(
        P2_U2847) );
  NAND2_X1 U19050 ( .A1(n15787), .A2(n15730), .ZN(n15732) );
  INV_X1 U19051 ( .A(n15730), .ZN(n19365) );
  AOI21_X1 U19052 ( .B1(n19344), .B2(n19365), .A(n19320), .ZN(n15731) );
  MUX2_X1 U19053 ( .A(n15732), .B(n15731), .S(n16252), .Z(n15740) );
  INV_X1 U19054 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20119) );
  OAI22_X1 U19055 ( .A1(n15733), .A2(n19356), .B1(n16250), .B2(n19375), .ZN(
        n15734) );
  INV_X1 U19056 ( .A(n15734), .ZN(n15735) );
  OAI211_X1 U19057 ( .C1(n20119), .C2(n19355), .A(n15735), .B(n19333), .ZN(
        n15736) );
  AOI21_X1 U19058 ( .B1(n19360), .B2(P2_EBX_REG_7__SCAN_IN), .A(n15736), .ZN(
        n15737) );
  OAI21_X1 U19059 ( .B1(n16566), .B2(n19368), .A(n15737), .ZN(n15738) );
  INV_X1 U19060 ( .A(n15738), .ZN(n15739) );
  OAI211_X1 U19061 ( .C1(n16572), .C2(n19366), .A(n15740), .B(n15739), .ZN(
        P2_U2848) );
  NOR2_X1 U19062 ( .A1(n15742), .A2(n15741), .ZN(n15743) );
  XNOR2_X1 U19063 ( .A(n15743), .B(n16271), .ZN(n15754) );
  XNOR2_X1 U19064 ( .A(n15744), .B(n15745), .ZN(n16589) );
  NOR2_X1 U19065 ( .A1(n16589), .A2(n19366), .ZN(n15753) );
  INV_X1 U19066 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15747) );
  NAND2_X1 U19067 ( .A1(n19360), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n15746) );
  OAI211_X1 U19068 ( .C1(n19355), .C2(n15747), .A(n19333), .B(n15746), .ZN(
        n15748) );
  AOI21_X1 U19069 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19337), .A(
        n15748), .ZN(n15751) );
  NAND2_X1 U19070 ( .A1(n15749), .A2(n16722), .ZN(n15750) );
  OAI211_X1 U19071 ( .C1(n16597), .C2(n19368), .A(n15751), .B(n15750), .ZN(
        n15752) );
  AOI211_X1 U19072 ( .C1(n15754), .C2(n19344), .A(n15753), .B(n15752), .ZN(
        n15755) );
  INV_X1 U19073 ( .A(n15755), .ZN(P2_U2850) );
  NAND2_X1 U19074 ( .A1(n15756), .A2(n15757), .ZN(n15758) );
  AND2_X1 U19075 ( .A1(n15744), .A2(n15758), .ZN(n19376) );
  INV_X1 U19076 ( .A(n16276), .ZN(n15762) );
  INV_X1 U19077 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n21249) );
  NAND2_X1 U19078 ( .A1(n19360), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n15760) );
  AOI22_X1 U19079 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19337), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19315), .ZN(n15759) );
  NAND3_X1 U19080 ( .A1(n15760), .A2(n15759), .A3(n19333), .ZN(n15761) );
  AOI21_X1 U19081 ( .B1(n15762), .B2(n16722), .A(n15761), .ZN(n15763) );
  OAI21_X1 U19082 ( .B1(n16607), .B2(n19368), .A(n15763), .ZN(n15769) );
  INV_X1 U19083 ( .A(n15765), .ZN(n15764) );
  NOR2_X1 U19084 ( .A1(n15816), .A2(n15764), .ZN(n15767) );
  OAI21_X1 U19085 ( .B1(n19364), .B2(n15765), .A(n16718), .ZN(n15766) );
  MUX2_X1 U19086 ( .A(n15767), .B(n15766), .S(n16285), .Z(n15768) );
  AOI211_X1 U19087 ( .C1(n19376), .C2(n19322), .A(n15769), .B(n15768), .ZN(
        n15770) );
  OAI21_X1 U19088 ( .B1(n19378), .B2(n15810), .A(n15770), .ZN(P2_U2851) );
  NAND2_X1 U19089 ( .A1(n15773), .A2(n15772), .ZN(n15774) );
  NAND2_X1 U19090 ( .A1(n15756), .A2(n15774), .ZN(n16021) );
  NOR2_X1 U19091 ( .A1(n15775), .A2(n19356), .ZN(n15777) );
  INV_X1 U19092 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20112) );
  OAI22_X1 U19093 ( .A1(n19354), .A2(n11032), .B1(n19355), .B2(n20112), .ZN(
        n15776) );
  AOI211_X1 U19094 ( .C1(n19337), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15777), .B(n15776), .ZN(n15778) );
  OAI21_X1 U19095 ( .B1(n16021), .B2(n19366), .A(n15778), .ZN(n15784) );
  INV_X1 U19096 ( .A(n15780), .ZN(n15779) );
  OAI21_X1 U19097 ( .B1(n19364), .B2(n15779), .A(n16718), .ZN(n15782) );
  NOR2_X1 U19098 ( .A1(n15816), .A2(n15780), .ZN(n15781) );
  MUX2_X1 U19099 ( .A(n15782), .B(n15781), .S(n16293), .Z(n15783) );
  AOI211_X1 U19100 ( .C1(n19324), .C2(n15771), .A(n15784), .B(n15783), .ZN(
        n15785) );
  OAI21_X1 U19101 ( .B1(n19807), .B2(n15810), .A(n15785), .ZN(P2_U2852) );
  AOI21_X1 U19102 ( .B1(n19344), .B2(n15798), .A(n19320), .ZN(n15789) );
  INV_X1 U19103 ( .A(n15798), .ZN(n15786) );
  NAND2_X1 U19104 ( .A1(n15787), .A2(n15786), .ZN(n15788) );
  MUX2_X1 U19105 ( .A(n15789), .B(n15788), .S(n19477), .Z(n15796) );
  NAND2_X1 U19106 ( .A1(n20194), .A2(n19322), .ZN(n15792) );
  INV_X1 U19107 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20110) );
  OAI22_X1 U19108 ( .A1(n10595), .A2(n19354), .B1(n20110), .B2(n19355), .ZN(
        n15790) );
  AOI21_X1 U19109 ( .B1(n19337), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15790), .ZN(n15791) );
  OAI211_X1 U19110 ( .C1(n15793), .C2(n19356), .A(n15792), .B(n15791), .ZN(
        n15794) );
  AOI21_X1 U19111 ( .B1(n19479), .B2(n19324), .A(n15794), .ZN(n15795) );
  OAI211_X1 U19112 ( .C1(n15810), .C2(n20190), .A(n15796), .B(n15795), .ZN(
        P2_U2853) );
  NOR2_X1 U19113 ( .A1(n15798), .A2(n10668), .ZN(n15799) );
  NAND2_X1 U19114 ( .A1(n11664), .A2(n15799), .ZN(n16653) );
  MUX2_X1 U19115 ( .A(n16718), .B(n19375), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15806) );
  INV_X1 U19116 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20108) );
  AOI22_X1 U19117 ( .A1(n16722), .A2(n15800), .B1(P2_EBX_REG_1__SCAN_IN), .B2(
        n19360), .ZN(n15802) );
  NAND2_X1 U19118 ( .A1(n19322), .A2(n20203), .ZN(n15801) );
  OAI211_X1 U19119 ( .C1(n19355), .C2(n20108), .A(n15802), .B(n15801), .ZN(
        n15804) );
  NOR2_X1 U19120 ( .A1(n19502), .A2(n15810), .ZN(n15803) );
  AOI211_X1 U19121 ( .C1(n19324), .C2(n19494), .A(n15804), .B(n15803), .ZN(
        n15805) );
  OAI211_X1 U19122 ( .C1(n16653), .C2(n19364), .A(n15806), .B(n15805), .ZN(
        P2_U2854) );
  INV_X1 U19123 ( .A(n16647), .ZN(n15817) );
  OAI21_X1 U19124 ( .B1(n19320), .B2(n19337), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15815) );
  AOI22_X1 U19125 ( .A1(n19322), .A2(n19400), .B1(P2_EBX_REG_0__SCAN_IN), .B2(
        n19360), .ZN(n15808) );
  NAND2_X1 U19126 ( .A1(n19315), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n15807) );
  OAI211_X1 U19127 ( .C1(n19356), .C2(n15809), .A(n15808), .B(n15807), .ZN(
        n15812) );
  NOR2_X1 U19128 ( .A1(n19501), .A2(n15810), .ZN(n15811) );
  AOI211_X1 U19129 ( .C1(n19324), .C2(n15813), .A(n15812), .B(n15811), .ZN(
        n15814) );
  OAI211_X1 U19130 ( .C1(n15817), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        P2_U2855) );
  NAND2_X1 U19131 ( .A1(n9733), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15818) );
  OAI21_X1 U19132 ( .B1(n12574), .B2(n9733), .A(n15818), .ZN(P2_U2856) );
  OR2_X1 U19133 ( .A1(n15821), .A2(n15820), .ZN(n15914) );
  NAND3_X1 U19134 ( .A1(n15819), .A2(n15914), .A3(n15904), .ZN(n15823) );
  NAND2_X1 U19135 ( .A1(n9733), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15822) );
  OAI211_X1 U19136 ( .C1(n15824), .C2(n16308), .A(n15823), .B(n15822), .ZN(
        P2_U2858) );
  INV_X1 U19137 ( .A(n15825), .ZN(n15826) );
  NAND2_X1 U19138 ( .A1(n15827), .A2(n15826), .ZN(n15829) );
  XNOR2_X1 U19139 ( .A(n15829), .B(n15828), .ZN(n15929) );
  NOR2_X1 U19140 ( .A1(n16321), .A2(n9733), .ZN(n15830) );
  AOI21_X1 U19141 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n9733), .A(n15830), .ZN(
        n15831) );
  OAI21_X1 U19142 ( .B1(n15929), .B2(n15897), .A(n15831), .ZN(P2_U2859) );
  NOR2_X1 U19143 ( .A1(n15832), .A2(n15842), .ZN(n15841) );
  NOR2_X1 U19144 ( .A1(n15841), .A2(n15833), .ZN(n15838) );
  NOR2_X1 U19145 ( .A1(n13063), .A2(n15834), .ZN(n15835) );
  XNOR2_X1 U19146 ( .A(n15836), .B(n15835), .ZN(n15837) );
  XNOR2_X1 U19147 ( .A(n15838), .B(n15837), .ZN(n15936) );
  MUX2_X1 U19148 ( .A(n16349), .B(n15839), .S(n9733), .Z(n15840) );
  OAI21_X1 U19149 ( .B1(n15936), .B2(n15897), .A(n15840), .ZN(P2_U2861) );
  AOI21_X1 U19150 ( .B1(n15832), .B2(n15842), .A(n15841), .ZN(n15937) );
  NAND2_X1 U19151 ( .A1(n15937), .A2(n15904), .ZN(n15844) );
  NAND2_X1 U19152 ( .A1(n9733), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15843) );
  OAI211_X1 U19153 ( .C1(n16078), .C2(n9733), .A(n15844), .B(n15843), .ZN(
        P2_U2862) );
  INV_X1 U19154 ( .A(n15845), .ZN(n15860) );
  XNOR2_X1 U19155 ( .A(n15845), .B(n15847), .ZN(n15856) );
  NOR2_X1 U19156 ( .A1(n13063), .A2(n15846), .ZN(n15855) );
  NAND2_X1 U19157 ( .A1(n15856), .A2(n15855), .ZN(n15854) );
  OAI21_X1 U19158 ( .B1(n15847), .B2(n15860), .A(n15854), .ZN(n15851) );
  XOR2_X1 U19159 ( .A(n15849), .B(n15848), .Z(n15850) );
  XNOR2_X1 U19160 ( .A(n15851), .B(n15850), .ZN(n15951) );
  NOR2_X1 U19161 ( .A1(n16362), .A2(n9733), .ZN(n15852) );
  AOI21_X1 U19162 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n9733), .A(n15852), .ZN(
        n15853) );
  OAI21_X1 U19163 ( .B1(n15951), .B2(n15897), .A(n15853), .ZN(P2_U2863) );
  OAI21_X1 U19164 ( .B1(n15856), .B2(n15855), .A(n15854), .ZN(n15957) );
  NOR2_X1 U19165 ( .A1(n16372), .A2(n9733), .ZN(n15857) );
  AOI21_X1 U19166 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n9733), .A(n15857), .ZN(
        n15858) );
  OAI21_X1 U19167 ( .B1(n15957), .B2(n15897), .A(n15858), .ZN(P2_U2864) );
  OAI21_X1 U19168 ( .B1(n15859), .B2(n15861), .A(n15860), .ZN(n15967) );
  INV_X1 U19169 ( .A(n15862), .ZN(n15865) );
  NAND2_X1 U19170 ( .A1(n11697), .A2(n15863), .ZN(n15864) );
  NAND2_X1 U19171 ( .A1(n15865), .A2(n15864), .ZN(n16710) );
  NOR2_X1 U19172 ( .A1(n16710), .A2(n9733), .ZN(n15866) );
  AOI21_X1 U19173 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n9733), .A(n15866), .ZN(
        n15867) );
  OAI21_X1 U19174 ( .B1(n15897), .B2(n15967), .A(n15867), .ZN(P2_U2865) );
  INV_X1 U19175 ( .A(n15859), .ZN(n15869) );
  OAI21_X1 U19176 ( .B1(n15868), .B2(n15870), .A(n15869), .ZN(n15972) );
  NOR2_X1 U19177 ( .A1(n19311), .A2(n9733), .ZN(n15871) );
  AOI21_X1 U19178 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n9733), .A(n15871), .ZN(
        n15872) );
  OAI21_X1 U19179 ( .B1(n15972), .B2(n15897), .A(n15872), .ZN(P2_U2866) );
  AOI21_X1 U19180 ( .B1(n15874), .B2(n15879), .A(n15868), .ZN(n15973) );
  NAND2_X1 U19181 ( .A1(n15973), .A2(n15904), .ZN(n15876) );
  NAND2_X1 U19182 ( .A1(n16400), .A2(n15887), .ZN(n15875) );
  OAI211_X1 U19183 ( .C1(n15887), .C2(n15877), .A(n15876), .B(n15875), .ZN(
        P2_U2867) );
  OAI21_X1 U19184 ( .B1(n15878), .B2(n15880), .A(n15879), .ZN(n15984) );
  NAND2_X1 U19185 ( .A1(n9733), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15882) );
  NAND2_X1 U19186 ( .A1(n16411), .A2(n15887), .ZN(n15881) );
  OAI211_X1 U19187 ( .C1(n15984), .C2(n15897), .A(n15882), .B(n15881), .ZN(
        P2_U2868) );
  INV_X1 U19188 ( .A(n15890), .ZN(n15886) );
  OAI21_X1 U19189 ( .B1(n15886), .B2(n15885), .A(n15884), .ZN(n15992) );
  NAND2_X1 U19190 ( .A1(n16425), .A2(n15887), .ZN(n15889) );
  NAND2_X1 U19191 ( .A1(n9733), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15888) );
  OAI211_X1 U19192 ( .C1(n15992), .C2(n15897), .A(n15889), .B(n15888), .ZN(
        P2_U2869) );
  OAI21_X1 U19193 ( .B1(n9813), .B2(n15891), .A(n15890), .ZN(n16001) );
  NAND2_X1 U19194 ( .A1(n15892), .A2(n15893), .ZN(n15894) );
  NAND2_X1 U19195 ( .A1(n15622), .A2(n15894), .ZN(n19321) );
  NOR2_X1 U19196 ( .A1(n19321), .A2(n9733), .ZN(n15895) );
  AOI21_X1 U19197 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n9733), .A(n15895), .ZN(
        n15896) );
  OAI21_X1 U19198 ( .B1(n15897), .B2(n16001), .A(n15896), .ZN(P2_U2870) );
  OR2_X1 U19199 ( .A1(n15639), .A2(n15898), .ZN(n15899) );
  NAND2_X1 U19200 ( .A1(n15892), .A2(n15899), .ZN(n19346) );
  INV_X1 U19201 ( .A(n15900), .ZN(n15901) );
  AOI21_X1 U19202 ( .B1(n15901), .B2(n9752), .A(n9813), .ZN(n16005) );
  NAND2_X1 U19203 ( .A1(n16005), .A2(n15904), .ZN(n15903) );
  NAND2_X1 U19204 ( .A1(n9733), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15902) );
  OAI211_X1 U19205 ( .C1(n19346), .C2(n9733), .A(n15903), .B(n15902), .ZN(
        P2_U2871) );
  INV_X1 U19206 ( .A(n13811), .ZN(n15906) );
  OAI211_X1 U19207 ( .C1(n15906), .C2(n15905), .A(n9752), .B(n15904), .ZN(
        n15908) );
  NAND2_X1 U19208 ( .A1(n9733), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n15907) );
  OAI211_X1 U19209 ( .C1(n15909), .C2(n9733), .A(n15908), .B(n15907), .ZN(
        P2_U2872) );
  INV_X1 U19210 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n15913) );
  NAND2_X1 U19211 ( .A1(n15910), .A2(n19397), .ZN(n15912) );
  AOI22_X1 U19212 ( .A1(n16011), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19396), .ZN(n15911) );
  OAI211_X1 U19213 ( .C1(n16007), .C2(n15913), .A(n15912), .B(n15911), .ZN(
        P2_U2888) );
  NAND3_X1 U19214 ( .A1(n15819), .A2(n15914), .A3(n19398), .ZN(n15921) );
  INV_X1 U19215 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n15917) );
  AOI22_X1 U19216 ( .A1(n15985), .A2(n15915), .B1(n19396), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15916) );
  OAI21_X1 U19217 ( .B1(n16007), .B2(n15917), .A(n15916), .ZN(n15919) );
  NOR2_X1 U19218 ( .A1(n16300), .A2(n16014), .ZN(n15918) );
  AOI211_X1 U19219 ( .C1(n16011), .C2(BUF1_REG_29__SCAN_IN), .A(n15919), .B(
        n15918), .ZN(n15920) );
  NAND2_X1 U19220 ( .A1(n15921), .A2(n15920), .ZN(P2_U2890) );
  INV_X1 U19221 ( .A(n15922), .ZN(n16322) );
  INV_X1 U19222 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n15926) );
  NAND2_X1 U19223 ( .A1(n16011), .A2(BUF1_REG_28__SCAN_IN), .ZN(n15925) );
  AOI22_X1 U19224 ( .A1(n15985), .A2(n15923), .B1(n19396), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15924) );
  OAI211_X1 U19225 ( .C1(n16007), .C2(n15926), .A(n15925), .B(n15924), .ZN(
        n15927) );
  AOI21_X1 U19226 ( .B1(n16322), .B2(n19397), .A(n15927), .ZN(n15928) );
  OAI21_X1 U19227 ( .B1(n15929), .B2(n16023), .A(n15928), .ZN(P2_U2891) );
  INV_X1 U19228 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n15932) );
  AOI22_X1 U19229 ( .A1(n15985), .A2(n15930), .B1(n19396), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15931) );
  OAI21_X1 U19230 ( .B1(n16007), .B2(n15932), .A(n15931), .ZN(n15934) );
  NOR2_X1 U19231 ( .A1(n16339), .A2(n16014), .ZN(n15933) );
  AOI211_X1 U19232 ( .C1(n16011), .C2(BUF1_REG_26__SCAN_IN), .A(n15934), .B(
        n15933), .ZN(n15935) );
  OAI21_X1 U19233 ( .B1(n15936), .B2(n16023), .A(n15935), .ZN(P2_U2893) );
  NAND2_X1 U19234 ( .A1(n15937), .A2(n19398), .ZN(n15943) );
  INV_X1 U19235 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n15940) );
  AOI22_X1 U19236 ( .A1(n15985), .A2(n15938), .B1(n19396), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15939) );
  OAI21_X1 U19237 ( .B1(n16007), .B2(n15940), .A(n15939), .ZN(n15941) );
  AOI21_X1 U19238 ( .B1(n16011), .B2(BUF1_REG_25__SCAN_IN), .A(n15941), .ZN(
        n15942) );
  OAI211_X1 U19239 ( .C1(n15944), .C2(n16014), .A(n15943), .B(n15942), .ZN(
        P2_U2894) );
  INV_X1 U19240 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n15948) );
  NAND2_X1 U19241 ( .A1(n16011), .A2(BUF1_REG_24__SCAN_IN), .ZN(n15947) );
  AOI22_X1 U19242 ( .A1(n15985), .A2(n15945), .B1(n19396), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15946) );
  OAI211_X1 U19243 ( .C1(n16007), .C2(n15948), .A(n15947), .B(n15946), .ZN(
        n15949) );
  AOI21_X1 U19244 ( .B1(n16359), .B2(n19397), .A(n15949), .ZN(n15950) );
  OAI21_X1 U19245 ( .B1(n15951), .B2(n16023), .A(n15950), .ZN(P2_U2895) );
  INV_X1 U19246 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15954) );
  NAND2_X1 U19247 ( .A1(n16011), .A2(BUF1_REG_23__SCAN_IN), .ZN(n15953) );
  AOI22_X1 U19248 ( .A1(n15985), .A2(n19552), .B1(n19396), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15952) );
  OAI211_X1 U19249 ( .C1(n15954), .C2(n16007), .A(n15953), .B(n15952), .ZN(
        n15955) );
  AOI21_X1 U19250 ( .B1(n16375), .B2(n19397), .A(n15955), .ZN(n15956) );
  OAI21_X1 U19251 ( .B1(n15957), .B2(n16023), .A(n15956), .ZN(P2_U2896) );
  OR2_X1 U19252 ( .A1(n15959), .A2(n15958), .ZN(n15960) );
  NAND2_X1 U19253 ( .A1(n15571), .A2(n15960), .ZN(n16709) );
  INV_X1 U19254 ( .A(n16709), .ZN(n15965) );
  INV_X1 U19255 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n15963) );
  NAND2_X1 U19256 ( .A1(n16011), .A2(BUF1_REG_22__SCAN_IN), .ZN(n15962) );
  AOI22_X1 U19257 ( .A1(n15985), .A2(n19543), .B1(n19396), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15961) );
  OAI211_X1 U19258 ( .C1(n15963), .C2(n16007), .A(n15962), .B(n15961), .ZN(
        n15964) );
  AOI21_X1 U19259 ( .B1(n15965), .B2(n19397), .A(n15964), .ZN(n15966) );
  OAI21_X1 U19260 ( .B1(n15967), .B2(n16023), .A(n15966), .ZN(P2_U2897) );
  NAND2_X1 U19261 ( .A1(n16011), .A2(BUF1_REG_21__SCAN_IN), .ZN(n15969) );
  AOI22_X1 U19262 ( .A1(n15985), .A2(n19535), .B1(n19396), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15968) );
  OAI211_X1 U19263 ( .C1(n18635), .C2(n16007), .A(n15969), .B(n15968), .ZN(
        n15970) );
  AOI21_X1 U19264 ( .B1(n19305), .B2(n19397), .A(n15970), .ZN(n15971) );
  OAI21_X1 U19265 ( .B1(n15972), .B2(n16023), .A(n15971), .ZN(P2_U2898) );
  NAND2_X1 U19266 ( .A1(n15973), .A2(n19398), .ZN(n15978) );
  INV_X1 U19267 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n15974) );
  NOR2_X1 U19268 ( .A1(n16007), .A2(n15974), .ZN(n15976) );
  INV_X1 U19269 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19429) );
  OAI22_X1 U19270 ( .A1(n16008), .A2(n19382), .B1(n16017), .B2(n19429), .ZN(
        n15975) );
  AOI211_X1 U19271 ( .C1(n16011), .C2(BUF1_REG_20__SCAN_IN), .A(n15976), .B(
        n15975), .ZN(n15977) );
  OAI211_X1 U19272 ( .C1(n16402), .C2(n16014), .A(n15978), .B(n15977), .ZN(
        P2_U2899) );
  INV_X1 U19273 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15981) );
  INV_X1 U19274 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19431) );
  OAI22_X1 U19275 ( .A1(n16008), .A2(n19389), .B1(n16017), .B2(n19431), .ZN(
        n15979) );
  AOI21_X1 U19276 ( .B1(n16011), .B2(BUF1_REG_19__SCAN_IN), .A(n15979), .ZN(
        n15980) );
  OAI21_X1 U19277 ( .B1(n16007), .B2(n15981), .A(n15980), .ZN(n15982) );
  AOI21_X1 U19278 ( .B1(n16412), .B2(n19397), .A(n15982), .ZN(n15983) );
  OAI21_X1 U19279 ( .B1(n15984), .B2(n16023), .A(n15983), .ZN(P2_U2900) );
  INV_X1 U19280 ( .A(n16422), .ZN(n15990) );
  INV_X1 U19281 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U19282 ( .A1(n16011), .A2(BUF1_REG_18__SCAN_IN), .ZN(n15987) );
  AOI22_X1 U19283 ( .A1(n15985), .A2(n19520), .B1(n19396), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15986) );
  OAI211_X1 U19284 ( .C1(n15988), .C2(n16007), .A(n15987), .B(n15986), .ZN(
        n15989) );
  AOI21_X1 U19285 ( .B1(n15990), .B2(n19397), .A(n15989), .ZN(n15991) );
  OAI21_X1 U19286 ( .B1(n15992), .B2(n16023), .A(n15991), .ZN(P2_U2901) );
  INV_X1 U19287 ( .A(n15994), .ZN(n16004) );
  AOI21_X1 U19288 ( .B1(n15995), .B2(n16004), .A(n10512), .ZN(n19323) );
  INV_X1 U19289 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n15998) );
  INV_X1 U19290 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n21396) );
  OAI22_X1 U19291 ( .A1(n16008), .A2(n19395), .B1(n16017), .B2(n21396), .ZN(
        n15996) );
  AOI21_X1 U19292 ( .B1(n16011), .B2(BUF1_REG_17__SCAN_IN), .A(n15996), .ZN(
        n15997) );
  OAI21_X1 U19293 ( .B1(n16007), .B2(n15998), .A(n15997), .ZN(n15999) );
  AOI21_X1 U19294 ( .B1(n19323), .B2(n19397), .A(n15999), .ZN(n16000) );
  OAI21_X1 U19295 ( .B1(n16001), .B2(n16023), .A(n16000), .ZN(P2_U2902) );
  NAND2_X1 U19296 ( .A1(n13737), .A2(n16002), .ZN(n16003) );
  NAND2_X1 U19297 ( .A1(n16004), .A2(n16003), .ZN(n19349) );
  NAND2_X1 U19298 ( .A1(n16005), .A2(n19398), .ZN(n16013) );
  INV_X1 U19299 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n16006) );
  NOR2_X1 U19300 ( .A1(n16007), .A2(n16006), .ZN(n16010) );
  INV_X1 U19301 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19438) );
  OAI22_X1 U19302 ( .A1(n16008), .A2(n19404), .B1(n16017), .B2(n19438), .ZN(
        n16009) );
  AOI211_X1 U19303 ( .C1(n16011), .C2(BUF1_REG_16__SCAN_IN), .A(n16010), .B(
        n16009), .ZN(n16012) );
  OAI211_X1 U19304 ( .C1(n19349), .C2(n16014), .A(n16013), .B(n16012), .ZN(
        P2_U2903) );
  INV_X1 U19305 ( .A(n16589), .ZN(n16027) );
  INV_X1 U19306 ( .A(n16015), .ZN(n16026) );
  INV_X1 U19307 ( .A(n19535), .ZN(n16018) );
  INV_X1 U19308 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n16016) );
  OAI22_X1 U19309 ( .A1(n19403), .A2(n16018), .B1(n16017), .B2(n16016), .ZN(
        n16025) );
  INV_X1 U19310 ( .A(n20190), .ZN(n16020) );
  OAI21_X1 U19311 ( .B1(n16020), .B2(n20194), .A(n16019), .ZN(n19384) );
  INV_X1 U19312 ( .A(n16021), .ZN(n20182) );
  XNOR2_X1 U19313 ( .A(n19807), .B(n20182), .ZN(n19385) );
  NAND2_X1 U19314 ( .A1(n19384), .A2(n19385), .ZN(n19383) );
  NAND2_X1 U19315 ( .A1(n19807), .A2(n16021), .ZN(n16022) );
  AOI21_X1 U19316 ( .B1(n19383), .B2(n16022), .A(n19376), .ZN(n19377) );
  NOR3_X1 U19317 ( .A1(n19377), .A2(n19378), .A3(n16023), .ZN(n16024) );
  AOI211_X1 U19318 ( .C1(n16027), .C2(n16026), .A(n16025), .B(n16024), .ZN(
        n16028) );
  INV_X1 U19319 ( .A(n16028), .ZN(P2_U2914) );
  NOR2_X1 U19320 ( .A1(n16030), .A2(n16029), .ZN(n16031) );
  AOI21_X1 U19321 ( .B1(n16303), .B2(n16039), .A(n16032), .ZN(n16311) );
  NAND2_X1 U19322 ( .A1(n16281), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16304) );
  OAI21_X1 U19323 ( .B1(n16283), .B2(n16033), .A(n16304), .ZN(n16034) );
  AOI21_X1 U19324 ( .B1(n16035), .B2(n19487), .A(n16034), .ZN(n16036) );
  OAI21_X1 U19325 ( .B1(n16308), .B2(n16287), .A(n16036), .ZN(n16037) );
  AOI21_X1 U19326 ( .B1(n19470), .B2(n16311), .A(n16037), .ZN(n16038) );
  OAI21_X1 U19327 ( .B1(n16313), .B2(n16299), .A(n16038), .ZN(P2_U2985) );
  NOR2_X1 U19328 ( .A1(n16055), .A2(n16315), .ZN(n16338) );
  INV_X1 U19329 ( .A(n16321), .ZN(n16043) );
  NAND2_X1 U19330 ( .A1(n16281), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16314) );
  NAND2_X1 U19331 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16040) );
  OAI211_X1 U19332 ( .C1(n16041), .C2(n19476), .A(n16314), .B(n16040), .ZN(
        n16042) );
  AOI21_X1 U19333 ( .B1(n16043), .B2(n19493), .A(n16042), .ZN(n16049) );
  INV_X1 U19334 ( .A(n16044), .ZN(n16046) );
  XOR2_X1 U19335 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n16047), .Z(
        n16048) );
  NAND2_X1 U19336 ( .A1(n16332), .A2(n19493), .ZN(n16060) );
  NOR2_X1 U19337 ( .A1(n19333), .A2(n20156), .ZN(n16326) );
  NOR2_X1 U19338 ( .A1(n16283), .A2(n16050), .ZN(n16051) );
  AOI211_X1 U19339 ( .C1(n16052), .C2(n19487), .A(n16326), .B(n16051), .ZN(
        n16059) );
  OR2_X1 U19340 ( .A1(n16053), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16334) );
  NAND3_X1 U19341 ( .A1(n16334), .A2(n19484), .A3(n16333), .ZN(n16058) );
  INV_X1 U19342 ( .A(n16338), .ZN(n16056) );
  NAND2_X1 U19343 ( .A1(n16055), .A2(n16315), .ZN(n16324) );
  NAND3_X1 U19344 ( .A1(n16056), .A2(n19470), .A3(n16324), .ZN(n16057) );
  NAND4_X1 U19345 ( .A1(n16060), .A2(n16059), .A3(n16058), .A4(n16057), .ZN(
        P2_U2987) );
  NAND2_X1 U19346 ( .A1(n16067), .A2(n16066), .ZN(n16354) );
  NOR2_X1 U19347 ( .A1(n16349), .A2(n16287), .ZN(n16072) );
  NAND2_X1 U19348 ( .A1(n16281), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16341) );
  NAND2_X1 U19349 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16069) );
  OAI211_X1 U19350 ( .C1(n16070), .C2(n19476), .A(n16341), .B(n16069), .ZN(
        n16071) );
  AOI211_X1 U19351 ( .C1(n16352), .C2(n19470), .A(n16072), .B(n16071), .ZN(
        n16073) );
  OAI21_X1 U19352 ( .B1(n16299), .B2(n16354), .A(n16073), .ZN(P2_U2988) );
  OAI21_X1 U19353 ( .B1(n16283), .B2(n10490), .A(n16074), .ZN(n16075) );
  AOI21_X1 U19354 ( .B1(n16076), .B2(n19487), .A(n16075), .ZN(n16077) );
  OAI21_X1 U19355 ( .B1(n16078), .B2(n16287), .A(n16077), .ZN(n16079) );
  AOI21_X1 U19356 ( .B1(n16080), .B2(n19484), .A(n16079), .ZN(n16081) );
  OAI21_X1 U19357 ( .B1(n19490), .B2(n16082), .A(n16081), .ZN(P2_U2989) );
  INV_X1 U19358 ( .A(n16100), .ZN(n16085) );
  INV_X1 U19359 ( .A(n16083), .ZN(n16084) );
  OAI21_X1 U19360 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16085), .A(
        n16084), .ZN(n16366) );
  XNOR2_X1 U19361 ( .A(n16086), .B(n21468), .ZN(n16087) );
  XNOR2_X1 U19362 ( .A(n16088), .B(n16087), .ZN(n16364) );
  AND2_X1 U19363 ( .A1(n19359), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16356) );
  NOR2_X1 U19364 ( .A1(n16089), .A2(n19476), .ZN(n16090) );
  AOI211_X1 U19365 ( .C1(n19483), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16356), .B(n16090), .ZN(n16091) );
  OAI21_X1 U19366 ( .B1(n16362), .B2(n16287), .A(n16091), .ZN(n16092) );
  AOI21_X1 U19367 ( .B1(n19484), .B2(n16364), .A(n16092), .ZN(n16093) );
  OAI21_X1 U19368 ( .B1(n16366), .B2(n19490), .A(n16093), .ZN(P2_U2990) );
  XNOR2_X1 U19369 ( .A(n16095), .B(n10350), .ZN(n16376) );
  NAND2_X1 U19370 ( .A1(n16281), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16369) );
  OAI21_X1 U19371 ( .B1(n16283), .B2(n16096), .A(n16369), .ZN(n16097) );
  AOI21_X1 U19372 ( .B1(n16098), .B2(n19487), .A(n16097), .ZN(n16099) );
  OAI21_X1 U19373 ( .B1(n16372), .B2(n16287), .A(n16099), .ZN(n16101) );
  OAI21_X1 U19374 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n10343), .A(
        n10268), .ZN(n16390) );
  INV_X1 U19375 ( .A(n16710), .ZN(n16105) );
  NAND2_X1 U19376 ( .A1(n16281), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16380) );
  NAND2_X1 U19377 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16103) );
  OAI211_X1 U19378 ( .C1(n16715), .C2(n19476), .A(n16380), .B(n16103), .ZN(
        n16104) );
  AOI21_X1 U19379 ( .B1(n16105), .B2(n19493), .A(n16104), .ZN(n16110) );
  OAI21_X1 U19380 ( .B1(n16108), .B2(n16107), .A(n16106), .ZN(n16388) );
  NAND2_X1 U19381 ( .A1(n16388), .A2(n19484), .ZN(n16109) );
  OAI211_X1 U19382 ( .C1(n16390), .C2(n19490), .A(n16110), .B(n16109), .ZN(
        P2_U2992) );
  NAND2_X1 U19383 ( .A1(n16112), .A2(n16111), .ZN(n16113) );
  XNOR2_X1 U19384 ( .A(n16114), .B(n16113), .ZN(n16406) );
  NAND2_X1 U19385 ( .A1(n16281), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n16396) );
  NAND2_X1 U19386 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16115) );
  OAI211_X1 U19387 ( .C1(n16116), .C2(n19476), .A(n16396), .B(n16115), .ZN(
        n16117) );
  AOI21_X1 U19388 ( .B1(n16400), .B2(n19493), .A(n16117), .ZN(n16120) );
  NAND2_X1 U19389 ( .A1(n16404), .A2(n19470), .ZN(n16119) );
  OAI211_X1 U19390 ( .C1(n16406), .C2(n16299), .A(n16120), .B(n16119), .ZN(
        P2_U2994) );
  NAND2_X1 U19391 ( .A1(n16122), .A2(n16121), .ZN(n16124) );
  XOR2_X1 U19392 ( .A(n16124), .B(n16123), .Z(n16428) );
  AOI21_X1 U19393 ( .B1(n16435), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16125) );
  NAND2_X1 U19394 ( .A1(n16417), .A2(n19470), .ZN(n16130) );
  NAND2_X1 U19395 ( .A1(n19359), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16419) );
  NAND2_X1 U19396 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16126) );
  OAI211_X1 U19397 ( .C1(n16127), .C2(n19476), .A(n16419), .B(n16126), .ZN(
        n16128) );
  AOI21_X1 U19398 ( .B1(n16425), .B2(n19493), .A(n16128), .ZN(n16129) );
  OAI211_X1 U19399 ( .C1(n16299), .C2(n16428), .A(n16130), .B(n16129), .ZN(
        P2_U2996) );
  XNOR2_X1 U19400 ( .A(n16435), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16136) );
  XNOR2_X1 U19401 ( .A(n9845), .B(n16131), .ZN(n16440) );
  NOR2_X1 U19402 ( .A1(n19321), .A2(n16287), .ZN(n16134) );
  INV_X1 U19403 ( .A(n19319), .ZN(n19327) );
  NAND2_X1 U19404 ( .A1(n19359), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16437) );
  NAND2_X1 U19405 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16132) );
  OAI211_X1 U19406 ( .C1(n19327), .C2(n19476), .A(n16437), .B(n16132), .ZN(
        n16133) );
  AOI211_X1 U19407 ( .C1(n16440), .C2(n19484), .A(n16134), .B(n16133), .ZN(
        n16135) );
  OAI21_X1 U19408 ( .B1(n16136), .B2(n19490), .A(n16135), .ZN(P2_U2997) );
  XNOR2_X1 U19409 ( .A(n16455), .B(n16436), .ZN(n16144) );
  XOR2_X1 U19410 ( .A(n16139), .B(n16138), .Z(n16451) );
  NOR2_X1 U19411 ( .A1(n19346), .A2(n16287), .ZN(n16142) );
  NAND2_X1 U19412 ( .A1(n19359), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16448) );
  NAND2_X1 U19413 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16140) );
  OAI211_X1 U19414 ( .C1(n19476), .C2(n19340), .A(n16448), .B(n16140), .ZN(
        n16141) );
  AOI211_X1 U19415 ( .C1(n16451), .C2(n19484), .A(n16142), .B(n16141), .ZN(
        n16143) );
  OAI21_X1 U19416 ( .B1(n16144), .B2(n19490), .A(n16143), .ZN(P2_U2998) );
  NAND2_X1 U19417 ( .A1(n16146), .A2(n16145), .ZN(n16149) );
  NAND2_X1 U19418 ( .A1(n16147), .A2(n16156), .ZN(n16148) );
  XOR2_X1 U19419 ( .A(n16149), .B(n16148), .Z(n16468) );
  NAND2_X1 U19420 ( .A1(n16150), .A2(n16461), .ZN(n16456) );
  NAND3_X1 U19421 ( .A1(n16456), .A2(n19470), .A3(n16455), .ZN(n16154) );
  NAND2_X1 U19422 ( .A1(n19359), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16459) );
  NAND2_X1 U19423 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16151) );
  OAI211_X1 U19424 ( .C1(n19476), .C2(n19338), .A(n16459), .B(n16151), .ZN(
        n16152) );
  AOI21_X1 U19425 ( .B1(n16465), .B2(n19493), .A(n16152), .ZN(n16153) );
  OAI211_X1 U19426 ( .C1(n16468), .C2(n16299), .A(n16154), .B(n16153), .ZN(
        P2_U2999) );
  NAND2_X1 U19427 ( .A1(n16156), .A2(n16155), .ZN(n16158) );
  XOR2_X1 U19428 ( .A(n16158), .B(n16157), .Z(n16481) );
  NAND2_X1 U19429 ( .A1(n16469), .A2(n19470), .ZN(n16164) );
  NAND2_X1 U19430 ( .A1(n19359), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n16472) );
  OAI21_X1 U19431 ( .B1(n16283), .B2(n16159), .A(n16472), .ZN(n16161) );
  NOR2_X1 U19432 ( .A1(n16470), .A2(n16287), .ZN(n16160) );
  AOI211_X1 U19433 ( .C1(n19487), .C2(n16162), .A(n16161), .B(n16160), .ZN(
        n16163) );
  OAI211_X1 U19434 ( .C1(n16299), .C2(n16481), .A(n16164), .B(n16163), .ZN(
        P2_U3000) );
  INV_X1 U19435 ( .A(n16201), .ZN(n16167) );
  NOR2_X1 U19436 ( .A1(n16166), .A2(n16167), .ZN(n16194) );
  AOI21_X1 U19437 ( .B1(n16194), .B2(n16195), .A(n16168), .ZN(n16182) );
  INV_X1 U19438 ( .A(n16180), .ZN(n16169) );
  AOI21_X1 U19439 ( .B1(n16182), .B2(n16179), .A(n16169), .ZN(n16173) );
  NAND2_X1 U19440 ( .A1(n16171), .A2(n16170), .ZN(n16172) );
  XNOR2_X1 U19441 ( .A(n16173), .B(n16172), .ZN(n16489) );
  NOR2_X1 U19442 ( .A1(n16485), .A2(n16287), .ZN(n16177) );
  NAND2_X1 U19443 ( .A1(n19359), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16484) );
  NAND2_X1 U19444 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16174) );
  OAI211_X1 U19445 ( .C1(n19476), .C2(n16175), .A(n16484), .B(n16174), .ZN(
        n16176) );
  AOI211_X1 U19446 ( .C1(n16489), .C2(n19484), .A(n16177), .B(n16176), .ZN(
        n16178) );
  OAI21_X1 U19447 ( .B1(n16492), .B2(n19490), .A(n16178), .ZN(P2_U3001) );
  NAND2_X1 U19448 ( .A1(n16180), .A2(n16179), .ZN(n16181) );
  XNOR2_X1 U19449 ( .A(n16182), .B(n16181), .ZN(n16503) );
  NAND2_X1 U19450 ( .A1(n16183), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16212) );
  NAND2_X1 U19451 ( .A1(n16204), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16189) );
  NAND2_X1 U19452 ( .A1(n16189), .A2(n21438), .ZN(n16493) );
  NAND2_X1 U19453 ( .A1(n19359), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n16494) );
  NAND2_X1 U19454 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16184) );
  OAI211_X1 U19455 ( .C1(n19476), .C2(n16185), .A(n16494), .B(n16184), .ZN(
        n16186) );
  AOI21_X1 U19456 ( .B1(n16500), .B2(n19493), .A(n16186), .ZN(n16187) );
  OAI211_X1 U19457 ( .C1(n16503), .C2(n16299), .A(n16188), .B(n16187), .ZN(
        P2_U3002) );
  OAI21_X1 U19458 ( .B1(n16204), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16189), .ZN(n16517) );
  NAND2_X1 U19459 ( .A1(n19487), .A2(n16190), .ZN(n16191) );
  NAND2_X1 U19460 ( .A1(n19359), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16505) );
  OAI211_X1 U19461 ( .C1(n16283), .C2(n21400), .A(n16191), .B(n16505), .ZN(
        n16199) );
  INV_X1 U19462 ( .A(n16192), .ZN(n16193) );
  NOR2_X1 U19463 ( .A1(n16194), .A2(n16193), .ZN(n16198) );
  NAND2_X1 U19464 ( .A1(n16196), .A2(n16195), .ZN(n16197) );
  NAND2_X1 U19465 ( .A1(n16201), .A2(n16200), .ZN(n16203) );
  NAND2_X1 U19466 ( .A1(n16166), .A2(n16216), .ZN(n16202) );
  XOR2_X1 U19467 ( .A(n16203), .B(n16202), .Z(n16530) );
  INV_X1 U19468 ( .A(n16204), .ZN(n16519) );
  NAND2_X1 U19469 ( .A1(n16212), .A2(n16205), .ZN(n16518) );
  NAND3_X1 U19470 ( .A1(n16519), .A2(n19470), .A3(n16518), .ZN(n16211) );
  NAND2_X1 U19471 ( .A1(n19359), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n16522) );
  OAI21_X1 U19472 ( .B1(n16283), .B2(n16206), .A(n16522), .ZN(n16208) );
  NOR2_X1 U19473 ( .A1(n16524), .A2(n16287), .ZN(n16207) );
  AOI211_X1 U19474 ( .C1(n16209), .C2(n19487), .A(n16208), .B(n16207), .ZN(
        n16210) );
  OAI211_X1 U19475 ( .C1(n16530), .C2(n16299), .A(n16211), .B(n16210), .ZN(
        P2_U3004) );
  OAI21_X1 U19476 ( .B1(n16183), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16212), .ZN(n16544) );
  INV_X1 U19477 ( .A(n16166), .ZN(n16217) );
  AOI21_X1 U19478 ( .B1(n16214), .B2(n16216), .A(n16213), .ZN(n16215) );
  AOI21_X1 U19479 ( .B1(n16217), .B2(n16216), .A(n16215), .ZN(n16542) );
  INV_X1 U19480 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20123) );
  NOR2_X1 U19481 ( .A1(n19333), .A2(n20123), .ZN(n16532) );
  NOR2_X1 U19482 ( .A1(n19476), .A2(n16218), .ZN(n16219) );
  AOI211_X1 U19483 ( .C1(n19483), .C2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16532), .B(n16219), .ZN(n16220) );
  OAI21_X1 U19484 ( .B1(n16531), .B2(n16287), .A(n16220), .ZN(n16221) );
  AOI21_X1 U19485 ( .B1(n16542), .B2(n19484), .A(n16221), .ZN(n16222) );
  OAI21_X1 U19486 ( .B1(n16544), .B2(n19490), .A(n16222), .ZN(P2_U3005) );
  NAND2_X1 U19487 ( .A1(n16224), .A2(n16223), .ZN(n16230) );
  XNOR2_X1 U19488 ( .A(n16226), .B(n16593), .ZN(n16264) );
  OAI22_X1 U19489 ( .A1(n16264), .A2(n16225), .B1(n16226), .B2(n16593), .ZN(
        n16256) );
  XOR2_X1 U19490 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16227), .Z(
        n16257) );
  AOI22_X1 U19491 ( .A1(n16256), .A2(n16257), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16227), .ZN(n16242) );
  INV_X1 U19492 ( .A(n16239), .ZN(n16228) );
  OAI21_X1 U19493 ( .B1(n16242), .B2(n16228), .A(n16240), .ZN(n16229) );
  XOR2_X1 U19494 ( .A(n16230), .B(n16229), .Z(n16564) );
  NAND2_X1 U19495 ( .A1(n19359), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16550) );
  OAI21_X1 U19496 ( .B1(n16283), .B2(n16231), .A(n16550), .ZN(n16233) );
  NOR2_X1 U19497 ( .A1(n16551), .A2(n16287), .ZN(n16232) );
  AOI211_X1 U19498 ( .C1(n16234), .C2(n19487), .A(n16233), .B(n16232), .ZN(
        n16238) );
  OR2_X1 U19499 ( .A1(n16236), .A2(n16235), .ZN(n16545) );
  NAND3_X1 U19500 ( .A1(n16545), .A2(n19470), .A3(n16546), .ZN(n16237) );
  OAI211_X1 U19501 ( .C1(n16564), .C2(n16299), .A(n16238), .B(n16237), .ZN(
        P2_U3006) );
  NAND2_X1 U19502 ( .A1(n16240), .A2(n16239), .ZN(n16241) );
  XNOR2_X1 U19503 ( .A(n16242), .B(n16241), .ZN(n16576) );
  NAND2_X1 U19504 ( .A1(n16258), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16245) );
  NAND2_X1 U19505 ( .A1(n16245), .A2(n16244), .ZN(n16249) );
  NAND2_X1 U19506 ( .A1(n16247), .A2(n16246), .ZN(n16248) );
  XNOR2_X1 U19507 ( .A(n16249), .B(n16248), .ZN(n16574) );
  OAI22_X1 U19508 ( .A1(n16283), .A2(n16250), .B1(n20119), .B2(n19333), .ZN(
        n16251) );
  AOI21_X1 U19509 ( .B1(n19487), .B2(n16252), .A(n16251), .ZN(n16253) );
  OAI21_X1 U19510 ( .B1(n16566), .B2(n16287), .A(n16253), .ZN(n16254) );
  AOI21_X1 U19511 ( .B1(n16574), .B2(n19470), .A(n16254), .ZN(n16255) );
  OAI21_X1 U19512 ( .B1(n16576), .B2(n16299), .A(n16255), .ZN(P2_U3007) );
  XNOR2_X1 U19513 ( .A(n16257), .B(n16256), .ZN(n16587) );
  XOR2_X1 U19514 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16258), .Z(
        n16585) );
  NAND2_X1 U19515 ( .A1(n19359), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n16582) );
  OAI21_X1 U19516 ( .B1(n16283), .B2(n16259), .A(n16582), .ZN(n16260) );
  AOI21_X1 U19517 ( .B1(n19487), .B2(n19363), .A(n16260), .ZN(n16261) );
  OAI21_X1 U19518 ( .B1(n19369), .B2(n16287), .A(n16261), .ZN(n16262) );
  AOI21_X1 U19519 ( .B1(n16585), .B2(n19470), .A(n16262), .ZN(n16263) );
  OAI21_X1 U19520 ( .B1(n16299), .B2(n16587), .A(n16263), .ZN(P2_U3008) );
  XNOR2_X1 U19521 ( .A(n16225), .B(n16264), .ZN(n16602) );
  AOI21_X1 U19522 ( .B1(n16268), .B2(n16266), .A(n16265), .ZN(n16267) );
  AOI21_X1 U19523 ( .B1(n16269), .B2(n16268), .A(n16267), .ZN(n16588) );
  NOR2_X1 U19524 ( .A1(n16597), .A2(n16287), .ZN(n16273) );
  NAND2_X1 U19525 ( .A1(n19359), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n16596) );
  NAND2_X1 U19526 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16270) );
  OAI211_X1 U19527 ( .C1(n19476), .C2(n16271), .A(n16596), .B(n16270), .ZN(
        n16272) );
  AOI211_X1 U19528 ( .C1(n16588), .C2(n19470), .A(n16273), .B(n16272), .ZN(
        n16274) );
  OAI21_X1 U19529 ( .B1(n16299), .B2(n16602), .A(n16274), .ZN(P2_U3009) );
  XNOR2_X1 U19530 ( .A(n16275), .B(n16617), .ZN(n16291) );
  AOI22_X1 U19531 ( .A1(n16291), .A2(n16290), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16275), .ZN(n16278) );
  XNOR2_X1 U19532 ( .A(n16276), .B(n16592), .ZN(n16277) );
  XNOR2_X1 U19533 ( .A(n16278), .B(n16277), .ZN(n16614) );
  XNOR2_X1 U19534 ( .A(n16280), .B(n16279), .ZN(n16611) );
  NAND2_X1 U19535 ( .A1(n16281), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n16603) );
  OAI21_X1 U19536 ( .B1(n16283), .B2(n16282), .A(n16603), .ZN(n16284) );
  AOI21_X1 U19537 ( .B1(n19487), .B2(n16285), .A(n16284), .ZN(n16286) );
  OAI21_X1 U19538 ( .B1(n16607), .B2(n16287), .A(n16286), .ZN(n16288) );
  AOI21_X1 U19539 ( .B1(n16611), .B2(n19470), .A(n16288), .ZN(n16289) );
  OAI21_X1 U19540 ( .B1(n16614), .B2(n16299), .A(n16289), .ZN(P2_U3010) );
  XNOR2_X1 U19541 ( .A(n16291), .B(n16290), .ZN(n16626) );
  AOI22_X1 U19542 ( .A1(n19483), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n19359), .ZN(n16292) );
  OAI21_X1 U19543 ( .B1(n19476), .B2(n16293), .A(n16292), .ZN(n16294) );
  AOI21_X1 U19544 ( .B1(n15771), .B2(n19493), .A(n16294), .ZN(n16298) );
  NAND3_X1 U19545 ( .A1(n16615), .A2(n19470), .A3(n16296), .ZN(n16297) );
  OAI211_X1 U19546 ( .C1(n16626), .C2(n16299), .A(n16298), .B(n16297), .ZN(
        P2_U3011) );
  NOR2_X1 U19547 ( .A1(n16300), .A2(n16590), .ZN(n16310) );
  OR2_X1 U19548 ( .A1(n16329), .A2(n16316), .ZN(n16302) );
  INV_X1 U19549 ( .A(n16327), .ZN(n16301) );
  NAND2_X1 U19550 ( .A1(n16302), .A2(n16301), .ZN(n16319) );
  NAND2_X1 U19551 ( .A1(n16316), .A2(n16303), .ZN(n16305) );
  OAI21_X1 U19552 ( .B1(n16329), .B2(n16305), .A(n16304), .ZN(n16306) );
  AOI21_X1 U19553 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16319), .A(
        n16306), .ZN(n16307) );
  OAI21_X1 U19554 ( .B1(n16308), .B2(n16836), .A(n16307), .ZN(n16309) );
  OAI21_X1 U19555 ( .B1(n16313), .B2(n16625), .A(n16312), .ZN(P2_U3017) );
  INV_X1 U19556 ( .A(n16314), .ZN(n16318) );
  NOR3_X1 U19557 ( .A1(n16329), .A2(n16316), .A3(n16315), .ZN(n16317) );
  AOI211_X1 U19558 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16319), .A(
        n16318), .B(n16317), .ZN(n16320) );
  NAND2_X1 U19559 ( .A1(n16324), .A2(n16640), .ZN(n16337) );
  NOR2_X1 U19560 ( .A1(n16325), .A2(n16590), .ZN(n16331) );
  AOI21_X1 U19561 ( .B1(n16327), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16326), .ZN(n16328) );
  OAI21_X1 U19562 ( .B1(n16329), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16328), .ZN(n16330) );
  AOI211_X1 U19563 ( .C1(n16332), .C2(n16633), .A(n16331), .B(n16330), .ZN(
        n16336) );
  NAND3_X1 U19564 ( .A1(n16334), .A2(n16832), .A3(n16333), .ZN(n16335) );
  OAI211_X1 U19565 ( .C1(n16338), .C2(n16337), .A(n16336), .B(n16335), .ZN(
        P2_U3019) );
  NOR2_X1 U19566 ( .A1(n16339), .A2(n16590), .ZN(n16351) );
  NAND2_X1 U19567 ( .A1(n16340), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16342) );
  OAI21_X1 U19568 ( .B1(n16355), .B2(n16342), .A(n16341), .ZN(n16343) );
  INV_X1 U19569 ( .A(n16343), .ZN(n16348) );
  INV_X1 U19570 ( .A(n16344), .ZN(n16345) );
  OAI211_X1 U19571 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n16346), .B(n16345), .ZN(
        n16347) );
  OAI211_X1 U19572 ( .C1(n16349), .C2(n16836), .A(n16348), .B(n16347), .ZN(
        n16350) );
  AOI211_X1 U19573 ( .C1(n16352), .C2(n16640), .A(n16351), .B(n16350), .ZN(
        n16353) );
  OAI21_X1 U19574 ( .B1(n16625), .B2(n16354), .A(n16353), .ZN(P2_U3020) );
  OAI21_X1 U19575 ( .B1(n16367), .B2(n16368), .A(n21468), .ZN(n16358) );
  INV_X1 U19576 ( .A(n16355), .ZN(n16357) );
  AOI21_X1 U19577 ( .B1(n16358), .B2(n16357), .A(n16356), .ZN(n16361) );
  NAND2_X1 U19578 ( .A1(n16359), .A2(n16838), .ZN(n16360) );
  OAI211_X1 U19579 ( .C1(n16362), .C2(n16836), .A(n16361), .B(n16360), .ZN(
        n16363) );
  AOI21_X1 U19580 ( .B1(n16832), .B2(n16364), .A(n16363), .ZN(n16365) );
  OAI21_X1 U19581 ( .B1(n16366), .B2(n16842), .A(n16365), .ZN(P2_U3022) );
  INV_X1 U19582 ( .A(n16367), .ZN(n16384) );
  OAI211_X1 U19583 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16384), .B(n16368), .ZN(
        n16370) );
  OAI211_X1 U19584 ( .C1(n16381), .C2(n16371), .A(n16370), .B(n16369), .ZN(
        n16374) );
  NOR2_X1 U19585 ( .A1(n16372), .A2(n16836), .ZN(n16373) );
  AOI211_X1 U19586 ( .C1(n16375), .C2(n16838), .A(n16374), .B(n16373), .ZN(
        n16378) );
  NAND2_X1 U19587 ( .A1(n16376), .A2(n16832), .ZN(n16377) );
  OAI211_X1 U19588 ( .C1(n16379), .C2(n16842), .A(n16378), .B(n16377), .ZN(
        P2_U3023) );
  NOR2_X1 U19589 ( .A1(n16709), .A2(n16590), .ZN(n16387) );
  OAI21_X1 U19590 ( .B1(n16381), .B2(n16383), .A(n16380), .ZN(n16382) );
  AOI21_X1 U19591 ( .B1(n16384), .B2(n16383), .A(n16382), .ZN(n16385) );
  OAI21_X1 U19592 ( .B1(n16710), .B2(n16836), .A(n16385), .ZN(n16386) );
  AOI211_X1 U19593 ( .C1(n16832), .C2(n16388), .A(n16387), .B(n16386), .ZN(
        n16389) );
  OAI21_X1 U19594 ( .B1(n16842), .B2(n16390), .A(n16389), .ZN(P2_U3024) );
  NAND2_X1 U19595 ( .A1(n16391), .A2(n16409), .ZN(n16408) );
  NAND2_X1 U19596 ( .A1(n16556), .A2(n16392), .ZN(n16393) );
  AND2_X1 U19597 ( .A1(n16462), .A2(n16393), .ZN(n16420) );
  AOI21_X1 U19598 ( .B1(n16408), .B2(n16420), .A(n16394), .ZN(n16399) );
  INV_X1 U19599 ( .A(n16441), .ZN(n16458) );
  NAND4_X1 U19600 ( .A1(n16458), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16395), .A4(n16394), .ZN(n16397) );
  NAND2_X1 U19601 ( .A1(n16397), .A2(n16396), .ZN(n16398) );
  AOI211_X1 U19602 ( .C1(n16400), .C2(n16633), .A(n16399), .B(n16398), .ZN(
        n16401) );
  OAI21_X1 U19603 ( .B1(n16590), .B2(n16402), .A(n16401), .ZN(n16403) );
  AOI21_X1 U19604 ( .B1(n16404), .B2(n16640), .A(n16403), .ZN(n16405) );
  OAI21_X1 U19605 ( .B1(n16406), .B2(n16625), .A(n16405), .ZN(P2_U3026) );
  OAI211_X1 U19606 ( .C1(n16420), .C2(n16409), .A(n16408), .B(n16407), .ZN(
        n16410) );
  AOI21_X1 U19607 ( .B1(n16411), .B2(n16633), .A(n16410), .ZN(n16414) );
  NAND2_X1 U19608 ( .A1(n16412), .A2(n16838), .ZN(n16413) );
  NAND2_X1 U19609 ( .A1(n16417), .A2(n16640), .ZN(n16427) );
  AOI21_X1 U19610 ( .B1(n16458), .B2(n16418), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16421) );
  OAI21_X1 U19611 ( .B1(n16421), .B2(n16420), .A(n16419), .ZN(n16424) );
  NOR2_X1 U19612 ( .A1(n16422), .A2(n16590), .ZN(n16423) );
  AOI211_X1 U19613 ( .C1(n16425), .C2(n16633), .A(n16424), .B(n16423), .ZN(
        n16426) );
  OAI211_X1 U19614 ( .C1(n16428), .C2(n16625), .A(n16427), .B(n16426), .ZN(
        P2_U3028) );
  INV_X1 U19615 ( .A(n16429), .ZN(n16642) );
  NOR2_X1 U19616 ( .A1(n16640), .A2(n16642), .ZN(n16434) );
  INV_X1 U19617 ( .A(n16462), .ZN(n16432) );
  AOI21_X1 U19618 ( .B1(n16436), .B2(n16556), .A(n16447), .ZN(n16445) );
  NAND2_X1 U19619 ( .A1(n19323), .A2(n16838), .ZN(n16438) );
  OAI211_X1 U19620 ( .C1(n19321), .C2(n16836), .A(n16438), .B(n16437), .ZN(
        n16439) );
  AOI21_X1 U19621 ( .B1(n16440), .B2(n16832), .A(n16439), .ZN(n16443) );
  NAND3_X1 U19622 ( .A1(n16446), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16444), .ZN(n16442) );
  OAI211_X1 U19623 ( .C1(n16445), .C2(n16444), .A(n16443), .B(n16442), .ZN(
        P2_U3029) );
  INV_X1 U19624 ( .A(n16446), .ZN(n16454) );
  NAND2_X1 U19625 ( .A1(n16447), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16453) );
  NOR2_X1 U19626 ( .A1(n19349), .A2(n16590), .ZN(n16450) );
  OAI21_X1 U19627 ( .B1(n19346), .B2(n16836), .A(n16448), .ZN(n16449) );
  AOI211_X1 U19628 ( .C1(n16451), .C2(n16832), .A(n16450), .B(n16449), .ZN(
        n16452) );
  OAI211_X1 U19629 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16454), .A(
        n16453), .B(n16452), .ZN(P2_U3030) );
  NAND3_X1 U19630 ( .A1(n16456), .A2(n16640), .A3(n16455), .ZN(n16467) );
  NOR2_X1 U19631 ( .A1(n16457), .A2(n16590), .ZN(n16464) );
  NAND2_X1 U19632 ( .A1(n16458), .A2(n16461), .ZN(n16460) );
  OAI211_X1 U19633 ( .C1(n16462), .C2(n16461), .A(n16460), .B(n16459), .ZN(
        n16463) );
  AOI211_X1 U19634 ( .C1(n16465), .C2(n16633), .A(n16464), .B(n16463), .ZN(
        n16466) );
  OAI211_X1 U19635 ( .C1(n16468), .C2(n16625), .A(n16467), .B(n16466), .ZN(
        P2_U3031) );
  NAND2_X1 U19636 ( .A1(n16469), .A2(n16640), .ZN(n16480) );
  INV_X1 U19637 ( .A(n16470), .ZN(n16478) );
  XNOR2_X1 U19638 ( .A(n21214), .B(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16471) );
  NAND2_X1 U19639 ( .A1(n16482), .A2(n16471), .ZN(n16473) );
  OAI211_X1 U19640 ( .C1(n16496), .C2(n16474), .A(n16473), .B(n16472), .ZN(
        n16477) );
  NOR2_X1 U19641 ( .A1(n16475), .A2(n16590), .ZN(n16476) );
  AOI211_X1 U19642 ( .C1(n16478), .C2(n16633), .A(n16477), .B(n16476), .ZN(
        n16479) );
  OAI211_X1 U19643 ( .C1(n16481), .C2(n16625), .A(n16480), .B(n16479), .ZN(
        P2_U3032) );
  NAND2_X1 U19644 ( .A1(n16482), .A2(n21438), .ZN(n16495) );
  AOI21_X1 U19645 ( .B1(n16495), .B2(n16496), .A(n21372), .ZN(n16487) );
  NAND3_X1 U19646 ( .A1(n16482), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n21372), .ZN(n16483) );
  OAI211_X1 U19647 ( .C1(n16485), .C2(n16836), .A(n16484), .B(n16483), .ZN(
        n16486) );
  AOI211_X1 U19648 ( .C1(n16488), .C2(n16838), .A(n16487), .B(n16486), .ZN(
        n16491) );
  NAND2_X1 U19649 ( .A1(n16489), .A2(n16832), .ZN(n16490) );
  OAI211_X1 U19650 ( .C1(n16492), .C2(n16842), .A(n16491), .B(n16490), .ZN(
        P2_U3033) );
  OAI211_X1 U19651 ( .C1(n16496), .C2(n21438), .A(n16495), .B(n16494), .ZN(
        n16499) );
  NOR2_X1 U19652 ( .A1(n16497), .A2(n16590), .ZN(n16498) );
  AOI211_X1 U19653 ( .C1(n16500), .C2(n16633), .A(n16499), .B(n16498), .ZN(
        n16501) );
  OAI211_X1 U19654 ( .C1(n16503), .C2(n16625), .A(n16502), .B(n16501), .ZN(
        P2_U3034) );
  INV_X1 U19655 ( .A(n16504), .ZN(n16515) );
  INV_X1 U19656 ( .A(n16505), .ZN(n16508) );
  INV_X1 U19657 ( .A(n16538), .ZN(n16510) );
  NOR3_X1 U19658 ( .A1(n16510), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16506), .ZN(n16507) );
  AOI211_X1 U19659 ( .C1(n16509), .C2(n16633), .A(n16508), .B(n16507), .ZN(
        n16512) );
  NOR3_X1 U19660 ( .A1(n16510), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n16537), .ZN(n16521) );
  OAI21_X1 U19661 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16846), .A(
        n16535), .ZN(n16527) );
  OAI21_X1 U19662 ( .B1(n16521), .B2(n16527), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16511) );
  OAI211_X1 U19663 ( .C1(n16513), .C2(n16590), .A(n16512), .B(n16511), .ZN(
        n16514) );
  AOI21_X1 U19664 ( .B1(n16515), .B2(n16832), .A(n16514), .ZN(n16516) );
  OAI21_X1 U19665 ( .B1(n16517), .B2(n16842), .A(n16516), .ZN(P2_U3035) );
  NAND3_X1 U19666 ( .A1(n16519), .A2(n16640), .A3(n16518), .ZN(n16529) );
  NOR2_X1 U19667 ( .A1(n16520), .A2(n16590), .ZN(n16526) );
  INV_X1 U19668 ( .A(n16521), .ZN(n16523) );
  OAI211_X1 U19669 ( .C1(n16524), .C2(n16836), .A(n16523), .B(n16522), .ZN(
        n16525) );
  AOI211_X1 U19670 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16527), .A(
        n16526), .B(n16525), .ZN(n16528) );
  OAI211_X1 U19671 ( .C1(n16530), .C2(n16625), .A(n16529), .B(n16528), .ZN(
        P2_U3036) );
  INV_X1 U19672 ( .A(n16531), .ZN(n16533) );
  AOI21_X1 U19673 ( .B1(n16533), .B2(n16633), .A(n16532), .ZN(n16534) );
  OAI21_X1 U19674 ( .B1(n16537), .B2(n16535), .A(n16534), .ZN(n16536) );
  AOI21_X1 U19675 ( .B1(n16538), .B2(n16537), .A(n16536), .ZN(n16539) );
  OAI21_X1 U19676 ( .B1(n16590), .B2(n16540), .A(n16539), .ZN(n16541) );
  AOI21_X1 U19677 ( .B1(n16542), .B2(n16832), .A(n16541), .ZN(n16543) );
  OAI21_X1 U19678 ( .B1(n16544), .B2(n16842), .A(n16543), .ZN(P2_U3037) );
  AND3_X1 U19679 ( .A1(n16546), .A2(n16640), .A3(n16545), .ZN(n16562) );
  AOI21_X1 U19680 ( .B1(n16558), .B2(n16569), .A(n16547), .ZN(n16548) );
  NAND2_X1 U19681 ( .A1(n16570), .A2(n16548), .ZN(n16549) );
  OAI211_X1 U19682 ( .C1(n16551), .C2(n16836), .A(n16550), .B(n16549), .ZN(
        n16561) );
  NAND2_X1 U19683 ( .A1(n16642), .A2(n16628), .ZN(n16552) );
  AND3_X1 U19684 ( .A1(n16553), .A2(n16552), .A3(n16627), .ZN(n16619) );
  INV_X1 U19685 ( .A(n16554), .ZN(n16555) );
  NAND2_X1 U19686 ( .A1(n16556), .A2(n16555), .ZN(n16557) );
  AND2_X1 U19687 ( .A1(n16619), .A2(n16557), .ZN(n16578) );
  OAI22_X1 U19688 ( .A1(n16559), .A2(n16590), .B1(n16578), .B2(n16558), .ZN(
        n16560) );
  NOR3_X1 U19689 ( .A1(n16562), .A2(n16561), .A3(n16560), .ZN(n16563) );
  OAI21_X1 U19690 ( .B1(n16564), .B2(n16625), .A(n16563), .ZN(P2_U3038) );
  NOR2_X1 U19691 ( .A1(n16578), .A2(n16569), .ZN(n16568) );
  NAND2_X1 U19692 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19359), .ZN(n16565) );
  OAI21_X1 U19693 ( .B1(n16566), .B2(n16836), .A(n16565), .ZN(n16567) );
  AOI211_X1 U19694 ( .C1(n16570), .C2(n16569), .A(n16568), .B(n16567), .ZN(
        n16571) );
  OAI21_X1 U19695 ( .B1(n16590), .B2(n16572), .A(n16571), .ZN(n16573) );
  AOI21_X1 U19696 ( .B1(n16574), .B2(n16640), .A(n16573), .ZN(n16575) );
  OAI21_X1 U19697 ( .B1(n16576), .B2(n16625), .A(n16575), .ZN(P2_U3039) );
  NAND2_X1 U19698 ( .A1(n16616), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16606) );
  INV_X1 U19699 ( .A(n16606), .ZN(n16577) );
  AOI21_X1 U19700 ( .B1(n16577), .B2(n16591), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16579) );
  NOR2_X1 U19701 ( .A1(n16579), .A2(n16578), .ZN(n16584) );
  NAND2_X1 U19702 ( .A1(n16580), .A2(n16838), .ZN(n16581) );
  OAI211_X1 U19703 ( .C1(n19369), .C2(n16836), .A(n16582), .B(n16581), .ZN(
        n16583) );
  AOI211_X1 U19704 ( .C1(n16585), .C2(n16640), .A(n16584), .B(n16583), .ZN(
        n16586) );
  OAI21_X1 U19705 ( .B1(n16625), .B2(n16587), .A(n16586), .ZN(P2_U3040) );
  NAND2_X1 U19706 ( .A1(n16588), .A2(n16640), .ZN(n16601) );
  OAI21_X1 U19707 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16846), .A(
        n16619), .ZN(n16610) );
  NOR2_X1 U19708 ( .A1(n16590), .A2(n16589), .ZN(n16599) );
  AOI211_X1 U19709 ( .C1(n16593), .C2(n16592), .A(n16591), .B(n16606), .ZN(
        n16594) );
  INV_X1 U19710 ( .A(n16594), .ZN(n16595) );
  OAI211_X1 U19711 ( .C1(n16597), .C2(n16836), .A(n16596), .B(n16595), .ZN(
        n16598) );
  AOI211_X1 U19712 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n16610), .A(
        n16599), .B(n16598), .ZN(n16600) );
  OAI211_X1 U19713 ( .C1(n16602), .C2(n16625), .A(n16601), .B(n16600), .ZN(
        P2_U3041) );
  INV_X1 U19714 ( .A(n16603), .ZN(n16604) );
  AOI21_X1 U19715 ( .B1(n19376), .B2(n16838), .A(n16604), .ZN(n16605) );
  OAI21_X1 U19716 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16606), .A(
        n16605), .ZN(n16609) );
  NOR2_X1 U19717 ( .A1(n16607), .A2(n16836), .ZN(n16608) );
  AOI211_X1 U19718 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n16610), .A(
        n16609), .B(n16608), .ZN(n16613) );
  NAND2_X1 U19719 ( .A1(n16611), .A2(n16640), .ZN(n16612) );
  OAI211_X1 U19720 ( .C1(n16614), .C2(n16625), .A(n16613), .B(n16612), .ZN(
        P2_U3042) );
  NAND3_X1 U19721 ( .A1(n16615), .A2(n16640), .A3(n16296), .ZN(n16623) );
  AOI22_X1 U19722 ( .A1(n16838), .A2(n20182), .B1(n19359), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n16622) );
  INV_X1 U19723 ( .A(n16616), .ZN(n16618) );
  MUX2_X1 U19724 ( .A(n16619), .B(n16618), .S(n16617), .Z(n16621) );
  NAND2_X1 U19725 ( .A1(n15771), .A2(n16633), .ZN(n16620) );
  AND4_X1 U19726 ( .A1(n16623), .A2(n16622), .A3(n16621), .A4(n16620), .ZN(
        n16624) );
  OAI21_X1 U19727 ( .B1(n16626), .B2(n16625), .A(n16624), .ZN(P2_U3043) );
  INV_X1 U19728 ( .A(n16627), .ZN(n16833) );
  INV_X1 U19729 ( .A(n16628), .ZN(n16630) );
  NAND2_X1 U19730 ( .A1(n16630), .A2(n16629), .ZN(n16641) );
  INV_X1 U19731 ( .A(n16641), .ZN(n16631) );
  AOI22_X1 U19732 ( .A1(n16833), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16632), .B2(n16631), .ZN(n16646) );
  AOI22_X1 U19733 ( .A1(n19479), .A2(n16633), .B1(n16838), .B2(n20194), .ZN(
        n16645) );
  OAI21_X1 U19734 ( .B1(n16636), .B2(n16635), .A(n16634), .ZN(n16637) );
  INV_X1 U19735 ( .A(n16637), .ZN(n19471) );
  XOR2_X1 U19736 ( .A(n16639), .B(n16638), .Z(n19472) );
  AOI22_X1 U19737 ( .A1(n19471), .A2(n16640), .B1(n16832), .B2(n19472), .ZN(
        n16644) );
  NOR2_X1 U19738 ( .A1(n19333), .A2(n20110), .ZN(n19473) );
  AOI21_X1 U19739 ( .B1(n16642), .B2(n16641), .A(n19473), .ZN(n16643) );
  NAND4_X1 U19740 ( .A1(n16646), .A2(n16645), .A3(n16644), .A4(n16643), .ZN(
        P2_U3044) );
  MUX2_X1 U19741 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16647), .S(
        n11664), .Z(n16652) );
  OAI222_X1 U19742 ( .A1(n16771), .A2(n16650), .B1(n16664), .B2(n16649), .C1(
        n16648), .C2(n16652), .ZN(n16651) );
  MUX2_X1 U19743 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n16651), .S(
        n16666), .Z(P2_U3601) );
  NAND2_X1 U19744 ( .A1(n16652), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16662) );
  OAI21_X1 U19745 ( .B1(n11664), .B2(n16654), .A(n16653), .ZN(n16659) );
  INV_X1 U19746 ( .A(n16771), .ZN(n16656) );
  AOI22_X1 U19747 ( .A1(n20199), .A2(n16656), .B1(n20179), .B2(n16655), .ZN(
        n16657) );
  OAI21_X1 U19748 ( .B1(n16662), .B2(n16659), .A(n16657), .ZN(n16658) );
  MUX2_X1 U19749 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16658), .S(
        n16666), .Z(P2_U3600) );
  INV_X1 U19750 ( .A(n16659), .ZN(n16661) );
  OAI222_X1 U19751 ( .A1(n20190), .A2(n16771), .B1(n16662), .B2(n16661), .C1(
        n16664), .C2(n16660), .ZN(n16663) );
  MUX2_X1 U19752 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16663), .S(
        n16666), .Z(P2_U3599) );
  OAI22_X1 U19753 ( .A1(n19807), .A2(n16771), .B1(n16665), .B2(n16664), .ZN(
        n16667) );
  MUX2_X1 U19754 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16667), .S(
        n16666), .Z(P2_U3596) );
  AOI22_X1 U19755 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16673) );
  AOI22_X1 U19756 ( .A1(n17580), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16672) );
  AOI22_X1 U19757 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16671) );
  AOI22_X1 U19758 ( .A1(n17596), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16670) );
  NAND4_X1 U19759 ( .A1(n16673), .A2(n16672), .A3(n16671), .A4(n16670), .ZN(
        n16680) );
  AOI22_X1 U19760 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16678) );
  AOI22_X1 U19761 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16677) );
  AOI22_X1 U19762 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16676) );
  AOI22_X1 U19763 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16675) );
  NAND4_X1 U19764 ( .A1(n16678), .A2(n16677), .A3(n16676), .A4(n16675), .ZN(
        n16679) );
  NOR2_X1 U19765 ( .A1(n16680), .A2(n16679), .ZN(n17755) );
  AOI22_X1 U19766 ( .A1(n16681), .A2(n17216), .B1(n9735), .B2(n17560), .ZN(
        n17547) );
  AND2_X1 U19767 ( .A1(n17216), .A2(n17560), .ZN(n16682) );
  OAI22_X1 U19768 ( .A1(n17755), .A2(n9735), .B1(n17547), .B2(n16682), .ZN(
        P3_U2690) );
  NAND2_X1 U19769 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18779) );
  AOI221_X1 U19770 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18779), .C1(n16684), 
        .C2(n18779), .A(n16683), .ZN(n18609) );
  NOR2_X1 U19771 ( .A1(n16685), .A2(n19067), .ZN(n16686) );
  OAI21_X1 U19772 ( .B1(n16686), .B2(n18964), .A(n18610), .ZN(n18607) );
  AOI22_X1 U19773 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18609), .B1(
        n18607), .B2(n18613), .ZN(P3_U2865) );
  NAND2_X1 U19774 ( .A1(n19054), .A2(n19254), .ZN(n16692) );
  NOR2_X1 U19775 ( .A1(n19260), .A2(n16690), .ZN(n19104) );
  OAI21_X1 U19776 ( .B1(n16691), .B2(n19104), .A(n19259), .ZN(n17814) );
  NOR2_X1 U19777 ( .A1(n16692), .A2(n17814), .ZN(n16694) );
  NOR2_X1 U19778 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19212), .ZN(n18616) );
  NOR2_X1 U19779 ( .A1(n17006), .A2(n19210), .ZN(n16696) );
  INV_X1 U19780 ( .A(n19240), .ZN(n19238) );
  AOI21_X1 U19781 ( .B1(n16698), .B2(n17317), .A(n16697), .ZN(n19062) );
  NAND3_X1 U19782 ( .A1(n19238), .A2(n19274), .A3(n19062), .ZN(n16699) );
  OAI21_X1 U19783 ( .B1(n19238), .B2(n17317), .A(n16699), .ZN(P3_U3284) );
  INV_X1 U19784 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16878) );
  NAND2_X1 U19785 ( .A1(n9780), .A2(n19088), .ZN(n18488) );
  AOI21_X1 U19786 ( .B1(n18307), .B2(n18488), .A(n16700), .ZN(n16893) );
  OAI21_X1 U19787 ( .B1(n9743), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16893), .ZN(n16703) );
  AOI21_X1 U19788 ( .B1(n18595), .B2(n16703), .A(n16702), .ZN(n16707) );
  NAND2_X1 U19789 ( .A1(n18199), .A2(n17939), .ZN(n16897) );
  NOR2_X1 U19790 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18117), .ZN(
        n16705) );
  OAI22_X1 U19791 ( .A1(n16710), .A2(n19368), .B1(n16709), .B2(n19366), .ZN(
        n16711) );
  INV_X1 U19792 ( .A(n16711), .ZN(n16724) );
  INV_X1 U19793 ( .A(n16712), .ZN(n16721) );
  AOI22_X1 U19794 ( .A1(n19315), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19360), .ZN(n16713) );
  OAI21_X1 U19795 ( .B1(n19375), .B2(n16714), .A(n16713), .ZN(n16720) );
  OAI21_X1 U19796 ( .B1(n19310), .B2(n16715), .A(n19344), .ZN(n16717) );
  AOI21_X1 U19797 ( .B1(n16718), .B2(n16717), .A(n16716), .ZN(n16719) );
  AOI211_X1 U19798 ( .C1(n16722), .C2(n16721), .A(n16720), .B(n16719), .ZN(
        n16723) );
  NAND2_X1 U19799 ( .A1(n16724), .A2(n16723), .ZN(P2_U2833) );
  INV_X1 U19800 ( .A(n16737), .ZN(n16740) );
  INV_X1 U19801 ( .A(n16725), .ZN(n16726) );
  OAI211_X1 U19802 ( .C1(n16728), .C2(n16727), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16726), .ZN(n16732) );
  INV_X1 U19803 ( .A(n16729), .ZN(n16731) );
  OAI211_X1 U19804 ( .C1(n20905), .C2(n16732), .A(n16731), .B(n16730), .ZN(
        n16734) );
  NAND2_X1 U19805 ( .A1(n20905), .A2(n16732), .ZN(n16733) );
  NAND2_X1 U19806 ( .A1(n16734), .A2(n16733), .ZN(n16738) );
  AND2_X1 U19807 ( .A1(n20830), .A2(n16738), .ZN(n16736) );
  OAI222_X1 U19808 ( .A1(n20830), .A2(n16738), .B1(n20834), .B2(n16737), .C1(
        n16736), .C2(n16735), .ZN(n16739) );
  OAI21_X1 U19809 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16740), .A(
        n16739), .ZN(n16748) );
  OAI21_X1 U19810 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16741), .ZN(n16742) );
  NAND4_X1 U19811 ( .A1(n16745), .A2(n16744), .A3(n16743), .A4(n16742), .ZN(
        n16746) );
  AOI211_X1 U19812 ( .C1(n20484), .C2(n16748), .A(n16747), .B(n16746), .ZN(
        n16763) );
  NAND3_X1 U19813 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21094), .A3(n21091), 
        .ZN(n16749) );
  AOI22_X1 U19814 ( .A1(n16752), .A2(n16751), .B1(n16750), .B2(n16749), .ZN(
        n16823) );
  OAI221_X1 U19815 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n16763), 
        .A(n16823), .ZN(n16830) );
  INV_X1 U19816 ( .A(n16753), .ZN(n16825) );
  NOR2_X1 U19817 ( .A1(n16825), .A2(n16754), .ZN(n16755) );
  NOR2_X1 U19818 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16755), .ZN(n16761) );
  INV_X1 U19819 ( .A(n16756), .ZN(n16757) );
  AOI211_X1 U19820 ( .C1(n21094), .C2(n13022), .A(n16758), .B(n16757), .ZN(
        n16759) );
  NAND2_X1 U19821 ( .A1(n16830), .A2(n16759), .ZN(n16760) );
  AOI22_X1 U19822 ( .A1(n16830), .A2(n16761), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16760), .ZN(n16762) );
  OAI21_X1 U19823 ( .B1(n16763), .B2(n20246), .A(n16762), .ZN(P1_U3161) );
  INV_X1 U19824 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20244) );
  NOR2_X1 U19825 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20244), .ZN(n21103) );
  INV_X1 U19826 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21101) );
  NOR2_X1 U19827 ( .A1(n21101), .A2(n21105), .ZN(n21100) );
  NAND2_X1 U19828 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n16764) );
  AOI22_X1 U19829 ( .A1(HOLD), .A2(n21103), .B1(n21100), .B2(n16764), .ZN(
        n16766) );
  OAI211_X1 U19830 ( .C1(n20244), .C2(n21102), .A(n16766), .B(n16765), .ZN(
        P1_U3195) );
  AND2_X1 U19831 ( .A1(n16767), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OR2_X1 U19832 ( .A1(n16769), .A2(n16768), .ZN(n16770) );
  AOI21_X4 U19833 ( .B1(n16771), .B2(n16770), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n20033) );
  OAI21_X1 U19834 ( .B1(n20216), .B2(n16773), .A(n16772), .ZN(n16774) );
  NOR2_X1 U19835 ( .A1(n20033), .A2(n16774), .ZN(n20214) );
  INV_X1 U19836 ( .A(n20214), .ZN(n20212) );
  NOR2_X1 U19837 ( .A1(n21284), .A2(n20212), .ZN(P2_U3047) );
  NOR3_X1 U19838 ( .A1(n16775), .A2(n17815), .A3(n19260), .ZN(n16776) );
  NOR2_X1 U19839 ( .A1(n17749), .A2(n17805), .ZN(n17706) );
  INV_X1 U19840 ( .A(n17706), .ZN(n17780) );
  INV_X1 U19841 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17885) );
  INV_X1 U19842 ( .A(n17805), .ZN(n16780) );
  NOR2_X1 U19843 ( .A1(n16778), .A2(n17806), .ZN(n17810) );
  NAND2_X1 U19844 ( .A1(n16778), .A2(n16780), .ZN(n17801) );
  AOI22_X1 U19845 ( .A1(n17810), .A2(BUF2_REG_0__SCAN_IN), .B1(n17809), .B2(
        n18288), .ZN(n16779) );
  OAI221_X1 U19846 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17780), .C1(n17885), 
        .C2(n16780), .A(n16779), .ZN(P3_U2735) );
  AOI21_X1 U19847 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n20272), .A(
        P1_REIP_REG_10__SCAN_IN), .ZN(n16789) );
  OAI22_X1 U19848 ( .A1(n21477), .A2(n16781), .B1(n20305), .B2(n21465), .ZN(
        n16782) );
  AOI211_X1 U19849 ( .C1(n16783), .C2(n20333), .A(n20296), .B(n16782), .ZN(
        n16788) );
  INV_X1 U19850 ( .A(n16784), .ZN(n16785) );
  AOI22_X1 U19851 ( .A1(n16786), .A2(n20298), .B1(n16785), .B2(n20344), .ZN(
        n16787) );
  OAI211_X1 U19852 ( .C1(n16790), .C2(n16789), .A(n16788), .B(n16787), .ZN(
        P1_U2830) );
  AOI22_X1 U19853 ( .A1(n20421), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20436), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16796) );
  NAND2_X1 U19854 ( .A1(n16793), .A2(n16792), .ZN(n16794) );
  XNOR2_X1 U19855 ( .A(n16791), .B(n16794), .ZN(n16808) );
  AOI22_X1 U19856 ( .A1(n20287), .A2(n20428), .B1(n16808), .B2(n20429), .ZN(
        n16795) );
  OAI211_X1 U19857 ( .C1(n20433), .C2(n20290), .A(n16796), .B(n16795), .ZN(
        P1_U2992) );
  AOI22_X1 U19858 ( .A1(n20421), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20436), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16801) );
  XNOR2_X1 U19859 ( .A(n16797), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16798) );
  XNOR2_X1 U19860 ( .A(n16799), .B(n16798), .ZN(n16817) );
  AOI22_X1 U19861 ( .A1(n20352), .A2(n20428), .B1(n16817), .B2(n20429), .ZN(
        n16800) );
  OAI211_X1 U19862 ( .C1(n20433), .C2(n20301), .A(n16801), .B(n16800), .ZN(
        P1_U2993) );
  AOI22_X1 U19863 ( .A1(n20421), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20436), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16806) );
  INV_X1 U19864 ( .A(n16802), .ZN(n16804) );
  INV_X1 U19865 ( .A(n16803), .ZN(n20311) );
  AOI22_X1 U19866 ( .A1(n20429), .A2(n16804), .B1(n20311), .B2(n20428), .ZN(
        n16805) );
  OAI211_X1 U19867 ( .C1(n20433), .C2(n20313), .A(n16806), .B(n16805), .ZN(
        P1_U2994) );
  INV_X1 U19868 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21122) );
  OAI22_X1 U19869 ( .A1(n20471), .A2(n20280), .B1(n21122), .B2(n20457), .ZN(
        n16807) );
  AOI21_X1 U19870 ( .B1(n16808), .B2(n20477), .A(n16807), .ZN(n16809) );
  OAI221_X1 U19871 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16812), .C1(
        n16811), .C2(n16810), .A(n16809), .ZN(P1_U3024) );
  INV_X1 U19872 ( .A(n16813), .ZN(n16815) );
  INV_X1 U19873 ( .A(n14256), .ZN(n16814) );
  AOI21_X1 U19874 ( .B1(n16815), .B2(n16814), .A(n9896), .ZN(n20349) );
  AOI22_X1 U19875 ( .A1(n20454), .A2(n20349), .B1(n20436), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16819) );
  AOI22_X1 U19876 ( .A1(n16817), .A2(n20477), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16816), .ZN(n16818) );
  OAI211_X1 U19877 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16820), .A(
        n16819), .B(n16818), .ZN(P1_U3025) );
  AOI21_X1 U19878 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16830), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16828) );
  NAND4_X1 U19879 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n13022), .A4(n21102), .ZN(n16821) );
  AND2_X1 U19880 ( .A1(n16822), .A2(n16821), .ZN(n21092) );
  AOI21_X1 U19881 ( .B1(n21092), .B2(n16824), .A(n16823), .ZN(n16827) );
  AOI21_X1 U19882 ( .B1(n20913), .B2(n21102), .A(n16825), .ZN(n16826) );
  NOR3_X1 U19883 ( .A1(n16828), .A2(n16827), .A3(n16826), .ZN(P1_U3162) );
  OAI221_X1 U19884 ( .B1(n20913), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20913), 
        .C2(n16830), .A(n16829), .ZN(P1_U3466) );
  AOI22_X1 U19885 ( .A1(n16833), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n16832), .B2(n16831), .ZN(n16845) );
  OAI21_X1 U19886 ( .B1(n16836), .B2(n16835), .A(n16834), .ZN(n16837) );
  INV_X1 U19887 ( .A(n16837), .ZN(n16840) );
  NAND2_X1 U19888 ( .A1(n16838), .A2(n19400), .ZN(n16839) );
  OAI211_X1 U19889 ( .C1(n16842), .C2(n16841), .A(n16840), .B(n16839), .ZN(
        n16843) );
  INV_X1 U19890 ( .A(n16843), .ZN(n16844) );
  OAI211_X1 U19891 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16846), .A(
        n16845), .B(n16844), .ZN(P2_U3046) );
  INV_X1 U19892 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19222) );
  NOR2_X1 U19893 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19222), .ZN(
        n16880) );
  NOR2_X1 U19894 ( .A1(n16847), .A2(n18117), .ZN(n16851) );
  NOR3_X1 U19895 ( .A1(n16880), .A2(n16851), .A3(n16848), .ZN(n16849) );
  AOI21_X1 U19896 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n19222), .A(
        n16849), .ZN(n16854) );
  AOI22_X1 U19897 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18199), .B1(
        n18117), .B2(n19222), .ZN(n16853) );
  OAI21_X1 U19898 ( .B1(n16851), .B2(n16850), .A(n16853), .ZN(n16852) );
  INV_X1 U19899 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19194) );
  NOR2_X1 U19900 ( .A1(n19194), .A2(n18481), .ZN(n16886) );
  XOR2_X1 U19901 ( .A(n10482), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16856) );
  OAI22_X1 U19902 ( .A1(n16857), .A2(n16856), .B1(n16855), .B2(n10482), .ZN(
        n16858) );
  AOI211_X1 U19903 ( .C1(n18145), .C2(n17362), .A(n16886), .B(n16858), .ZN(
        n16864) );
  NAND3_X1 U19904 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n19222), .ZN(n16881) );
  OAI21_X1 U19905 ( .B1(n16861), .B2(n16859), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16860) );
  OAI21_X1 U19906 ( .B1(n16867), .B2(n16881), .A(n16860), .ZN(n16888) );
  OAI21_X1 U19907 ( .B1(n16861), .B2(n16865), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16862) );
  OAI21_X1 U19908 ( .B1(n16881), .B2(n16896), .A(n16862), .ZN(n16889) );
  AOI22_X1 U19909 ( .A1(n18261), .A2(n16888), .B1(n18202), .B2(n16889), .ZN(
        n16863) );
  OAI211_X1 U19910 ( .C1(n16892), .C2(n18164), .A(n16864), .B(n16863), .ZN(
        P3_U2799) );
  NAND2_X1 U19911 ( .A1(n18202), .A2(n16865), .ZN(n16879) );
  AOI211_X1 U19912 ( .C1(n16867), .C2(n16878), .A(n16866), .B(n18293), .ZN(
        n16876) );
  AOI22_X1 U19913 ( .A1(n9732), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16868), .ZN(n16872) );
  INV_X1 U19914 ( .A(n17022), .ZN(n16869) );
  AOI21_X1 U19915 ( .B1(n10481), .B2(n16869), .A(n9894), .ZN(n17047) );
  OAI21_X1 U19916 ( .B1(n16870), .B2(n18145), .A(n17047), .ZN(n16871) );
  OAI211_X1 U19917 ( .C1(n16874), .C2(n16873), .A(n16872), .B(n16871), .ZN(
        n16875) );
  OAI221_X1 U19918 ( .B1(n16879), .B2(n16878), .C1(n16879), .C2(n16896), .A(
        n16877), .ZN(P3_U2801) );
  INV_X1 U19919 ( .A(n16880), .ZN(n16883) );
  OAI22_X1 U19920 ( .A1(n9743), .A2(n16883), .B1(n16882), .B2(n16881), .ZN(
        n16887) );
  AOI21_X1 U19921 ( .B1(n18581), .B2(n16884), .A(n19222), .ZN(n16885) );
  AOI211_X1 U19922 ( .C1(n18595), .C2(n16887), .A(n16886), .B(n16885), .ZN(
        n16891) );
  AOI22_X1 U19923 ( .A1(n18318), .A2(n16889), .B1(n18598), .B2(n16888), .ZN(
        n16890) );
  OAI211_X1 U19924 ( .C1(n16892), .C2(n18485), .A(n16891), .B(n16890), .ZN(
        P3_U2831) );
  OR4_X1 U19925 ( .A1(n18307), .A2(n18117), .A3(n16704), .A4(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16910) );
  NOR2_X1 U19926 ( .A1(n19055), .A2(n18586), .ZN(n18583) );
  INV_X1 U19927 ( .A(n18583), .ZN(n18602) );
  OAI211_X1 U19928 ( .C1(n16894), .C2(n18574), .A(n16893), .B(n18581), .ZN(
        n16895) );
  AOI21_X1 U19929 ( .B1(n18452), .B2(n16896), .A(n16895), .ZN(n16899) );
  INV_X1 U19930 ( .A(n17940), .ZN(n16907) );
  AOI22_X1 U19931 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18199), .B1(
        n18117), .B2(n17921), .ZN(n17934) );
  NAND2_X1 U19932 ( .A1(n17935), .A2(n17934), .ZN(n17933) );
  NAND3_X1 U19933 ( .A1(n18514), .A2(n16897), .A3(n17933), .ZN(n16898) );
  AOI21_X1 U19934 ( .B1(n16899), .B2(n16898), .A(n17921), .ZN(n16906) );
  INV_X1 U19935 ( .A(n16900), .ZN(n16904) );
  INV_X1 U19936 ( .A(n16901), .ZN(n18473) );
  INV_X1 U19937 ( .A(n18475), .ZN(n18160) );
  OAI22_X1 U19938 ( .A1(n18473), .A2(n18574), .B1(n18160), .B2(n18508), .ZN(
        n18399) );
  AOI21_X1 U19939 ( .B1(n16902), .B2(n18399), .A(n18320), .ZN(n18345) );
  NOR2_X2 U19940 ( .A1(n18345), .A2(n18586), .ZN(n18365) );
  NAND2_X1 U19941 ( .A1(n16903), .A2(n18365), .ZN(n18351) );
  NOR4_X1 U19942 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18307), .A3(
        n16904), .A4(n18351), .ZN(n16905) );
  AOI221_X2 U19943 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n9732), .C1(n16906), 
        .C2(n18481), .A(n16905), .ZN(n16909) );
  OR3_X1 U19944 ( .A1(n16907), .A2(n18485), .A3(n17934), .ZN(n16908) );
  OAI211_X1 U19945 ( .C1(n16910), .C2(n18602), .A(n16909), .B(n16908), .ZN(
        P3_U2834) );
  NOR3_X1 U19946 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16912) );
  NOR4_X1 U19947 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16911) );
  NAND4_X1 U19948 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16912), .A3(n16911), .A4(
        U215), .ZN(U213) );
  NOR2_X1 U19949 ( .A1(n16957), .A2(n16913), .ZN(n16958) );
  AOI222_X1 U19950 ( .A1(n16947), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(n16958), 
        .B2(BUF1_REG_31__SCAN_IN), .C1(n16957), .C2(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n16914) );
  INV_X1 U19951 ( .A(n16914), .ZN(U216) );
  INV_X1 U19952 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19540) );
  AOI22_X1 U19953 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16947), .ZN(n16915) );
  OAI21_X1 U19954 ( .B1(n19540), .B2(n16954), .A(n16915), .ZN(U217) );
  INV_X1 U19955 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n19533) );
  AOI22_X1 U19956 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16947), .ZN(n16916) );
  OAI21_X1 U19957 ( .B1(n19533), .B2(n16954), .A(n16916), .ZN(U218) );
  INV_X1 U19958 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19528) );
  AOI22_X1 U19959 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16947), .ZN(n16917) );
  OAI21_X1 U19960 ( .B1(n19528), .B2(n16954), .A(n16917), .ZN(U219) );
  INV_X1 U19961 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U19962 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16947), .ZN(n16918) );
  OAI21_X1 U19963 ( .B1(n16919), .B2(n16954), .A(n16918), .ZN(U220) );
  AOI222_X1 U19964 ( .A1(n16947), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(n16958), 
        .B2(BUF1_REG_26__SCAN_IN), .C1(n16957), .C2(P1_DATAO_REG_26__SCAN_IN), 
        .ZN(n16920) );
  INV_X1 U19965 ( .A(n16920), .ZN(U221) );
  INV_X1 U19966 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n21320) );
  AOI22_X1 U19967 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16947), .ZN(n16921) );
  OAI21_X1 U19968 ( .B1(n21320), .B2(n16954), .A(n16921), .ZN(U222) );
  INV_X1 U19969 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n19500) );
  AOI22_X1 U19970 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16947), .ZN(n16922) );
  OAI21_X1 U19971 ( .B1(n19500), .B2(n16954), .A(n16922), .ZN(U223) );
  INV_X1 U19972 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n21421) );
  AOI22_X1 U19973 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16947), .ZN(n16923) );
  OAI21_X1 U19974 ( .B1(n21421), .B2(n16954), .A(n16923), .ZN(U224) );
  INV_X1 U19975 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n21300) );
  AOI22_X1 U19976 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16947), .ZN(n16924) );
  OAI21_X1 U19977 ( .B1(n21300), .B2(n16954), .A(n16924), .ZN(U225) );
  AOI222_X1 U19978 ( .A1(n16947), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(n16958), 
        .B2(BUF1_REG_21__SCAN_IN), .C1(n16957), .C2(P1_DATAO_REG_21__SCAN_IN), 
        .ZN(n16925) );
  INV_X1 U19979 ( .A(n16925), .ZN(U226) );
  INV_X1 U19980 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U19981 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16947), .ZN(n16926) );
  OAI21_X1 U19982 ( .B1(n16927), .B2(n16954), .A(n16926), .ZN(U227) );
  INV_X1 U19983 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U19984 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16947), .ZN(n16928) );
  OAI21_X1 U19985 ( .B1(n16929), .B2(n16954), .A(n16928), .ZN(U228) );
  INV_X1 U19986 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U19987 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16947), .ZN(n16930) );
  OAI21_X1 U19988 ( .B1(n16931), .B2(n16954), .A(n16930), .ZN(U229) );
  INV_X1 U19989 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19512) );
  AOI22_X1 U19990 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16947), .ZN(n16932) );
  OAI21_X1 U19991 ( .B1(n19512), .B2(n16954), .A(n16932), .ZN(U230) );
  INV_X1 U19992 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U19993 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16947), .ZN(n16933) );
  OAI21_X1 U19994 ( .B1(n16934), .B2(n16954), .A(n16933), .ZN(U231) );
  AOI22_X1 U19995 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16947), .ZN(n16935) );
  OAI21_X1 U19996 ( .B1(n13117), .B2(n16954), .A(n16935), .ZN(U232) );
  AOI22_X1 U19997 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16947), .ZN(n16936) );
  OAI21_X1 U19998 ( .B1(n13270), .B2(n16954), .A(n16936), .ZN(U233) );
  AOI22_X1 U19999 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16947), .ZN(n16937) );
  OAI21_X1 U20000 ( .B1(n14937), .B2(n16954), .A(n16937), .ZN(U234) );
  AOI22_X1 U20001 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16947), .ZN(n16938) );
  OAI21_X1 U20002 ( .B1(n14247), .B2(n16954), .A(n16938), .ZN(U235) );
  AOI22_X1 U20003 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16947), .ZN(n16939) );
  OAI21_X1 U20004 ( .B1(n16940), .B2(n16954), .A(n16939), .ZN(U236) );
  AOI22_X1 U20005 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16947), .ZN(n16941) );
  OAI21_X1 U20006 ( .B1(n16942), .B2(n16954), .A(n16941), .ZN(U237) );
  AOI22_X1 U20007 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16947), .ZN(n16943) );
  OAI21_X1 U20008 ( .B1(n14953), .B2(n16954), .A(n16943), .ZN(U238) );
  AOI22_X1 U20009 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16947), .ZN(n16944) );
  OAI21_X1 U20010 ( .B1(n16945), .B2(n16954), .A(n16944), .ZN(U239) );
  INV_X1 U20011 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n21281) );
  AOI22_X1 U20012 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16958), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16947), .ZN(n16946) );
  OAI21_X1 U20013 ( .B1(n21281), .B2(U214), .A(n16946), .ZN(U240) );
  AOI22_X1 U20014 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16947), .ZN(n16948) );
  OAI21_X1 U20015 ( .B1(n16949), .B2(n16954), .A(n16948), .ZN(U241) );
  INV_X1 U20016 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20017 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16958), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16957), .ZN(n16950) );
  OAI21_X1 U20018 ( .B1(n16964), .B2(U212), .A(n16950), .ZN(U242) );
  INV_X1 U20019 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16963) );
  INV_X1 U20020 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16951) );
  INV_X1 U20021 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n21287) );
  OAI222_X1 U20022 ( .A1(U212), .A2(n16963), .B1(n16954), .B2(n16951), .C1(
        U214), .C2(n21287), .ZN(U243) );
  INV_X1 U20023 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20024 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16958), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16957), .ZN(n16952) );
  OAI21_X1 U20025 ( .B1(n16962), .B2(U212), .A(n16952), .ZN(U244) );
  INV_X1 U20026 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16955) );
  AOI22_X1 U20027 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16957), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16947), .ZN(n16953) );
  OAI21_X1 U20028 ( .B1(n16955), .B2(n16954), .A(n16953), .ZN(U245) );
  INV_X1 U20029 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n21402) );
  AOI22_X1 U20030 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16958), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16957), .ZN(n16956) );
  OAI21_X1 U20031 ( .B1(n21402), .B2(U212), .A(n16956), .ZN(U246) );
  INV_X1 U20032 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20033 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16958), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16957), .ZN(n16959) );
  OAI21_X1 U20034 ( .B1(n16960), .B2(U212), .A(n16959), .ZN(U247) );
  INV_X1 U20035 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18612) );
  AOI22_X1 U20036 ( .A1(n16990), .A2(n16960), .B1(n18612), .B2(U215), .ZN(U251) );
  INV_X1 U20037 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18620) );
  AOI22_X1 U20038 ( .A1(n16990), .A2(n21402), .B1(n18620), .B2(U215), .ZN(U252) );
  INV_X1 U20039 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U20040 ( .A1(n16990), .A2(n16961), .B1(n18624), .B2(U215), .ZN(U253) );
  INV_X1 U20041 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18628) );
  AOI22_X1 U20042 ( .A1(n16990), .A2(n16962), .B1(n18628), .B2(U215), .ZN(U254) );
  INV_X1 U20043 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21290) );
  AOI22_X1 U20044 ( .A1(n16990), .A2(n16963), .B1(n21290), .B2(U215), .ZN(U255) );
  AOI22_X1 U20045 ( .A1(n16989), .A2(n16964), .B1(n13138), .B2(U215), .ZN(U256) );
  INV_X1 U20046 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20047 ( .A1(n16989), .A2(n16965), .B1(n12944), .B2(U215), .ZN(U257) );
  INV_X1 U20048 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20049 ( .A1(n16990), .A2(n16966), .B1(n13056), .B2(U215), .ZN(U258) );
  INV_X1 U20050 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U20051 ( .A1(n16989), .A2(n16967), .B1(n17778), .B2(U215), .ZN(U259) );
  INV_X1 U20052 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20053 ( .A1(n16990), .A2(n16968), .B1(n13132), .B2(U215), .ZN(U260) );
  INV_X1 U20054 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20055 ( .A1(n16989), .A2(n16969), .B1(n17768), .B2(U215), .ZN(U261) );
  OAI22_X1 U20056 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16990), .ZN(n16970) );
  INV_X1 U20057 ( .A(n16970), .ZN(U262) );
  INV_X1 U20058 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20059 ( .A1(n16989), .A2(n16971), .B1(n13126), .B2(U215), .ZN(U263) );
  INV_X1 U20060 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20061 ( .A1(n16990), .A2(n16972), .B1(n13123), .B2(U215), .ZN(U264) );
  OAI22_X1 U20062 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16990), .ZN(n16973) );
  INV_X1 U20063 ( .A(n16973), .ZN(U265) );
  OAI22_X1 U20064 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16990), .ZN(n16974) );
  INV_X1 U20065 ( .A(n16974), .ZN(U266) );
  OAI22_X1 U20066 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16990), .ZN(n16975) );
  INV_X1 U20067 ( .A(n16975), .ZN(U267) );
  INV_X1 U20068 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20069 ( .A1(n16990), .A2(n16976), .B1(n15998), .B2(U215), .ZN(U268) );
  OAI22_X1 U20070 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16990), .ZN(n16977) );
  INV_X1 U20071 ( .A(n16977), .ZN(U269) );
  OAI22_X1 U20072 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16989), .ZN(n16978) );
  INV_X1 U20073 ( .A(n16978), .ZN(U270) );
  OAI22_X1 U20074 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16989), .ZN(n16979) );
  INV_X1 U20075 ( .A(n16979), .ZN(U271) );
  INV_X1 U20076 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16980) );
  INV_X1 U20077 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18635) );
  AOI22_X1 U20078 ( .A1(n16990), .A2(n16980), .B1(n18635), .B2(U215), .ZN(U272) );
  INV_X1 U20079 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20080 ( .A1(n16990), .A2(n16981), .B1(n15963), .B2(U215), .ZN(U273) );
  OAI22_X1 U20081 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16989), .ZN(n16982) );
  INV_X1 U20082 ( .A(n16982), .ZN(U274) );
  INV_X1 U20083 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20084 ( .A1(n16990), .A2(n16983), .B1(n15948), .B2(U215), .ZN(U275) );
  OAI22_X1 U20085 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16990), .ZN(n16984) );
  INV_X1 U20086 ( .A(n16984), .ZN(U276) );
  OAI22_X1 U20087 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16990), .ZN(n16985) );
  INV_X1 U20088 ( .A(n16985), .ZN(U277) );
  OAI22_X1 U20089 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16990), .ZN(n16986) );
  INV_X1 U20090 ( .A(n16986), .ZN(U278) );
  INV_X1 U20091 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20092 ( .A1(n16989), .A2(n16987), .B1(n15926), .B2(U215), .ZN(U279) );
  INV_X1 U20093 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20094 ( .A1(n16990), .A2(n16988), .B1(n15917), .B2(U215), .ZN(U280) );
  INV_X1 U20095 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20096 ( .A1(n16989), .A2(n16993), .B1(n12431), .B2(U215), .ZN(U281) );
  OAI22_X1 U20097 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16990), .ZN(n16991) );
  INV_X1 U20098 ( .A(n16991), .ZN(U282) );
  INV_X1 U20099 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16994) );
  INV_X1 U20100 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16992) );
  OAI222_X1 U20101 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n16994), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n16993), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n16992), .ZN(n16995) );
  INV_X2 U20102 ( .A(n21188), .ZN(n21189) );
  INV_X1 U20103 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n21381) );
  INV_X1 U20104 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20126) );
  AOI22_X1 U20105 ( .A1(n21189), .A2(n21381), .B1(n20126), .B2(n21188), .ZN(
        U347) );
  INV_X1 U20106 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19154) );
  INV_X1 U20107 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20124) );
  AOI22_X1 U20108 ( .A1(n21189), .A2(n19154), .B1(n20124), .B2(n21188), .ZN(
        U348) );
  INV_X1 U20109 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19151) );
  INV_X1 U20110 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U20111 ( .A1(n21189), .A2(n19151), .B1(n20122), .B2(n21188), .ZN(
        U349) );
  INV_X1 U20112 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19150) );
  INV_X1 U20113 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20120) );
  AOI22_X1 U20114 ( .A1(n21189), .A2(n19150), .B1(n20120), .B2(n21188), .ZN(
        U350) );
  INV_X1 U20115 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19145) );
  INV_X1 U20116 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20116) );
  AOI22_X1 U20117 ( .A1(n21189), .A2(n19145), .B1(n20116), .B2(n21188), .ZN(
        U352) );
  INV_X1 U20118 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19144) );
  INV_X1 U20119 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20115) );
  AOI22_X1 U20120 ( .A1(n21189), .A2(n19144), .B1(n20115), .B2(n21188), .ZN(
        U353) );
  INV_X1 U20121 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19142) );
  AOI22_X1 U20122 ( .A1(n21189), .A2(n19142), .B1(n20113), .B2(n21188), .ZN(
        U354) );
  INV_X1 U20123 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19195) );
  INV_X1 U20124 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20164) );
  AOI22_X1 U20125 ( .A1(n21189), .A2(n19195), .B1(n20164), .B2(n21188), .ZN(
        U355) );
  INV_X1 U20126 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19191) );
  INV_X1 U20127 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20160) );
  AOI22_X1 U20128 ( .A1(n21189), .A2(n19191), .B1(n20160), .B2(n21188), .ZN(
        U356) );
  INV_X1 U20129 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19188) );
  INV_X1 U20130 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n21240) );
  AOI22_X1 U20131 ( .A1(n21189), .A2(n19188), .B1(n21240), .B2(n16995), .ZN(
        U357) );
  INV_X1 U20132 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19187) );
  INV_X1 U20133 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20155) );
  AOI22_X1 U20134 ( .A1(n21189), .A2(n19187), .B1(n20155), .B2(n21188), .ZN(
        U358) );
  INV_X1 U20135 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19185) );
  INV_X1 U20136 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20154) );
  AOI22_X1 U20137 ( .A1(n21189), .A2(n19185), .B1(n20154), .B2(n16995), .ZN(
        U359) );
  INV_X1 U20138 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19183) );
  INV_X1 U20139 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20152) );
  AOI22_X1 U20140 ( .A1(n21189), .A2(n19183), .B1(n20152), .B2(n21188), .ZN(
        U360) );
  INV_X1 U20141 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19181) );
  INV_X1 U20142 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U20143 ( .A1(n21189), .A2(n19181), .B1(n20150), .B2(n21188), .ZN(
        U361) );
  INV_X1 U20144 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19179) );
  INV_X1 U20145 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n21337) );
  AOI22_X1 U20146 ( .A1(n21189), .A2(n19179), .B1(n21337), .B2(n21188), .ZN(
        U362) );
  INV_X1 U20147 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19177) );
  INV_X1 U20148 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20148) );
  AOI22_X1 U20149 ( .A1(n21189), .A2(n19177), .B1(n20148), .B2(n21188), .ZN(
        U363) );
  INV_X1 U20150 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19176) );
  INV_X1 U20151 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20146) );
  AOI22_X1 U20152 ( .A1(n21189), .A2(n19176), .B1(n20146), .B2(n21188), .ZN(
        U364) );
  INV_X1 U20153 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19140) );
  INV_X1 U20154 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20111) );
  AOI22_X1 U20155 ( .A1(n21189), .A2(n19140), .B1(n20111), .B2(n21188), .ZN(
        U365) );
  INV_X1 U20156 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19174) );
  INV_X1 U20157 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20144) );
  AOI22_X1 U20158 ( .A1(n21189), .A2(n19174), .B1(n20144), .B2(n21188), .ZN(
        U366) );
  INV_X1 U20159 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19172) );
  INV_X1 U20160 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20142) );
  AOI22_X1 U20161 ( .A1(n21189), .A2(n19172), .B1(n20142), .B2(n16995), .ZN(
        U367) );
  INV_X1 U20162 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19170) );
  INV_X1 U20163 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n21316) );
  AOI22_X1 U20164 ( .A1(n21189), .A2(n19170), .B1(n21316), .B2(n16995), .ZN(
        U368) );
  INV_X1 U20165 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19167) );
  INV_X1 U20166 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U20167 ( .A1(n21189), .A2(n19167), .B1(n20139), .B2(n16995), .ZN(
        U369) );
  INV_X1 U20168 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19166) );
  INV_X1 U20169 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20137) );
  AOI22_X1 U20170 ( .A1(n21189), .A2(n19166), .B1(n20137), .B2(n16995), .ZN(
        U370) );
  INV_X1 U20171 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19164) );
  INV_X1 U20172 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20135) );
  AOI22_X1 U20173 ( .A1(n21189), .A2(n19164), .B1(n20135), .B2(n16995), .ZN(
        U371) );
  INV_X1 U20174 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19162) );
  INV_X1 U20175 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20133) );
  AOI22_X1 U20176 ( .A1(n21189), .A2(n19162), .B1(n20133), .B2(n16995), .ZN(
        U372) );
  INV_X1 U20177 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19161) );
  INV_X1 U20178 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20131) );
  AOI22_X1 U20179 ( .A1(n21189), .A2(n19161), .B1(n20131), .B2(n21188), .ZN(
        U373) );
  INV_X1 U20180 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19159) );
  INV_X1 U20181 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U20182 ( .A1(n21189), .A2(n19159), .B1(n20130), .B2(n21188), .ZN(
        U374) );
  INV_X1 U20183 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19157) );
  INV_X1 U20184 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20128) );
  AOI22_X1 U20185 ( .A1(n21189), .A2(n19157), .B1(n20128), .B2(n21188), .ZN(
        U375) );
  INV_X1 U20186 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19138) );
  INV_X1 U20187 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20109) );
  AOI22_X1 U20188 ( .A1(n21189), .A2(n19138), .B1(n20109), .B2(n21188), .ZN(
        U376) );
  INV_X1 U20189 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16996) );
  INV_X1 U20190 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19137) );
  NAND2_X1 U20191 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19137), .ZN(n19129) );
  AOI21_X1 U20192 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n19129), .A(n19272), 
        .ZN(n19208) );
  INV_X1 U20193 ( .A(n19208), .ZN(n19204) );
  OAI21_X1 U20194 ( .B1(n16996), .B2(n19134), .A(n19204), .ZN(P3_U2633) );
  OAI21_X1 U20195 ( .B1(n17004), .B2(n17853), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16997) );
  OAI21_X1 U20196 ( .B1(n16998), .B2(n19105), .A(n16997), .ZN(P3_U2634) );
  AOI21_X1 U20197 ( .B1(n19134), .B2(n19137), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16999) );
  AOI22_X1 U20198 ( .A1(n19272), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16999), 
        .B2(n19270), .ZN(P3_U2635) );
  OAI21_X1 U20199 ( .B1(n17000), .B2(BS16), .A(n19208), .ZN(n19206) );
  OAI21_X1 U20200 ( .B1(n19208), .B2(n17001), .A(n19206), .ZN(P3_U2636) );
  NOR3_X1 U20201 ( .A1(n17004), .A2(n17003), .A3(n17002), .ZN(n19098) );
  NOR2_X1 U20202 ( .A1(n19098), .A2(n19102), .ZN(n19250) );
  OAI21_X1 U20203 ( .B1(n19250), .B2(n17006), .A(n17005), .ZN(P3_U2637) );
  NOR4_X1 U20204 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17010) );
  NOR4_X1 U20205 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17009) );
  NOR4_X1 U20206 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17008) );
  NOR4_X1 U20207 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17007) );
  NAND4_X1 U20208 ( .A1(n17010), .A2(n17009), .A3(n17008), .A4(n17007), .ZN(
        n17016) );
  NOR4_X1 U20209 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17014) );
  AOI211_X1 U20210 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_10__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17013) );
  NOR4_X1 U20211 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17012) );
  NOR4_X1 U20212 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n17011) );
  NAND4_X1 U20213 ( .A1(n17014), .A2(n17013), .A3(n17012), .A4(n17011), .ZN(
        n17015) );
  NOR2_X1 U20214 ( .A1(n17016), .A2(n17015), .ZN(n19245) );
  INV_X1 U20215 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19201) );
  NOR3_X1 U20216 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17018) );
  OAI21_X1 U20217 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17018), .A(n19245), .ZN(
        n17017) );
  OAI21_X1 U20218 ( .B1(n19245), .B2(n19201), .A(n17017), .ZN(P3_U2638) );
  INV_X1 U20219 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19241) );
  INV_X1 U20220 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19207) );
  AOI21_X1 U20221 ( .B1(n19241), .B2(n19207), .A(n17018), .ZN(n17019) );
  INV_X1 U20222 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19198) );
  INV_X1 U20223 ( .A(n19245), .ZN(n19247) );
  AOI22_X1 U20224 ( .A1(n19245), .A2(n17019), .B1(n19198), .B2(n19247), .ZN(
        P3_U2639) );
  INV_X1 U20225 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19196) );
  NOR2_X1 U20226 ( .A1(n19184), .A2(n17020), .ZN(n17056) );
  NAND4_X1 U20227 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17056), .ZN(n17029) );
  NOR3_X1 U20228 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19196), .A3(n17029), 
        .ZN(n17021) );
  AOI21_X1 U20229 ( .B1(n17377), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17021), .ZN(
        n17038) );
  NAND3_X1 U20230 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n12629), .A3(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17023) );
  AOI21_X1 U20231 ( .B1(n17922), .B2(n17023), .A(n17022), .ZN(n17932) );
  OAI21_X1 U20232 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17024), .A(
        n17023), .ZN(n17025) );
  INV_X1 U20233 ( .A(n17025), .ZN(n17942) );
  NOR2_X1 U20234 ( .A1(n17026), .A2(n17294), .ZN(n17068) );
  NOR2_X1 U20235 ( .A1(n17942), .A2(n17068), .ZN(n17067) );
  NOR2_X1 U20236 ( .A1(n17067), .A2(n17294), .ZN(n17060) );
  NOR2_X1 U20237 ( .A1(n17932), .A2(n17060), .ZN(n17059) );
  NOR2_X1 U20238 ( .A1(n17059), .A2(n17294), .ZN(n17046) );
  NOR2_X1 U20239 ( .A1(n17047), .A2(n17046), .ZN(n17045) );
  INV_X1 U20240 ( .A(n17040), .ZN(n17036) );
  OR2_X1 U20241 ( .A1(n17041), .A2(n19118), .ZN(n17027) );
  INV_X1 U20242 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17411) );
  NAND2_X1 U20243 ( .A1(n17058), .A2(n17384), .ZN(n17039) );
  INV_X1 U20244 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17390) );
  NAND2_X1 U20245 ( .A1(n17372), .A2(n17366), .ZN(n17375) );
  NAND3_X1 U20246 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n17028) );
  AOI21_X1 U20247 ( .B1(n17375), .B2(n17028), .A(n17072), .ZN(n17055) );
  NOR2_X1 U20248 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17029), .ZN(n17043) );
  INV_X1 U20249 ( .A(n17043), .ZN(n17030) );
  AOI21_X1 U20250 ( .B1(n17055), .B2(n17030), .A(n19194), .ZN(n17031) );
  INV_X1 U20251 ( .A(n17031), .ZN(n17032) );
  OAI211_X1 U20252 ( .C1(n10482), .C2(n17363), .A(n17038), .B(n17037), .ZN(
        P3_U2640) );
  NAND2_X1 U20253 ( .A1(n17376), .A2(n17039), .ZN(n17051) );
  OAI22_X1 U20254 ( .A1(n17055), .A2(n19196), .B1(n10483), .B2(n17363), .ZN(
        n17042) );
  INV_X1 U20255 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21459) );
  AOI211_X1 U20256 ( .C1(n17047), .C2(n17046), .A(n17045), .B(n19118), .ZN(
        n17050) );
  NAND3_X1 U20257 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17056), .ZN(n17048) );
  OAI22_X1 U20258 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17048), .B1(n10481), 
        .B2(n17363), .ZN(n17049) );
  AOI211_X1 U20259 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17377), .A(n17050), .B(
        n17049), .ZN(n17054) );
  INV_X1 U20260 ( .A(n17051), .ZN(n17052) );
  OAI21_X1 U20261 ( .B1(n17058), .B2(n17384), .A(n17052), .ZN(n17053) );
  OAI211_X1 U20262 ( .C1(n17055), .C2(n21459), .A(n17054), .B(n17053), .ZN(
        P3_U2642) );
  NAND2_X1 U20263 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17056), .ZN(n17066) );
  AOI22_X1 U20264 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17345), .B1(
        n17377), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17065) );
  INV_X1 U20265 ( .A(n17056), .ZN(n17077) );
  OAI21_X1 U20266 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n17077), .A(n17057), 
        .ZN(n17063) );
  AOI211_X1 U20267 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17073), .A(n17058), .B(
        n17365), .ZN(n17062) );
  AOI211_X1 U20268 ( .C1(n17932), .C2(n17060), .A(n17059), .B(n19118), .ZN(
        n17061) );
  OAI211_X1 U20269 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17066), .A(n17065), 
        .B(n17064), .ZN(P3_U2643) );
  AOI211_X1 U20270 ( .C1(n17942), .C2(n17068), .A(n17067), .B(n19118), .ZN(
        n17071) );
  AOI22_X1 U20271 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17345), .B1(
        n17377), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n17069) );
  INV_X1 U20272 ( .A(n17069), .ZN(n17070) );
  AOI211_X1 U20273 ( .C1(n17072), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17071), 
        .B(n17070), .ZN(n17076) );
  OAI211_X1 U20274 ( .C1(n17074), .C2(n17411), .A(n17376), .B(n17073), .ZN(
        n17075) );
  OAI211_X1 U20275 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17077), .A(n17076), 
        .B(n17075), .ZN(P3_U2644) );
  INV_X1 U20276 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19180) );
  OAI21_X1 U20277 ( .B1(n17089), .B2(n17366), .A(n17372), .ZN(n17102) );
  AOI21_X1 U20278 ( .B1(n17353), .B2(n19180), .A(n17102), .ZN(n17087) );
  AOI211_X1 U20279 ( .C1(n17968), .C2(n17079), .A(n17078), .B(n19118), .ZN(
        n17083) );
  NOR3_X1 U20280 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17366), .A3(n17080), 
        .ZN(n17082) );
  OAI22_X1 U20281 ( .A1(n17965), .A2(n17363), .B1(n17334), .B2(n17383), .ZN(
        n17081) );
  NOR3_X1 U20282 ( .A1(n17083), .A2(n17082), .A3(n17081), .ZN(n17086) );
  OAI211_X1 U20283 ( .C1(n17090), .C2(n17383), .A(n17376), .B(n17084), .ZN(
        n17085) );
  OAI211_X1 U20284 ( .C1(n17087), .C2(n19182), .A(n17086), .B(n17085), .ZN(
        P3_U2646) );
  NOR2_X1 U20285 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17366), .ZN(n17088) );
  AOI22_X1 U20286 ( .A1(n17377), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17089), 
        .B2(n17088), .ZN(n17096) );
  AOI211_X1 U20287 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17103), .A(n17090), .B(
        n17365), .ZN(n17094) );
  AOI211_X1 U20288 ( .C1(n17981), .C2(n17092), .A(n17091), .B(n19118), .ZN(
        n17093) );
  AOI211_X1 U20289 ( .C1(n17102), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17094), 
        .B(n17093), .ZN(n17095) );
  OAI211_X1 U20290 ( .C1(n17978), .C2(n17363), .A(n17096), .B(n17095), .ZN(
        P3_U2647) );
  OAI21_X1 U20291 ( .B1(n17366), .B2(n17097), .A(n19178), .ZN(n17101) );
  AOI211_X1 U20292 ( .C1(n17997), .C2(n10485), .A(n17098), .B(n19118), .ZN(
        n17100) );
  OAI22_X1 U20293 ( .A1(n17993), .A2(n17363), .B1(n17334), .B2(n17104), .ZN(
        n17099) );
  AOI211_X1 U20294 ( .C1(n17102), .C2(n17101), .A(n17100), .B(n17099), .ZN(
        n17106) );
  OAI211_X1 U20295 ( .C1(n17109), .C2(n17104), .A(n17376), .B(n17103), .ZN(
        n17105) );
  NAND2_X1 U20296 ( .A1(n17106), .A2(n17105), .ZN(P3_U2648) );
  NOR2_X1 U20297 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17366), .ZN(n17107) );
  AOI22_X1 U20298 ( .A1(n17377), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n17108), 
        .B2(n17107), .ZN(n17116) );
  AOI21_X1 U20299 ( .B1(n17353), .B2(n17127), .A(n17373), .ZN(n17118) );
  OAI21_X1 U20300 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n17366), .A(n17118), 
        .ZN(n17114) );
  AOI211_X1 U20301 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17123), .A(n17109), .B(
        n17365), .ZN(n17113) );
  AOI211_X1 U20302 ( .C1(n18009), .C2(n17111), .A(n17110), .B(n19118), .ZN(
        n17112) );
  AOI211_X1 U20303 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17114), .A(n17113), 
        .B(n17112), .ZN(n17115) );
  OAI211_X1 U20304 ( .C1(n17117), .C2(n17363), .A(n17116), .B(n17115), .ZN(
        P3_U2649) );
  NAND2_X1 U20305 ( .A1(n17353), .A2(n19175), .ZN(n17128) );
  INV_X1 U20306 ( .A(n17118), .ZN(n17134) );
  AOI211_X1 U20307 ( .C1(n18022), .C2(n17120), .A(n17119), .B(n19118), .ZN(
        n17122) );
  INV_X1 U20308 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18025) );
  OAI22_X1 U20309 ( .A1(n18025), .A2(n17363), .B1(n17334), .B2(n17124), .ZN(
        n17121) );
  AOI211_X1 U20310 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n17134), .A(n17122), 
        .B(n17121), .ZN(n17126) );
  OAI211_X1 U20311 ( .C1(n17131), .C2(n17124), .A(n17376), .B(n17123), .ZN(
        n17125) );
  OAI211_X1 U20312 ( .C1(n17128), .C2(n17127), .A(n17126), .B(n17125), .ZN(
        P3_U2650) );
  AOI211_X1 U20313 ( .C1(n18035), .C2(n17130), .A(n17129), .B(n19118), .ZN(
        n17133) );
  AOI211_X1 U20314 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17148), .A(n17131), .B(
        n17365), .ZN(n17132) );
  AOI211_X1 U20315 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17377), .A(n17133), .B(
        n17132), .ZN(n17137) );
  OAI221_X1 U20316 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n17353), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(n17135), .A(n17134), .ZN(n17136) );
  OAI211_X1 U20317 ( .C1(n17363), .C2(n17138), .A(n17137), .B(n17136), .ZN(
        P3_U2651) );
  INV_X1 U20318 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18052) );
  AOI21_X1 U20319 ( .B1(n17143), .B2(n17353), .A(n17373), .ZN(n17168) );
  INV_X1 U20320 ( .A(n17168), .ZN(n17158) );
  INV_X1 U20321 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18061) );
  NOR2_X1 U20322 ( .A1(n18285), .A2(n17139), .ZN(n17164) );
  NAND2_X1 U20323 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17164), .ZN(
        n18050) );
  NOR2_X1 U20324 ( .A1(n18061), .A2(n18050), .ZN(n17155) );
  OAI21_X1 U20325 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17155), .A(
        n18007), .ZN(n18048) );
  INV_X1 U20326 ( .A(n17155), .ZN(n17140) );
  NAND2_X1 U20327 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9917), .ZN(
        n17186) );
  INV_X1 U20328 ( .A(n17186), .ZN(n18083) );
  INV_X1 U20329 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21451) );
  NAND3_X1 U20330 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18083), .A3(
        n21451), .ZN(n17176) );
  OAI21_X1 U20331 ( .B1(n17140), .B2(n17176), .A(n17362), .ZN(n17142) );
  OAI21_X1 U20332 ( .B1(n18048), .B2(n17142), .A(n17338), .ZN(n17141) );
  AOI21_X1 U20333 ( .B1(n18048), .B2(n17142), .A(n17141), .ZN(n17147) );
  NOR2_X1 U20334 ( .A1(n17366), .A2(n17143), .ZN(n17154) );
  OAI211_X1 U20335 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n17154), .B(n17144), .ZN(n17145) );
  OAI211_X1 U20336 ( .C1(n17334), .C2(n17149), .A(n18481), .B(n17145), .ZN(
        n17146) );
  AOI211_X1 U20337 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n17158), .A(n17147), 
        .B(n17146), .ZN(n17151) );
  OAI211_X1 U20338 ( .C1(n17152), .C2(n17149), .A(n17376), .B(n17148), .ZN(
        n17150) );
  OAI211_X1 U20339 ( .C1(n17363), .C2(n18052), .A(n17151), .B(n17150), .ZN(
        P3_U2652) );
  AOI22_X1 U20340 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17345), .B1(
        n17377), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n17162) );
  INV_X1 U20341 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19169) );
  AOI211_X1 U20342 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17170), .A(n17152), .B(
        n17365), .ZN(n17153) );
  AOI211_X1 U20343 ( .C1(n17154), .C2(n19169), .A(n9732), .B(n17153), .ZN(
        n17161) );
  AOI21_X1 U20344 ( .B1(n18061), .B2(n18050), .A(n17155), .ZN(n18064) );
  AOI21_X1 U20345 ( .B1(n17156), .B2(n17199), .A(n17294), .ZN(n17157) );
  XOR2_X1 U20346 ( .A(n18064), .B(n17157), .Z(n17159) );
  AOI22_X1 U20347 ( .A1(n17338), .A2(n17159), .B1(P3_REIP_REG_18__SCAN_IN), 
        .B2(n17158), .ZN(n17160) );
  NAND3_X1 U20348 ( .A1(n17162), .A2(n17161), .A3(n17160), .ZN(P3_U2653) );
  AOI21_X1 U20349 ( .B1(n17353), .B2(n17163), .A(P3_REIP_REG_17__SCAN_IN), 
        .ZN(n17167) );
  OAI21_X1 U20350 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17164), .A(
        n18050), .ZN(n18081) );
  INV_X1 U20351 ( .A(n17164), .ZN(n17174) );
  OAI21_X1 U20352 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17174), .A(
        n17362), .ZN(n17165) );
  XNOR2_X1 U20353 ( .A(n18081), .B(n17165), .ZN(n17166) );
  OAI22_X1 U20354 ( .A1(n17168), .A2(n17167), .B1(n19118), .B2(n17166), .ZN(
        n17169) );
  AOI211_X1 U20355 ( .C1(n17377), .C2(P3_EBX_REG_17__SCAN_IN), .A(n9732), .B(
        n17169), .ZN(n17173) );
  OAI211_X1 U20356 ( .C1(n17178), .C2(n17171), .A(n17376), .B(n17170), .ZN(
        n17172) );
  OAI211_X1 U20357 ( .C1(n17363), .C2(n18072), .A(n17173), .B(n17172), .ZN(
        P3_U2654) );
  AOI21_X1 U20358 ( .B1(n17353), .B2(n17203), .A(n17373), .ZN(n17204) );
  INV_X1 U20359 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19165) );
  INV_X1 U20360 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18085) );
  NOR2_X1 U20361 ( .A1(n18085), .A2(n17186), .ZN(n17175) );
  OAI21_X1 U20362 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17175), .A(
        n17174), .ZN(n18086) );
  NAND2_X1 U20363 ( .A1(n17362), .A2(n17176), .ZN(n17189) );
  OAI21_X1 U20364 ( .B1(n18086), .B2(n17189), .A(n17338), .ZN(n17177) );
  AOI21_X1 U20365 ( .B1(n18086), .B2(n17189), .A(n17177), .ZN(n17182) );
  AOI211_X1 U20366 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17193), .A(n17178), .B(
        n17365), .ZN(n17181) );
  INV_X1 U20367 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18084) );
  INV_X1 U20368 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17179) );
  OAI22_X1 U20369 ( .A1(n18084), .A2(n17363), .B1(n17334), .B2(n17179), .ZN(
        n17180) );
  NOR4_X1 U20370 ( .A1(n9732), .A2(n17182), .A3(n17181), .A4(n17180), .ZN(
        n17185) );
  INV_X1 U20371 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n21405) );
  NAND3_X1 U20372 ( .A1(n17353), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n17214), 
        .ZN(n17205) );
  NOR2_X1 U20373 ( .A1(n21405), .A2(n17205), .ZN(n17191) );
  OAI211_X1 U20374 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17191), .B(n17183), .ZN(n17184) );
  OAI211_X1 U20375 ( .C1(n17204), .C2(n19165), .A(n17185), .B(n17184), .ZN(
        P3_U2655) );
  AOI22_X1 U20376 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17345), .B1(
        n17377), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n17197) );
  INV_X1 U20377 ( .A(n17204), .ZN(n17192) );
  INV_X1 U20378 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19163) );
  AOI22_X1 U20379 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17186), .B1(
        n18083), .B2(n18085), .ZN(n18096) );
  NAND2_X1 U20380 ( .A1(n17338), .A2(n17294), .ZN(n17360) );
  NOR2_X1 U20381 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17186), .ZN(
        n17187) );
  OAI21_X1 U20382 ( .B1(n17187), .B2(n18096), .A(n17338), .ZN(n17188) );
  AOI22_X1 U20383 ( .A1(n18096), .A2(n17189), .B1(n17360), .B2(n17188), .ZN(
        n17190) );
  AOI221_X1 U20384 ( .B1(n17192), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n17191), 
        .C2(n19163), .A(n17190), .ZN(n17196) );
  OAI211_X1 U20385 ( .C1(n17202), .C2(n17194), .A(n17376), .B(n17193), .ZN(
        n17195) );
  NAND4_X1 U20386 ( .A1(n17197), .A2(n17196), .A3(n18481), .A4(n17195), .ZN(
        P3_U2656) );
  INV_X1 U20387 ( .A(n17199), .ZN(n17347) );
  NOR2_X1 U20388 ( .A1(n17198), .A2(n17347), .ZN(n17286) );
  INV_X1 U20389 ( .A(n17286), .ZN(n17283) );
  NOR2_X1 U20390 ( .A1(n18123), .A2(n17283), .ZN(n17227) );
  AOI21_X1 U20391 ( .B1(n18128), .B2(n17227), .A(n17294), .ZN(n17201) );
  NAND2_X1 U20392 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17200), .ZN(
        n17226) );
  INV_X1 U20393 ( .A(n17226), .ZN(n18126) );
  NAND2_X1 U20394 ( .A1(n18128), .A2(n18126), .ZN(n17212) );
  AOI21_X1 U20395 ( .B1(n18112), .B2(n17212), .A(n18083), .ZN(n18114) );
  XNOR2_X1 U20396 ( .A(n17201), .B(n18114), .ZN(n17211) );
  AOI211_X1 U20397 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17215), .A(n17202), .B(
        n17365), .ZN(n17209) );
  INV_X1 U20398 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17546) );
  OAI22_X1 U20399 ( .A1(n18112), .A2(n17363), .B1(n17334), .B2(n17546), .ZN(
        n17208) );
  INV_X1 U20400 ( .A(n17203), .ZN(n17206) );
  OAI22_X1 U20401 ( .A1(n17206), .A2(n17205), .B1(n21405), .B2(n17204), .ZN(
        n17207) );
  NOR4_X1 U20402 ( .A1(n9732), .A2(n17209), .A3(n17208), .A4(n17207), .ZN(
        n17210) );
  OAI21_X1 U20403 ( .B1(n19118), .B2(n17211), .A(n17210), .ZN(P3_U2657) );
  INV_X1 U20404 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19160) );
  AOI21_X1 U20405 ( .B1(n17353), .B2(n17230), .A(n17373), .ZN(n17240) );
  NAND2_X1 U20406 ( .A1(n17353), .A2(n19158), .ZN(n17229) );
  AOI21_X1 U20407 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17227), .A(
        n17294), .ZN(n17213) );
  NOR2_X1 U20408 ( .A1(n18130), .A2(n17226), .ZN(n17225) );
  OAI21_X1 U20409 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17225), .A(
        n17212), .ZN(n18139) );
  XNOR2_X1 U20410 ( .A(n17213), .B(n18139), .ZN(n17221) );
  OAI22_X1 U20411 ( .A1(n18129), .A2(n17363), .B1(n17334), .B2(n17216), .ZN(
        n17220) );
  NAND2_X1 U20412 ( .A1(n17353), .A2(n17214), .ZN(n17218) );
  OAI211_X1 U20413 ( .C1(n17223), .C2(n17216), .A(n17376), .B(n17215), .ZN(
        n17217) );
  OAI211_X1 U20414 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17218), .A(n18481), 
        .B(n17217), .ZN(n17219) );
  AOI211_X1 U20415 ( .C1(n17338), .C2(n17221), .A(n17220), .B(n17219), .ZN(
        n17222) );
  OAI221_X1 U20416 ( .B1(n19160), .B2(n17240), .C1(n19160), .C2(n17229), .A(
        n17222), .ZN(P3_U2658) );
  AOI211_X1 U20417 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17242), .A(n17223), .B(
        n17365), .ZN(n17224) );
  AOI21_X1 U20418 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17377), .A(n17224), .ZN(
        n17234) );
  AOI21_X1 U20419 ( .B1(n18130), .B2(n17226), .A(n17225), .ZN(n18144) );
  NOR2_X1 U20420 ( .A1(n17227), .A2(n17294), .ZN(n17228) );
  XOR2_X1 U20421 ( .A(n18144), .B(n17228), .Z(n17232) );
  OAI22_X1 U20422 ( .A1(n18130), .A2(n17363), .B1(n17230), .B2(n17229), .ZN(
        n17231) );
  AOI211_X1 U20423 ( .C1(n17338), .C2(n17232), .A(n9732), .B(n17231), .ZN(
        n17233) );
  OAI211_X1 U20424 ( .C1(n17240), .C2(n19158), .A(n17234), .B(n17233), .ZN(
        P3_U2659) );
  INV_X1 U20425 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17246) );
  INV_X1 U20426 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19155) );
  INV_X1 U20427 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19153) );
  NOR2_X1 U20428 ( .A1(n19155), .A2(n19153), .ZN(n17236) );
  INV_X1 U20429 ( .A(n17235), .ZN(n17250) );
  NOR2_X1 U20430 ( .A1(n17366), .A2(n17250), .ZN(n17251) );
  AOI21_X1 U20431 ( .B1(n17236), .B2(n17251), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17239) );
  INV_X1 U20432 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18178) );
  NOR3_X1 U20433 ( .A1(n18285), .A2(n17198), .A3(n21384), .ZN(n17282) );
  NAND2_X1 U20434 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17282), .ZN(
        n17271) );
  NOR2_X1 U20435 ( .A1(n18178), .A2(n17271), .ZN(n17259) );
  NAND2_X1 U20436 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17259), .ZN(
        n17248) );
  AOI21_X1 U20437 ( .B1(n17246), .B2(n17248), .A(n18126), .ZN(n18159) );
  AND3_X1 U20438 ( .A1(n18192), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17286), .ZN(n17247) );
  AOI21_X1 U20439 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17247), .A(
        n17294), .ZN(n17237) );
  XNOR2_X1 U20440 ( .A(n18159), .B(n17237), .ZN(n17238) );
  OAI22_X1 U20441 ( .A1(n17240), .A2(n17239), .B1(n19118), .B2(n17238), .ZN(
        n17241) );
  AOI211_X1 U20442 ( .C1(n17377), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9732), .B(
        n17241), .ZN(n17245) );
  OAI211_X1 U20443 ( .C1(n17252), .C2(n17243), .A(n17376), .B(n17242), .ZN(
        n17244) );
  OAI211_X1 U20444 ( .C1(n17363), .C2(n17246), .A(n17245), .B(n17244), .ZN(
        P3_U2660) );
  OR2_X1 U20445 ( .A1(n17247), .A2(n17294), .ZN(n17261) );
  OAI21_X1 U20446 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17259), .A(
        n17248), .ZN(n18173) );
  XNOR2_X1 U20447 ( .A(n17261), .B(n18173), .ZN(n17257) );
  AND3_X1 U20448 ( .A1(n19155), .A2(P3_REIP_REG_9__SCAN_IN), .A3(n17251), .ZN(
        n17249) );
  AOI211_X1 U20449 ( .C1(n17377), .C2(P3_EBX_REG_10__SCAN_IN), .A(n9732), .B(
        n17249), .ZN(n17256) );
  AOI21_X1 U20450 ( .B1(n17353), .B2(n17250), .A(n17373), .ZN(n17274) );
  NAND2_X1 U20451 ( .A1(n17251), .A2(n19153), .ZN(n17258) );
  AOI21_X1 U20452 ( .B1(n17274), .B2(n17258), .A(n19155), .ZN(n17254) );
  AOI211_X1 U20453 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17267), .A(n17252), .B(
        n17365), .ZN(n17253) );
  AOI211_X1 U20454 ( .C1(n17345), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17254), .B(n17253), .ZN(n17255) );
  OAI211_X1 U20455 ( .C1(n19118), .C2(n17257), .A(n17256), .B(n17255), .ZN(
        P3_U2661) );
  INV_X1 U20456 ( .A(n17258), .ZN(n17266) );
  AOI21_X1 U20457 ( .B1(n18178), .B2(n17271), .A(n17259), .ZN(n18182) );
  NAND2_X1 U20458 ( .A1(n18192), .A2(n17286), .ZN(n17260) );
  OAI22_X1 U20459 ( .A1(n18182), .A2(n17261), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17260), .ZN(n17262) );
  AOI211_X1 U20460 ( .C1(n18182), .C2(n17294), .A(n9732), .B(n17262), .ZN(
        n17263) );
  OAI22_X1 U20461 ( .A1(n17264), .A2(n17263), .B1(n17274), .B2(n19153), .ZN(
        n17265) );
  AOI211_X1 U20462 ( .C1(n17345), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17266), .B(n17265), .ZN(n17269) );
  OAI211_X1 U20463 ( .C1(n17276), .C2(n17270), .A(n17376), .B(n17267), .ZN(
        n17268) );
  OAI211_X1 U20464 ( .C1(n17270), .C2(n17334), .A(n17269), .B(n17268), .ZN(
        P3_U2662) );
  AOI21_X1 U20465 ( .B1(n17282), .B2(n21451), .A(n17294), .ZN(n17272) );
  OAI21_X1 U20466 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17282), .A(
        n17271), .ZN(n18195) );
  XOR2_X1 U20467 ( .A(n17272), .B(n18195), .Z(n17281) );
  AOI21_X1 U20468 ( .B1(n17377), .B2(P3_EBX_REG_8__SCAN_IN), .A(n9732), .ZN(
        n17280) );
  INV_X1 U20469 ( .A(n17273), .ZN(n17305) );
  NAND2_X1 U20470 ( .A1(n17353), .A2(n17305), .ZN(n17285) );
  AOI221_X1 U20471 ( .B1(n17275), .B2(n19152), .C1(n17285), .C2(n19152), .A(
        n17274), .ZN(n17278) );
  AOI211_X1 U20472 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17287), .A(n17276), .B(
        n17365), .ZN(n17277) );
  AOI211_X1 U20473 ( .C1(n17345), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17278), .B(n17277), .ZN(n17279) );
  OAI211_X1 U20474 ( .C1(n19118), .C2(n17281), .A(n17280), .B(n17279), .ZN(
        P3_U2663) );
  AND2_X1 U20475 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18209), .ZN(
        n17304) );
  NAND2_X1 U20476 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17304), .ZN(
        n17293) );
  AOI21_X1 U20477 ( .B1(n21384), .B2(n17293), .A(n17282), .ZN(n18215) );
  NAND3_X1 U20478 ( .A1(n17338), .A2(n17362), .A3(n17283), .ZN(n17302) );
  INV_X1 U20479 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19147) );
  NOR3_X1 U20480 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n19147), .A3(n17285), .ZN(
        n17284) );
  AOI211_X1 U20481 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n17345), .A(
        n9732), .B(n17284), .ZN(n17292) );
  NOR2_X1 U20482 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17285), .ZN(n17299) );
  OAI21_X1 U20483 ( .B1(n17305), .B2(n17366), .A(n17372), .ZN(n17311) );
  OAI211_X1 U20484 ( .C1(n17286), .C2(n17294), .A(n17338), .B(n18215), .ZN(
        n17289) );
  OAI211_X1 U20485 ( .C1(n17295), .C2(n17631), .A(n17376), .B(n17287), .ZN(
        n17288) );
  OAI211_X1 U20486 ( .C1(n17631), .C2(n17334), .A(n17289), .B(n17288), .ZN(
        n17290) );
  AOI221_X1 U20487 ( .B1(n17299), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n17311), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n17290), .ZN(n17291) );
  OAI211_X1 U20488 ( .C1(n18215), .C2(n17302), .A(n17292), .B(n17291), .ZN(
        P3_U2664) );
  OAI21_X1 U20489 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17304), .A(
        n17293), .ZN(n18225) );
  INV_X1 U20490 ( .A(n18225), .ZN(n17303) );
  OAI221_X1 U20491 ( .B1(n17294), .B2(n17304), .C1(n17294), .C2(n21451), .A(
        n17338), .ZN(n17301) );
  AOI211_X1 U20492 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17312), .A(n17295), .B(
        n17365), .ZN(n17298) );
  AOI22_X1 U20493 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17345), .B1(
        P3_REIP_REG_6__SCAN_IN), .B2(n17311), .ZN(n17296) );
  OAI21_X1 U20494 ( .B1(n17334), .B2(n21399), .A(n17296), .ZN(n17297) );
  NOR4_X1 U20495 ( .A1(n9732), .A2(n17299), .A3(n17298), .A4(n17297), .ZN(
        n17300) );
  OAI221_X1 U20496 ( .B1(n17303), .B2(n17302), .C1(n18225), .C2(n17301), .A(
        n17300), .ZN(P3_U2665) );
  OR2_X1 U20497 ( .A1(n18285), .A2(n18237), .ZN(n17320) );
  AOI21_X1 U20498 ( .B1(n18238), .B2(n17320), .A(n17304), .ZN(n18240) );
  OAI21_X1 U20499 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17320), .A(
        n17362), .ZN(n17321) );
  XOR2_X1 U20500 ( .A(n18240), .B(n17321), .Z(n17309) );
  NOR2_X1 U20501 ( .A1(n17305), .A2(n17366), .ZN(n17306) );
  AOI22_X1 U20502 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17345), .B1(
        n17307), .B2(n17306), .ZN(n17308) );
  OAI211_X1 U20503 ( .C1(n19118), .C2(n17309), .A(n17308), .B(n18481), .ZN(
        n17310) );
  AOI21_X1 U20504 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n17311), .A(n17310), .ZN(
        n17314) );
  OAI211_X1 U20505 ( .C1(n17323), .C2(n17315), .A(n17376), .B(n17312), .ZN(
        n17313) );
  OAI211_X1 U20506 ( .C1(n17315), .C2(n17334), .A(n17314), .B(n17313), .ZN(
        P3_U2666) );
  AOI21_X1 U20507 ( .B1(n17353), .B2(n17316), .A(n17373), .ZN(n17331) );
  NOR3_X1 U20508 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17366), .A3(n17316), .ZN(
        n17319) );
  NAND2_X1 U20509 ( .A1(n18617), .A2(n19276), .ZN(n17380) );
  OAI221_X1 U20510 ( .B1(n17380), .B2(n17333), .C1(n17380), .C2(n17317), .A(
        n18481), .ZN(n17318) );
  AOI211_X1 U20511 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17377), .A(n17319), .B(
        n17318), .ZN(n17329) );
  AND2_X1 U20512 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18252), .ZN(
        n17330) );
  OAI21_X1 U20513 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17330), .A(
        n17320), .ZN(n18255) );
  INV_X1 U20514 ( .A(n18255), .ZN(n17322) );
  INV_X1 U20515 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17324) );
  NAND2_X1 U20516 ( .A1(n18252), .A2(n17324), .ZN(n18245) );
  OAI22_X1 U20517 ( .A1(n17322), .A2(n17321), .B1(n17347), .B2(n18245), .ZN(
        n17327) );
  AOI211_X1 U20518 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17339), .A(n17323), .B(
        n17365), .ZN(n17326) );
  OAI22_X1 U20519 ( .A1(n17324), .A2(n17363), .B1(n18255), .B2(n17360), .ZN(
        n17325) );
  AOI211_X1 U20520 ( .C1(n17338), .C2(n17327), .A(n17326), .B(n17325), .ZN(
        n17328) );
  OAI211_X1 U20521 ( .C1(n19143), .C2(n17331), .A(n17329), .B(n17328), .ZN(
        P3_U2667) );
  NAND2_X1 U20522 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17344) );
  AOI21_X1 U20523 ( .B1(n17343), .B2(n17344), .A(n17330), .ZN(n18258) );
  OAI21_X1 U20524 ( .B1(n18275), .B2(n17347), .A(n17362), .ZN(n17346) );
  XNOR2_X1 U20525 ( .A(n18258), .B(n17346), .ZN(n17337) );
  INV_X1 U20526 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19141) );
  NAND2_X1 U20527 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17352) );
  AOI221_X1 U20528 ( .B1(n17366), .B2(n19141), .C1(n17352), .C2(n19141), .A(
        n17331), .ZN(n17336) );
  NAND2_X1 U20529 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19086) );
  NOR2_X1 U20530 ( .A1(n17332), .A2(n19086), .ZN(n19083) );
  OAI21_X1 U20531 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19083), .A(
        n17333), .ZN(n19213) );
  OAI22_X1 U20532 ( .A1(n17334), .A2(n17340), .B1(n17380), .B2(n19213), .ZN(
        n17335) );
  AOI211_X1 U20533 ( .C1(n17338), .C2(n17337), .A(n17336), .B(n17335), .ZN(
        n17342) );
  OAI211_X1 U20534 ( .C1(n17349), .C2(n17340), .A(n17376), .B(n17339), .ZN(
        n17341) );
  OAI211_X1 U20535 ( .C1(n17363), .C2(n17343), .A(n17342), .B(n17341), .ZN(
        P3_U2668) );
  OAI21_X1 U20536 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17344), .ZN(n18271) );
  AOI22_X1 U20537 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17345), .B1(
        n17377), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n17359) );
  INV_X1 U20538 ( .A(n17380), .ZN(n19278) );
  AOI21_X1 U20539 ( .B1(n19226), .B2(n19081), .A(n19083), .ZN(n19223) );
  INV_X1 U20540 ( .A(n18271), .ZN(n17348) );
  AOI211_X1 U20541 ( .C1(n17348), .C2(n17347), .A(n19118), .B(n17346), .ZN(
        n17357) );
  INV_X1 U20542 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19139) );
  NOR2_X1 U20543 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17351) );
  INV_X1 U20544 ( .A(n17349), .ZN(n17350) );
  OAI211_X1 U20545 ( .C1(n17351), .C2(n9996), .A(n17376), .B(n17350), .ZN(
        n17355) );
  OAI211_X1 U20546 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17353), .B(n17352), .ZN(n17354) );
  OAI211_X1 U20547 ( .C1(n19139), .C2(n17372), .A(n17355), .B(n17354), .ZN(
        n17356) );
  AOI211_X1 U20548 ( .C1(n19278), .C2(n19223), .A(n17357), .B(n17356), .ZN(
        n17358) );
  OAI211_X1 U20549 ( .C1(n18271), .C2(n17360), .A(n17359), .B(n17358), .ZN(
        P3_U2669) );
  AND2_X1 U20550 ( .A1(n17361), .A2(n19081), .ZN(n19231) );
  AOI22_X1 U20551 ( .A1(n17377), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n19231), .B2(
        n19278), .ZN(n17371) );
  AOI21_X1 U20552 ( .B1(n17362), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n19118), .ZN(n17369) );
  NAND2_X1 U20553 ( .A1(n17362), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17364) );
  OAI21_X1 U20554 ( .B1(n19118), .B2(n17364), .A(n17363), .ZN(n17368) );
  NAND2_X1 U20555 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17649) );
  OAI21_X1 U20556 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17649), .ZN(n17656) );
  OAI22_X1 U20557 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17366), .B1(n17365), 
        .B2(n17656), .ZN(n17367) );
  AOI221_X1 U20558 ( .B1(n17369), .B2(n18285), .C1(n17368), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n17367), .ZN(n17370) );
  OAI211_X1 U20559 ( .C1(n17372), .C2(n19241), .A(n17371), .B(n17370), .ZN(
        P3_U2670) );
  NOR3_X1 U20560 ( .A1(n19274), .A2(n17373), .A3(n21451), .ZN(n17374) );
  AOI21_X1 U20561 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n17375), .A(n17374), .ZN(
        n17379) );
  OAI21_X1 U20562 ( .B1(n17377), .B2(n17376), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17378) );
  OAI211_X1 U20563 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17380), .A(
        n17379), .B(n17378), .ZN(P3_U2671) );
  NOR4_X1 U20564 ( .A1(n17384), .A2(n17383), .A3(n17382), .A4(n17381), .ZN(
        n17385) );
  NAND4_X1 U20565 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17452), .A3(n17386), 
        .A4(n17385), .ZN(n17389) );
  NAND2_X1 U20566 ( .A1(n9735), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17388) );
  NAND2_X1 U20567 ( .A1(n17408), .A2(n18645), .ZN(n17387) );
  OAI22_X1 U20568 ( .A1(n17408), .A2(n17388), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17387), .ZN(P3_U2672) );
  NAND2_X1 U20569 ( .A1(n17390), .A2(n17389), .ZN(n17391) );
  NAND2_X1 U20570 ( .A1(n17391), .A2(n9735), .ZN(n17407) );
  AOI22_X1 U20571 ( .A1(n17612), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20572 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U20573 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20574 ( .B1(n17533), .B2(n17393), .A(n17392), .ZN(n17399) );
  AOI22_X1 U20575 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20576 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20577 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20578 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17394) );
  NAND4_X1 U20579 ( .A1(n17397), .A2(n17396), .A3(n17395), .A4(n17394), .ZN(
        n17398) );
  AOI211_X1 U20580 ( .C1(n17613), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n17399), .B(n17398), .ZN(n17400) );
  NAND3_X1 U20581 ( .A1(n17402), .A2(n17401), .A3(n17400), .ZN(n17406) );
  NOR3_X1 U20582 ( .A1(n17404), .A2(n17403), .A3(n17681), .ZN(n17405) );
  XNOR2_X1 U20583 ( .A(n17406), .B(n17405), .ZN(n17671) );
  OAI22_X1 U20584 ( .A1(n17408), .A2(n17407), .B1(n17671), .B2(n9735), .ZN(
        P3_U2673) );
  OAI211_X1 U20585 ( .C1(n17683), .C2(n17682), .A(n17658), .B(n17681), .ZN(
        n17409) );
  OAI221_X1 U20586 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17412), .C1(n17411), 
        .C2(n17410), .A(n17409), .ZN(P3_U2676) );
  AOI21_X1 U20587 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n9735), .A(n17420), .ZN(
        n17414) );
  XNOR2_X1 U20588 ( .A(n17413), .B(n17416), .ZN(n17691) );
  OAI22_X1 U20589 ( .A1(n17415), .A2(n17414), .B1(n9735), .B2(n17691), .ZN(
        P3_U2677) );
  AOI21_X1 U20590 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n9735), .A(n9863), .ZN(
        n17419) );
  OAI21_X1 U20591 ( .B1(n17418), .B2(n17417), .A(n17416), .ZN(n17695) );
  OAI22_X1 U20592 ( .A1(n17420), .A2(n17419), .B1(n9735), .B2(n17695), .ZN(
        P3_U2678) );
  AOI22_X1 U20593 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n9735), .B1(
        P3_EBX_REG_23__SCAN_IN), .B2(n17423), .ZN(n17422) );
  XNOR2_X1 U20594 ( .A(n17421), .B(n17424), .ZN(n17701) );
  OAI22_X1 U20595 ( .A1(n9863), .A2(n17422), .B1(n9735), .B2(n17701), .ZN(
        P3_U2679) );
  OAI21_X1 U20596 ( .B1(n17426), .B2(n17425), .A(n17424), .ZN(n17705) );
  NAND3_X1 U20597 ( .A1(n10218), .A2(P3_EBX_REG_23__SCAN_IN), .A3(n9735), .ZN(
        n17427) );
  OAI221_X1 U20598 ( .B1(n10218), .B2(P3_EBX_REG_23__SCAN_IN), .C1(n9735), 
        .C2(n17705), .A(n17427), .ZN(P3_U2680) );
  AOI22_X1 U20599 ( .A1(n9724), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20600 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20601 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17429) );
  AOI22_X1 U20602 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17428) );
  NAND4_X1 U20603 ( .A1(n17431), .A2(n17430), .A3(n17429), .A4(n17428), .ZN(
        n17437) );
  AOI22_X1 U20604 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U20605 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17434) );
  AOI22_X1 U20606 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U20607 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17432) );
  NAND4_X1 U20608 ( .A1(n17435), .A2(n17434), .A3(n17433), .A4(n17432), .ZN(
        n17436) );
  NOR2_X1 U20609 ( .A1(n17437), .A2(n17436), .ZN(n17708) );
  NAND3_X1 U20610 ( .A1(n17439), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n9735), .ZN(
        n17438) );
  OAI221_X1 U20611 ( .B1(n17439), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n9735), 
        .C2(n17708), .A(n17438), .ZN(P3_U2681) );
  OAI21_X1 U20612 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n10205), .A(n9735), .ZN(
        n17451) );
  AOI22_X1 U20613 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20614 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20615 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20616 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17441) );
  NAND4_X1 U20617 ( .A1(n17444), .A2(n17443), .A3(n17442), .A4(n17441), .ZN(
        n17450) );
  AOI22_X1 U20618 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20619 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U20620 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U20621 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17445) );
  NAND4_X1 U20622 ( .A1(n17448), .A2(n17447), .A3(n17446), .A4(n17445), .ZN(
        n17449) );
  NOR2_X1 U20623 ( .A1(n17450), .A2(n17449), .ZN(n17714) );
  OAI22_X1 U20624 ( .A1(n17452), .A2(n17451), .B1(n17714), .B2(n9735), .ZN(
        P3_U2682) );
  AOI22_X1 U20625 ( .A1(n18645), .A2(n17476), .B1(P3_EBX_REG_20__SCAN_IN), 
        .B2(n9735), .ZN(n17464) );
  AOI22_X1 U20626 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20627 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U20628 ( .A1(n17596), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20629 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17453) );
  NAND4_X1 U20630 ( .A1(n17456), .A2(n17455), .A3(n17454), .A4(n17453), .ZN(
        n17463) );
  AOI22_X1 U20631 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17461) );
  AOI22_X1 U20632 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20633 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9723), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U20634 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17458) );
  NAND4_X1 U20635 ( .A1(n17461), .A2(n17460), .A3(n17459), .A4(n17458), .ZN(
        n17462) );
  NOR2_X1 U20636 ( .A1(n17463), .A2(n17462), .ZN(n17718) );
  OAI22_X1 U20637 ( .A1(n10205), .A2(n17464), .B1(n17718), .B2(n9735), .ZN(
        P3_U2683) );
  OAI21_X1 U20638 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n10207), .A(n9735), .ZN(
        n17475) );
  AOI22_X1 U20639 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20640 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U20641 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U20642 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9724), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17465) );
  NAND4_X1 U20643 ( .A1(n17468), .A2(n17467), .A3(n17466), .A4(n17465), .ZN(
        n17474) );
  AOI22_X1 U20644 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U20645 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U20646 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U20647 ( .A1(n17594), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17469) );
  NAND4_X1 U20648 ( .A1(n17472), .A2(n17471), .A3(n17470), .A4(n17469), .ZN(
        n17473) );
  NOR2_X1 U20649 ( .A1(n17474), .A2(n17473), .ZN(n17726) );
  OAI22_X1 U20650 ( .A1(n17476), .A2(n17475), .B1(n17726), .B2(n9735), .ZN(
        P3_U2684) );
  AOI22_X1 U20651 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17480) );
  AOI22_X1 U20652 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U20653 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U20654 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17477) );
  NAND4_X1 U20655 ( .A1(n17480), .A2(n17479), .A3(n17478), .A4(n17477), .ZN(
        n17486) );
  AOI22_X1 U20656 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U20657 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U20658 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U20659 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17481) );
  NAND4_X1 U20660 ( .A1(n17484), .A2(n17483), .A3(n17482), .A4(n17481), .ZN(
        n17485) );
  NOR2_X1 U20661 ( .A1(n17486), .A2(n17485), .ZN(n17731) );
  OAI21_X1 U20662 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17502), .A(n17487), .ZN(
        n17488) );
  AOI22_X1 U20663 ( .A1(n17658), .A2(n17731), .B1(n17488), .B2(n9735), .ZN(
        P3_U2685) );
  INV_X1 U20664 ( .A(n17489), .ZN(n17490) );
  OAI21_X1 U20665 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17490), .A(n9735), .ZN(
        n17501) );
  AOI22_X1 U20666 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17553), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17494) );
  AOI22_X1 U20667 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U20668 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17597), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9728), .ZN(n17492) );
  AOI22_X1 U20669 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17596), .ZN(n17491) );
  NAND4_X1 U20670 ( .A1(n17494), .A2(n17493), .A3(n17492), .A4(n17491), .ZN(
        n17500) );
  AOI22_X1 U20671 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U20672 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n16674), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9737), .ZN(n17497) );
  AOI22_X1 U20673 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U20674 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17594), .ZN(n17495) );
  NAND4_X1 U20675 ( .A1(n17498), .A2(n17497), .A3(n17496), .A4(n17495), .ZN(
        n17499) );
  NOR2_X1 U20676 ( .A1(n17500), .A2(n17499), .ZN(n17737) );
  OAI22_X1 U20677 ( .A1(n17502), .A2(n17501), .B1(n17737), .B2(n9735), .ZN(
        P3_U2686) );
  NAND2_X1 U20678 ( .A1(n18645), .A2(n17503), .ZN(n17516) );
  NOR2_X1 U20679 ( .A1(n17658), .A2(n17503), .ZN(n17529) );
  AOI22_X1 U20680 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U20681 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U20682 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12500), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17504) );
  OAI21_X1 U20683 ( .B1(n17505), .B2(n21458), .A(n17504), .ZN(n17511) );
  AOI22_X1 U20684 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U20685 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17508) );
  AOI22_X1 U20686 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U20687 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17506) );
  NAND4_X1 U20688 ( .A1(n17509), .A2(n17508), .A3(n17507), .A4(n17506), .ZN(
        n17510) );
  AOI211_X1 U20689 ( .C1(n17613), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17511), .B(n17510), .ZN(n17512) );
  NAND3_X1 U20690 ( .A1(n17514), .A2(n17513), .A3(n17512), .ZN(n17738) );
  AOI22_X1 U20691 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17529), .B1(n17658), 
        .B2(n17738), .ZN(n17515) );
  OAI21_X1 U20692 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17516), .A(n17515), .ZN(
        P3_U2687) );
  AOI22_X1 U20693 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17520) );
  AOI22_X1 U20694 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U20695 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9723), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17518) );
  AOI22_X1 U20696 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17517) );
  NAND4_X1 U20697 ( .A1(n17520), .A2(n17519), .A3(n17518), .A4(n17517), .ZN(
        n17527) );
  AOI22_X1 U20698 ( .A1(n9728), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U20699 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U20700 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17523) );
  AOI22_X1 U20701 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17522) );
  NAND4_X1 U20702 ( .A1(n17525), .A2(n17524), .A3(n17523), .A4(n17522), .ZN(
        n17526) );
  NOR2_X1 U20703 ( .A1(n17527), .A2(n17526), .ZN(n17747) );
  INV_X1 U20704 ( .A(n17528), .ZN(n17530) );
  OAI21_X1 U20705 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17530), .A(n17529), .ZN(
        n17531) );
  OAI21_X1 U20706 ( .B1(n17747), .B2(n9735), .A(n17531), .ZN(P3_U2688) );
  AOI22_X1 U20707 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17542) );
  AOI22_X1 U20708 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U20709 ( .A1(n17596), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17532) );
  OAI21_X1 U20710 ( .B1(n17533), .B2(n21397), .A(n17532), .ZN(n17539) );
  AOI22_X1 U20711 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U20712 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17536) );
  AOI22_X1 U20713 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17535) );
  AOI22_X1 U20714 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17534) );
  NAND4_X1 U20715 ( .A1(n17537), .A2(n17536), .A3(n17535), .A4(n17534), .ZN(
        n17538) );
  AOI211_X1 U20716 ( .C1(n17580), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17539), .B(n17538), .ZN(n17540) );
  NAND3_X1 U20717 ( .A1(n17542), .A2(n17541), .A3(n17540), .ZN(n17748) );
  NOR2_X1 U20718 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17749), .ZN(n17543) );
  AOI22_X1 U20719 ( .A1(n17658), .A2(n17748), .B1(n17544), .B2(n17543), .ZN(
        n17545) );
  OAI21_X1 U20720 ( .B1(n17547), .B2(n17546), .A(n17545), .ZN(P3_U2689) );
  AOI22_X1 U20721 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17552) );
  AOI22_X1 U20722 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17551) );
  AOI22_X1 U20723 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U20724 ( .A1(n17548), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17549) );
  NAND4_X1 U20725 ( .A1(n17552), .A2(n17551), .A3(n17550), .A4(n17549), .ZN(
        n17559) );
  AOI22_X1 U20726 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17557) );
  AOI22_X1 U20727 ( .A1(n17553), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U20728 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17555) );
  AOI22_X1 U20729 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17554) );
  NAND4_X1 U20730 ( .A1(n17557), .A2(n17556), .A3(n17555), .A4(n17554), .ZN(
        n17558) );
  NOR2_X1 U20731 ( .A1(n17559), .A2(n17558), .ZN(n17759) );
  OAI211_X1 U20732 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17579), .A(n17560), .B(
        n9735), .ZN(n17561) );
  OAI21_X1 U20733 ( .B1(n17759), .B2(n9735), .A(n17561), .ZN(P3_U2691) );
  INV_X1 U20734 ( .A(n17591), .ZN(n17562) );
  OAI21_X1 U20735 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17562), .A(n9735), .ZN(
        n17578) );
  AOI22_X1 U20736 ( .A1(n17563), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17613), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17576) );
  AOI22_X1 U20737 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9728), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17575) );
  INV_X1 U20738 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n21437) );
  AOI22_X1 U20739 ( .A1(n17564), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17565) );
  OAI21_X1 U20740 ( .B1(n17566), .B2(n21437), .A(n17565), .ZN(n17573) );
  AOI22_X1 U20741 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17571) );
  AOI22_X1 U20742 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9725), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17570) );
  AOI22_X1 U20743 ( .A1(n17567), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17569) );
  AOI22_X1 U20744 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17596), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17568) );
  NAND4_X1 U20745 ( .A1(n17571), .A2(n17570), .A3(n17569), .A4(n17568), .ZN(
        n17572) );
  AOI211_X1 U20746 ( .C1(n17615), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17573), .B(n17572), .ZN(n17574) );
  NAND3_X1 U20747 ( .A1(n17576), .A2(n17575), .A3(n17574), .ZN(n17762) );
  INV_X1 U20748 ( .A(n17762), .ZN(n17577) );
  OAI22_X1 U20749 ( .A1(n17579), .A2(n17578), .B1(n17577), .B2(n9735), .ZN(
        P3_U2692) );
  AOI22_X1 U20750 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17584) );
  AOI22_X1 U20751 ( .A1(n17616), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16674), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17583) );
  AOI22_X1 U20752 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17582) );
  AOI22_X1 U20753 ( .A1(n17596), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17581) );
  NAND4_X1 U20754 ( .A1(n17584), .A2(n17583), .A3(n17582), .A4(n17581), .ZN(
        n17590) );
  AOI22_X1 U20755 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U20756 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9741), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17587) );
  AOI22_X1 U20757 ( .A1(n9725), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17521), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17586) );
  AOI22_X1 U20758 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9737), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17585) );
  NAND4_X1 U20759 ( .A1(n17588), .A2(n17587), .A3(n17586), .A4(n17585), .ZN(
        n17589) );
  NOR2_X1 U20760 ( .A1(n17590), .A2(n17589), .ZN(n17765) );
  OAI21_X1 U20761 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17610), .A(n17591), .ZN(
        n17592) );
  AOI22_X1 U20762 ( .A1(n17658), .A2(n17765), .B1(n17592), .B2(n9735), .ZN(
        P3_U2693) );
  INV_X1 U20763 ( .A(n17593), .ZN(n17630) );
  OAI21_X1 U20764 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17630), .A(n9735), .ZN(
        n17609) );
  AOI22_X1 U20765 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17616), .B1(
        n17580), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17601) );
  AOI22_X1 U20766 ( .A1(n17595), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17594), .ZN(n17600) );
  AOI22_X1 U20767 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17596), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9737), .ZN(n17599) );
  AOI22_X1 U20768 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17597), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n16674), .ZN(n17598) );
  NAND4_X1 U20769 ( .A1(n17601), .A2(n17600), .A3(n17599), .A4(n17598), .ZN(
        n17608) );
  AOI22_X1 U20770 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9724), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17606) );
  AOI22_X1 U20771 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9729), .B1(
        n17602), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17605) );
  AOI22_X1 U20772 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17613), .ZN(n17604) );
  AOI22_X1 U20773 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17603) );
  NAND4_X1 U20774 ( .A1(n17606), .A2(n17605), .A3(n17604), .A4(n17603), .ZN(
        n17607) );
  NOR2_X1 U20775 ( .A1(n17608), .A2(n17607), .ZN(n17770) );
  OAI22_X1 U20776 ( .A1(n17610), .A2(n17609), .B1(n17770), .B2(n9735), .ZN(
        P3_U2694) );
  NOR2_X1 U20777 ( .A1(n17611), .A2(n17660), .ZN(n17648) );
  NAND3_X1 U20778 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .A3(n17648), .ZN(n17638) );
  NOR2_X1 U20779 ( .A1(n21399), .A2(n17638), .ZN(n17632) );
  AOI22_X1 U20780 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n9735), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17632), .ZN(n17629) );
  AOI22_X1 U20781 ( .A1(n9721), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17564), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17627) );
  AOI22_X1 U20782 ( .A1(n17602), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17626) );
  AOI22_X1 U20783 ( .A1(n17613), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17594), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17614) );
  OAI21_X1 U20784 ( .B1(n9720), .B2(n21458), .A(n17614), .ZN(n17624) );
  AOI22_X1 U20785 ( .A1(n17615), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17548), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17622) );
  AOI22_X1 U20786 ( .A1(n17617), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17616), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17621) );
  AOI22_X1 U20787 ( .A1(n9741), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17618), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U20788 ( .A1(n17596), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9728), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17619) );
  NAND4_X1 U20789 ( .A1(n17622), .A2(n17621), .A3(n17620), .A4(n17619), .ZN(
        n17623) );
  AOI211_X1 U20790 ( .C1(n9725), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17624), .B(n17623), .ZN(n17625) );
  NAND3_X1 U20791 ( .A1(n17627), .A2(n17626), .A3(n17625), .ZN(n17776) );
  INV_X1 U20792 ( .A(n17776), .ZN(n17628) );
  OAI22_X1 U20793 ( .A1(n17630), .A2(n17629), .B1(n17628), .B2(n9735), .ZN(
        P3_U2695) );
  NAND2_X1 U20794 ( .A1(n9735), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U20795 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17658), .B1(
        n17632), .B2(n17631), .ZN(n17633) );
  OAI21_X1 U20796 ( .B1(n17635), .B2(n17634), .A(n17633), .ZN(P3_U2696) );
  INV_X1 U20797 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17637) );
  NAND3_X1 U20798 ( .A1(n17638), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n9735), .ZN(
        n17636) );
  OAI221_X1 U20799 ( .B1(n17638), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n9735), .C2(
        n17637), .A(n17636), .ZN(P3_U2697) );
  INV_X1 U20800 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17641) );
  INV_X1 U20801 ( .A(n17642), .ZN(n17639) );
  OAI211_X1 U20802 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17639), .A(n17638), .B(
        n9735), .ZN(n17640) );
  OAI21_X1 U20803 ( .B1(n9735), .B2(n17641), .A(n17640), .ZN(P3_U2698) );
  OAI21_X1 U20804 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17643), .A(n17642), .ZN(
        n17644) );
  AOI22_X1 U20805 ( .A1(n17658), .A2(n17645), .B1(n17644), .B2(n9735), .ZN(
        P3_U2699) );
  NOR3_X1 U20806 ( .A1(n9996), .A2(n17649), .A3(n17660), .ZN(n17653) );
  AOI21_X1 U20807 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n9735), .A(n17653), .ZN(
        n17647) );
  INV_X1 U20808 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17646) );
  OAI22_X1 U20809 ( .A1(n17648), .A2(n17647), .B1(n17646), .B2(n9735), .ZN(
        P3_U2700) );
  NOR2_X1 U20810 ( .A1(n17649), .A2(n17660), .ZN(n17650) );
  AOI21_X1 U20811 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n9735), .A(n17650), .ZN(
        n17652) );
  INV_X1 U20812 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17651) );
  OAI22_X1 U20813 ( .A1(n17653), .A2(n17652), .B1(n17651), .B2(n9735), .ZN(
        P3_U2701) );
  OAI222_X1 U20814 ( .A1(n17656), .A2(n17660), .B1(n9997), .B2(n17655), .C1(
        n17654), .C2(n9735), .ZN(P3_U2702) );
  AOI22_X1 U20815 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17658), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17657), .ZN(n17659) );
  OAI21_X1 U20816 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17660), .A(n17659), .ZN(
        P3_U2703) );
  INV_X1 U20817 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n21310) );
  INV_X1 U20818 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17876) );
  INV_X1 U20819 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17920) );
  NAND3_X1 U20820 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .ZN(n17782) );
  INV_X1 U20821 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17889) );
  NAND2_X1 U20822 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17781) );
  INV_X1 U20823 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17901) );
  INV_X1 U20824 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17911) );
  INV_X1 U20825 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17907) );
  INV_X1 U20826 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17905) );
  INV_X1 U20827 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17903) );
  NOR4_X1 U20828 ( .A1(n17911), .A2(n17907), .A3(n17905), .A4(n17903), .ZN(
        n17750) );
  NOR2_X4 U20829 ( .A1(n17920), .A2(n17751), .ZN(n17744) );
  INV_X1 U20830 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17867) );
  INV_X1 U20831 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17865) );
  NOR2_X1 U20832 ( .A1(n17867), .A2(n17865), .ZN(n17662) );
  NAND4_X1 U20833 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17662), .ZN(n17707) );
  INV_X1 U20834 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17869) );
  NAND2_X1 U20835 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17677), .ZN(n17673) );
  NAND2_X1 U20836 ( .A1(n17668), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17664) );
  NOR2_X2 U20837 ( .A1(n18640), .A2(n17806), .ZN(n17739) );
  NAND2_X1 U20838 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17739), .ZN(n17663) );
  OAI221_X1 U20839 ( .B1(n17668), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17664), 
        .C2(n17774), .A(n17663), .ZN(P3_U2704) );
  NAND2_X1 U20840 ( .A1(n18636), .A2(n17774), .ZN(n17743) );
  AOI22_X1 U20841 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17739), .ZN(n17670) );
  NAND2_X1 U20842 ( .A1(n17668), .A2(n17667), .ZN(n17669) );
  OAI211_X1 U20843 ( .C1(n17671), .C2(n17801), .A(n17670), .B(n17669), .ZN(
        P3_U2705) );
  INV_X1 U20844 ( .A(n17739), .ZN(n17713) );
  AOI22_X1 U20845 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17732), .B1(n17672), .B2(
        n17809), .ZN(n17675) );
  OAI211_X1 U20846 ( .C1(n17677), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17806), .B(
        n17673), .ZN(n17674) );
  OAI211_X1 U20847 ( .C1(n17713), .C2(n15917), .A(n17675), .B(n17674), .ZN(
        P3_U2706) );
  AOI22_X1 U20848 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17732), .B1(n17676), .B2(
        n17809), .ZN(n17680) );
  AOI211_X1 U20849 ( .C1(n21310), .C2(n17684), .A(n17677), .B(n17774), .ZN(
        n17678) );
  INV_X1 U20850 ( .A(n17678), .ZN(n17679) );
  OAI211_X1 U20851 ( .C1(n17713), .C2(n15926), .A(n17680), .B(n17679), .ZN(
        P3_U2707) );
  OAI21_X1 U20852 ( .B1(n17683), .B2(n17682), .A(n17681), .ZN(n17687) );
  AOI22_X1 U20853 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17739), .ZN(n17686) );
  OAI211_X1 U20854 ( .C1(n9788), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17806), .B(
        n17684), .ZN(n17685) );
  OAI211_X1 U20855 ( .C1(n17801), .C2(n17687), .A(n17686), .B(n17685), .ZN(
        P3_U2708) );
  AOI22_X1 U20856 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17739), .ZN(n17690) );
  AOI211_X1 U20857 ( .C1(n17876), .C2(n17692), .A(n9788), .B(n17774), .ZN(
        n17688) );
  INV_X1 U20858 ( .A(n17688), .ZN(n17689) );
  OAI211_X1 U20859 ( .C1(n17801), .C2(n17691), .A(n17690), .B(n17689), .ZN(
        P3_U2709) );
  AOI22_X1 U20860 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17739), .ZN(n17694) );
  OAI211_X1 U20861 ( .C1(n17696), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17806), .B(
        n17692), .ZN(n17693) );
  OAI211_X1 U20862 ( .C1(n17801), .C2(n17695), .A(n17694), .B(n17693), .ZN(
        P3_U2710) );
  AOI22_X1 U20863 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17739), .ZN(n17700) );
  OAI211_X1 U20864 ( .C1(n17698), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17806), .B(
        n17697), .ZN(n17699) );
  OAI211_X1 U20865 ( .C1(n17801), .C2(n17701), .A(n17700), .B(n17699), .ZN(
        P3_U2711) );
  AOI22_X1 U20866 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17739), .ZN(n17704) );
  OAI211_X1 U20867 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n9884), .A(n17806), .B(
        n17702), .ZN(n17703) );
  OAI211_X1 U20868 ( .C1(n17801), .C2(n17705), .A(n17704), .B(n17703), .ZN(
        P3_U2712) );
  INV_X1 U20869 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17861) );
  NAND2_X1 U20870 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17727), .ZN(n17723) );
  NOR2_X1 U20871 ( .A1(n17865), .A2(n17723), .ZN(n17716) );
  NOR2_X1 U20872 ( .A1(n17774), .A2(n17716), .ZN(n17720) );
  AOI21_X1 U20873 ( .B1(n17706), .B2(n17867), .A(n17720), .ZN(n17712) );
  NOR4_X1 U20874 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17749), .A3(n17740), .A4(
        n17707), .ZN(n17710) );
  OAI22_X1 U20875 ( .A1(n17708), .A2(n17801), .B1(n15963), .B2(n17713), .ZN(
        n17709) );
  AOI211_X1 U20876 ( .C1(n17732), .C2(BUF2_REG_6__SCAN_IN), .A(n17710), .B(
        n17709), .ZN(n17711) );
  OAI21_X1 U20877 ( .B1(n17712), .B2(n17869), .A(n17711), .ZN(P3_U2713) );
  OAI22_X1 U20878 ( .A1(n17714), .A2(n17801), .B1(n18635), .B2(n17713), .ZN(
        n17715) );
  AOI221_X1 U20879 ( .B1(n17720), .B2(P3_EAX_REG_21__SCAN_IN), .C1(n17716), 
        .C2(n17867), .A(n17715), .ZN(n17717) );
  OAI21_X1 U20880 ( .B1(n13138), .B2(n17743), .A(n17717), .ZN(P3_U2714) );
  INV_X1 U20881 ( .A(n17718), .ZN(n17719) );
  AOI22_X1 U20882 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17739), .B1(n17809), .B2(
        n17719), .ZN(n17722) );
  AOI22_X1 U20883 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17732), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n17720), .ZN(n17721) );
  OAI211_X1 U20884 ( .C1(P3_EAX_REG_20__SCAN_IN), .C2(n17723), .A(n17722), .B(
        n17721), .ZN(P3_U2715) );
  AOI22_X1 U20885 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17739), .ZN(n17725) );
  OAI211_X1 U20886 ( .C1(n17727), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17806), .B(
        n17723), .ZN(n17724) );
  OAI211_X1 U20887 ( .C1(n17726), .C2(n17801), .A(n17725), .B(n17724), .ZN(
        P3_U2716) );
  AOI22_X1 U20888 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17739), .ZN(n17730) );
  AOI211_X1 U20889 ( .C1(n17861), .C2(n17733), .A(n17727), .B(n17774), .ZN(
        n17728) );
  INV_X1 U20890 ( .A(n17728), .ZN(n17729) );
  OAI211_X1 U20891 ( .C1(n17731), .C2(n17801), .A(n17730), .B(n17729), .ZN(
        P3_U2717) );
  AOI22_X1 U20892 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17732), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17739), .ZN(n17736) );
  OAI211_X1 U20893 ( .C1(n17734), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17806), .B(
        n17733), .ZN(n17735) );
  OAI211_X1 U20894 ( .C1(n17737), .C2(n17801), .A(n17736), .B(n17735), .ZN(
        P3_U2718) );
  AOI22_X1 U20895 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17739), .B1(n17809), .B2(
        n17738), .ZN(n17742) );
  OAI211_X1 U20896 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17744), .A(n17806), .B(
        n17740), .ZN(n17741) );
  OAI211_X1 U20897 ( .C1(n17743), .C2(n18612), .A(n17742), .B(n17741), .ZN(
        P3_U2719) );
  AOI211_X1 U20898 ( .C1(n17920), .C2(n17751), .A(n17774), .B(n17744), .ZN(
        n17745) );
  AOI21_X1 U20899 ( .B1(n17810), .B2(BUF2_REG_15__SCAN_IN), .A(n17745), .ZN(
        n17746) );
  OAI21_X1 U20900 ( .B1(n17747), .B2(n17801), .A(n17746), .ZN(P3_U2720) );
  AOI22_X1 U20901 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17810), .B1(n17809), .B2(
        n17748), .ZN(n17753) );
  INV_X1 U20902 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17913) );
  NOR3_X1 U20903 ( .A1(n17749), .A2(n17901), .A3(n17779), .ZN(n17769) );
  NAND2_X1 U20904 ( .A1(n17750), .A2(n17769), .ZN(n17754) );
  NOR2_X1 U20905 ( .A1(n17913), .A2(n17754), .ZN(n17757) );
  OAI211_X1 U20906 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17757), .A(n17806), .B(
        n17751), .ZN(n17752) );
  NAND2_X1 U20907 ( .A1(n17753), .A2(n17752), .ZN(P3_U2721) );
  INV_X1 U20908 ( .A(n17754), .ZN(n17761) );
  AOI21_X1 U20909 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17806), .A(n17761), .ZN(
        n17756) );
  OAI222_X1 U20910 ( .A1(n17804), .A2(n13123), .B1(n17757), .B2(n17756), .C1(
        n17801), .C2(n17755), .ZN(P3_U2722) );
  NAND3_X1 U20911 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n17769), .ZN(n17764) );
  INV_X1 U20912 ( .A(n17764), .ZN(n17758) );
  AOI22_X1 U20913 ( .A1(n17758), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17806), .ZN(n17760) );
  OAI222_X1 U20914 ( .A1(n17804), .A2(n13126), .B1(n17761), .B2(n17760), .C1(
        n17801), .C2(n17759), .ZN(P3_U2723) );
  NAND2_X1 U20915 ( .A1(n17806), .A2(n17764), .ZN(n17767) );
  AOI22_X1 U20916 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17810), .B1(n17809), .B2(
        n17762), .ZN(n17763) );
  OAI221_X1 U20917 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17764), .C1(n17907), 
        .C2(n17767), .A(n17763), .ZN(P3_U2724) );
  AOI21_X1 U20918 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17769), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n17766) );
  OAI222_X1 U20919 ( .A1(n17804), .A2(n17768), .B1(n17767), .B2(n17766), .C1(
        n17801), .C2(n17765), .ZN(P3_U2725) );
  AND2_X1 U20920 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17769), .ZN(n17772) );
  AOI21_X1 U20921 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17806), .A(n17769), .ZN(
        n17771) );
  OAI222_X1 U20922 ( .A1(n17804), .A2(n13132), .B1(n17772), .B2(n17771), .C1(
        n17801), .C2(n17770), .ZN(P3_U2726) );
  AOI211_X1 U20923 ( .C1(n17901), .C2(n17779), .A(n17774), .B(n17773), .ZN(
        n17775) );
  AOI21_X1 U20924 ( .B1(n17809), .B2(n17776), .A(n17775), .ZN(n17777) );
  OAI21_X1 U20925 ( .B1(n17778), .B2(n17804), .A(n17777), .ZN(P3_U2727) );
  INV_X1 U20926 ( .A(n17779), .ZN(n17785) );
  NAND2_X1 U20927 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17813), .ZN(n17796) );
  NOR2_X1 U20928 ( .A1(n17782), .A2(n17796), .ZN(n17792) );
  AOI22_X1 U20929 ( .A1(n17792), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17806), .ZN(n17784) );
  OAI222_X1 U20930 ( .A1(n17804), .A2(n13056), .B1(n17785), .B2(n17784), .C1(
        n17801), .C2(n17783), .ZN(P3_U2728) );
  AOI21_X1 U20931 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17806), .A(n17792), .ZN(
        n17788) );
  AND2_X1 U20932 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17792), .ZN(n17787) );
  OAI222_X1 U20933 ( .A1(n17804), .A2(n12944), .B1(n17788), .B2(n17787), .C1(
        n17801), .C2(n17786), .ZN(P3_U2729) );
  NAND2_X1 U20934 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n17789) );
  NOR2_X1 U20935 ( .A1(n17789), .A2(n17796), .ZN(n17795) );
  AOI21_X1 U20936 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17806), .A(n17795), .ZN(
        n17791) );
  OAI222_X1 U20937 ( .A1(n13138), .A2(n17804), .B1(n17792), .B2(n17791), .C1(
        n17801), .C2(n17790), .ZN(P3_U2730) );
  INV_X1 U20938 ( .A(n17796), .ZN(n17803) );
  AOI22_X1 U20939 ( .A1(n17803), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17806), .ZN(n17794) );
  OAI222_X1 U20940 ( .A1(n21290), .A2(n17804), .B1(n17795), .B2(n17794), .C1(
        n17801), .C2(n17793), .ZN(P3_U2731) );
  INV_X1 U20941 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17891) );
  NOR2_X1 U20942 ( .A1(n17891), .A2(n17796), .ZN(n17799) );
  AOI21_X1 U20943 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17806), .A(n17803), .ZN(
        n17798) );
  OAI222_X1 U20944 ( .A1(n18628), .A2(n17804), .B1(n17799), .B2(n17798), .C1(
        n17801), .C2(n17797), .ZN(P3_U2732) );
  AOI21_X1 U20945 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17806), .A(n17813), .ZN(
        n17802) );
  OAI222_X1 U20946 ( .A1(n18624), .A2(n17804), .B1(n17803), .B2(n17802), .C1(
        n17801), .C2(n17800), .ZN(P3_U2733) );
  NOR2_X1 U20947 ( .A1(n17805), .A2(n17885), .ZN(n17807) );
  OAI21_X1 U20948 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17807), .A(n17806), .ZN(
        n17812) );
  AOI22_X1 U20949 ( .A1(n17810), .A2(BUF2_REG_1__SCAN_IN), .B1(n17809), .B2(
        n17808), .ZN(n17811) );
  OAI21_X1 U20950 ( .B1(n17813), .B2(n17812), .A(n17811), .ZN(P3_U2734) );
  NOR2_X1 U20951 ( .A1(n19221), .A2(n19123), .ZN(n17842) );
  AND2_X1 U20952 ( .A1(n17850), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20953 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17883) );
  NAND2_X1 U20954 ( .A1(n17832), .A2(n17815), .ZN(n17831) );
  AOI22_X1 U20955 ( .A1(n19255), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17848), .ZN(n17816) );
  OAI21_X1 U20956 ( .B1(n17883), .B2(n17831), .A(n17816), .ZN(P3_U2737) );
  INV_X1 U20957 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17881) );
  AOI22_X1 U20958 ( .A1(n19255), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17817) );
  OAI21_X1 U20959 ( .B1(n17881), .B2(n17831), .A(n17817), .ZN(P3_U2738) );
  AOI22_X1 U20960 ( .A1(n19255), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17818) );
  OAI21_X1 U20961 ( .B1(n21310), .B2(n17831), .A(n17818), .ZN(P3_U2739) );
  INV_X1 U20962 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17878) );
  AOI22_X1 U20963 ( .A1(n19255), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17819) );
  OAI21_X1 U20964 ( .B1(n17878), .B2(n17831), .A(n17819), .ZN(P3_U2740) );
  AOI22_X1 U20965 ( .A1(n19255), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17820) );
  OAI21_X1 U20966 ( .B1(n17876), .B2(n17831), .A(n17820), .ZN(P3_U2741) );
  INV_X1 U20967 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17874) );
  AOI22_X1 U20968 ( .A1(n19255), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17821) );
  OAI21_X1 U20969 ( .B1(n17874), .B2(n17831), .A(n17821), .ZN(P3_U2742) );
  INV_X1 U20970 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17872) );
  AOI22_X1 U20971 ( .A1(n19255), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17822) );
  OAI21_X1 U20972 ( .B1(n17872), .B2(n17831), .A(n17822), .ZN(P3_U2743) );
  AOI22_X1 U20973 ( .A1(n19255), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17823) );
  OAI21_X1 U20974 ( .B1(n10263), .B2(n17831), .A(n17823), .ZN(P3_U2744) );
  AOI22_X1 U20975 ( .A1(n19255), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17824) );
  OAI21_X1 U20976 ( .B1(n17869), .B2(n17831), .A(n17824), .ZN(P3_U2745) );
  AOI22_X1 U20977 ( .A1(n17842), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17825) );
  OAI21_X1 U20978 ( .B1(n17867), .B2(n17831), .A(n17825), .ZN(P3_U2746) );
  AOI22_X1 U20979 ( .A1(n17842), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17826) );
  OAI21_X1 U20980 ( .B1(n17865), .B2(n17831), .A(n17826), .ZN(P3_U2747) );
  INV_X1 U20981 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17863) );
  AOI22_X1 U20982 ( .A1(n17842), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17827) );
  OAI21_X1 U20983 ( .B1(n17863), .B2(n17831), .A(n17827), .ZN(P3_U2748) );
  AOI22_X1 U20984 ( .A1(n17842), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17828) );
  OAI21_X1 U20985 ( .B1(n17861), .B2(n17831), .A(n17828), .ZN(P3_U2749) );
  INV_X1 U20986 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17859) );
  AOI22_X1 U20987 ( .A1(n17842), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17829) );
  OAI21_X1 U20988 ( .B1(n17859), .B2(n17831), .A(n17829), .ZN(P3_U2750) );
  INV_X1 U20989 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17857) );
  AOI22_X1 U20990 ( .A1(n17842), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17830) );
  OAI21_X1 U20991 ( .B1(n17857), .B2(n17831), .A(n17830), .ZN(P3_U2751) );
  AOI22_X1 U20992 ( .A1(n17842), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17833) );
  OAI21_X1 U20993 ( .B1(n17920), .B2(n17852), .A(n17833), .ZN(P3_U2752) );
  INV_X1 U20994 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17915) );
  AOI22_X1 U20995 ( .A1(n17842), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17834) );
  OAI21_X1 U20996 ( .B1(n17915), .B2(n17852), .A(n17834), .ZN(P3_U2753) );
  AOI22_X1 U20997 ( .A1(n17842), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17835) );
  OAI21_X1 U20998 ( .B1(n17913), .B2(n17852), .A(n17835), .ZN(P3_U2754) );
  AOI22_X1 U20999 ( .A1(n17842), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17836) );
  OAI21_X1 U21000 ( .B1(n17911), .B2(n17852), .A(n17836), .ZN(P3_U2755) );
  AOI22_X1 U21001 ( .A1(n19255), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17837) );
  OAI21_X1 U21002 ( .B1(n17907), .B2(n17852), .A(n17837), .ZN(P3_U2756) );
  AOI22_X1 U21003 ( .A1(n19255), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17838) );
  OAI21_X1 U21004 ( .B1(n17905), .B2(n17852), .A(n17838), .ZN(P3_U2757) );
  AOI22_X1 U21005 ( .A1(n19255), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17839) );
  OAI21_X1 U21006 ( .B1(n17903), .B2(n17852), .A(n17839), .ZN(P3_U2758) );
  AOI22_X1 U21007 ( .A1(n19255), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17840) );
  OAI21_X1 U21008 ( .B1(n17901), .B2(n17852), .A(n17840), .ZN(P3_U2759) );
  INV_X1 U21009 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17899) );
  AOI22_X1 U21010 ( .A1(n19255), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17841) );
  OAI21_X1 U21011 ( .B1(n17899), .B2(n17852), .A(n17841), .ZN(P3_U2760) );
  INV_X1 U21012 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17897) );
  AOI22_X1 U21013 ( .A1(n17842), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17843) );
  OAI21_X1 U21014 ( .B1(n17897), .B2(n17852), .A(n17843), .ZN(P3_U2761) );
  INV_X1 U21015 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17895) );
  AOI22_X1 U21016 ( .A1(n19255), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17844) );
  OAI21_X1 U21017 ( .B1(n17895), .B2(n17852), .A(n17844), .ZN(P3_U2762) );
  INV_X1 U21018 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17893) );
  AOI22_X1 U21019 ( .A1(n19255), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17845) );
  OAI21_X1 U21020 ( .B1(n17893), .B2(n17852), .A(n17845), .ZN(P3_U2763) );
  AOI22_X1 U21021 ( .A1(n19255), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17846) );
  OAI21_X1 U21022 ( .B1(n17891), .B2(n17852), .A(n17846), .ZN(P3_U2764) );
  AOI22_X1 U21023 ( .A1(n19255), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17847) );
  OAI21_X1 U21024 ( .B1(n17889), .B2(n17852), .A(n17847), .ZN(P3_U2765) );
  INV_X1 U21025 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17887) );
  AOI22_X1 U21026 ( .A1(n19255), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17848), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17849) );
  OAI21_X1 U21027 ( .B1(n17887), .B2(n17852), .A(n17849), .ZN(P3_U2766) );
  AOI22_X1 U21028 ( .A1(n19255), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17850), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17851) );
  OAI21_X1 U21029 ( .B1(n17885), .B2(n17852), .A(n17851), .ZN(P3_U2767) );
  INV_X1 U21030 ( .A(n17853), .ZN(n17854) );
  AOI22_X1 U21031 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17917), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17908), .ZN(n17856) );
  OAI21_X1 U21032 ( .B1(n17857), .B2(n17919), .A(n17856), .ZN(P3_U2768) );
  AOI22_X1 U21033 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17917), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17908), .ZN(n17858) );
  OAI21_X1 U21034 ( .B1(n17859), .B2(n17919), .A(n17858), .ZN(P3_U2769) );
  AOI22_X1 U21035 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17917), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17908), .ZN(n17860) );
  OAI21_X1 U21036 ( .B1(n17861), .B2(n17919), .A(n17860), .ZN(P3_U2770) );
  AOI22_X1 U21037 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17908), .ZN(n17862) );
  OAI21_X1 U21038 ( .B1(n17863), .B2(n17919), .A(n17862), .ZN(P3_U2771) );
  AOI22_X1 U21039 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17908), .ZN(n17864) );
  OAI21_X1 U21040 ( .B1(n17865), .B2(n17919), .A(n17864), .ZN(P3_U2772) );
  AOI22_X1 U21041 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17908), .ZN(n17866) );
  OAI21_X1 U21042 ( .B1(n17867), .B2(n17919), .A(n17866), .ZN(P3_U2773) );
  AOI22_X1 U21043 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17908), .ZN(n17868) );
  OAI21_X1 U21044 ( .B1(n17869), .B2(n17919), .A(n17868), .ZN(P3_U2774) );
  AOI22_X1 U21045 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17908), .ZN(n17870) );
  OAI21_X1 U21046 ( .B1(n10263), .B2(n17919), .A(n17870), .ZN(P3_U2775) );
  AOI22_X1 U21047 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17908), .ZN(n17871) );
  OAI21_X1 U21048 ( .B1(n17872), .B2(n17919), .A(n17871), .ZN(P3_U2776) );
  AOI22_X1 U21049 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17908), .ZN(n17873) );
  OAI21_X1 U21050 ( .B1(n17874), .B2(n17919), .A(n17873), .ZN(P3_U2777) );
  AOI22_X1 U21051 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17908), .ZN(n17875) );
  OAI21_X1 U21052 ( .B1(n17876), .B2(n17919), .A(n17875), .ZN(P3_U2778) );
  AOI22_X1 U21053 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17909), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17908), .ZN(n17877) );
  OAI21_X1 U21054 ( .B1(n17878), .B2(n17919), .A(n17877), .ZN(P3_U2779) );
  AOI22_X1 U21055 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17917), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17908), .ZN(n17879) );
  OAI21_X1 U21056 ( .B1(n21310), .B2(n17919), .A(n17879), .ZN(P3_U2780) );
  AOI22_X1 U21057 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17917), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17908), .ZN(n17880) );
  OAI21_X1 U21058 ( .B1(n17881), .B2(n17919), .A(n17880), .ZN(P3_U2781) );
  AOI22_X1 U21059 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17917), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17908), .ZN(n17882) );
  OAI21_X1 U21060 ( .B1(n17883), .B2(n17919), .A(n17882), .ZN(P3_U2782) );
  AOI22_X1 U21061 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17908), .ZN(n17884) );
  OAI21_X1 U21062 ( .B1(n17885), .B2(n17919), .A(n17884), .ZN(P3_U2783) );
  AOI22_X1 U21063 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17908), .ZN(n17886) );
  OAI21_X1 U21064 ( .B1(n17887), .B2(n17919), .A(n17886), .ZN(P3_U2784) );
  AOI22_X1 U21065 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17908), .ZN(n17888) );
  OAI21_X1 U21066 ( .B1(n17889), .B2(n17919), .A(n17888), .ZN(P3_U2785) );
  AOI22_X1 U21067 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17908), .ZN(n17890) );
  OAI21_X1 U21068 ( .B1(n17891), .B2(n17919), .A(n17890), .ZN(P3_U2786) );
  AOI22_X1 U21069 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17916), .ZN(n17892) );
  OAI21_X1 U21070 ( .B1(n17893), .B2(n17919), .A(n17892), .ZN(P3_U2787) );
  AOI22_X1 U21071 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17916), .ZN(n17894) );
  OAI21_X1 U21072 ( .B1(n17895), .B2(n17919), .A(n17894), .ZN(P3_U2788) );
  AOI22_X1 U21073 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17916), .ZN(n17896) );
  OAI21_X1 U21074 ( .B1(n17897), .B2(n17919), .A(n17896), .ZN(P3_U2789) );
  AOI22_X1 U21075 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17916), .ZN(n17898) );
  OAI21_X1 U21076 ( .B1(n17899), .B2(n17919), .A(n17898), .ZN(P3_U2790) );
  AOI22_X1 U21077 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17916), .ZN(n17900) );
  OAI21_X1 U21078 ( .B1(n17901), .B2(n17919), .A(n17900), .ZN(P3_U2791) );
  AOI22_X1 U21079 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17916), .ZN(n17902) );
  OAI21_X1 U21080 ( .B1(n17903), .B2(n17919), .A(n17902), .ZN(P3_U2792) );
  AOI22_X1 U21081 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17909), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17908), .ZN(n17904) );
  OAI21_X1 U21082 ( .B1(n17905), .B2(n17919), .A(n17904), .ZN(P3_U2793) );
  AOI22_X1 U21083 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17916), .ZN(n17906) );
  OAI21_X1 U21084 ( .B1(n17907), .B2(n17919), .A(n17906), .ZN(P3_U2794) );
  AOI22_X1 U21085 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17909), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17908), .ZN(n17910) );
  OAI21_X1 U21086 ( .B1(n17911), .B2(n17919), .A(n17910), .ZN(P3_U2795) );
  AOI22_X1 U21087 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17916), .ZN(n17912) );
  OAI21_X1 U21088 ( .B1(n17913), .B2(n17919), .A(n17912), .ZN(P3_U2796) );
  AOI22_X1 U21089 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17916), .ZN(n17914) );
  OAI21_X1 U21090 ( .B1(n17915), .B2(n17919), .A(n17914), .ZN(P3_U2797) );
  AOI22_X1 U21091 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17917), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17916), .ZN(n17918) );
  OAI21_X1 U21092 ( .B1(n17920), .B2(n17919), .A(n17918), .ZN(P3_U2798) );
  NAND4_X1 U21093 ( .A1(n18321), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(n18068), .ZN(n17944) );
  NAND2_X1 U21094 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17921), .ZN(
        n17938) );
  NOR2_X1 U21095 ( .A1(n18261), .A2(n18202), .ZN(n18015) );
  OAI22_X1 U21096 ( .A1(n18303), .A2(n18293), .B1(n18302), .B2(n18122), .ZN(
        n17957) );
  NOR2_X1 U21097 ( .A1(n18307), .A2(n17957), .ZN(n17943) );
  NOR3_X1 U21098 ( .A1(n18015), .A2(n17943), .A3(n17921), .ZN(n17931) );
  NAND2_X1 U21099 ( .A1(n18127), .A2(n17922), .ZN(n17928) );
  NOR3_X1 U21100 ( .A1(n18018), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17923), .ZN(n17946) );
  OAI21_X1 U21101 ( .B1(n12629), .B2(n18251), .A(n18289), .ZN(n17924) );
  AOI21_X1 U21102 ( .B1(n18051), .B2(n17925), .A(n17924), .ZN(n17950) );
  OAI21_X1 U21103 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18008), .A(
        n17950), .ZN(n17947) );
  OAI21_X1 U21104 ( .B1(n17946), .B2(n17947), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17927) );
  NAND2_X1 U21105 ( .A1(n9732), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17926) );
  OAI211_X1 U21106 ( .C1(n17929), .C2(n17928), .A(n17927), .B(n17926), .ZN(
        n17930) );
  AOI211_X1 U21107 ( .C1(n18145), .C2(n17932), .A(n17931), .B(n17930), .ZN(
        n17937) );
  OAI211_X1 U21108 ( .C1(n17935), .C2(n17934), .A(n18200), .B(n17933), .ZN(
        n17936) );
  OAI211_X1 U21109 ( .C1(n17944), .C2(n17938), .A(n17937), .B(n17936), .ZN(
        P3_U2802) );
  NOR2_X1 U21110 ( .A1(n17940), .A2(n17939), .ZN(n17941) );
  XNOR2_X1 U21111 ( .A(n17941), .B(n18117), .ZN(n18311) );
  AOI22_X1 U21112 ( .A1(n9732), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n18145), 
        .B2(n17942), .ZN(n17949) );
  AOI21_X1 U21113 ( .B1(n18307), .B2(n17944), .A(n17943), .ZN(n17945) );
  AOI211_X1 U21114 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17947), .A(
        n17946), .B(n17945), .ZN(n17948) );
  OAI211_X1 U21115 ( .C1(n18311), .C2(n18164), .A(n17949), .B(n17948), .ZN(
        P3_U2803) );
  NAND3_X1 U21116 ( .A1(n18321), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n18068), .ZN(n17960) );
  INV_X1 U21117 ( .A(n18008), .ZN(n17992) );
  NOR2_X1 U21118 ( .A1(n18481), .A2(n19184), .ZN(n18315) );
  AOI221_X1 U21119 ( .B1(n18639), .B2(n17952), .C1(n17951), .C2(n17952), .A(
        n17950), .ZN(n17953) );
  AOI211_X1 U21120 ( .C1(n17954), .C2(n18281), .A(n18315), .B(n17953), .ZN(
        n17959) );
  OAI21_X1 U21121 ( .B1(n17956), .B2(n18317), .A(n17955), .ZN(n18316) );
  AOI22_X1 U21122 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17957), .B1(
        n18200), .B2(n18316), .ZN(n17958) );
  OAI211_X1 U21123 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17960), .A(
        n17959), .B(n17958), .ZN(P3_U2804) );
  OAI21_X1 U21124 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17962), .A(
        n17961), .ZN(n18331) );
  NAND2_X1 U21125 ( .A1(n12628), .A2(n18127), .ZN(n17979) );
  AOI221_X1 U21126 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C1(n17978), .C2(n17965), .A(
        n17979), .ZN(n17967) );
  OAI22_X1 U21127 ( .A1(n18639), .A2(n12628), .B1(n19123), .B2(n17963), .ZN(
        n17964) );
  INV_X1 U21128 ( .A(n18289), .ZN(n18259) );
  OR2_X1 U21129 ( .A1(n17964), .A2(n18259), .ZN(n17996) );
  AOI21_X1 U21130 ( .B1(n17992), .B2(n17993), .A(n17996), .ZN(n17977) );
  OAI22_X1 U21131 ( .A1(n17977), .A2(n17965), .B1(n18481), .B2(n19182), .ZN(
        n17966) );
  AOI211_X1 U21132 ( .C1(n17968), .C2(n18145), .A(n17967), .B(n17966), .ZN(
        n17974) );
  XNOR2_X1 U21133 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17969), .ZN(
        n18328) );
  OAI21_X1 U21134 ( .B1(n18199), .B2(n17970), .A(n17971), .ZN(n17972) );
  XNOR2_X1 U21135 ( .A(n17972), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18327) );
  AOI22_X1 U21136 ( .A1(n18261), .A2(n18328), .B1(n18200), .B2(n18327), .ZN(
        n17973) );
  OAI211_X1 U21137 ( .C1(n18122), .C2(n18331), .A(n17974), .B(n17973), .ZN(
        P3_U2805) );
  OAI21_X1 U21138 ( .B1(n9849), .B2(n18296), .A(n17975), .ZN(n18333) );
  INV_X1 U21139 ( .A(n18333), .ZN(n17987) );
  NAND2_X1 U21140 ( .A1(n9732), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17976) );
  OAI221_X1 U21141 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17979), .C1(
        n17978), .C2(n17977), .A(n17976), .ZN(n17980) );
  AOI21_X1 U21142 ( .B1(n18145), .B2(n17981), .A(n17980), .ZN(n17986) );
  NAND2_X1 U21143 ( .A1(n18016), .A2(n17982), .ZN(n18335) );
  AOI22_X1 U21144 ( .A1(n18334), .A2(n18202), .B1(n18335), .B2(n18261), .ZN(
        n17983) );
  INV_X1 U21145 ( .A(n17983), .ZN(n18002) );
  NOR2_X1 U21146 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17984), .ZN(
        n18332) );
  AOI22_X1 U21147 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18002), .B1(
        n18068), .B2(n18332), .ZN(n17985) );
  OAI211_X1 U21148 ( .C1(n17987), .C2(n18164), .A(n17986), .B(n17985), .ZN(
        P3_U2806) );
  OAI22_X1 U21149 ( .A1(n18199), .A2(n21331), .B1(n17988), .B2(n18010), .ZN(
        n17990) );
  NOR2_X1 U21150 ( .A1(n17990), .A2(n18011), .ZN(n17991) );
  XNOR2_X1 U21151 ( .A(n17991), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18350) );
  NAND2_X1 U21152 ( .A1(n17992), .A2(n17993), .ZN(n18000) );
  OAI21_X1 U21153 ( .B1(n18639), .B2(n17994), .A(n17993), .ZN(n17995) );
  AOI22_X1 U21154 ( .A1(n18145), .A2(n17997), .B1(n17996), .B2(n17995), .ZN(
        n17998) );
  NAND2_X1 U21155 ( .A1(n9732), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18348) );
  OAI211_X1 U21156 ( .C1(n18000), .C2(n17999), .A(n17998), .B(n18348), .ZN(
        n18001) );
  AOI21_X1 U21157 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18002), .A(
        n18001), .ZN(n18004) );
  INV_X1 U21158 ( .A(n18068), .ZN(n18095) );
  OAI211_X1 U21159 ( .C1(n18350), .C2(n18164), .A(n18004), .B(n18003), .ZN(
        P3_U2807) );
  OAI21_X1 U21160 ( .B1(n18005), .B2(n18251), .A(n18289), .ZN(n18006) );
  AOI21_X1 U21161 ( .B1(n18051), .B2(n18007), .A(n18006), .ZN(n18045) );
  OAI21_X1 U21162 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18008), .A(
        n18045), .ZN(n18024) );
  AOI22_X1 U21163 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18024), .B1(
        n18145), .B2(n18009), .ZN(n18021) );
  INV_X1 U21164 ( .A(n18010), .ZN(n18013) );
  AOI21_X1 U21165 ( .B1(n18013), .B2(n18012), .A(n18011), .ZN(n18014) );
  XNOR2_X1 U21166 ( .A(n18014), .B(n21331), .ZN(n18362) );
  INV_X1 U21167 ( .A(n18015), .ZN(n18039) );
  OAI22_X1 U21168 ( .A1(n18016), .A2(n18293), .B1(n18352), .B2(n18122), .ZN(
        n18092) );
  NAND2_X1 U21169 ( .A1(n9732), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18363) );
  NOR2_X1 U21170 ( .A1(n18018), .A2(n18017), .ZN(n18026) );
  OAI211_X1 U21171 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18026), .B(n18019), .ZN(n18020) );
  INV_X1 U21172 ( .A(n18022), .ZN(n18034) );
  NOR2_X1 U21173 ( .A1(n18481), .A2(n19175), .ZN(n18023) );
  AOI221_X1 U21174 ( .B1(n18026), .B2(n18025), .C1(n18024), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18023), .ZN(n18033) );
  NOR3_X1 U21175 ( .A1(n18071), .A2(n18117), .A3(n18027), .ZN(n18036) );
  INV_X1 U21176 ( .A(n18036), .ZN(n18046) );
  OAI22_X1 U21177 ( .A1(n18031), .A2(n18046), .B1(n18028), .B2(n18029), .ZN(
        n18030) );
  XNOR2_X1 U21178 ( .A(n18357), .B(n18030), .ZN(n18367) );
  INV_X1 U21179 ( .A(n18031), .ZN(n18369) );
  NAND2_X1 U21180 ( .A1(n18369), .A2(n18357), .ZN(n18374) );
  AOI21_X1 U21181 ( .B1(n12635), .B2(n18998), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18044) );
  AOI22_X1 U21182 ( .A1(n9732), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18035), 
        .B2(n18281), .ZN(n18043) );
  OAI221_X1 U21183 ( .B1(n18037), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), 
        .C1(n18037), .C2(n18036), .A(n17989), .ZN(n18038) );
  XNOR2_X1 U21184 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18038), .ZN(
        n18375) );
  NAND2_X1 U21185 ( .A1(n18366), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18377) );
  AOI21_X1 U21186 ( .B1(n18039), .B2(n18377), .A(n18092), .ZN(n18056) );
  NAND2_X1 U21187 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18040), .ZN(
        n18383) );
  OAI22_X1 U21188 ( .A1(n18056), .A2(n18040), .B1(n18383), .B2(n18058), .ZN(
        n18041) );
  AOI21_X1 U21189 ( .B1(n18200), .B2(n18375), .A(n18041), .ZN(n18042) );
  OAI211_X1 U21190 ( .C1(n18045), .C2(n18044), .A(n18043), .B(n18042), .ZN(
        P3_U2810) );
  INV_X1 U21191 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18057) );
  OAI21_X1 U21192 ( .B1(n18065), .B2(n18028), .A(n18046), .ZN(n18047) );
  XOR2_X1 U21193 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n18047), .Z(
        n18384) );
  OAI211_X1 U21194 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17156), .B(n18127), .ZN(n18049) );
  OAI22_X1 U21195 ( .A1(n10643), .A2(n18049), .B1(n18048), .B2(n18140), .ZN(
        n18054) );
  OAI21_X1 U21196 ( .B1(n17156), .B2(n18251), .A(n18289), .ZN(n18074) );
  AOI21_X1 U21197 ( .B1(n18051), .B2(n18050), .A(n18074), .ZN(n18060) );
  NAND2_X1 U21198 ( .A1(n9732), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18386) );
  OAI21_X1 U21199 ( .B1(n18060), .B2(n18052), .A(n18386), .ZN(n18053) );
  AOI211_X1 U21200 ( .C1(n18200), .C2(n18384), .A(n18054), .B(n18053), .ZN(
        n18055) );
  OAI221_X1 U21201 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18058), 
        .C1(n18057), .C2(n18056), .A(n18055), .ZN(P3_U2811) );
  AOI21_X1 U21202 ( .B1(n18068), .B2(n18067), .A(n18092), .ZN(n18077) );
  NAND2_X1 U21203 ( .A1(n17156), .A2(n18127), .ZN(n18062) );
  NAND2_X1 U21204 ( .A1(n9732), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18059) );
  OAI221_X1 U21205 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18062), .C1(
        n18061), .C2(n18060), .A(n18059), .ZN(n18063) );
  AOI21_X1 U21206 ( .B1(n18145), .B2(n18064), .A(n18063), .ZN(n18070) );
  OAI21_X1 U21207 ( .B1(n18071), .B2(n18117), .A(n18065), .ZN(n18066) );
  XOR2_X1 U21208 ( .A(n18028), .B(n18066), .Z(n18402) );
  NOR2_X1 U21209 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18067), .ZN(
        n18401) );
  AOI22_X1 U21210 ( .A1(n18200), .A2(n18402), .B1(n18068), .B2(n18401), .ZN(
        n18069) );
  OAI211_X1 U21211 ( .C1(n18077), .C2(n18071), .A(n18070), .B(n18069), .ZN(
        P3_U2812) );
  OAI21_X1 U21212 ( .B1(n17139), .B2(n18639), .A(n18072), .ZN(n18073) );
  AOI22_X1 U21213 ( .A1(n9732), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18074), 
        .B2(n18073), .ZN(n18080) );
  OAI21_X1 U21214 ( .B1(n18076), .B2(n18396), .A(n18075), .ZN(n18405) );
  NAND2_X1 U21215 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18396), .ZN(
        n18410) );
  OAI22_X1 U21216 ( .A1(n18077), .A2(n18396), .B1(n18095), .B2(n18410), .ZN(
        n18078) );
  AOI21_X1 U21217 ( .B1(n18200), .B2(n18405), .A(n18078), .ZN(n18079) );
  OAI211_X1 U21218 ( .C1(n18272), .C2(n18081), .A(n18080), .B(n18079), .ZN(
        P3_U2813) );
  OAI21_X1 U21219 ( .B1(n18251), .B2(n9917), .A(n18289), .ZN(n18082) );
  INV_X1 U21220 ( .A(n18082), .ZN(n18110) );
  OAI21_X1 U21221 ( .B1(n18083), .B2(n19123), .A(n18110), .ZN(n18100) );
  NAND2_X1 U21222 ( .A1(n9917), .A2(n18127), .ZN(n18097) );
  AOI221_X1 U21223 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n18085), .C2(n18084), .A(
        n18097), .ZN(n18088) );
  OAI22_X1 U21224 ( .A1(n18481), .A2(n19165), .B1(n18140), .B2(n18086), .ZN(
        n18087) );
  AOI211_X1 U21225 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n18100), .A(
        n18088), .B(n18087), .ZN(n18094) );
  AOI21_X1 U21226 ( .B1(n18199), .B2(n18090), .A(n18089), .ZN(n18091) );
  XNOR2_X1 U21227 ( .A(n18091), .B(n18417), .ZN(n18419) );
  AOI22_X1 U21228 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18092), .B1(
        n18200), .B2(n18419), .ZN(n18093) );
  OAI211_X1 U21229 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18095), .A(
        n18094), .B(n18093), .ZN(P3_U2814) );
  NOR2_X1 U21230 ( .A1(n18429), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18108) );
  NAND2_X1 U21231 ( .A1(n18261), .A2(n18428), .ZN(n18107) );
  NOR2_X1 U21232 ( .A1(n18481), .A2(n19163), .ZN(n18099) );
  OAI22_X1 U21233 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18097), .B1(
        n18096), .B2(n18140), .ZN(n18098) );
  AOI211_X1 U21234 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18100), .A(
        n18099), .B(n18098), .ZN(n18106) );
  INV_X1 U21235 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18460) );
  NOR4_X1 U21236 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n18199), .A4(n18165), .ZN(
        n18153) );
  NAND2_X1 U21237 ( .A1(n18153), .A2(n18154), .ZN(n18141) );
  AOI22_X1 U21238 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18101), .B1(
        n18141), .B2(n18135), .ZN(n18102) );
  OAI221_X1 U21239 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18441), 
        .C1(n18460), .C2(n18199), .A(n18102), .ZN(n18103) );
  XNOR2_X1 U21240 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18103), .ZN(
        n18432) );
  NOR2_X1 U21241 ( .A1(n18352), .A2(n18122), .ZN(n18104) );
  NAND2_X1 U21242 ( .A1(n18423), .A2(n18109), .ZN(n18426) );
  AOI22_X1 U21243 ( .A1(n18200), .A2(n18432), .B1(n18104), .B2(n18426), .ZN(
        n18105) );
  OAI211_X1 U21244 ( .C1(n18108), .C2(n18107), .A(n18106), .B(n18105), .ZN(
        P3_U2815) );
  OAI221_X1 U21245 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18475), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n9770), .A(n18109), .ZN(
        n18448) );
  AOI221_X1 U21246 ( .B1(n18639), .B2(n18112), .C1(n18111), .C2(n18112), .A(
        n18110), .ZN(n18113) );
  NOR2_X1 U21247 ( .A1(n18481), .A2(n21405), .ZN(n18443) );
  AOI211_X1 U21248 ( .C1(n18114), .C2(n18281), .A(n18113), .B(n18443), .ZN(
        n18121) );
  AOI21_X1 U21249 ( .B1(n18441), .B2(n18115), .A(n18429), .ZN(n18445) );
  NOR2_X1 U21250 ( .A1(n18117), .A2(n18116), .ZN(n18184) );
  NAND2_X1 U21251 ( .A1(n18436), .A2(n18184), .ZN(n18133) );
  NAND2_X1 U21252 ( .A1(n18460), .A2(n18135), .ZN(n18118) );
  OAI22_X1 U21253 ( .A1(n18135), .A2(n18133), .B1(n18118), .B2(n18141), .ZN(
        n18119) );
  XNOR2_X1 U21254 ( .A(n18441), .B(n18119), .ZN(n18444) );
  AOI22_X1 U21255 ( .A1(n18261), .A2(n18445), .B1(n18200), .B2(n18444), .ZN(
        n18120) );
  OAI211_X1 U21256 ( .C1(n18122), .C2(n18448), .A(n18121), .B(n18120), .ZN(
        P3_U2816) );
  AOI21_X1 U21257 ( .B1(n18124), .B2(n17198), .A(n18259), .ZN(n18210) );
  NAND2_X1 U21258 ( .A1(n18124), .A2(n18123), .ZN(n18125) );
  OAI211_X1 U21259 ( .C1(n18126), .C2(n19123), .A(n18210), .B(n18125), .ZN(
        n18146) );
  NAND2_X1 U21260 ( .A1(n17200), .A2(n18127), .ZN(n18148) );
  AOI211_X1 U21261 ( .C1(n18130), .C2(n18129), .A(n18128), .B(n18148), .ZN(
        n18132) );
  NOR2_X1 U21262 ( .A1(n18481), .A2(n19160), .ZN(n18131) );
  AOI211_X1 U21263 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18146), .A(
        n18132), .B(n18131), .ZN(n18138) );
  OAI21_X1 U21264 ( .B1(n18141), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18133), .ZN(n18134) );
  XNOR2_X1 U21265 ( .A(n18134), .B(n18135), .ZN(n18450) );
  NAND2_X1 U21266 ( .A1(n18436), .A2(n18135), .ZN(n18459) );
  NAND2_X1 U21267 ( .A1(n18436), .A2(n18475), .ZN(n18451) );
  AOI22_X1 U21268 ( .A1(n18261), .A2(n18453), .B1(n18202), .B2(n18451), .ZN(
        n18151) );
  OAI22_X1 U21269 ( .A1(n18167), .A2(n18459), .B1(n18151), .B2(n18135), .ZN(
        n18136) );
  AOI21_X1 U21270 ( .B1(n18200), .B2(n18450), .A(n18136), .ZN(n18137) );
  OAI211_X1 U21271 ( .C1(n18140), .C2(n18139), .A(n18138), .B(n18137), .ZN(
        P3_U2817) );
  INV_X1 U21272 ( .A(n18167), .ZN(n18186) );
  NAND2_X1 U21273 ( .A1(n18480), .A2(n18186), .ZN(n18152) );
  INV_X1 U21274 ( .A(n18477), .ZN(n18169) );
  NAND2_X1 U21275 ( .A1(n18169), .A2(n18184), .ZN(n18142) );
  OAI21_X1 U21276 ( .B1(n18154), .B2(n18142), .A(n18141), .ZN(n18143) );
  XNOR2_X1 U21277 ( .A(n18143), .B(n18460), .ZN(n18464) );
  AOI22_X1 U21278 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18146), .B1(
        n18145), .B2(n18144), .ZN(n18147) );
  NAND2_X1 U21279 ( .A1(n9732), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18465) );
  OAI211_X1 U21280 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n18148), .A(
        n18147), .B(n18465), .ZN(n18149) );
  AOI21_X1 U21281 ( .B1(n18200), .B2(n18464), .A(n18149), .ZN(n18150) );
  OAI221_X1 U21282 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18152), 
        .C1(n18460), .C2(n18151), .A(n18150), .ZN(P3_U2818) );
  AOI21_X1 U21283 ( .B1(n18184), .B2(n18169), .A(n18153), .ZN(n18155) );
  XNOR2_X1 U21284 ( .A(n18155), .B(n18154), .ZN(n18486) );
  NAND4_X1 U21285 ( .A1(n18209), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18998), .A4(n18192), .ZN(n18179) );
  NOR2_X1 U21286 ( .A1(n18178), .A2(n18179), .ZN(n18177) );
  NAND2_X1 U21287 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18177), .ZN(
        n18170) );
  NAND2_X1 U21288 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18218), .ZN(
        n18156) );
  AOI22_X1 U21289 ( .A1(n18998), .A2(n17200), .B1(n18170), .B2(n18156), .ZN(
        n18158) );
  INV_X1 U21290 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19156) );
  NOR2_X1 U21291 ( .A1(n18481), .A2(n19156), .ZN(n18157) );
  AOI211_X1 U21292 ( .C1(n18159), .C2(n18281), .A(n18158), .B(n18157), .ZN(
        n18163) );
  AOI22_X1 U21293 ( .A1(n18261), .A2(n18473), .B1(n18202), .B2(n18160), .ZN(
        n18189) );
  OAI21_X1 U21294 ( .B1(n18169), .B2(n18167), .A(n18189), .ZN(n18161) );
  NOR2_X1 U21295 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18477), .ZN(
        n18469) );
  AOI22_X1 U21296 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18161), .B1(
        n18469), .B2(n18186), .ZN(n18162) );
  OAI211_X1 U21297 ( .C1(n18486), .C2(n18164), .A(n18163), .B(n18162), .ZN(
        P3_U2819) );
  NOR2_X1 U21298 ( .A1(n18199), .A2(n18165), .ZN(n18183) );
  AOI22_X1 U21299 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18184), .B1(
        n18183), .B2(n12119), .ZN(n18166) );
  XNOR2_X1 U21300 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18166), .ZN(
        n18490) );
  NOR2_X1 U21301 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18168) );
  NOR3_X1 U21302 ( .A1(n18169), .A2(n18168), .A3(n18167), .ZN(n18175) );
  OAI211_X1 U21303 ( .C1(n18177), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18218), .B(n18170), .ZN(n18172) );
  NAND2_X1 U21304 ( .A1(n9732), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18171) );
  OAI211_X1 U21305 ( .C1(n18272), .C2(n18173), .A(n18172), .B(n18171), .ZN(
        n18174) );
  AOI211_X1 U21306 ( .C1(n18200), .C2(n18490), .A(n18175), .B(n18174), .ZN(
        n18176) );
  OAI21_X1 U21307 ( .B1(n18189), .B2(n12120), .A(n18176), .ZN(P3_U2820) );
  INV_X1 U21308 ( .A(n18218), .ZN(n18286) );
  AOI211_X1 U21309 ( .C1(n18179), .C2(n18178), .A(n18286), .B(n18177), .ZN(
        n18181) );
  NOR2_X1 U21310 ( .A1(n18481), .A2(n19153), .ZN(n18180) );
  AOI211_X1 U21311 ( .C1(n18182), .C2(n18281), .A(n18181), .B(n18180), .ZN(
        n18188) );
  NOR2_X1 U21312 ( .A1(n18184), .A2(n18183), .ZN(n18185) );
  XNOR2_X1 U21313 ( .A(n18185), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18495) );
  AOI22_X1 U21314 ( .A1(n18200), .A2(n18495), .B1(n12119), .B2(n18186), .ZN(
        n18187) );
  OAI211_X1 U21315 ( .C1(n18189), .C2(n12119), .A(n18188), .B(n18187), .ZN(
        P3_U2821) );
  OAI21_X1 U21316 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18191), .A(
        n18190), .ZN(n18510) );
  OR2_X1 U21317 ( .A1(n17198), .A2(n21384), .ZN(n18193) );
  AOI211_X1 U21318 ( .C1(n18194), .C2(n18193), .A(n18192), .B(n18639), .ZN(
        n18197) );
  OAI22_X1 U21319 ( .A1(n18272), .A2(n18195), .B1(n18210), .B2(n18194), .ZN(
        n18196) );
  AOI211_X1 U21320 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n9732), .A(n18197), .B(
        n18196), .ZN(n18204) );
  INV_X1 U21321 ( .A(n18509), .ZN(n18201) );
  AOI21_X1 U21322 ( .B1(n18199), .B2(n18509), .A(n18198), .ZN(n18513) );
  AOI22_X1 U21323 ( .A1(n18202), .A2(n18201), .B1(n18200), .B2(n18513), .ZN(
        n18203) );
  OAI211_X1 U21324 ( .C1(n18293), .C2(n18510), .A(n18204), .B(n18203), .ZN(
        P3_U2822) );
  OAI21_X1 U21325 ( .B1(n18207), .B2(n18206), .A(n18205), .ZN(n18208) );
  XNOR2_X1 U21326 ( .A(n18208), .B(n18504), .ZN(n18519) );
  INV_X1 U21327 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21271) );
  NAND2_X1 U21328 ( .A1(n18998), .A2(n18209), .ZN(n18222) );
  NOR2_X1 U21329 ( .A1(n21271), .A2(n18222), .ZN(n18212) );
  INV_X1 U21330 ( .A(n18210), .ZN(n18211) );
  INV_X1 U21331 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19149) );
  NOR2_X1 U21332 ( .A1(n18481), .A2(n19149), .ZN(n18523) );
  AOI221_X1 U21333 ( .B1(n18212), .B2(n21384), .C1(n18211), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18523), .ZN(n18217) );
  AOI21_X1 U21334 ( .B1(n18504), .B2(n18214), .A(n18213), .ZN(n18517) );
  AOI22_X1 U21335 ( .A1(n18282), .A2(n18517), .B1(n18215), .B2(n18281), .ZN(
        n18216) );
  OAI211_X1 U21336 ( .C1(n18293), .C2(n18519), .A(n18217), .B(n18216), .ZN(
        P3_U2823) );
  NAND2_X1 U21337 ( .A1(n18218), .A2(n18222), .ZN(n18236) );
  AOI21_X1 U21338 ( .B1(n18221), .B2(n18220), .A(n18219), .ZN(n18530) );
  OAI22_X1 U21339 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18222), .B1(
        n18481), .B2(n19147), .ZN(n18227) );
  OAI21_X1 U21340 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18224), .A(
        n18223), .ZN(n18533) );
  OAI22_X1 U21341 ( .A1(n18272), .A2(n18225), .B1(n18293), .B2(n18533), .ZN(
        n18226) );
  AOI211_X1 U21342 ( .C1(n18282), .C2(n18530), .A(n18227), .B(n18226), .ZN(
        n18228) );
  OAI21_X1 U21343 ( .B1(n21271), .B2(n18236), .A(n18228), .ZN(P3_U2824) );
  OAI21_X1 U21344 ( .B1(n18231), .B2(n18230), .A(n18229), .ZN(n18540) );
  AOI21_X1 U21345 ( .B1(n18232), .B2(n18234), .A(n18233), .ZN(n18235) );
  XNOR2_X1 U21346 ( .A(n18235), .B(n10560), .ZN(n18537) );
  AOI22_X1 U21347 ( .A1(n18282), .A2(n18537), .B1(n9732), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18242) );
  AOI221_X1 U21348 ( .B1(n18259), .B2(n18238), .C1(n18237), .C2(n18238), .A(
        n18236), .ZN(n18239) );
  AOI21_X1 U21349 ( .B1(n18240), .B2(n18281), .A(n18239), .ZN(n18241) );
  OAI211_X1 U21350 ( .C1(n18293), .C2(n18540), .A(n18242), .B(n18241), .ZN(
        P3_U2825) );
  OAI21_X1 U21351 ( .B1(n18244), .B2(n18544), .A(n18243), .ZN(n18541) );
  OAI22_X1 U21352 ( .A1(n18481), .A2(n19143), .B1(n18639), .B2(n18245), .ZN(
        n18246) );
  AOI21_X1 U21353 ( .B1(n18282), .B2(n18541), .A(n18246), .ZN(n18254) );
  AOI21_X1 U21354 ( .B1(n18249), .B2(n18248), .A(n18247), .ZN(n18250) );
  XNOR2_X1 U21355 ( .A(n18250), .B(n18544), .ZN(n18547) );
  OAI21_X1 U21356 ( .B1(n18252), .B2(n18251), .A(n18289), .ZN(n18260) );
  AOI22_X1 U21357 ( .A1(n18261), .A2(n18547), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18260), .ZN(n18253) );
  OAI211_X1 U21358 ( .C1(n18272), .C2(n18255), .A(n18254), .B(n18253), .ZN(
        P3_U2826) );
  AOI21_X1 U21359 ( .B1(n9897), .B2(n18257), .A(n18256), .ZN(n18551) );
  AOI22_X1 U21360 ( .A1(n18282), .A2(n18551), .B1(n18258), .B2(n18281), .ZN(
        n18264) );
  NOR2_X1 U21361 ( .A1(n18259), .A2(n18275), .ZN(n18276) );
  OAI21_X1 U21362 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18276), .A(
        n18260), .ZN(n18263) );
  NAND2_X1 U21363 ( .A1(n9732), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18561) );
  OAI211_X1 U21364 ( .C1(n18554), .C2(n18553), .A(n18261), .B(n18552), .ZN(
        n18262) );
  NAND4_X1 U21365 ( .A1(n18264), .A2(n18263), .A3(n18561), .A4(n18262), .ZN(
        P3_U2827) );
  AOI21_X1 U21366 ( .B1(n18267), .B2(n18266), .A(n18265), .ZN(n18575) );
  NOR2_X1 U21367 ( .A1(n18481), .A2(n19139), .ZN(n18577) );
  OAI21_X1 U21368 ( .B1(n18270), .B2(n18269), .A(n18268), .ZN(n18573) );
  OAI22_X1 U21369 ( .A1(n18272), .A2(n18271), .B1(n18293), .B2(n18573), .ZN(
        n18273) );
  AOI211_X1 U21370 ( .C1(n18282), .C2(n18575), .A(n18577), .B(n18273), .ZN(
        n18274) );
  OAI221_X1 U21371 ( .B1(n18276), .B2(n18639), .C1(n18276), .C2(n18275), .A(
        n18274), .ZN(P3_U2828) );
  NOR2_X1 U21372 ( .A1(n18288), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18277) );
  XOR2_X1 U21373 ( .A(n18277), .B(n18280), .Z(n18594) );
  OAI22_X1 U21374 ( .A1(n18293), .A2(n18594), .B1(n18481), .B2(n19241), .ZN(
        n18278) );
  INV_X1 U21375 ( .A(n18278), .ZN(n18284) );
  AOI21_X1 U21376 ( .B1(n18280), .B2(n18287), .A(n18279), .ZN(n18582) );
  AOI22_X1 U21377 ( .A1(n18282), .A2(n18582), .B1(n18285), .B2(n18281), .ZN(
        n18283) );
  OAI211_X1 U21378 ( .C1(n18286), .C2(n18285), .A(n18284), .B(n18283), .ZN(
        P3_U2829) );
  OAI21_X1 U21379 ( .B1(n18288), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18287), .ZN(n18601) );
  INV_X1 U21380 ( .A(n18601), .ZN(n18294) );
  NAND3_X1 U21381 ( .A1(n19221), .A2(n19123), .A3(n18289), .ZN(n18290) );
  AOI22_X1 U21382 ( .A1(n9732), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18290), .ZN(n18291) );
  OAI221_X1 U21383 ( .B1(n18294), .B2(n18293), .C1(n18601), .C2(n18292), .A(
        n18291), .ZN(P3_U2830) );
  AOI22_X1 U21384 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18588), .B1(
        n9732), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n18310) );
  NOR3_X1 U21385 ( .A1(n18345), .A2(n18295), .A3(n18344), .ZN(n18308) );
  NOR2_X1 U21386 ( .A1(n18338), .A2(n18296), .ZN(n18300) );
  INV_X1 U21387 ( .A(n18297), .ZN(n18356) );
  AOI21_X1 U21388 ( .B1(n18502), .B2(n18298), .A(n18356), .ZN(n18337) );
  OAI211_X1 U21389 ( .C1(n9743), .C2(n18300), .A(n18337), .B(n18299), .ZN(
        n18319) );
  OAI22_X1 U21390 ( .A1(n9780), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18301), .B2(n18587), .ZN(n18305) );
  OAI22_X1 U21391 ( .A1(n18303), .A2(n18574), .B1(n18302), .B2(n18508), .ZN(
        n18304) );
  OAI21_X1 U21392 ( .B1(n9780), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n18314), .ZN(n18306) );
  OAI221_X1 U21393 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18308), 
        .C1(n18307), .C2(n18306), .A(n18595), .ZN(n18309) );
  OAI211_X1 U21394 ( .C1(n18311), .C2(n18485), .A(n18310), .B(n18309), .ZN(
        P3_U2835) );
  AND2_X1 U21395 ( .A1(n18321), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18312) );
  AOI22_X1 U21396 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18595), .B1(
        n18365), .B2(n18312), .ZN(n18313) );
  INV_X1 U21397 ( .A(n18318), .ZN(n18449) );
  NOR2_X1 U21398 ( .A1(n18481), .A2(n19182), .ZN(n18326) );
  INV_X1 U21399 ( .A(n18319), .ZN(n18324) );
  NAND2_X1 U21400 ( .A1(n18321), .A2(n18320), .ZN(n18323) );
  AOI221_X1 U21401 ( .B1(n18324), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n18323), .C2(n18322), .A(n18586), .ZN(n18325) );
  AOI211_X1 U21402 ( .C1(n18588), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18326), .B(n18325), .ZN(n18330) );
  AOI22_X1 U21403 ( .A1(n18598), .A2(n18328), .B1(n18496), .B2(n18327), .ZN(
        n18329) );
  OAI211_X1 U21404 ( .C1(n18449), .C2(n18331), .A(n18330), .B(n18329), .ZN(
        P3_U2837) );
  AOI22_X1 U21405 ( .A1(n18496), .A2(n18333), .B1(n18365), .B2(n18332), .ZN(
        n18343) );
  INV_X1 U21406 ( .A(n18574), .ZN(n19058) );
  AOI22_X1 U21407 ( .A1(n19058), .A2(n18335), .B1(n18452), .B2(n18334), .ZN(
        n18336) );
  NAND3_X1 U21408 ( .A1(n18337), .A2(n18336), .A3(n18581), .ZN(n18341) );
  NOR3_X1 U21409 ( .A1(n18339), .A2(n18338), .A3(n18341), .ZN(n18340) );
  NOR2_X1 U21410 ( .A1(n9732), .A2(n18340), .ZN(n18346) );
  OAI211_X1 U21411 ( .C1(n18505), .C2(n18341), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18346), .ZN(n18342) );
  OAI211_X1 U21412 ( .C1(n19180), .C2(n18481), .A(n18343), .B(n18342), .ZN(
        P3_U2838) );
  NOR2_X1 U21413 ( .A1(n18345), .A2(n18344), .ZN(n18347) );
  OAI221_X1 U21414 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18347), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18581), .A(n18346), .ZN(
        n18349) );
  OAI211_X1 U21415 ( .C1(n18485), .C2(n18350), .A(n18349), .B(n18348), .ZN(
        P3_U2839) );
  OAI21_X1 U21416 ( .B1(n18586), .B2(n21331), .A(n18351), .ZN(n18361) );
  NOR2_X1 U21417 ( .A1(n18352), .A2(n18508), .ZN(n18427) );
  AOI21_X1 U21418 ( .B1(n19058), .B2(n18428), .A(n18427), .ZN(n18394) );
  NAND2_X1 U21419 ( .A1(n18574), .A2(n18508), .ZN(n18476) );
  OAI21_X1 U21420 ( .B1(n18389), .B2(n18377), .A(n19080), .ZN(n18353) );
  OAI221_X1 U21421 ( .B1(n19088), .B2(n18366), .C1(n19088), .C2(n18391), .A(
        n18353), .ZN(n18376) );
  AOI21_X1 U21422 ( .B1(n18354), .B2(n18476), .A(n18376), .ZN(n18355) );
  OAI211_X1 U21423 ( .C1(n9780), .C2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n18394), .B(n18355), .ZN(n18371) );
  AOI211_X1 U21424 ( .C1(n19080), .C2(n18357), .A(n18356), .B(n18371), .ZN(
        n18358) );
  OAI211_X1 U21425 ( .C1(n18359), .C2(n19088), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18358), .ZN(n18360) );
  AOI22_X1 U21426 ( .A1(n18496), .A2(n18362), .B1(n18361), .B2(n18360), .ZN(
        n18364) );
  OAI211_X1 U21427 ( .C1(n18581), .C2(n21331), .A(n18364), .B(n18363), .ZN(
        P3_U2840) );
  NAND2_X1 U21428 ( .A1(n18366), .A2(n18365), .ZN(n18388) );
  AOI22_X1 U21429 ( .A1(n9732), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18496), 
        .B2(n18367), .ZN(n18373) );
  OAI21_X1 U21430 ( .B1(n18368), .B2(n18413), .A(n18462), .ZN(n18378) );
  OAI211_X1 U21431 ( .C1(n18587), .C2(n18369), .A(n18378), .B(n18595), .ZN(
        n18370) );
  OAI211_X1 U21432 ( .C1(n18371), .C2(n18370), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18481), .ZN(n18372) );
  OAI211_X1 U21433 ( .C1(n18388), .C2(n18374), .A(n18373), .B(n18372), .ZN(
        P3_U2841) );
  AOI22_X1 U21434 ( .A1(n9732), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18496), 
        .B2(n18375), .ZN(n18382) );
  NAND2_X1 U21435 ( .A1(n18394), .A2(n18581), .ZN(n18416) );
  AOI211_X1 U21436 ( .C1(n18377), .C2(n18476), .A(n18416), .B(n18376), .ZN(
        n18379) );
  AOI21_X1 U21437 ( .B1(n18379), .B2(n18378), .A(n9732), .ZN(n18385) );
  NOR3_X1 U21438 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18587), .A3(
        n19273), .ZN(n18380) );
  OAI21_X1 U21439 ( .B1(n18385), .B2(n18380), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18381) );
  OAI211_X1 U21440 ( .C1(n18383), .C2(n18388), .A(n18382), .B(n18381), .ZN(
        P3_U2842) );
  AOI22_X1 U21441 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18385), .B1(
        n18496), .B2(n18384), .ZN(n18387) );
  OAI211_X1 U21442 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18388), .A(
        n18387), .B(n18386), .ZN(P3_U2843) );
  INV_X1 U21443 ( .A(n18502), .ZN(n18566) );
  NOR2_X1 U21444 ( .A1(n19064), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18568) );
  NOR3_X1 U21445 ( .A1(n18568), .A2(n18389), .A3(n18417), .ZN(n18395) );
  OAI21_X1 U21446 ( .B1(n18391), .B2(n19088), .A(n18390), .ZN(n18392) );
  AOI221_X1 U21447 ( .B1(n19060), .B2(n18392), .C1(n18476), .C2(n18392), .A(
        n18586), .ZN(n18393) );
  OAI211_X1 U21448 ( .C1(n18566), .C2(n18395), .A(n18394), .B(n18393), .ZN(
        n18406) );
  OAI221_X1 U21449 ( .B1(n18406), .B2(n18502), .C1(n18406), .C2(n18396), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18404) );
  INV_X1 U21450 ( .A(n18397), .ZN(n18398) );
  OAI22_X1 U21451 ( .A1(n18500), .A2(n19088), .B1(n18564), .B2(n18501), .ZN(
        n18559) );
  NAND2_X1 U21452 ( .A1(n18503), .A2(n18559), .ZN(n18526) );
  NOR2_X1 U21453 ( .A1(n18398), .A2(n18526), .ZN(n18422) );
  OAI21_X1 U21454 ( .B1(n18422), .B2(n18399), .A(n18595), .ZN(n18499) );
  NOR2_X1 U21455 ( .A1(n18400), .A2(n18499), .ZN(n18418) );
  AOI22_X1 U21456 ( .A1(n18496), .A2(n18402), .B1(n18418), .B2(n18401), .ZN(
        n18403) );
  OAI221_X1 U21457 ( .B1(n9732), .B2(n18404), .C1(n18481), .C2(n19169), .A(
        n18403), .ZN(P3_U2844) );
  INV_X1 U21458 ( .A(n18418), .ZN(n18409) );
  AOI22_X1 U21459 ( .A1(n9732), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18496), 
        .B2(n18405), .ZN(n18408) );
  NAND3_X1 U21460 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18481), .A3(
        n18406), .ZN(n18407) );
  OAI211_X1 U21461 ( .C1(n18410), .C2(n18409), .A(n18408), .B(n18407), .ZN(
        P3_U2845) );
  INV_X1 U21462 ( .A(n18488), .ZN(n18479) );
  AOI22_X1 U21463 ( .A1(n19060), .A2(n18412), .B1(n19080), .B2(n18411), .ZN(
        n18470) );
  OAI21_X1 U21464 ( .B1(n18423), .B2(n18462), .A(n18413), .ZN(n18414) );
  OAI211_X1 U21465 ( .C1(n18415), .C2(n18479), .A(n18470), .B(n18414), .ZN(
        n18425) );
  OAI221_X1 U21466 ( .B1(n18416), .B2(n18505), .C1(n18416), .C2(n18425), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18421) );
  AOI22_X1 U21467 ( .A1(n18419), .A2(n18496), .B1(n18418), .B2(n18417), .ZN(
        n18420) );
  OAI221_X1 U21468 ( .B1(n9732), .B2(n18421), .C1(n18481), .C2(n19165), .A(
        n18420), .ZN(P3_U2846) );
  NAND2_X1 U21469 ( .A1(n9770), .A2(n18422), .ZN(n18440) );
  OAI21_X1 U21470 ( .B1(n18441), .B2(n18440), .A(n18423), .ZN(n18424) );
  AOI22_X1 U21471 ( .A1(n18427), .A2(n18426), .B1(n18425), .B2(n18424), .ZN(
        n18435) );
  AOI22_X1 U21472 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18588), .B1(
        n9732), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18434) );
  OAI211_X1 U21473 ( .C1(n18429), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18428), .B(n18598), .ZN(n18430) );
  INV_X1 U21474 ( .A(n18430), .ZN(n18431) );
  AOI21_X1 U21475 ( .B1(n18432), .B2(n18496), .A(n18431), .ZN(n18433) );
  OAI211_X1 U21476 ( .C1(n18435), .C2(n18586), .A(n18434), .B(n18433), .ZN(
        P3_U2847) );
  NAND2_X1 U21477 ( .A1(n18436), .A2(n18471), .ZN(n18463) );
  NAND2_X1 U21478 ( .A1(n18462), .A2(n18463), .ZN(n18455) );
  OAI211_X1 U21479 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18587), .A(
        n18470), .B(n18455), .ZN(n18437) );
  AOI211_X1 U21480 ( .C1(n18438), .C2(n18488), .A(n18441), .B(n18437), .ZN(
        n18439) );
  AOI211_X1 U21481 ( .C1(n18441), .C2(n18440), .A(n18439), .B(n18586), .ZN(
        n18442) );
  AOI211_X1 U21482 ( .C1(n18588), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18443), .B(n18442), .ZN(n18447) );
  AOI22_X1 U21483 ( .A1(n18598), .A2(n18445), .B1(n18496), .B2(n18444), .ZN(
        n18446) );
  OAI211_X1 U21484 ( .C1(n18449), .C2(n18448), .A(n18447), .B(n18446), .ZN(
        P3_U2848) );
  AOI22_X1 U21485 ( .A1(n9732), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18496), 
        .B2(n18450), .ZN(n18458) );
  AOI22_X1 U21486 ( .A1(n19058), .A2(n18453), .B1(n18452), .B2(n18451), .ZN(
        n18454) );
  OAI211_X1 U21487 ( .C1(n18480), .C2(n18479), .A(n18470), .B(n18454), .ZN(
        n18461) );
  OAI211_X1 U21488 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18479), .A(
        n18595), .B(n18455), .ZN(n18456) );
  OAI211_X1 U21489 ( .C1(n18461), .C2(n18456), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18481), .ZN(n18457) );
  OAI211_X1 U21490 ( .C1(n18459), .C2(n18499), .A(n18458), .B(n18457), .ZN(
        P3_U2849) );
  AOI211_X1 U21491 ( .C1(n18463), .C2(n18462), .A(n18461), .B(n18460), .ZN(
        n18468) );
  INV_X1 U21492 ( .A(n18499), .ZN(n18487) );
  AOI22_X1 U21493 ( .A1(n18480), .A2(n18487), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18595), .ZN(n18467) );
  AOI22_X1 U21494 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18588), .B1(
        n18496), .B2(n18464), .ZN(n18466) );
  OAI211_X1 U21495 ( .C1(n18468), .C2(n18467), .A(n18466), .B(n18465), .ZN(
        P3_U2850) );
  AOI22_X1 U21496 ( .A1(n9732), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18487), 
        .B2(n18469), .ZN(n18484) );
  OAI211_X1 U21497 ( .C1(n19064), .C2(n18471), .A(n18595), .B(n18470), .ZN(
        n18472) );
  AOI21_X1 U21498 ( .B1(n19058), .B2(n18473), .A(n18472), .ZN(n18474) );
  OAI21_X1 U21499 ( .B1(n18475), .B2(n18508), .A(n18474), .ZN(n18494) );
  AOI21_X1 U21500 ( .B1(n18477), .B2(n18476), .A(n18494), .ZN(n18478) );
  OAI21_X1 U21501 ( .B1(n19064), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18478), .ZN(n18489) );
  OAI22_X1 U21502 ( .A1(n19064), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18480), .B2(n18479), .ZN(n18482) );
  OAI211_X1 U21503 ( .C1(n18489), .C2(n18482), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18481), .ZN(n18483) );
  OAI211_X1 U21504 ( .C1(n18486), .C2(n18485), .A(n18484), .B(n18483), .ZN(
        P3_U2851) );
  NAND2_X1 U21505 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18487), .ZN(
        n18493) );
  OAI221_X1 U21506 ( .B1(n18489), .B2(n12119), .C1(n18489), .C2(n18488), .A(
        n18481), .ZN(n18492) );
  AOI22_X1 U21507 ( .A1(n9732), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18496), 
        .B2(n18490), .ZN(n18491) );
  OAI221_X1 U21508 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18493), 
        .C1(n12120), .C2(n18492), .A(n18491), .ZN(P3_U2852) );
  NAND2_X1 U21509 ( .A1(n18481), .A2(n18494), .ZN(n18498) );
  AOI22_X1 U21510 ( .A1(n9732), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18496), .B2(
        n18495), .ZN(n18497) );
  OAI221_X1 U21511 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18499), .C1(
        n12119), .C2(n18498), .A(n18497), .ZN(P3_U2853) );
  NOR2_X1 U21512 ( .A1(n10171), .A2(n18526), .ZN(n18518) );
  AND2_X1 U21513 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18518), .ZN(
        n18507) );
  NAND2_X1 U21514 ( .A1(n19060), .A2(n18500), .ZN(n18571) );
  AOI21_X1 U21515 ( .B1(n18502), .B2(n18501), .A(n18568), .ZN(n18542) );
  OAI211_X1 U21516 ( .C1(n9743), .C2(n18503), .A(n18571), .B(n18542), .ZN(
        n18528) );
  AOI211_X1 U21517 ( .C1(n18505), .C2(n10171), .A(n18504), .B(n18528), .ZN(
        n18521) );
  NOR2_X1 U21518 ( .A1(n9743), .A2(n18521), .ZN(n18506) );
  MUX2_X1 U21519 ( .A(n18507), .B(n18506), .S(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(n18512) );
  OAI22_X1 U21520 ( .A1(n18574), .A2(n18510), .B1(n18509), .B2(n18508), .ZN(
        n18511) );
  AOI211_X1 U21521 ( .C1(n18514), .C2(n18513), .A(n18512), .B(n18511), .ZN(
        n18516) );
  AOI22_X1 U21522 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18588), .B1(
        n9732), .B2(P3_REIP_REG_8__SCAN_IN), .ZN(n18515) );
  OAI21_X1 U21523 ( .B1(n18516), .B2(n18586), .A(n18515), .ZN(P3_U2854) );
  INV_X1 U21524 ( .A(n18517), .ZN(n18525) );
  OAI21_X1 U21525 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18518), .A(
        n18595), .ZN(n18520) );
  OAI22_X1 U21526 ( .A1(n18521), .A2(n18520), .B1(n18593), .B2(n18519), .ZN(
        n18522) );
  AOI211_X1 U21527 ( .C1(n18588), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18523), .B(n18522), .ZN(n18524) );
  OAI21_X1 U21528 ( .B1(n18602), .B2(n18525), .A(n18524), .ZN(P3_U2855) );
  NOR3_X1 U21529 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18586), .A3(
        n18526), .ZN(n18527) );
  AOI21_X1 U21530 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n9732), .A(n18527), .ZN(
        n18532) );
  AOI21_X1 U21531 ( .B1(n18528), .B2(n18595), .A(n18588), .ZN(n18529) );
  INV_X1 U21532 ( .A(n18529), .ZN(n18534) );
  AOI22_X1 U21533 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18534), .B1(
        n18583), .B2(n18530), .ZN(n18531) );
  OAI211_X1 U21534 ( .C1(n18593), .C2(n18533), .A(n18532), .B(n18531), .ZN(
        P3_U2856) );
  NAND3_X1 U21535 ( .A1(n18595), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18559), .ZN(n18550) );
  NOR2_X1 U21536 ( .A1(n18544), .A2(n18550), .ZN(n18535) );
  MUX2_X1 U21537 ( .A(n18535), .B(n18534), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18536) );
  AOI21_X1 U21538 ( .B1(n18583), .B2(n18537), .A(n18536), .ZN(n18539) );
  NAND2_X1 U21539 ( .A1(n9732), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18538) );
  OAI211_X1 U21540 ( .C1(n18540), .C2(n18593), .A(n18539), .B(n18538), .ZN(
        P3_U2857) );
  AOI22_X1 U21541 ( .A1(n9732), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18583), .B2(
        n18541), .ZN(n18549) );
  AND2_X1 U21542 ( .A1(n18571), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18543) );
  AOI21_X1 U21543 ( .B1(n18543), .B2(n18542), .A(n18586), .ZN(n18560) );
  NOR2_X1 U21544 ( .A1(n18588), .A2(n18560), .ZN(n18557) );
  NOR2_X1 U21545 ( .A1(n18557), .A2(n18544), .ZN(n18546) );
  AOI22_X1 U21546 ( .A1(n18547), .A2(n18598), .B1(n18546), .B2(n18545), .ZN(
        n18548) );
  OAI211_X1 U21547 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18550), .A(
        n18549), .B(n18548), .ZN(P3_U2858) );
  INV_X1 U21548 ( .A(n18551), .ZN(n18563) );
  OAI21_X1 U21549 ( .B1(n18554), .B2(n18553), .A(n18552), .ZN(n18555) );
  OAI22_X1 U21550 ( .A1(n18557), .A2(n18556), .B1(n18593), .B2(n18555), .ZN(
        n18558) );
  AOI21_X1 U21551 ( .B1(n18560), .B2(n18559), .A(n18558), .ZN(n18562) );
  OAI211_X1 U21552 ( .C1(n18563), .C2(n18602), .A(n18562), .B(n18561), .ZN(
        P3_U2859) );
  OR2_X1 U21553 ( .A1(n21317), .A2(n18564), .ZN(n18570) );
  NAND2_X1 U21554 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18565) );
  OAI22_X1 U21555 ( .A1(n18566), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19088), .B2(n18565), .ZN(n18567) );
  NOR2_X1 U21556 ( .A1(n18568), .A2(n18567), .ZN(n18569) );
  MUX2_X1 U21557 ( .A(n18570), .B(n18569), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18572) );
  OAI211_X1 U21558 ( .C1(n18574), .C2(n18573), .A(n18572), .B(n18571), .ZN(
        n18576) );
  AOI22_X1 U21559 ( .A1(n18595), .A2(n18576), .B1(n18583), .B2(n18575), .ZN(
        n18579) );
  INV_X1 U21560 ( .A(n18577), .ZN(n18578) );
  OAI211_X1 U21561 ( .C1(n18581), .C2(n18580), .A(n18579), .B(n18578), .ZN(
        P3_U2860) );
  AOI22_X1 U21562 ( .A1(n9732), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18583), .B2(
        n18582), .ZN(n18592) );
  AOI211_X1 U21563 ( .C1(n9780), .C2(n19237), .A(n9743), .B(n18586), .ZN(
        n18585) );
  INV_X1 U21564 ( .A(n18585), .ZN(n18590) );
  NOR3_X1 U21565 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18587), .A3(
        n18586), .ZN(n18597) );
  NOR2_X1 U21566 ( .A1(n18588), .A2(n18597), .ZN(n18589) );
  MUX2_X1 U21567 ( .A(n18590), .B(n18589), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n18591) );
  OAI211_X1 U21568 ( .C1(n18594), .C2(n18593), .A(n18592), .B(n18591), .ZN(
        P3_U2861) );
  AOI211_X1 U21569 ( .C1(n9780), .C2(n18595), .A(n9732), .B(n19237), .ZN(
        n18596) );
  AOI211_X1 U21570 ( .C1(n18598), .C2(n18601), .A(n18597), .B(n18596), .ZN(
        n18600) );
  NAND2_X1 U21571 ( .A1(n9732), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18599) );
  OAI211_X1 U21572 ( .C1(n18602), .C2(n18601), .A(n18600), .B(n18599), .ZN(
        P3_U2862) );
  OAI211_X1 U21573 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18603), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n19111)
         );
  OAI21_X1 U21574 ( .B1(n18606), .B2(n18604), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18605) );
  OAI221_X1 U21575 ( .B1(n18606), .B2(n19111), .C1(n18606), .C2(n18649), .A(
        n18605), .ZN(P3_U2863) );
  INV_X1 U21576 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19095) );
  NOR2_X1 U21577 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18613), .ZN(
        n18780) );
  INV_X1 U21578 ( .A(n18780), .ZN(n18756) );
  NAND2_X1 U21579 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18613), .ZN(
        n18852) );
  INV_X1 U21580 ( .A(n18852), .ZN(n18877) );
  NAND2_X1 U21581 ( .A1(n18964), .A2(n18877), .ZN(n18902) );
  AND2_X1 U21582 ( .A1(n18756), .A2(n18902), .ZN(n18608) );
  OAI22_X1 U21583 ( .A1(n18609), .A2(n19095), .B1(n18608), .B2(n18607), .ZN(
        P3_U2866) );
  NOR2_X1 U21584 ( .A1(n18611), .A2(n18610), .ZN(P3_U2867) );
  NAND2_X1 U21585 ( .A1(n18998), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18909) );
  NAND2_X1 U21586 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18614) );
  NAND2_X1 U21587 ( .A1(n19066), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18853) );
  NOR2_X1 U21588 ( .A1(n18614), .A2(n18853), .ZN(n18662) );
  INV_X1 U21589 ( .A(n18662), .ZN(n18992) );
  NOR2_X1 U21590 ( .A1(n18614), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18997) );
  INV_X1 U21591 ( .A(n18997), .ZN(n18931) );
  NOR2_X2 U21592 ( .A1(n19066), .A2(n18931), .ZN(n19036) );
  NOR2_X2 U21593 ( .A1(n15948), .A2(n18639), .ZN(n18999) );
  NOR2_X2 U21594 ( .A1(n18690), .A2(n18612), .ZN(n18993) );
  NOR2_X1 U21595 ( .A1(n19095), .A2(n18779), .ZN(n18996) );
  NAND2_X1 U21596 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18996), .ZN(
        n19041) );
  NOR2_X1 U21597 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19070) );
  INV_X1 U21598 ( .A(n19070), .ZN(n18803) );
  NAND2_X1 U21599 ( .A1(n18613), .A2(n19095), .ZN(n18689) );
  NOR2_X2 U21600 ( .A1(n18803), .A2(n18689), .ZN(n18702) );
  INV_X1 U21601 ( .A(n18702), .ZN(n18711) );
  NAND2_X1 U21602 ( .A1(n19041), .A2(n18711), .ZN(n18669) );
  AND2_X1 U21603 ( .A1(n19113), .A2(n18669), .ZN(n18643) );
  AOI22_X1 U21604 ( .A1(n19036), .A2(n18999), .B1(n18993), .B2(n18643), .ZN(
        n18619) );
  NAND2_X1 U21605 ( .A1(n19067), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18829) );
  AND2_X1 U21606 ( .A1(n18853), .A2(n18829), .ZN(n18903) );
  NOR2_X1 U21607 ( .A1(n18903), .A2(n18614), .ZN(n18965) );
  AOI21_X1 U21608 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18690), .ZN(n18962) );
  AOI22_X1 U21609 ( .A1(n18998), .A2(n18965), .B1(n18962), .B2(n18669), .ZN(
        n18646) );
  NAND2_X1 U21610 ( .A1(n18616), .A2(n18615), .ZN(n18644) );
  NOR2_X1 U21611 ( .A1(n18617), .A2(n18644), .ZN(n18906) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18646), .B1(
        n18702), .B2(n18906), .ZN(n18618) );
  OAI211_X1 U21613 ( .C1(n18909), .C2(n18992), .A(n18619), .B(n18618), .ZN(
        P3_U2868) );
  INV_X1 U21614 ( .A(n19036), .ZN(n19052) );
  NAND2_X1 U21615 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18998), .ZN(n18939) );
  NOR2_X2 U21616 ( .A1(n18639), .A2(n15998), .ZN(n19005) );
  NOR2_X2 U21617 ( .A1(n18690), .A2(n18620), .ZN(n19003) );
  AOI22_X1 U21618 ( .A1(n18662), .A2(n19005), .B1(n18643), .B2(n19003), .ZN(
        n18623) );
  NOR2_X1 U21619 ( .A1(n18621), .A2(n18644), .ZN(n18936) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18646), .B1(
        n18702), .B2(n18936), .ZN(n18622) );
  OAI211_X1 U21621 ( .C1(n19052), .C2(n18939), .A(n18623), .B(n18622), .ZN(
        P3_U2869) );
  NAND2_X1 U21622 ( .A1(n18998), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19014) );
  AND2_X1 U21623 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18998), .ZN(n19009) );
  NOR2_X2 U21624 ( .A1(n18690), .A2(n18624), .ZN(n19010) );
  AOI22_X1 U21625 ( .A1(n19036), .A2(n19009), .B1(n18643), .B2(n19010), .ZN(
        n18627) );
  NOR2_X1 U21626 ( .A1(n18625), .A2(n18644), .ZN(n19011) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18646), .B1(
        n18702), .B2(n19011), .ZN(n18626) );
  OAI211_X1 U21628 ( .C1(n18992), .C2(n19014), .A(n18627), .B(n18626), .ZN(
        P3_U2870) );
  NAND2_X1 U21629 ( .A1(n18998), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19020) );
  NAND2_X1 U21630 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18998), .ZN(n18916) );
  INV_X1 U21631 ( .A(n18916), .ZN(n19016) );
  NOR2_X2 U21632 ( .A1(n18690), .A2(n18628), .ZN(n19015) );
  AOI22_X1 U21633 ( .A1(n19036), .A2(n19016), .B1(n18643), .B2(n19015), .ZN(
        n18631) );
  NOR2_X2 U21634 ( .A1(n18629), .A2(n18644), .ZN(n19017) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18646), .B1(
        n18702), .B2(n19017), .ZN(n18630) );
  OAI211_X1 U21636 ( .C1(n18992), .C2(n19020), .A(n18631), .B(n18630), .ZN(
        P3_U2871) );
  NAND2_X1 U21637 ( .A1(n18998), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18891) );
  NOR2_X1 U21638 ( .A1(n15926), .A2(n18639), .ZN(n19023) );
  NOR2_X2 U21639 ( .A1(n18690), .A2(n21290), .ZN(n19021) );
  AOI22_X1 U21640 ( .A1(n19036), .A2(n19023), .B1(n18643), .B2(n19021), .ZN(
        n18634) );
  NOR2_X2 U21641 ( .A1(n18632), .A2(n18644), .ZN(n18944) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18646), .B1(
        n18702), .B2(n18944), .ZN(n18633) );
  OAI211_X1 U21643 ( .C1(n18992), .C2(n18891), .A(n18634), .B(n18633), .ZN(
        P3_U2872) );
  NAND2_X1 U21644 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18998), .ZN(n18951) );
  NOR2_X1 U21645 ( .A1(n18639), .A2(n18635), .ZN(n19028) );
  NOR2_X2 U21646 ( .A1(n18690), .A2(n13138), .ZN(n19027) );
  AOI22_X1 U21647 ( .A1(n18662), .A2(n19028), .B1(n18643), .B2(n19027), .ZN(
        n18638) );
  NOR2_X2 U21648 ( .A1(n18636), .A2(n18644), .ZN(n18948) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18646), .B1(
        n18702), .B2(n18948), .ZN(n18637) );
  OAI211_X1 U21650 ( .C1(n19052), .C2(n18951), .A(n18638), .B(n18637), .ZN(
        P3_U2873) );
  NAND2_X1 U21651 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18998), .ZN(n18925) );
  NOR2_X2 U21652 ( .A1(n12431), .A2(n18639), .ZN(n19037) );
  NOR2_X2 U21653 ( .A1(n12944), .A2(n18690), .ZN(n19034) );
  AOI22_X1 U21654 ( .A1(n19036), .A2(n19037), .B1(n18643), .B2(n19034), .ZN(
        n18642) );
  NOR2_X1 U21655 ( .A1(n18640), .A2(n18644), .ZN(n18922) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18646), .B1(
        n18702), .B2(n18922), .ZN(n18641) );
  OAI211_X1 U21657 ( .C1(n18992), .C2(n18925), .A(n18642), .B(n18641), .ZN(
        P3_U2874) );
  NAND2_X1 U21658 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18998), .ZN(n18960) );
  NAND2_X1 U21659 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18998), .ZN(n19051) );
  INV_X1 U21660 ( .A(n19051), .ZN(n18987) );
  NOR2_X2 U21661 ( .A1(n13056), .A2(n18690), .ZN(n19043) );
  AOI22_X1 U21662 ( .A1(n18662), .A2(n18987), .B1(n18643), .B2(n19043), .ZN(
        n18648) );
  NOR2_X2 U21663 ( .A1(n18645), .A2(n18644), .ZN(n19046) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18646), .B1(
        n18702), .B2(n19046), .ZN(n18647) );
  OAI211_X1 U21665 ( .C1(n19052), .C2(n18960), .A(n18648), .B(n18647), .ZN(
        P3_U2875) );
  NAND2_X1 U21666 ( .A1(n19067), .A2(n19113), .ZN(n18830) );
  NOR2_X1 U21667 ( .A1(n18689), .A2(n18830), .ZN(n18665) );
  AOI22_X1 U21668 ( .A1(n18662), .A2(n18999), .B1(n18993), .B2(n18665), .ZN(
        n18651) );
  INV_X1 U21669 ( .A(n18689), .ZN(n18691) );
  NAND2_X1 U21670 ( .A1(n18905), .A2(n18649), .ZN(n18831) );
  NOR2_X1 U21671 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18831), .ZN(
        n18734) );
  AOI22_X1 U21672 ( .A1(n18998), .A2(n18996), .B1(n18691), .B2(n18734), .ZN(
        n18666) );
  NOR2_X2 U21673 ( .A1(n18689), .A2(n18829), .ZN(n18730) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18666), .B1(
        n18906), .B2(n18730), .ZN(n18650) );
  OAI211_X1 U21675 ( .C1(n19041), .C2(n18909), .A(n18651), .B(n18650), .ZN(
        P3_U2876) );
  INV_X1 U21676 ( .A(n19041), .ZN(n19047) );
  AOI22_X1 U21677 ( .A1(n19047), .A2(n19005), .B1(n19003), .B2(n18665), .ZN(
        n18653) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18666), .B1(
        n18936), .B2(n18730), .ZN(n18652) );
  OAI211_X1 U21679 ( .C1(n18992), .C2(n18939), .A(n18653), .B(n18652), .ZN(
        P3_U2877) );
  AOI22_X1 U21680 ( .A1(n18662), .A2(n19009), .B1(n19010), .B2(n18665), .ZN(
        n18655) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18666), .B1(
        n19011), .B2(n18730), .ZN(n18654) );
  OAI211_X1 U21682 ( .C1(n19041), .C2(n19014), .A(n18655), .B(n18654), .ZN(
        P3_U2878) );
  INV_X1 U21683 ( .A(n19020), .ZN(n18974) );
  AOI22_X1 U21684 ( .A1(n19047), .A2(n18974), .B1(n19015), .B2(n18665), .ZN(
        n18657) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18666), .B1(
        n19017), .B2(n18730), .ZN(n18656) );
  OAI211_X1 U21686 ( .C1(n18992), .C2(n18916), .A(n18657), .B(n18656), .ZN(
        P3_U2879) );
  INV_X1 U21687 ( .A(n19023), .ZN(n18947) );
  INV_X1 U21688 ( .A(n18891), .ZN(n19022) );
  AOI22_X1 U21689 ( .A1(n19047), .A2(n19022), .B1(n19021), .B2(n18665), .ZN(
        n18659) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18666), .B1(
        n18944), .B2(n18730), .ZN(n18658) );
  OAI211_X1 U21691 ( .C1(n18992), .C2(n18947), .A(n18659), .B(n18658), .ZN(
        P3_U2880) );
  INV_X1 U21692 ( .A(n19028), .ZN(n18894) );
  INV_X1 U21693 ( .A(n18951), .ZN(n19030) );
  AOI22_X1 U21694 ( .A1(n18662), .A2(n19030), .B1(n19027), .B2(n18665), .ZN(
        n18661) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18666), .B1(
        n18948), .B2(n18730), .ZN(n18660) );
  OAI211_X1 U21696 ( .C1(n19041), .C2(n18894), .A(n18661), .B(n18660), .ZN(
        P3_U2881) );
  AOI22_X1 U21697 ( .A1(n18662), .A2(n19037), .B1(n19034), .B2(n18665), .ZN(
        n18664) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18666), .B1(
        n18922), .B2(n18730), .ZN(n18663) );
  OAI211_X1 U21699 ( .C1(n19041), .C2(n18925), .A(n18664), .B(n18663), .ZN(
        P3_U2882) );
  AOI22_X1 U21700 ( .A1(n19047), .A2(n18987), .B1(n19043), .B2(n18665), .ZN(
        n18668) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18666), .B1(
        n19046), .B2(n18730), .ZN(n18667) );
  OAI211_X1 U21702 ( .C1(n18992), .C2(n18960), .A(n18668), .B(n18667), .ZN(
        P3_U2883) );
  INV_X1 U21703 ( .A(n18906), .ZN(n19002) );
  NOR2_X2 U21704 ( .A1(n18689), .A2(n18853), .ZN(n18748) );
  INV_X1 U21705 ( .A(n18748), .ZN(n18755) );
  INV_X1 U21706 ( .A(n18909), .ZN(n18994) );
  NOR2_X1 U21707 ( .A1(n18730), .A2(n18748), .ZN(n18712) );
  NOR2_X1 U21708 ( .A1(n18932), .A2(n18712), .ZN(n18685) );
  AOI22_X1 U21709 ( .A1(n18702), .A2(n18994), .B1(n18993), .B2(n18685), .ZN(
        n18672) );
  INV_X1 U21710 ( .A(n18712), .ZN(n18670) );
  OAI221_X1 U21711 ( .B1(n18670), .B2(n18964), .C1(n18670), .C2(n18669), .A(
        n18962), .ZN(n18686) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18686), .B1(
        n19047), .B2(n18999), .ZN(n18671) );
  OAI211_X1 U21713 ( .C1(n19002), .C2(n18755), .A(n18672), .B(n18671), .ZN(
        P3_U2884) );
  INV_X1 U21714 ( .A(n18936), .ZN(n19008) );
  INV_X1 U21715 ( .A(n18939), .ZN(n19004) );
  AOI22_X1 U21716 ( .A1(n19047), .A2(n19004), .B1(n19003), .B2(n18685), .ZN(
        n18674) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18686), .B1(
        n18702), .B2(n19005), .ZN(n18673) );
  OAI211_X1 U21718 ( .C1(n19008), .C2(n18755), .A(n18674), .B(n18673), .ZN(
        P3_U2885) );
  AOI22_X1 U21719 ( .A1(n19047), .A2(n19009), .B1(n19010), .B2(n18685), .ZN(
        n18676) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18686), .B1(
        n19011), .B2(n18748), .ZN(n18675) );
  OAI211_X1 U21721 ( .C1(n18711), .C2(n19014), .A(n18676), .B(n18675), .ZN(
        P3_U2886) );
  AOI22_X1 U21722 ( .A1(n19047), .A2(n19016), .B1(n19015), .B2(n18685), .ZN(
        n18678) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18686), .B1(
        n19017), .B2(n18748), .ZN(n18677) );
  OAI211_X1 U21724 ( .C1(n18711), .C2(n19020), .A(n18678), .B(n18677), .ZN(
        P3_U2887) );
  AOI22_X1 U21725 ( .A1(n19047), .A2(n19023), .B1(n19021), .B2(n18685), .ZN(
        n18680) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18686), .B1(
        n18944), .B2(n18748), .ZN(n18679) );
  OAI211_X1 U21727 ( .C1(n18711), .C2(n18891), .A(n18680), .B(n18679), .ZN(
        P3_U2888) );
  AOI22_X1 U21728 ( .A1(n19047), .A2(n19030), .B1(n19027), .B2(n18685), .ZN(
        n18682) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18686), .B1(
        n18948), .B2(n18748), .ZN(n18681) );
  OAI211_X1 U21730 ( .C1(n18711), .C2(n18894), .A(n18682), .B(n18681), .ZN(
        P3_U2889) );
  INV_X1 U21731 ( .A(n19037), .ZN(n18822) );
  INV_X1 U21732 ( .A(n18925), .ZN(n19035) );
  AOI22_X1 U21733 ( .A1(n18702), .A2(n19035), .B1(n19034), .B2(n18685), .ZN(
        n18684) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18686), .B1(
        n18922), .B2(n18748), .ZN(n18683) );
  OAI211_X1 U21735 ( .C1(n19041), .C2(n18822), .A(n18684), .B(n18683), .ZN(
        P3_U2890) );
  INV_X1 U21736 ( .A(n18960), .ZN(n19045) );
  AOI22_X1 U21737 ( .A1(n19047), .A2(n19045), .B1(n19043), .B2(n18685), .ZN(
        n18688) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18686), .B1(
        n19046), .B2(n18748), .ZN(n18687) );
  OAI211_X1 U21739 ( .C1(n18711), .C2(n19051), .A(n18688), .B(n18687), .ZN(
        P3_U2891) );
  NOR2_X1 U21740 ( .A1(n19067), .A2(n18689), .ZN(n18735) );
  NAND2_X1 U21741 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18735), .ZN(
        n18778) );
  INV_X1 U21742 ( .A(n18778), .ZN(n18771) );
  INV_X1 U21743 ( .A(n18964), .ZN(n18854) );
  AOI21_X1 U21744 ( .B1(n19067), .B2(n18854), .A(n18690), .ZN(n18781) );
  OAI211_X1 U21745 ( .C1(n18771), .C2(n19212), .A(n18691), .B(n18781), .ZN(
        n18708) );
  AND2_X1 U21746 ( .A1(n19113), .A2(n18735), .ZN(n18707) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18708), .B1(
        n18993), .B2(n18707), .ZN(n18693) );
  AOI22_X1 U21748 ( .A1(n18702), .A2(n18999), .B1(n18994), .B2(n18730), .ZN(
        n18692) );
  OAI211_X1 U21749 ( .C1(n19002), .C2(n18778), .A(n18693), .B(n18692), .ZN(
        P3_U2892) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18708), .B1(
        n19003), .B2(n18707), .ZN(n18695) );
  AOI22_X1 U21751 ( .A1(n18936), .A2(n18771), .B1(n19005), .B2(n18730), .ZN(
        n18694) );
  OAI211_X1 U21752 ( .C1(n18711), .C2(n18939), .A(n18695), .B(n18694), .ZN(
        P3_U2893) );
  INV_X1 U21753 ( .A(n18730), .ZN(n18726) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18708), .B1(
        n19010), .B2(n18707), .ZN(n18697) );
  AOI22_X1 U21755 ( .A1(n18702), .A2(n19009), .B1(n19011), .B2(n18771), .ZN(
        n18696) );
  OAI211_X1 U21756 ( .C1(n19014), .C2(n18726), .A(n18697), .B(n18696), .ZN(
        P3_U2894) );
  AOI22_X1 U21757 ( .A1(n18702), .A2(n19016), .B1(n19015), .B2(n18707), .ZN(
        n18699) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18708), .B1(
        n19017), .B2(n18771), .ZN(n18698) );
  OAI211_X1 U21759 ( .C1(n19020), .C2(n18726), .A(n18699), .B(n18698), .ZN(
        P3_U2895) );
  AOI22_X1 U21760 ( .A1(n18702), .A2(n19023), .B1(n19021), .B2(n18707), .ZN(
        n18701) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18708), .B1(
        n18944), .B2(n18771), .ZN(n18700) );
  OAI211_X1 U21762 ( .C1(n18891), .C2(n18726), .A(n18701), .B(n18700), .ZN(
        P3_U2896) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18708), .B1(
        n19027), .B2(n18707), .ZN(n18704) );
  AOI22_X1 U21764 ( .A1(n18702), .A2(n19030), .B1(n18948), .B2(n18771), .ZN(
        n18703) );
  OAI211_X1 U21765 ( .C1(n18894), .C2(n18726), .A(n18704), .B(n18703), .ZN(
        P3_U2897) );
  AOI22_X1 U21766 ( .A1(n19035), .A2(n18730), .B1(n19034), .B2(n18707), .ZN(
        n18706) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18708), .B1(
        n18922), .B2(n18771), .ZN(n18705) );
  OAI211_X1 U21768 ( .C1(n18711), .C2(n18822), .A(n18706), .B(n18705), .ZN(
        P3_U2898) );
  AOI22_X1 U21769 ( .A1(n18987), .A2(n18730), .B1(n19043), .B2(n18707), .ZN(
        n18710) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18708), .B1(
        n19046), .B2(n18771), .ZN(n18709) );
  OAI211_X1 U21771 ( .C1(n18711), .C2(n18960), .A(n18710), .B(n18709), .ZN(
        P3_U2899) );
  NAND2_X1 U21772 ( .A1(n19070), .A2(n18780), .ZN(n18802) );
  INV_X1 U21773 ( .A(n18802), .ZN(n18795) );
  NOR2_X1 U21774 ( .A1(n18771), .A2(n18795), .ZN(n18757) );
  NOR2_X1 U21775 ( .A1(n18932), .A2(n18757), .ZN(n18729) );
  AOI22_X1 U21776 ( .A1(n18994), .A2(n18748), .B1(n18993), .B2(n18729), .ZN(
        n18715) );
  OAI21_X1 U21777 ( .B1(n18712), .B2(n18854), .A(n18757), .ZN(n18713) );
  OAI211_X1 U21778 ( .C1(n18795), .C2(n19212), .A(n18905), .B(n18713), .ZN(
        n18731) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18731), .B1(
        n18999), .B2(n18730), .ZN(n18714) );
  OAI211_X1 U21780 ( .C1(n19002), .C2(n18802), .A(n18715), .B(n18714), .ZN(
        P3_U2900) );
  AOI22_X1 U21781 ( .A1(n19005), .A2(n18748), .B1(n19003), .B2(n18729), .ZN(
        n18717) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18731), .B1(
        n18936), .B2(n18795), .ZN(n18716) );
  OAI211_X1 U21783 ( .C1(n18939), .C2(n18726), .A(n18717), .B(n18716), .ZN(
        P3_U2901) );
  AOI22_X1 U21784 ( .A1(n19010), .A2(n18729), .B1(n19009), .B2(n18730), .ZN(
        n18719) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18731), .B1(
        n19011), .B2(n18795), .ZN(n18718) );
  OAI211_X1 U21786 ( .C1(n19014), .C2(n18755), .A(n18719), .B(n18718), .ZN(
        P3_U2902) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18731), .B1(
        n19015), .B2(n18729), .ZN(n18721) );
  AOI22_X1 U21788 ( .A1(n19017), .A2(n18795), .B1(n19016), .B2(n18730), .ZN(
        n18720) );
  OAI211_X1 U21789 ( .C1(n19020), .C2(n18755), .A(n18721), .B(n18720), .ZN(
        P3_U2903) );
  AOI22_X1 U21790 ( .A1(n19021), .A2(n18729), .B1(n19023), .B2(n18730), .ZN(
        n18723) );
  AOI22_X1 U21791 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18731), .B1(
        n18944), .B2(n18795), .ZN(n18722) );
  OAI211_X1 U21792 ( .C1(n18891), .C2(n18755), .A(n18723), .B(n18722), .ZN(
        P3_U2904) );
  AOI22_X1 U21793 ( .A1(n19028), .A2(n18748), .B1(n19027), .B2(n18729), .ZN(
        n18725) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18731), .B1(
        n18948), .B2(n18795), .ZN(n18724) );
  OAI211_X1 U21795 ( .C1(n18951), .C2(n18726), .A(n18725), .B(n18724), .ZN(
        P3_U2905) );
  AOI22_X1 U21796 ( .A1(n19037), .A2(n18730), .B1(n19034), .B2(n18729), .ZN(
        n18728) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18731), .B1(
        n18922), .B2(n18795), .ZN(n18727) );
  OAI211_X1 U21798 ( .C1(n18925), .C2(n18755), .A(n18728), .B(n18727), .ZN(
        P3_U2906) );
  AOI22_X1 U21799 ( .A1(n19045), .A2(n18730), .B1(n19043), .B2(n18729), .ZN(
        n18733) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18731), .B1(
        n19046), .B2(n18795), .ZN(n18732) );
  OAI211_X1 U21801 ( .C1(n19051), .C2(n18755), .A(n18733), .B(n18732), .ZN(
        P3_U2907) );
  NOR2_X2 U21802 ( .A1(n18829), .A2(n18756), .ZN(n18824) );
  INV_X1 U21803 ( .A(n18824), .ZN(n18821) );
  NOR2_X1 U21804 ( .A1(n18830), .A2(n18756), .ZN(n18751) );
  AOI22_X1 U21805 ( .A1(n18994), .A2(n18771), .B1(n18993), .B2(n18751), .ZN(
        n18737) );
  AOI22_X1 U21806 ( .A1(n18998), .A2(n18735), .B1(n18734), .B2(n18780), .ZN(
        n18752) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18752), .B1(
        n18999), .B2(n18748), .ZN(n18736) );
  OAI211_X1 U21808 ( .C1(n19002), .C2(n18821), .A(n18737), .B(n18736), .ZN(
        P3_U2908) );
  AOI22_X1 U21809 ( .A1(n19004), .A2(n18748), .B1(n19003), .B2(n18751), .ZN(
        n18739) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18752), .B1(
        n19005), .B2(n18771), .ZN(n18738) );
  OAI211_X1 U21811 ( .C1(n19008), .C2(n18821), .A(n18739), .B(n18738), .ZN(
        P3_U2909) );
  INV_X1 U21812 ( .A(n19011), .ZN(n18973) );
  INV_X1 U21813 ( .A(n19014), .ZN(n18970) );
  AOI22_X1 U21814 ( .A1(n18970), .A2(n18771), .B1(n19010), .B2(n18751), .ZN(
        n18741) );
  AOI22_X1 U21815 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18752), .B1(
        n19009), .B2(n18748), .ZN(n18740) );
  OAI211_X1 U21816 ( .C1(n18973), .C2(n18821), .A(n18741), .B(n18740), .ZN(
        P3_U2910) );
  AOI22_X1 U21817 ( .A1(n18974), .A2(n18771), .B1(n19015), .B2(n18751), .ZN(
        n18743) );
  AOI22_X1 U21818 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18752), .B1(
        n19017), .B2(n18824), .ZN(n18742) );
  OAI211_X1 U21819 ( .C1(n18916), .C2(n18755), .A(n18743), .B(n18742), .ZN(
        P3_U2911) );
  AOI22_X1 U21820 ( .A1(n19022), .A2(n18771), .B1(n19021), .B2(n18751), .ZN(
        n18745) );
  AOI22_X1 U21821 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18752), .B1(
        n18944), .B2(n18824), .ZN(n18744) );
  OAI211_X1 U21822 ( .C1(n18947), .C2(n18755), .A(n18745), .B(n18744), .ZN(
        P3_U2912) );
  AOI22_X1 U21823 ( .A1(n19028), .A2(n18771), .B1(n19027), .B2(n18751), .ZN(
        n18747) );
  AOI22_X1 U21824 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18752), .B1(
        n18948), .B2(n18824), .ZN(n18746) );
  OAI211_X1 U21825 ( .C1(n18951), .C2(n18755), .A(n18747), .B(n18746), .ZN(
        P3_U2913) );
  AOI22_X1 U21826 ( .A1(n19037), .A2(n18748), .B1(n19034), .B2(n18751), .ZN(
        n18750) );
  AOI22_X1 U21827 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18752), .B1(
        n18922), .B2(n18824), .ZN(n18749) );
  OAI211_X1 U21828 ( .C1(n18925), .C2(n18778), .A(n18750), .B(n18749), .ZN(
        P3_U2914) );
  AOI22_X1 U21829 ( .A1(n18987), .A2(n18771), .B1(n19043), .B2(n18751), .ZN(
        n18754) );
  AOI22_X1 U21830 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18752), .B1(
        n19046), .B2(n18824), .ZN(n18753) );
  OAI211_X1 U21831 ( .C1(n18960), .C2(n18755), .A(n18754), .B(n18753), .ZN(
        P3_U2915) );
  INV_X1 U21832 ( .A(n18843), .ZN(n18828) );
  NOR2_X1 U21833 ( .A1(n18824), .A2(n18843), .ZN(n18805) );
  NOR2_X1 U21834 ( .A1(n18932), .A2(n18805), .ZN(n18774) );
  AOI22_X1 U21835 ( .A1(n18999), .A2(n18771), .B1(n18993), .B2(n18774), .ZN(
        n18760) );
  OAI21_X1 U21836 ( .B1(n18757), .B2(n18854), .A(n18805), .ZN(n18758) );
  OAI211_X1 U21837 ( .C1(n18843), .C2(n19212), .A(n18905), .B(n18758), .ZN(
        n18775) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18775), .B1(
        n18994), .B2(n18795), .ZN(n18759) );
  OAI211_X1 U21839 ( .C1(n19002), .C2(n18828), .A(n18760), .B(n18759), .ZN(
        P3_U2916) );
  AOI22_X1 U21840 ( .A1(n19005), .A2(n18795), .B1(n19003), .B2(n18774), .ZN(
        n18762) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18775), .B1(
        n18936), .B2(n18843), .ZN(n18761) );
  OAI211_X1 U21842 ( .C1(n18939), .C2(n18778), .A(n18762), .B(n18761), .ZN(
        P3_U2917) );
  AOI22_X1 U21843 ( .A1(n19010), .A2(n18774), .B1(n19009), .B2(n18771), .ZN(
        n18764) );
  AOI22_X1 U21844 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18775), .B1(
        n19011), .B2(n18843), .ZN(n18763) );
  OAI211_X1 U21845 ( .C1(n19014), .C2(n18802), .A(n18764), .B(n18763), .ZN(
        P3_U2918) );
  AOI22_X1 U21846 ( .A1(n19016), .A2(n18771), .B1(n19015), .B2(n18774), .ZN(
        n18766) );
  AOI22_X1 U21847 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18775), .B1(
        n19017), .B2(n18843), .ZN(n18765) );
  OAI211_X1 U21848 ( .C1(n19020), .C2(n18802), .A(n18766), .B(n18765), .ZN(
        P3_U2919) );
  AOI22_X1 U21849 ( .A1(n19021), .A2(n18774), .B1(n19023), .B2(n18771), .ZN(
        n18768) );
  AOI22_X1 U21850 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18775), .B1(
        n18944), .B2(n18843), .ZN(n18767) );
  OAI211_X1 U21851 ( .C1(n18891), .C2(n18802), .A(n18768), .B(n18767), .ZN(
        P3_U2920) );
  AOI22_X1 U21852 ( .A1(n19030), .A2(n18771), .B1(n19027), .B2(n18774), .ZN(
        n18770) );
  AOI22_X1 U21853 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18775), .B1(
        n18948), .B2(n18843), .ZN(n18769) );
  OAI211_X1 U21854 ( .C1(n18894), .C2(n18802), .A(n18770), .B(n18769), .ZN(
        P3_U2921) );
  AOI22_X1 U21855 ( .A1(n19037), .A2(n18771), .B1(n19034), .B2(n18774), .ZN(
        n18773) );
  AOI22_X1 U21856 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18775), .B1(
        n18922), .B2(n18843), .ZN(n18772) );
  OAI211_X1 U21857 ( .C1(n18925), .C2(n18802), .A(n18773), .B(n18772), .ZN(
        P3_U2922) );
  AOI22_X1 U21858 ( .A1(n18987), .A2(n18795), .B1(n19043), .B2(n18774), .ZN(
        n18777) );
  AOI22_X1 U21859 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18775), .B1(
        n19046), .B2(n18843), .ZN(n18776) );
  OAI211_X1 U21860 ( .C1(n18960), .C2(n18778), .A(n18777), .B(n18776), .ZN(
        P3_U2923) );
  NOR2_X1 U21861 ( .A1(n18779), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18832) );
  INV_X1 U21862 ( .A(n18832), .ZN(n18782) );
  NOR2_X1 U21863 ( .A1(n19066), .A2(n18782), .ZN(n18867) );
  CLKBUF_X1 U21864 ( .A(n18867), .Z(n18873) );
  OAI211_X1 U21865 ( .C1(n18873), .C2(n19212), .A(n18781), .B(n18780), .ZN(
        n18799) );
  NOR2_X1 U21866 ( .A1(n18932), .A2(n18782), .ZN(n18798) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18799), .B1(
        n18993), .B2(n18798), .ZN(n18784) );
  AOI22_X1 U21868 ( .A1(n18906), .A2(n18873), .B1(n18999), .B2(n18795), .ZN(
        n18783) );
  OAI211_X1 U21869 ( .C1(n18909), .C2(n18821), .A(n18784), .B(n18783), .ZN(
        P3_U2924) );
  AOI22_X1 U21870 ( .A1(n19005), .A2(n18824), .B1(n19003), .B2(n18798), .ZN(
        n18786) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18799), .B1(
        n18936), .B2(n18867), .ZN(n18785) );
  OAI211_X1 U21872 ( .C1(n18939), .C2(n18802), .A(n18786), .B(n18785), .ZN(
        P3_U2925) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18799), .B1(
        n19010), .B2(n18798), .ZN(n18788) );
  AOI22_X1 U21874 ( .A1(n19011), .A2(n18873), .B1(n19009), .B2(n18795), .ZN(
        n18787) );
  OAI211_X1 U21875 ( .C1(n19014), .C2(n18821), .A(n18788), .B(n18787), .ZN(
        P3_U2926) );
  AOI22_X1 U21876 ( .A1(n18974), .A2(n18824), .B1(n19015), .B2(n18798), .ZN(
        n18790) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18799), .B1(
        n19017), .B2(n18867), .ZN(n18789) );
  OAI211_X1 U21878 ( .C1(n18916), .C2(n18802), .A(n18790), .B(n18789), .ZN(
        P3_U2927) );
  AOI22_X1 U21879 ( .A1(n19022), .A2(n18824), .B1(n19021), .B2(n18798), .ZN(
        n18792) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18799), .B1(
        n18944), .B2(n18873), .ZN(n18791) );
  OAI211_X1 U21881 ( .C1(n18947), .C2(n18802), .A(n18792), .B(n18791), .ZN(
        P3_U2928) );
  AOI22_X1 U21882 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18799), .B1(
        n19027), .B2(n18798), .ZN(n18794) );
  AOI22_X1 U21883 ( .A1(n18948), .A2(n18873), .B1(n19028), .B2(n18824), .ZN(
        n18793) );
  OAI211_X1 U21884 ( .C1(n18951), .C2(n18802), .A(n18794), .B(n18793), .ZN(
        P3_U2929) );
  AOI22_X1 U21885 ( .A1(n19037), .A2(n18795), .B1(n19034), .B2(n18798), .ZN(
        n18797) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18799), .B1(
        n18922), .B2(n18873), .ZN(n18796) );
  OAI211_X1 U21887 ( .C1(n18925), .C2(n18821), .A(n18797), .B(n18796), .ZN(
        P3_U2930) );
  AOI22_X1 U21888 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18799), .B1(
        n19043), .B2(n18798), .ZN(n18801) );
  AOI22_X1 U21889 ( .A1(n19046), .A2(n18873), .B1(n18987), .B2(n18824), .ZN(
        n18800) );
  OAI211_X1 U21890 ( .C1(n18960), .C2(n18802), .A(n18801), .B(n18800), .ZN(
        P3_U2931) );
  OR2_X1 U21891 ( .A1(n18803), .A2(n18852), .ZN(n18888) );
  INV_X1 U21892 ( .A(n18888), .ZN(n18898) );
  NOR2_X1 U21893 ( .A1(n18873), .A2(n18898), .ZN(n18855) );
  NOR2_X1 U21894 ( .A1(n18932), .A2(n18855), .ZN(n18823) );
  AOI22_X1 U21895 ( .A1(n18999), .A2(n18824), .B1(n18993), .B2(n18823), .ZN(
        n18808) );
  INV_X1 U21896 ( .A(n18962), .ZN(n18804) );
  AOI221_X1 U21897 ( .B1(n18855), .B2(n18854), .C1(n18855), .C2(n18805), .A(
        n18804), .ZN(n18806) );
  INV_X1 U21898 ( .A(n18806), .ZN(n18825) );
  AOI22_X1 U21899 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18825), .B1(
        n18906), .B2(n18898), .ZN(n18807) );
  OAI211_X1 U21900 ( .C1(n18909), .C2(n18828), .A(n18808), .B(n18807), .ZN(
        P3_U2932) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18825), .B1(
        n19003), .B2(n18823), .ZN(n18810) );
  AOI22_X1 U21902 ( .A1(n18936), .A2(n18898), .B1(n19005), .B2(n18843), .ZN(
        n18809) );
  OAI211_X1 U21903 ( .C1(n18939), .C2(n18821), .A(n18810), .B(n18809), .ZN(
        P3_U2933) );
  AOI22_X1 U21904 ( .A1(n19010), .A2(n18823), .B1(n19009), .B2(n18824), .ZN(
        n18812) );
  AOI22_X1 U21905 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18825), .B1(
        n19011), .B2(n18898), .ZN(n18811) );
  OAI211_X1 U21906 ( .C1(n19014), .C2(n18828), .A(n18812), .B(n18811), .ZN(
        P3_U2934) );
  AOI22_X1 U21907 ( .A1(n18974), .A2(n18843), .B1(n19015), .B2(n18823), .ZN(
        n18814) );
  AOI22_X1 U21908 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18825), .B1(
        n19017), .B2(n18898), .ZN(n18813) );
  OAI211_X1 U21909 ( .C1(n18916), .C2(n18821), .A(n18814), .B(n18813), .ZN(
        P3_U2935) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18825), .B1(
        n19021), .B2(n18823), .ZN(n18816) );
  AOI22_X1 U21911 ( .A1(n18944), .A2(n18898), .B1(n19023), .B2(n18824), .ZN(
        n18815) );
  OAI211_X1 U21912 ( .C1(n18891), .C2(n18828), .A(n18816), .B(n18815), .ZN(
        P3_U2936) );
  AOI22_X1 U21913 ( .A1(n19028), .A2(n18843), .B1(n19027), .B2(n18823), .ZN(
        n18818) );
  AOI22_X1 U21914 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18825), .B1(
        n18948), .B2(n18898), .ZN(n18817) );
  OAI211_X1 U21915 ( .C1(n18951), .C2(n18821), .A(n18818), .B(n18817), .ZN(
        P3_U2937) );
  AOI22_X1 U21916 ( .A1(n19035), .A2(n18843), .B1(n19034), .B2(n18823), .ZN(
        n18820) );
  AOI22_X1 U21917 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18825), .B1(
        n18922), .B2(n18898), .ZN(n18819) );
  OAI211_X1 U21918 ( .C1(n18822), .C2(n18821), .A(n18820), .B(n18819), .ZN(
        P3_U2938) );
  AOI22_X1 U21919 ( .A1(n19045), .A2(n18824), .B1(n19043), .B2(n18823), .ZN(
        n18827) );
  AOI22_X1 U21920 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18825), .B1(
        n19046), .B2(n18898), .ZN(n18826) );
  OAI211_X1 U21921 ( .C1(n19051), .C2(n18828), .A(n18827), .B(n18826), .ZN(
        P3_U2939) );
  NOR2_X1 U21922 ( .A1(n18829), .A2(n18852), .ZN(n18928) );
  INV_X1 U21923 ( .A(n18928), .ZN(n18921) );
  NOR2_X1 U21924 ( .A1(n18830), .A2(n18852), .ZN(n18848) );
  AOI22_X1 U21925 ( .A1(n18999), .A2(n18843), .B1(n18993), .B2(n18848), .ZN(
        n18834) );
  INV_X1 U21926 ( .A(n18831), .ZN(n18995) );
  NOR2_X1 U21927 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18852), .ZN(
        n18878) );
  AOI22_X1 U21928 ( .A1(n18998), .A2(n18832), .B1(n18995), .B2(n18878), .ZN(
        n18849) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18849), .B1(
        n18994), .B2(n18873), .ZN(n18833) );
  OAI211_X1 U21930 ( .C1(n19002), .C2(n18921), .A(n18834), .B(n18833), .ZN(
        P3_U2940) );
  AOI22_X1 U21931 ( .A1(n19004), .A2(n18843), .B1(n19003), .B2(n18848), .ZN(
        n18836) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18849), .B1(
        n19005), .B2(n18873), .ZN(n18835) );
  OAI211_X1 U21933 ( .C1(n19008), .C2(n18921), .A(n18836), .B(n18835), .ZN(
        P3_U2941) );
  AOI22_X1 U21934 ( .A1(n18970), .A2(n18873), .B1(n19010), .B2(n18848), .ZN(
        n18838) );
  AOI22_X1 U21935 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18849), .B1(
        n19009), .B2(n18843), .ZN(n18837) );
  OAI211_X1 U21936 ( .C1(n18973), .C2(n18921), .A(n18838), .B(n18837), .ZN(
        P3_U2942) );
  INV_X1 U21937 ( .A(n19017), .ZN(n18977) );
  AOI22_X1 U21938 ( .A1(n19016), .A2(n18843), .B1(n19015), .B2(n18848), .ZN(
        n18840) );
  AOI22_X1 U21939 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18849), .B1(
        n18974), .B2(n18867), .ZN(n18839) );
  OAI211_X1 U21940 ( .C1(n18977), .C2(n18921), .A(n18840), .B(n18839), .ZN(
        P3_U2943) );
  INV_X1 U21941 ( .A(n18944), .ZN(n19026) );
  AOI22_X1 U21942 ( .A1(n19021), .A2(n18848), .B1(n19023), .B2(n18843), .ZN(
        n18842) );
  AOI22_X1 U21943 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18849), .B1(
        n19022), .B2(n18867), .ZN(n18841) );
  OAI211_X1 U21944 ( .C1(n19026), .C2(n18921), .A(n18842), .B(n18841), .ZN(
        P3_U2944) );
  INV_X1 U21945 ( .A(n18948), .ZN(n19033) );
  AOI22_X1 U21946 ( .A1(n19030), .A2(n18843), .B1(n19027), .B2(n18848), .ZN(
        n18845) );
  AOI22_X1 U21947 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18849), .B1(
        n19028), .B2(n18867), .ZN(n18844) );
  OAI211_X1 U21948 ( .C1(n19033), .C2(n18921), .A(n18845), .B(n18844), .ZN(
        P3_U2945) );
  INV_X1 U21949 ( .A(n18922), .ZN(n19040) );
  AOI22_X1 U21950 ( .A1(n19037), .A2(n18843), .B1(n19034), .B2(n18848), .ZN(
        n18847) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18849), .B1(
        n19035), .B2(n18873), .ZN(n18846) );
  OAI211_X1 U21952 ( .C1(n19040), .C2(n18921), .A(n18847), .B(n18846), .ZN(
        P3_U2946) );
  INV_X1 U21953 ( .A(n19046), .ZN(n18991) );
  AOI22_X1 U21954 ( .A1(n19045), .A2(n18843), .B1(n19043), .B2(n18848), .ZN(
        n18851) );
  AOI22_X1 U21955 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18849), .B1(
        n18987), .B2(n18873), .ZN(n18850) );
  OAI211_X1 U21956 ( .C1(n18991), .C2(n18921), .A(n18851), .B(n18850), .ZN(
        P3_U2947) );
  NOR2_X1 U21957 ( .A1(n18853), .A2(n18852), .ZN(n18952) );
  INV_X1 U21958 ( .A(n18952), .ZN(n18959) );
  AOI21_X1 U21959 ( .B1(n18921), .B2(n18959), .A(n18932), .ZN(n18872) );
  AOI22_X1 U21960 ( .A1(n18994), .A2(n18898), .B1(n18993), .B2(n18872), .ZN(
        n18858) );
  OAI211_X1 U21961 ( .C1(n18855), .C2(n18854), .A(n18921), .B(n18959), .ZN(
        n18856) );
  OAI211_X1 U21962 ( .C1(n18952), .C2(n19212), .A(n18905), .B(n18856), .ZN(
        n18874) );
  AOI22_X1 U21963 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18874), .B1(
        n18999), .B2(n18867), .ZN(n18857) );
  OAI211_X1 U21964 ( .C1(n19002), .C2(n18959), .A(n18858), .B(n18857), .ZN(
        P3_U2948) );
  AOI22_X1 U21965 ( .A1(n19005), .A2(n18898), .B1(n19003), .B2(n18872), .ZN(
        n18860) );
  AOI22_X1 U21966 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18874), .B1(
        n19004), .B2(n18867), .ZN(n18859) );
  OAI211_X1 U21967 ( .C1(n19008), .C2(n18959), .A(n18860), .B(n18859), .ZN(
        P3_U2949) );
  AOI22_X1 U21968 ( .A1(n19010), .A2(n18872), .B1(n19009), .B2(n18867), .ZN(
        n18862) );
  AOI22_X1 U21969 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18874), .B1(
        n18970), .B2(n18898), .ZN(n18861) );
  OAI211_X1 U21970 ( .C1(n18973), .C2(n18959), .A(n18862), .B(n18861), .ZN(
        P3_U2950) );
  AOI22_X1 U21971 ( .A1(n19016), .A2(n18873), .B1(n19015), .B2(n18872), .ZN(
        n18864) );
  AOI22_X1 U21972 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18874), .B1(
        n18974), .B2(n18898), .ZN(n18863) );
  OAI211_X1 U21973 ( .C1(n18977), .C2(n18959), .A(n18864), .B(n18863), .ZN(
        P3_U2951) );
  AOI22_X1 U21974 ( .A1(n19021), .A2(n18872), .B1(n19023), .B2(n18867), .ZN(
        n18866) );
  AOI22_X1 U21975 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18874), .B1(
        n19022), .B2(n18898), .ZN(n18865) );
  OAI211_X1 U21976 ( .C1(n19026), .C2(n18959), .A(n18866), .B(n18865), .ZN(
        P3_U2952) );
  AOI22_X1 U21977 ( .A1(n19028), .A2(n18898), .B1(n19027), .B2(n18872), .ZN(
        n18869) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18874), .B1(
        n19030), .B2(n18867), .ZN(n18868) );
  OAI211_X1 U21979 ( .C1(n19033), .C2(n18959), .A(n18869), .B(n18868), .ZN(
        P3_U2953) );
  AOI22_X1 U21980 ( .A1(n19035), .A2(n18898), .B1(n19034), .B2(n18872), .ZN(
        n18871) );
  AOI22_X1 U21981 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18874), .B1(
        n19037), .B2(n18873), .ZN(n18870) );
  OAI211_X1 U21982 ( .C1(n19040), .C2(n18959), .A(n18871), .B(n18870), .ZN(
        P3_U2954) );
  AOI22_X1 U21983 ( .A1(n19045), .A2(n18873), .B1(n19043), .B2(n18872), .ZN(
        n18876) );
  AOI22_X1 U21984 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18874), .B1(
        n18987), .B2(n18898), .ZN(n18875) );
  OAI211_X1 U21985 ( .C1(n18991), .C2(n18959), .A(n18876), .B(n18875), .ZN(
        P3_U2955) );
  NAND2_X1 U21986 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18877), .ZN(
        n18879) );
  NOR2_X1 U21987 ( .A1(n18932), .A2(n18879), .ZN(n18897) );
  AOI22_X1 U21988 ( .A1(n18999), .A2(n18898), .B1(n18993), .B2(n18897), .ZN(
        n18881) );
  INV_X1 U21989 ( .A(n18879), .ZN(n18933) );
  AOI22_X1 U21990 ( .A1(n18998), .A2(n18878), .B1(n18995), .B2(n18933), .ZN(
        n18899) );
  NOR2_X1 U21991 ( .A1(n19066), .A2(n18879), .ZN(n18980) );
  AOI22_X1 U21992 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18899), .B1(
        n18906), .B2(n18980), .ZN(n18880) );
  OAI211_X1 U21993 ( .C1(n18909), .C2(n18921), .A(n18881), .B(n18880), .ZN(
        P3_U2956) );
  AOI22_X1 U21994 ( .A1(n19005), .A2(n18928), .B1(n19003), .B2(n18897), .ZN(
        n18883) );
  CLKBUF_X1 U21995 ( .A(n18980), .Z(n18986) );
  AOI22_X1 U21996 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18899), .B1(
        n18936), .B2(n18986), .ZN(n18882) );
  OAI211_X1 U21997 ( .C1(n18939), .C2(n18888), .A(n18883), .B(n18882), .ZN(
        P3_U2957) );
  AOI22_X1 U21998 ( .A1(n19010), .A2(n18897), .B1(n19009), .B2(n18898), .ZN(
        n18885) );
  AOI22_X1 U21999 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18899), .B1(
        n19011), .B2(n18986), .ZN(n18884) );
  OAI211_X1 U22000 ( .C1(n19014), .C2(n18921), .A(n18885), .B(n18884), .ZN(
        P3_U2958) );
  AOI22_X1 U22001 ( .A1(n18974), .A2(n18928), .B1(n19015), .B2(n18897), .ZN(
        n18887) );
  AOI22_X1 U22002 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18899), .B1(
        n19017), .B2(n18980), .ZN(n18886) );
  OAI211_X1 U22003 ( .C1(n18916), .C2(n18888), .A(n18887), .B(n18886), .ZN(
        P3_U2959) );
  AOI22_X1 U22004 ( .A1(n19021), .A2(n18897), .B1(n19023), .B2(n18898), .ZN(
        n18890) );
  AOI22_X1 U22005 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18899), .B1(
        n18944), .B2(n18980), .ZN(n18889) );
  OAI211_X1 U22006 ( .C1(n18891), .C2(n18921), .A(n18890), .B(n18889), .ZN(
        P3_U2960) );
  AOI22_X1 U22007 ( .A1(n19030), .A2(n18898), .B1(n19027), .B2(n18897), .ZN(
        n18893) );
  AOI22_X1 U22008 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18899), .B1(
        n18948), .B2(n18980), .ZN(n18892) );
  OAI211_X1 U22009 ( .C1(n18894), .C2(n18921), .A(n18893), .B(n18892), .ZN(
        P3_U2961) );
  AOI22_X1 U22010 ( .A1(n19037), .A2(n18898), .B1(n19034), .B2(n18897), .ZN(
        n18896) );
  AOI22_X1 U22011 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18899), .B1(
        n18922), .B2(n18980), .ZN(n18895) );
  OAI211_X1 U22012 ( .C1(n18925), .C2(n18921), .A(n18896), .B(n18895), .ZN(
        P3_U2962) );
  AOI22_X1 U22013 ( .A1(n19045), .A2(n18898), .B1(n19043), .B2(n18897), .ZN(
        n18901) );
  AOI22_X1 U22014 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18899), .B1(
        n19046), .B2(n18980), .ZN(n18900) );
  OAI211_X1 U22015 ( .C1(n19051), .C2(n18921), .A(n18901), .B(n18900), .ZN(
        P3_U2963) );
  NOR2_X1 U22016 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18931), .ZN(
        n19029) );
  CLKBUF_X1 U22017 ( .A(n19029), .Z(n19044) );
  NOR2_X1 U22018 ( .A1(n18986), .A2(n19044), .ZN(n18961) );
  OAI21_X1 U22019 ( .B1(n18903), .B2(n18902), .A(n18961), .ZN(n18904) );
  OAI211_X1 U22020 ( .C1(n19029), .C2(n19212), .A(n18905), .B(n18904), .ZN(
        n18927) );
  NOR2_X1 U22021 ( .A1(n18932), .A2(n18961), .ZN(n18926) );
  AOI22_X1 U22022 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18927), .B1(
        n18993), .B2(n18926), .ZN(n18908) );
  AOI22_X1 U22023 ( .A1(n18906), .A2(n19044), .B1(n18999), .B2(n18928), .ZN(
        n18907) );
  OAI211_X1 U22024 ( .C1(n18909), .C2(n18959), .A(n18908), .B(n18907), .ZN(
        P3_U2964) );
  AOI22_X1 U22025 ( .A1(n19005), .A2(n18952), .B1(n19003), .B2(n18926), .ZN(
        n18911) );
  AOI22_X1 U22026 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18927), .B1(
        n18936), .B2(n19044), .ZN(n18910) );
  OAI211_X1 U22027 ( .C1(n18939), .C2(n18921), .A(n18911), .B(n18910), .ZN(
        P3_U2965) );
  AOI22_X1 U22028 ( .A1(n19010), .A2(n18926), .B1(n19009), .B2(n18928), .ZN(
        n18913) );
  AOI22_X1 U22029 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18927), .B1(
        n19011), .B2(n19029), .ZN(n18912) );
  OAI211_X1 U22030 ( .C1(n19014), .C2(n18959), .A(n18913), .B(n18912), .ZN(
        P3_U2966) );
  AOI22_X1 U22031 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18927), .B1(
        n19015), .B2(n18926), .ZN(n18915) );
  AOI22_X1 U22032 ( .A1(n18974), .A2(n18952), .B1(n19017), .B2(n19029), .ZN(
        n18914) );
  OAI211_X1 U22033 ( .C1(n18916), .C2(n18921), .A(n18915), .B(n18914), .ZN(
        P3_U2967) );
  AOI22_X1 U22034 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18927), .B1(
        n19021), .B2(n18926), .ZN(n18918) );
  AOI22_X1 U22035 ( .A1(n19022), .A2(n18952), .B1(n18944), .B2(n19044), .ZN(
        n18917) );
  OAI211_X1 U22036 ( .C1(n18947), .C2(n18921), .A(n18918), .B(n18917), .ZN(
        P3_U2968) );
  AOI22_X1 U22037 ( .A1(n19028), .A2(n18952), .B1(n19027), .B2(n18926), .ZN(
        n18920) );
  AOI22_X1 U22038 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18927), .B1(
        n18948), .B2(n19029), .ZN(n18919) );
  OAI211_X1 U22039 ( .C1(n18951), .C2(n18921), .A(n18920), .B(n18919), .ZN(
        P3_U2969) );
  AOI22_X1 U22040 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18927), .B1(
        n19034), .B2(n18926), .ZN(n18924) );
  AOI22_X1 U22041 ( .A1(n18922), .A2(n19044), .B1(n19037), .B2(n18928), .ZN(
        n18923) );
  OAI211_X1 U22042 ( .C1(n18925), .C2(n18959), .A(n18924), .B(n18923), .ZN(
        P3_U2970) );
  AOI22_X1 U22043 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18927), .B1(
        n19043), .B2(n18926), .ZN(n18930) );
  AOI22_X1 U22044 ( .A1(n19045), .A2(n18928), .B1(n19046), .B2(n19044), .ZN(
        n18929) );
  OAI211_X1 U22045 ( .C1(n19051), .C2(n18959), .A(n18930), .B(n18929), .ZN(
        P3_U2971) );
  NOR2_X1 U22046 ( .A1(n18932), .A2(n18931), .ZN(n18955) );
  AOI22_X1 U22047 ( .A1(n18994), .A2(n18986), .B1(n18993), .B2(n18955), .ZN(
        n18935) );
  AOI22_X1 U22048 ( .A1(n18998), .A2(n18933), .B1(n18997), .B2(n18995), .ZN(
        n18956) );
  AOI22_X1 U22049 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18956), .B1(
        n18999), .B2(n18952), .ZN(n18934) );
  OAI211_X1 U22050 ( .C1(n19002), .C2(n19052), .A(n18935), .B(n18934), .ZN(
        P3_U2972) );
  AOI22_X1 U22051 ( .A1(n19005), .A2(n18986), .B1(n19003), .B2(n18955), .ZN(
        n18938) );
  AOI22_X1 U22052 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18956), .B1(
        n19036), .B2(n18936), .ZN(n18937) );
  OAI211_X1 U22053 ( .C1(n18939), .C2(n18959), .A(n18938), .B(n18937), .ZN(
        P3_U2973) );
  AOI22_X1 U22054 ( .A1(n19010), .A2(n18955), .B1(n19009), .B2(n18952), .ZN(
        n18941) );
  AOI22_X1 U22055 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18956), .B1(
        n18970), .B2(n18980), .ZN(n18940) );
  OAI211_X1 U22056 ( .C1(n19052), .C2(n18973), .A(n18941), .B(n18940), .ZN(
        P3_U2974) );
  AOI22_X1 U22057 ( .A1(n19016), .A2(n18952), .B1(n19015), .B2(n18955), .ZN(
        n18943) );
  AOI22_X1 U22058 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18956), .B1(
        n18974), .B2(n18980), .ZN(n18942) );
  OAI211_X1 U22059 ( .C1(n19052), .C2(n18977), .A(n18943), .B(n18942), .ZN(
        P3_U2975) );
  AOI22_X1 U22060 ( .A1(n19022), .A2(n18986), .B1(n19021), .B2(n18955), .ZN(
        n18946) );
  AOI22_X1 U22061 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18956), .B1(
        n19036), .B2(n18944), .ZN(n18945) );
  OAI211_X1 U22062 ( .C1(n18947), .C2(n18959), .A(n18946), .B(n18945), .ZN(
        P3_U2976) );
  AOI22_X1 U22063 ( .A1(n19028), .A2(n18986), .B1(n19027), .B2(n18955), .ZN(
        n18950) );
  AOI22_X1 U22064 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18956), .B1(
        n19036), .B2(n18948), .ZN(n18949) );
  OAI211_X1 U22065 ( .C1(n18951), .C2(n18959), .A(n18950), .B(n18949), .ZN(
        P3_U2977) );
  AOI22_X1 U22066 ( .A1(n19037), .A2(n18952), .B1(n19034), .B2(n18955), .ZN(
        n18954) );
  AOI22_X1 U22067 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18956), .B1(
        n19035), .B2(n18980), .ZN(n18953) );
  OAI211_X1 U22068 ( .C1(n19052), .C2(n19040), .A(n18954), .B(n18953), .ZN(
        P3_U2978) );
  AOI22_X1 U22069 ( .A1(n18987), .A2(n18986), .B1(n19043), .B2(n18955), .ZN(
        n18958) );
  AOI22_X1 U22070 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18956), .B1(
        n19036), .B2(n19046), .ZN(n18957) );
  OAI211_X1 U22071 ( .C1(n18960), .C2(n18959), .A(n18958), .B(n18957), .ZN(
        P3_U2979) );
  AND2_X1 U22072 ( .A1(n19113), .A2(n18965), .ZN(n18985) );
  AOI22_X1 U22073 ( .A1(n18999), .A2(n18986), .B1(n18993), .B2(n18985), .ZN(
        n18967) );
  INV_X1 U22074 ( .A(n18961), .ZN(n18963) );
  OAI221_X1 U22075 ( .B1(n18965), .B2(n18964), .C1(n18965), .C2(n18963), .A(
        n18962), .ZN(n18988) );
  AOI22_X1 U22076 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18988), .B1(
        n18994), .B2(n19029), .ZN(n18966) );
  OAI211_X1 U22077 ( .C1(n18992), .C2(n19002), .A(n18967), .B(n18966), .ZN(
        P3_U2980) );
  AOI22_X1 U22078 ( .A1(n19004), .A2(n18986), .B1(n19003), .B2(n18985), .ZN(
        n18969) );
  AOI22_X1 U22079 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18988), .B1(
        n19005), .B2(n19029), .ZN(n18968) );
  OAI211_X1 U22080 ( .C1(n18992), .C2(n19008), .A(n18969), .B(n18968), .ZN(
        P3_U2981) );
  AOI22_X1 U22081 ( .A1(n19010), .A2(n18985), .B1(n19009), .B2(n18986), .ZN(
        n18972) );
  AOI22_X1 U22082 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18988), .B1(
        n18970), .B2(n19029), .ZN(n18971) );
  OAI211_X1 U22083 ( .C1(n18992), .C2(n18973), .A(n18972), .B(n18971), .ZN(
        P3_U2982) );
  AOI22_X1 U22084 ( .A1(n19016), .A2(n18986), .B1(n19015), .B2(n18985), .ZN(
        n18976) );
  AOI22_X1 U22085 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18988), .B1(
        n18974), .B2(n19029), .ZN(n18975) );
  OAI211_X1 U22086 ( .C1(n18992), .C2(n18977), .A(n18976), .B(n18975), .ZN(
        P3_U2983) );
  AOI22_X1 U22087 ( .A1(n19021), .A2(n18985), .B1(n19023), .B2(n18986), .ZN(
        n18979) );
  AOI22_X1 U22088 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18988), .B1(
        n19022), .B2(n19029), .ZN(n18978) );
  OAI211_X1 U22089 ( .C1(n18992), .C2(n19026), .A(n18979), .B(n18978), .ZN(
        P3_U2984) );
  AOI22_X1 U22090 ( .A1(n19028), .A2(n19044), .B1(n19027), .B2(n18985), .ZN(
        n18982) );
  AOI22_X1 U22091 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18988), .B1(
        n19030), .B2(n18980), .ZN(n18981) );
  OAI211_X1 U22092 ( .C1(n18992), .C2(n19033), .A(n18982), .B(n18981), .ZN(
        P3_U2985) );
  AOI22_X1 U22093 ( .A1(n19037), .A2(n18986), .B1(n19034), .B2(n18985), .ZN(
        n18984) );
  AOI22_X1 U22094 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18988), .B1(
        n19035), .B2(n19029), .ZN(n18983) );
  OAI211_X1 U22095 ( .C1(n18992), .C2(n19040), .A(n18984), .B(n18983), .ZN(
        P3_U2986) );
  AOI22_X1 U22096 ( .A1(n19045), .A2(n18986), .B1(n19043), .B2(n18985), .ZN(
        n18990) );
  AOI22_X1 U22097 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18988), .B1(
        n18987), .B2(n19044), .ZN(n18989) );
  OAI211_X1 U22098 ( .C1(n18992), .C2(n18991), .A(n18990), .B(n18989), .ZN(
        P3_U2987) );
  AND2_X1 U22099 ( .A1(n19113), .A2(n18996), .ZN(n19042) );
  AOI22_X1 U22100 ( .A1(n18994), .A2(n19036), .B1(n18993), .B2(n19042), .ZN(
        n19001) );
  AOI22_X1 U22101 ( .A1(n18998), .A2(n18997), .B1(n18996), .B2(n18995), .ZN(
        n19048) );
  AOI22_X1 U22102 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19048), .B1(
        n18999), .B2(n19044), .ZN(n19000) );
  OAI211_X1 U22103 ( .C1(n19041), .C2(n19002), .A(n19001), .B(n19000), .ZN(
        P3_U2988) );
  AOI22_X1 U22104 ( .A1(n19004), .A2(n19044), .B1(n19003), .B2(n19042), .ZN(
        n19007) );
  AOI22_X1 U22105 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19048), .B1(
        n19036), .B2(n19005), .ZN(n19006) );
  OAI211_X1 U22106 ( .C1(n19041), .C2(n19008), .A(n19007), .B(n19006), .ZN(
        P3_U2989) );
  AOI22_X1 U22107 ( .A1(n19010), .A2(n19042), .B1(n19009), .B2(n19044), .ZN(
        n19013) );
  AOI22_X1 U22108 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n19011), .ZN(n19012) );
  OAI211_X1 U22109 ( .C1(n19052), .C2(n19014), .A(n19013), .B(n19012), .ZN(
        P3_U2990) );
  AOI22_X1 U22110 ( .A1(n19016), .A2(n19044), .B1(n19015), .B2(n19042), .ZN(
        n19019) );
  AOI22_X1 U22111 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n19017), .ZN(n19018) );
  OAI211_X1 U22112 ( .C1(n19052), .C2(n19020), .A(n19019), .B(n19018), .ZN(
        P3_U2991) );
  AOI22_X1 U22113 ( .A1(n19036), .A2(n19022), .B1(n19021), .B2(n19042), .ZN(
        n19025) );
  AOI22_X1 U22114 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19048), .B1(
        n19023), .B2(n19044), .ZN(n19024) );
  OAI211_X1 U22115 ( .C1(n19041), .C2(n19026), .A(n19025), .B(n19024), .ZN(
        P3_U2992) );
  AOI22_X1 U22116 ( .A1(n19036), .A2(n19028), .B1(n19027), .B2(n19042), .ZN(
        n19032) );
  AOI22_X1 U22117 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19048), .B1(
        n19030), .B2(n19029), .ZN(n19031) );
  OAI211_X1 U22118 ( .C1(n19041), .C2(n19033), .A(n19032), .B(n19031), .ZN(
        P3_U2993) );
  AOI22_X1 U22119 ( .A1(n19036), .A2(n19035), .B1(n19034), .B2(n19042), .ZN(
        n19039) );
  AOI22_X1 U22120 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19048), .B1(
        n19037), .B2(n19044), .ZN(n19038) );
  OAI211_X1 U22121 ( .C1(n19041), .C2(n19040), .A(n19039), .B(n19038), .ZN(
        P3_U2994) );
  AOI22_X1 U22122 ( .A1(n19045), .A2(n19044), .B1(n19043), .B2(n19042), .ZN(
        n19050) );
  AOI22_X1 U22123 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n19046), .ZN(n19049) );
  OAI211_X1 U22124 ( .C1(n19052), .C2(n19051), .A(n19050), .B(n19049), .ZN(
        P3_U2995) );
  OAI22_X1 U22125 ( .A1(n19056), .A2(n19055), .B1(n19054), .B2(n19053), .ZN(
        n19057) );
  AOI221_X1 U22126 ( .B1(n19060), .B2(n19059), .C1(n19058), .C2(n19059), .A(
        n19057), .ZN(n19252) );
  AOI211_X1 U22127 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19091), .A(
        n19062), .B(n19061), .ZN(n19101) );
  NAND2_X1 U22128 ( .A1(n19064), .A2(n19063), .ZN(n19065) );
  OAI21_X1 U22129 ( .B1(n19064), .B2(n17332), .A(n9780), .ZN(n19085) );
  AOI22_X1 U22130 ( .A1(n19231), .A2(n19065), .B1(n19234), .B2(n19085), .ZN(
        n19227) );
  AOI22_X1 U22131 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19080), .B1(
        n19065), .B2(n17332), .ZN(n19068) );
  INV_X1 U22132 ( .A(n19068), .ZN(n19236) );
  NOR3_X1 U22133 ( .A1(n19067), .A2(n19066), .A3(n19236), .ZN(n19069) );
  OAI22_X1 U22134 ( .A1(n19227), .A2(n19069), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19068), .ZN(n19071) );
  AOI21_X1 U22135 ( .B1(n19071), .B2(n10333), .A(n19070), .ZN(n19078) );
  AOI21_X1 U22136 ( .B1(n19074), .B2(n19073), .A(n19072), .ZN(n19084) );
  OR3_X1 U22137 ( .A1(n19226), .A2(n11865), .A3(n19084), .ZN(n19076) );
  OAI211_X1 U22138 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n19085), .B(n19086), .ZN(
        n19075) );
  OAI211_X1 U22139 ( .C1(n19223), .C2(n19088), .A(n19076), .B(n19075), .ZN(
        n19224) );
  AOI22_X1 U22140 ( .A1(n19091), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19224), .B2(n10333), .ZN(n19093) );
  OR2_X1 U22141 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19093), .ZN(
        n19077) );
  AOI221_X1 U22142 ( .B1(n19078), .B2(n19077), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n19093), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19097) );
  AOI22_X1 U22143 ( .A1(n19226), .A2(n19081), .B1(n19080), .B2(n19086), .ZN(
        n19082) );
  OAI21_X1 U22144 ( .B1(n19084), .B2(n19083), .A(n19082), .ZN(n19218) );
  NOR2_X1 U22145 ( .A1(n19218), .A2(n19091), .ZN(n19092) );
  NOR2_X1 U22146 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11865), .ZN(
        n19089) );
  INV_X1 U22147 ( .A(n19085), .ZN(n19087) );
  OAI22_X1 U22148 ( .A1(n19089), .A2(n19088), .B1(n19087), .B2(n19086), .ZN(
        n19090) );
  NAND2_X1 U22149 ( .A1(n19079), .A2(n19090), .ZN(n19215) );
  OAI22_X1 U22150 ( .A1(n19079), .A2(n19092), .B1(n19091), .B2(n19215), .ZN(
        n19096) );
  OAI21_X1 U22151 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n19093), .ZN(n19094) );
  AOI222_X1 U22152 ( .A1(n19097), .A2(n19096), .B1(n19097), .B2(n19095), .C1(
        n19096), .C2(n19094), .ZN(n19100) );
  OAI21_X1 U22153 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19098), .ZN(n19099) );
  NOR2_X1 U22154 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19254), .ZN(n19112) );
  NOR2_X1 U22155 ( .A1(n19105), .A2(n19113), .ZN(n19108) );
  NAND2_X1 U22156 ( .A1(n19261), .A2(n19255), .ZN(n19117) );
  INV_X1 U22157 ( .A(n19117), .ZN(n19106) );
  AOI211_X1 U22158 ( .C1(n19235), .C2(n19266), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n19106), .ZN(n19107) );
  AOI211_X1 U22159 ( .C1(n19258), .C2(n19109), .A(n19108), .B(n19107), .ZN(
        n19110) );
  NAND3_X1 U22160 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n19112), .ZN(n19120) );
  NAND3_X1 U22161 ( .A1(n19115), .A2(n19114), .A3(n19113), .ZN(n19116) );
  NAND4_X1 U22162 ( .A1(n19118), .A2(n19117), .A3(n19120), .A4(n19116), .ZN(
        P3_U2997) );
  OAI21_X1 U22163 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n19119), .ZN(n19122) );
  INV_X1 U22164 ( .A(n19120), .ZN(n19121) );
  AOI21_X1 U22165 ( .B1(n19123), .B2(n19122), .A(n19121), .ZN(P3_U2998) );
  AND2_X1 U22166 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19204), .ZN(
        P3_U2999) );
  AND2_X1 U22167 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19204), .ZN(
        P3_U3000) );
  AND2_X1 U22168 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19204), .ZN(
        P3_U3001) );
  AND2_X1 U22169 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19204), .ZN(
        P3_U3002) );
  AND2_X1 U22170 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19204), .ZN(
        P3_U3003) );
  AND2_X1 U22171 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19204), .ZN(
        P3_U3004) );
  AND2_X1 U22172 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19204), .ZN(
        P3_U3005) );
  AND2_X1 U22173 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19204), .ZN(
        P3_U3006) );
  AND2_X1 U22174 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19204), .ZN(
        P3_U3007) );
  AND2_X1 U22175 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19204), .ZN(
        P3_U3008) );
  AND2_X1 U22176 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19204), .ZN(
        P3_U3009) );
  AND2_X1 U22177 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19204), .ZN(
        P3_U3010) );
  AND2_X1 U22178 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19204), .ZN(
        P3_U3011) );
  AND2_X1 U22179 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19204), .ZN(
        P3_U3012) );
  AND2_X1 U22180 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19204), .ZN(
        P3_U3013) );
  AND2_X1 U22181 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19204), .ZN(
        P3_U3014) );
  AND2_X1 U22182 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19204), .ZN(
        P3_U3015) );
  AND2_X1 U22183 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19204), .ZN(
        P3_U3016) );
  AND2_X1 U22184 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19204), .ZN(
        P3_U3017) );
  AND2_X1 U22185 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19204), .ZN(
        P3_U3018) );
  AND2_X1 U22186 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19204), .ZN(
        P3_U3019) );
  INV_X1 U22187 ( .A(P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21307) );
  NOR2_X1 U22188 ( .A1(n19208), .A2(n21307), .ZN(P3_U3020) );
  AND2_X1 U22189 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19204), .ZN(P3_U3021) );
  AND2_X1 U22190 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19204), .ZN(P3_U3022) );
  AND2_X1 U22191 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19204), .ZN(P3_U3023) );
  AND2_X1 U22192 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19204), .ZN(P3_U3024) );
  AND2_X1 U22193 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19204), .ZN(P3_U3025) );
  AND2_X1 U22194 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19204), .ZN(P3_U3026) );
  AND2_X1 U22195 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19204), .ZN(P3_U3027) );
  AND2_X1 U22196 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19204), .ZN(P3_U3028) );
  INV_X1 U22197 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19268) );
  AOI21_X1 U22198 ( .B1(HOLD), .B2(n19124), .A(n19268), .ZN(n19126) );
  AOI21_X1 U22199 ( .B1(n19261), .B2(P3_STATE_REG_1__SCAN_IN), .A(n19134), 
        .ZN(n19136) );
  INV_X1 U22200 ( .A(NA), .ZN(n21099) );
  OAI21_X1 U22201 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n21099), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n19135) );
  INV_X1 U22202 ( .A(n19135), .ZN(n19125) );
  OAI22_X1 U22203 ( .A1(n19272), .A2(n19126), .B1(n19136), .B2(n19125), .ZN(
        P3_U3029) );
  INV_X1 U22204 ( .A(HOLD), .ZN(n21095) );
  NOR2_X1 U22205 ( .A1(n19137), .A2(n21095), .ZN(n19132) );
  NOR3_X1 U22206 ( .A1(n19132), .A2(n19134), .A3(n19268), .ZN(n19127) );
  NOR2_X1 U22207 ( .A1(n19127), .A2(n19259), .ZN(n19128) );
  NAND2_X1 U22208 ( .A1(n19261), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19130) );
  OAI211_X1 U22209 ( .C1(n21095), .C2(n19129), .A(n19128), .B(n19130), .ZN(
        P3_U3030) );
  OAI22_X1 U22210 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19130), .ZN(n19131) );
  OAI22_X1 U22211 ( .A1(n19132), .A2(n19131), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19133) );
  OAI22_X1 U22212 ( .A1(n19136), .A2(n19135), .B1(n19134), .B2(n19133), .ZN(
        P3_U3031) );
  NAND2_X1 U22213 ( .A1(n19272), .A2(n19137), .ZN(n19192) );
  CLKBUF_X1 U22214 ( .A(n19192), .Z(n19193) );
  OAI222_X1 U22215 ( .A1(n19241), .A2(n19189), .B1(n19138), .B2(n19272), .C1(
        n19139), .C2(n19193), .ZN(P3_U3032) );
  OAI222_X1 U22216 ( .A1(n19193), .A2(n19141), .B1(n19140), .B2(n19272), .C1(
        n19139), .C2(n19189), .ZN(P3_U3033) );
  OAI222_X1 U22217 ( .A1(n19192), .A2(n19143), .B1(n19142), .B2(n19272), .C1(
        n19141), .C2(n19189), .ZN(P3_U3034) );
  INV_X1 U22218 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19146) );
  OAI222_X1 U22219 ( .A1(n19192), .A2(n19146), .B1(n19144), .B2(n19272), .C1(
        n19143), .C2(n19189), .ZN(P3_U3035) );
  OAI222_X1 U22220 ( .A1(n19146), .A2(n19189), .B1(n19145), .B2(n19272), .C1(
        n19147), .C2(n19193), .ZN(P3_U3036) );
  INV_X1 U22221 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19148) );
  OAI222_X1 U22222 ( .A1(n19192), .A2(n19149), .B1(n19148), .B2(n19272), .C1(
        n19147), .C2(n19189), .ZN(P3_U3037) );
  OAI222_X1 U22223 ( .A1(n19192), .A2(n19152), .B1(n19150), .B2(n19272), .C1(
        n19149), .C2(n19189), .ZN(P3_U3038) );
  OAI222_X1 U22224 ( .A1(n19152), .A2(n19189), .B1(n19151), .B2(n19272), .C1(
        n19153), .C2(n19193), .ZN(P3_U3039) );
  OAI222_X1 U22225 ( .A1(n19192), .A2(n19155), .B1(n19154), .B2(n19272), .C1(
        n19153), .C2(n19189), .ZN(P3_U3040) );
  OAI222_X1 U22226 ( .A1(n19193), .A2(n19156), .B1(n21381), .B2(n19272), .C1(
        n19155), .C2(n19189), .ZN(P3_U3041) );
  OAI222_X1 U22227 ( .A1(n19193), .A2(n19158), .B1(n19157), .B2(n19272), .C1(
        n19156), .C2(n19189), .ZN(P3_U3042) );
  OAI222_X1 U22228 ( .A1(n19193), .A2(n19160), .B1(n19159), .B2(n19272), .C1(
        n19158), .C2(n19189), .ZN(P3_U3043) );
  OAI222_X1 U22229 ( .A1(n19193), .A2(n21405), .B1(n19161), .B2(n19272), .C1(
        n19160), .C2(n19189), .ZN(P3_U3044) );
  OAI222_X1 U22230 ( .A1(n21405), .A2(n19189), .B1(n19162), .B2(n19272), .C1(
        n19163), .C2(n19193), .ZN(P3_U3045) );
  OAI222_X1 U22231 ( .A1(n19193), .A2(n19165), .B1(n19164), .B2(n19272), .C1(
        n19163), .C2(n19189), .ZN(P3_U3046) );
  INV_X1 U22232 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19168) );
  OAI222_X1 U22233 ( .A1(n19193), .A2(n19168), .B1(n19166), .B2(n19272), .C1(
        n19165), .C2(n19189), .ZN(P3_U3047) );
  OAI222_X1 U22234 ( .A1(n19168), .A2(n19189), .B1(n19167), .B2(n19272), .C1(
        n19169), .C2(n19193), .ZN(P3_U3048) );
  INV_X1 U22235 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19171) );
  OAI222_X1 U22236 ( .A1(n19192), .A2(n19171), .B1(n19170), .B2(n19272), .C1(
        n19169), .C2(n19189), .ZN(P3_U3049) );
  INV_X1 U22237 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19173) );
  OAI222_X1 U22238 ( .A1(n19192), .A2(n19173), .B1(n19172), .B2(n19272), .C1(
        n19171), .C2(n19189), .ZN(P3_U3050) );
  OAI222_X1 U22239 ( .A1(n19192), .A2(n19175), .B1(n19174), .B2(n19272), .C1(
        n19173), .C2(n19189), .ZN(P3_U3051) );
  INV_X1 U22240 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21373) );
  OAI222_X1 U22241 ( .A1(n19192), .A2(n21373), .B1(n19176), .B2(n19272), .C1(
        n19175), .C2(n19189), .ZN(P3_U3052) );
  OAI222_X1 U22242 ( .A1(n19193), .A2(n19178), .B1(n19177), .B2(n19272), .C1(
        n21373), .C2(n19189), .ZN(P3_U3053) );
  OAI222_X1 U22243 ( .A1(n19192), .A2(n19180), .B1(n19179), .B2(n19272), .C1(
        n19178), .C2(n19189), .ZN(P3_U3054) );
  OAI222_X1 U22244 ( .A1(n19192), .A2(n19182), .B1(n19181), .B2(n19272), .C1(
        n19180), .C2(n19189), .ZN(P3_U3055) );
  OAI222_X1 U22245 ( .A1(n19193), .A2(n19184), .B1(n19183), .B2(n19272), .C1(
        n19182), .C2(n19189), .ZN(P3_U3056) );
  INV_X1 U22246 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19186) );
  OAI222_X1 U22247 ( .A1(n19193), .A2(n19186), .B1(n19185), .B2(n19272), .C1(
        n19184), .C2(n19189), .ZN(P3_U3057) );
  INV_X1 U22248 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19190) );
  OAI222_X1 U22249 ( .A1(n19193), .A2(n19190), .B1(n19187), .B2(n19272), .C1(
        n19186), .C2(n19189), .ZN(P3_U3058) );
  OAI222_X1 U22250 ( .A1(n19190), .A2(n19189), .B1(n19188), .B2(n19272), .C1(
        n21459), .C2(n19193), .ZN(P3_U3059) );
  OAI222_X1 U22251 ( .A1(n19192), .A2(n19196), .B1(n19191), .B2(n19272), .C1(
        n21459), .C2(n19189), .ZN(P3_U3060) );
  OAI222_X1 U22252 ( .A1(n19189), .A2(n19196), .B1(n19195), .B2(n19272), .C1(
        n19194), .C2(n19193), .ZN(P3_U3061) );
  INV_X1 U22253 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19197) );
  AOI22_X1 U22254 ( .A1(n19272), .A2(n19198), .B1(n19197), .B2(n19270), .ZN(
        P3_U3274) );
  INV_X1 U22255 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19243) );
  INV_X1 U22256 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19199) );
  AOI22_X1 U22257 ( .A1(n19272), .A2(n19243), .B1(n19199), .B2(n19270), .ZN(
        P3_U3275) );
  INV_X1 U22258 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19200) );
  AOI22_X1 U22259 ( .A1(n19272), .A2(n19201), .B1(n19200), .B2(n19270), .ZN(
        P3_U3276) );
  INV_X1 U22260 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19248) );
  INV_X1 U22261 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19202) );
  AOI22_X1 U22262 ( .A1(n19272), .A2(n19248), .B1(n19202), .B2(n19270), .ZN(
        P3_U3277) );
  INV_X1 U22263 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19205) );
  INV_X1 U22264 ( .A(n19206), .ZN(n19203) );
  AOI21_X1 U22265 ( .B1(n19205), .B2(n19204), .A(n19203), .ZN(P3_U3280) );
  OAI21_X1 U22266 ( .B1(n19208), .B2(n19207), .A(n19206), .ZN(P3_U3281) );
  INV_X1 U22267 ( .A(n19209), .ZN(n19211) );
  OAI221_X1 U22268 ( .B1(n19212), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19212), 
        .C2(n19211), .A(n19210), .ZN(P3_U3282) );
  OAI22_X1 U22269 ( .A1(n19216), .A2(n19215), .B1(n19214), .B2(n19213), .ZN(
        n19217) );
  INV_X1 U22270 ( .A(n19217), .ZN(n19220) );
  AOI21_X1 U22271 ( .B1(n19274), .B2(n19218), .A(n19240), .ZN(n19219) );
  OAI22_X1 U22272 ( .A1(n19240), .A2(n19220), .B1(n19219), .B2(n19079), .ZN(
        P3_U3285) );
  NOR2_X1 U22273 ( .A1(n19221), .A2(n19237), .ZN(n19229) );
  AOI22_X1 U22274 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n21317), .B2(n19222), .ZN(
        n19228) );
  AOI222_X1 U22275 ( .A1(n19224), .A2(n19274), .B1(n19229), .B2(n19228), .C1(
        n19235), .C2(n19223), .ZN(n19225) );
  AOI22_X1 U22276 ( .A1(n19240), .A2(n19226), .B1(n19225), .B2(n19238), .ZN(
        P3_U3288) );
  INV_X1 U22277 ( .A(n19227), .ZN(n19232) );
  INV_X1 U22278 ( .A(n19228), .ZN(n19230) );
  AOI222_X1 U22279 ( .A1(n19232), .A2(n19274), .B1(n19235), .B2(n19231), .C1(
        n19230), .C2(n19229), .ZN(n19233) );
  AOI22_X1 U22280 ( .A1(n19240), .A2(n19234), .B1(n19233), .B2(n19238), .ZN(
        P3_U3289) );
  AOI222_X1 U22281 ( .A1(n19237), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19274), 
        .B2(n19236), .C1(n17332), .C2(n19235), .ZN(n19239) );
  AOI22_X1 U22282 ( .A1(n19240), .A2(n17332), .B1(n19239), .B2(n19238), .ZN(
        P3_U3290) );
  AOI21_X1 U22283 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19242) );
  AOI22_X1 U22284 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19242), .B2(n19241), .ZN(n19244) );
  AOI22_X1 U22285 ( .A1(n19245), .A2(n19244), .B1(n19243), .B2(n19247), .ZN(
        P3_U3292) );
  INV_X1 U22286 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n21367) );
  NOR2_X1 U22287 ( .A1(n19247), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19246) );
  AOI22_X1 U22288 ( .A1(n19248), .A2(n19247), .B1(n21367), .B2(n19246), .ZN(
        P3_U3293) );
  INV_X1 U22289 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19249) );
  AOI22_X1 U22290 ( .A1(n19272), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19249), 
        .B2(n19270), .ZN(P3_U3294) );
  INV_X1 U22291 ( .A(n19250), .ZN(n19253) );
  NAND2_X1 U22292 ( .A1(n19253), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19251) );
  OAI21_X1 U22293 ( .B1(n19253), .B2(n19252), .A(n19251), .ZN(P3_U3295) );
  AOI21_X1 U22294 ( .B1(n19255), .B2(n19254), .A(n19276), .ZN(n19256) );
  OAI21_X1 U22295 ( .B1(n19258), .B2(n19257), .A(n19256), .ZN(n19269) );
  OAI21_X1 U22296 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19260), .A(n19259), 
        .ZN(n19262) );
  AOI211_X1 U22297 ( .C1(n19275), .C2(n19262), .A(n19261), .B(n19273), .ZN(
        n19264) );
  NOR2_X1 U22298 ( .A1(n19264), .A2(n19263), .ZN(n19265) );
  OAI21_X1 U22299 ( .B1(n19266), .B2(n19265), .A(n19269), .ZN(n19267) );
  OAI21_X1 U22300 ( .B1(n19269), .B2(n19268), .A(n19267), .ZN(P3_U3296) );
  INV_X1 U22301 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19279) );
  INV_X1 U22302 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19271) );
  AOI22_X1 U22303 ( .A1(n19272), .A2(n19279), .B1(n19271), .B2(n19270), .ZN(
        P3_U3297) );
  AOI21_X1 U22304 ( .B1(n19274), .B2(n19273), .A(n19276), .ZN(n19280) );
  INV_X1 U22305 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19277) );
  AOI22_X1 U22306 ( .A1(n19280), .A2(n19277), .B1(n19276), .B2(n19275), .ZN(
        P3_U3298) );
  AOI21_X1 U22307 ( .B1(n19280), .B2(n19279), .A(n19278), .ZN(P3_U3299) );
  INV_X1 U22308 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19281) );
  NAND2_X1 U22309 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21283), .ZN(n20096) );
  AOI22_X1 U22310 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20096), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20089), .ZN(n20175) );
  INV_X1 U22311 ( .A(n20175), .ZN(n20088) );
  OAI21_X1 U22312 ( .B1(n20089), .B2(n19281), .A(n20088), .ZN(P2_U2815) );
  NAND2_X1 U22313 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20089), .ZN(n20241) );
  INV_X2 U22314 ( .A(n20241), .ZN(n20158) );
  AOI21_X1 U22315 ( .B1(n20089), .B2(n21283), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19282) );
  AOI22_X1 U22316 ( .A1(n20158), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19282), 
        .B2(n20241), .ZN(P2_U2817) );
  OAI21_X1 U22317 ( .B1(n20099), .B2(BS16), .A(n20175), .ZN(n20173) );
  OAI21_X1 U22318 ( .B1(n20175), .B2(n20227), .A(n20173), .ZN(P2_U2818) );
  NOR4_X1 U22319 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_10__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19292) );
  NOR4_X1 U22320 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19291) );
  AOI211_X1 U22321 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_3__SCAN_IN), .B(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19283) );
  INV_X1 U22322 ( .A(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(n21431) );
  INV_X1 U22323 ( .A(P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21482) );
  NAND3_X1 U22324 ( .A1(n19283), .A2(n21431), .A3(n21482), .ZN(n19289) );
  NOR4_X1 U22325 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19287) );
  NOR4_X1 U22326 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19286) );
  NOR4_X1 U22327 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19285) );
  NOR4_X1 U22328 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19284) );
  NAND4_X1 U22329 ( .A1(n19287), .A2(n19286), .A3(n19285), .A4(n19284), .ZN(
        n19288) );
  NOR4_X1 U22330 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(n19289), .A4(n19288), .ZN(n19290) );
  NAND3_X1 U22331 ( .A1(n19292), .A2(n19291), .A3(n19290), .ZN(n19299) );
  NOR2_X1 U22332 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19299), .ZN(n19293) );
  INV_X1 U22333 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20171) );
  AOI22_X1 U22334 ( .A1(n19293), .A2(n19294), .B1(n19299), .B2(n20171), .ZN(
        P2_U2820) );
  OR3_X1 U22335 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19298) );
  INV_X1 U22336 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20169) );
  AOI22_X1 U22337 ( .A1(n19293), .A2(n19298), .B1(n19299), .B2(n20169), .ZN(
        P2_U2821) );
  INV_X1 U22338 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20174) );
  NAND2_X1 U22339 ( .A1(n19293), .A2(n20174), .ZN(n19297) );
  INV_X1 U22340 ( .A(n19299), .ZN(n19300) );
  OAI21_X1 U22341 ( .B1(n20108), .B2(n19294), .A(n19300), .ZN(n19295) );
  OAI21_X1 U22342 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19300), .A(n19295), 
        .ZN(n19296) );
  OAI221_X1 U22343 ( .B1(n19297), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19297), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19296), .ZN(P2_U2822) );
  INV_X1 U22344 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20167) );
  OAI221_X1 U22345 ( .B1(n19300), .B2(n20167), .C1(n19299), .C2(n19298), .A(
        n19297), .ZN(P2_U2823) );
  INV_X1 U22346 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20145) );
  OAI22_X1 U22347 ( .A1(n19354), .A2(n10096), .B1(n19355), .B2(n20145), .ZN(
        n19301) );
  AOI21_X1 U22348 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19337), .A(
        n19301), .ZN(n19302) );
  OAI21_X1 U22349 ( .B1(n19303), .B2(n19356), .A(n19302), .ZN(n19304) );
  AOI21_X1 U22350 ( .B1(n19305), .B2(n19322), .A(n19304), .ZN(n19314) );
  NAND2_X1 U22351 ( .A1(n19307), .A2(n19306), .ZN(n19308) );
  AOI21_X1 U22352 ( .B1(n19308), .B2(n19344), .A(n19320), .ZN(n19309) );
  OAI22_X1 U22353 ( .A1(n19311), .A2(n19368), .B1(n19310), .B2(n19309), .ZN(
        n19312) );
  INV_X1 U22354 ( .A(n19312), .ZN(n19313) );
  NAND2_X1 U22355 ( .A1(n19314), .A2(n19313), .ZN(P2_U2834) );
  AOI22_X1 U22356 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19337), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19315), .ZN(n19332) );
  AOI21_X1 U22357 ( .B1(n19360), .B2(P2_EBX_REG_17__SCAN_IN), .A(n19359), .ZN(
        n19316) );
  OAI21_X1 U22358 ( .B1(n19317), .B2(n19356), .A(n19316), .ZN(n19318) );
  AOI21_X1 U22359 ( .B1(n19320), .B2(n19319), .A(n19318), .ZN(n19331) );
  INV_X1 U22360 ( .A(n19321), .ZN(n19325) );
  AOI22_X1 U22361 ( .A1(n19325), .A2(n19324), .B1(n19323), .B2(n19322), .ZN(
        n19330) );
  INV_X1 U22362 ( .A(n19343), .ZN(n19328) );
  OAI21_X1 U22363 ( .B1(n19328), .B2(n19327), .A(n19326), .ZN(n19329) );
  NAND4_X1 U22364 ( .A1(n19332), .A2(n19331), .A3(n19330), .A4(n19329), .ZN(
        P2_U2838) );
  INV_X1 U22365 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20136) );
  OAI21_X1 U22366 ( .B1(n19355), .B2(n20136), .A(n19333), .ZN(n19336) );
  NOR2_X1 U22367 ( .A1(n19334), .A2(n19356), .ZN(n19335) );
  AOI211_X1 U22368 ( .C1(n19337), .C2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19336), .B(n19335), .ZN(n19353) );
  NOR2_X1 U22369 ( .A1(n19340), .A2(n19338), .ZN(n19339) );
  MUX2_X1 U22370 ( .A(n19340), .B(n19339), .S(n11664), .Z(n19348) );
  INV_X1 U22371 ( .A(n19340), .ZN(n19342) );
  NAND3_X1 U22372 ( .A1(n11664), .A2(n19342), .A3(n19341), .ZN(n19345) );
  NAND3_X1 U22373 ( .A1(n19345), .A2(n19344), .A3(n19343), .ZN(n19347) );
  OAI22_X1 U22374 ( .A1(n19348), .A2(n19347), .B1(n19346), .B2(n19368), .ZN(
        n19351) );
  NOR2_X1 U22375 ( .A1(n19349), .A2(n19366), .ZN(n19350) );
  NOR2_X1 U22376 ( .A1(n19351), .A2(n19350), .ZN(n19352) );
  OAI211_X1 U22377 ( .C1(n11094), .C2(n19354), .A(n19353), .B(n19352), .ZN(
        P2_U2839) );
  INV_X1 U22378 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20117) );
  OAI22_X1 U22379 ( .A1(n19357), .A2(n19356), .B1(n20117), .B2(n19355), .ZN(
        n19358) );
  AOI211_X1 U22380 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19360), .A(n19359), .B(
        n19358), .ZN(n19374) );
  NAND2_X1 U22381 ( .A1(n19361), .A2(n19363), .ZN(n19362) );
  MUX2_X1 U22382 ( .A(n19363), .B(n19362), .S(n11664), .Z(n19372) );
  NOR2_X1 U22383 ( .A1(n19365), .A2(n19364), .ZN(n19371) );
  OAI22_X1 U22384 ( .A1(n19369), .A2(n19368), .B1(n19367), .B2(n19366), .ZN(
        n19370) );
  AOI21_X1 U22385 ( .B1(n19372), .B2(n19371), .A(n19370), .ZN(n19373) );
  OAI211_X1 U22386 ( .C1(n16259), .C2(n19375), .A(n19374), .B(n19373), .ZN(
        P2_U2849) );
  AOI22_X1 U22387 ( .A1(n19376), .A2(n19397), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19396), .ZN(n19381) );
  XOR2_X1 U22388 ( .A(n19378), .B(n19377), .Z(n19379) );
  NAND2_X1 U22389 ( .A1(n19379), .A2(n19398), .ZN(n19380) );
  OAI211_X1 U22390 ( .C1(n19382), .C2(n19403), .A(n19381), .B(n19380), .ZN(
        P2_U2915) );
  AOI22_X1 U22391 ( .A1(n20182), .A2(n19397), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19396), .ZN(n19388) );
  OAI21_X1 U22392 ( .B1(n19385), .B2(n19384), .A(n19383), .ZN(n19386) );
  NAND2_X1 U22393 ( .A1(n19386), .A2(n19398), .ZN(n19387) );
  OAI211_X1 U22394 ( .C1(n19389), .C2(n19403), .A(n19388), .B(n19387), .ZN(
        P2_U2916) );
  AOI22_X1 U22395 ( .A1(n19397), .A2(n20203), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19396), .ZN(n19394) );
  OAI21_X1 U22396 ( .B1(n19391), .B2(n19399), .A(n19390), .ZN(n19392) );
  NAND2_X1 U22397 ( .A1(n19392), .A2(n19398), .ZN(n19393) );
  OAI211_X1 U22398 ( .C1(n19395), .C2(n19403), .A(n19394), .B(n19393), .ZN(
        P2_U2918) );
  AOI22_X1 U22399 ( .A1(n19397), .A2(n19400), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19396), .ZN(n19402) );
  OAI211_X1 U22400 ( .C1(n20211), .C2(n19400), .A(n19399), .B(n19398), .ZN(
        n19401) );
  OAI211_X1 U22401 ( .C1(n19404), .C2(n19403), .A(n19402), .B(n19401), .ZN(
        P2_U2919) );
  INV_X1 U22402 ( .A(n19405), .ZN(n19407) );
  NAND2_X1 U22403 ( .A1(n19407), .A2(n19406), .ZN(n19409) );
  NOR2_X1 U22404 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19410), .ZN(n19460) );
  AND2_X1 U22405 ( .A1(n19435), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NAND2_X1 U22406 ( .A1(n19439), .A2(n19411), .ZN(n19437) );
  AOI22_X1 U22407 ( .A1(n20237), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n19467), .ZN(n19412) );
  OAI21_X1 U22408 ( .B1(n21272), .B2(n19437), .A(n19412), .ZN(P2_U2921) );
  INV_X1 U22409 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19414) );
  AOI22_X1 U22410 ( .A1(n20237), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19413) );
  OAI21_X1 U22411 ( .B1(n19414), .B2(n19437), .A(n19413), .ZN(P2_U2922) );
  INV_X1 U22412 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n21370) );
  AOI22_X1 U22413 ( .A1(n20237), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19415) );
  OAI21_X1 U22414 ( .B1(n21370), .B2(n19437), .A(n19415), .ZN(P2_U2923) );
  INV_X1 U22415 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19417) );
  AOI22_X1 U22416 ( .A1(n20237), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19416) );
  OAI21_X1 U22417 ( .B1(n19417), .B2(n19437), .A(n19416), .ZN(P2_U2924) );
  AOI22_X1 U22418 ( .A1(n20237), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19418) );
  OAI21_X1 U22419 ( .B1(n19419), .B2(n19437), .A(n19418), .ZN(P2_U2925) );
  INV_X1 U22420 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n21239) );
  AOI22_X1 U22421 ( .A1(n20237), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19420) );
  OAI21_X1 U22422 ( .B1(n21239), .B2(n19437), .A(n19420), .ZN(P2_U2926) );
  AOI22_X1 U22423 ( .A1(n20237), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19421) );
  OAI21_X1 U22424 ( .B1(n21340), .B2(n19437), .A(n19421), .ZN(P2_U2927) );
  INV_X1 U22425 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19423) );
  AOI22_X1 U22426 ( .A1(n20237), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19422) );
  OAI21_X1 U22427 ( .B1(n19423), .B2(n19437), .A(n19422), .ZN(P2_U2928) );
  INV_X1 U22428 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19425) );
  AOI22_X1 U22429 ( .A1(n20237), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19424) );
  OAI21_X1 U22430 ( .B1(n19425), .B2(n19437), .A(n19424), .ZN(P2_U2929) );
  INV_X1 U22431 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19427) );
  AOI22_X1 U22432 ( .A1(n20237), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19426) );
  OAI21_X1 U22433 ( .B1(n19427), .B2(n19437), .A(n19426), .ZN(P2_U2930) );
  AOI22_X1 U22434 ( .A1(n20237), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19428) );
  OAI21_X1 U22435 ( .B1(n19429), .B2(n19437), .A(n19428), .ZN(P2_U2931) );
  AOI22_X1 U22436 ( .A1(n20237), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19430) );
  OAI21_X1 U22437 ( .B1(n19431), .B2(n19437), .A(n19430), .ZN(P2_U2932) );
  INV_X1 U22438 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19433) );
  AOI22_X1 U22439 ( .A1(n20237), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19432) );
  OAI21_X1 U22440 ( .B1(n19433), .B2(n19437), .A(n19432), .ZN(P2_U2933) );
  AOI22_X1 U22441 ( .A1(n20237), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19434) );
  OAI21_X1 U22442 ( .B1(n21396), .B2(n19437), .A(n19434), .ZN(P2_U2934) );
  AOI22_X1 U22443 ( .A1(n20237), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19435), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19436) );
  OAI21_X1 U22444 ( .B1(n19438), .B2(n19437), .A(n19436), .ZN(P2_U2935) );
  AOI22_X1 U22445 ( .A1(n20237), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19440) );
  OAI21_X1 U22446 ( .B1(n13119), .B2(n19469), .A(n19440), .ZN(P2_U2936) );
  AOI22_X1 U22447 ( .A1(n20237), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19441) );
  OAI21_X1 U22448 ( .B1(n19442), .B2(n19469), .A(n19441), .ZN(P2_U2937) );
  AOI22_X1 U22449 ( .A1(n20237), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19443) );
  OAI21_X1 U22450 ( .B1(n19444), .B2(n19469), .A(n19443), .ZN(P2_U2938) );
  AOI22_X1 U22451 ( .A1(n19460), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19445) );
  OAI21_X1 U22452 ( .B1(n19446), .B2(n19469), .A(n19445), .ZN(P2_U2939) );
  AOI22_X1 U22453 ( .A1(n19460), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19447) );
  OAI21_X1 U22454 ( .B1(n19448), .B2(n19469), .A(n19447), .ZN(P2_U2940) );
  AOI22_X1 U22455 ( .A1(n19460), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19449) );
  OAI21_X1 U22456 ( .B1(n19450), .B2(n19469), .A(n19449), .ZN(P2_U2941) );
  AOI22_X1 U22457 ( .A1(n19460), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19451) );
  OAI21_X1 U22458 ( .B1(n21406), .B2(n19469), .A(n19451), .ZN(P2_U2942) );
  AOI22_X1 U22459 ( .A1(n19460), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19452) );
  OAI21_X1 U22460 ( .B1(n19453), .B2(n19469), .A(n19452), .ZN(P2_U2943) );
  AOI22_X1 U22461 ( .A1(n19460), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19454) );
  OAI21_X1 U22462 ( .B1(n19455), .B2(n19469), .A(n19454), .ZN(P2_U2944) );
  AOI22_X1 U22463 ( .A1(n19460), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19456) );
  OAI21_X1 U22464 ( .B1(n21457), .B2(n19469), .A(n19456), .ZN(P2_U2945) );
  AOI22_X1 U22465 ( .A1(n19460), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19457) );
  OAI21_X1 U22466 ( .B1(n16016), .B2(n19469), .A(n19457), .ZN(P2_U2946) );
  INV_X1 U22467 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19459) );
  AOI22_X1 U22468 ( .A1(n19460), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19458) );
  OAI21_X1 U22469 ( .B1(n19459), .B2(n19469), .A(n19458), .ZN(P2_U2947) );
  INV_X1 U22470 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19462) );
  AOI22_X1 U22471 ( .A1(n19460), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19461) );
  OAI21_X1 U22472 ( .B1(n19462), .B2(n19469), .A(n19461), .ZN(P2_U2948) );
  INV_X1 U22473 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19464) );
  AOI22_X1 U22474 ( .A1(n20237), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19463) );
  OAI21_X1 U22475 ( .B1(n19464), .B2(n19469), .A(n19463), .ZN(P2_U2949) );
  INV_X1 U22476 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19466) );
  AOI22_X1 U22477 ( .A1(n20237), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19465) );
  OAI21_X1 U22478 ( .B1(n19466), .B2(n19469), .A(n19465), .ZN(P2_U2950) );
  AOI22_X1 U22479 ( .A1(n20237), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19467), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19468) );
  OAI21_X1 U22480 ( .B1(n11393), .B2(n19469), .A(n19468), .ZN(P2_U2951) );
  AOI22_X1 U22481 ( .A1(n19471), .A2(n19470), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19483), .ZN(n19481) );
  NAND2_X1 U22482 ( .A1(n19472), .A2(n19484), .ZN(n19475) );
  INV_X1 U22483 ( .A(n19473), .ZN(n19474) );
  OAI211_X1 U22484 ( .C1(n19477), .C2(n19476), .A(n19475), .B(n19474), .ZN(
        n19478) );
  AOI21_X1 U22485 ( .B1(n19479), .B2(n19493), .A(n19478), .ZN(n19480) );
  NAND2_X1 U22486 ( .A1(n19481), .A2(n19480), .ZN(P2_U3012) );
  INV_X1 U22487 ( .A(n19482), .ZN(n19485) );
  AOI22_X1 U22488 ( .A1(n19485), .A2(n19484), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19483), .ZN(n19496) );
  NAND2_X1 U22489 ( .A1(n19487), .A2(n19486), .ZN(n19489) );
  OAI211_X1 U22490 ( .C1(n19491), .C2(n19490), .A(n19489), .B(n19488), .ZN(
        n19492) );
  AOI21_X1 U22491 ( .B1(n19494), .B2(n19493), .A(n19492), .ZN(n19495) );
  NAND2_X1 U22492 ( .A1(n19496), .A2(n19495), .ZN(P2_U3013) );
  AND2_X1 U22493 ( .A1(n20180), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20201) );
  AOI22_X2 U22494 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19546), .ZN(n20038) );
  OAI22_X2 U22495 ( .A1(n19500), .A2(n19539), .B1(n15948), .B2(n19538), .ZN(
        n20035) );
  NOR2_X2 U22496 ( .A1(n19549), .A2(n20229), .ZN(n20025) );
  NAND2_X1 U22497 ( .A1(n20188), .A2(n20196), .ZN(n19619) );
  OR2_X1 U22498 ( .A1(n19619), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19561) );
  NOR2_X1 U22499 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19561), .ZN(
        n19542) );
  AOI22_X1 U22500 ( .A1(n20035), .A2(n20082), .B1(n20025), .B2(n19542), .ZN(
        n19511) );
  AOI21_X1 U22501 ( .B1(n20075), .B2(n19576), .A(n20227), .ZN(n19503) );
  NOR2_X1 U22502 ( .A1(n19503), .A2(n20176), .ZN(n19507) );
  OAI21_X1 U22503 ( .B1(n10950), .B2(n20207), .A(n19977), .ZN(n19504) );
  AOI21_X1 U22504 ( .B1(n19507), .B2(n20030), .A(n19504), .ZN(n19505) );
  INV_X1 U22505 ( .A(n20030), .ZN(n20078) );
  OAI21_X1 U22506 ( .B1(n20078), .B2(n19542), .A(n19507), .ZN(n19509) );
  OAI21_X1 U22507 ( .B1(n10950), .B2(n19542), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19508) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19554), .B1(
        n20026), .B2(n19553), .ZN(n19510) );
  OAI211_X1 U22509 ( .C1(n20038), .C2(n19576), .A(n19511), .B(n19510), .ZN(
        P2_U3048) );
  AOI22_X1 U22510 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19546), .ZN(n19991) );
  NOR2_X2 U22511 ( .A1(n19549), .A2(n19513), .ZN(n20039) );
  INV_X1 U22512 ( .A(n20039), .ZN(n19818) );
  INV_X1 U22513 ( .A(n19542), .ZN(n19550) );
  OAI22_X1 U22514 ( .A1(n20075), .A2(n19991), .B1(n19818), .B2(n19550), .ZN(
        n19514) );
  INV_X1 U22515 ( .A(n19514), .ZN(n19517) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19554), .B1(
        n20040), .B2(n19553), .ZN(n19516) );
  OAI211_X1 U22517 ( .C1(n20044), .C2(n19576), .A(n19517), .B(n19516), .ZN(
        P2_U3049) );
  AOI22_X1 U22518 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19546), .ZN(n20050) );
  NOR2_X2 U22519 ( .A1(n19549), .A2(n19518), .ZN(n20045) );
  INV_X1 U22520 ( .A(n20045), .ZN(n19992) );
  OAI22_X1 U22521 ( .A1(n20075), .A2(n20050), .B1(n19992), .B2(n19550), .ZN(
        n19519) );
  INV_X1 U22522 ( .A(n19519), .ZN(n19522) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19554), .B1(
        n20046), .B2(n19553), .ZN(n19521) );
  OAI211_X1 U22524 ( .C1(n19996), .C2(n19576), .A(n19522), .B(n19521), .ZN(
        P2_U3050) );
  AOI22_X2 U22525 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19546), .ZN(n20001) );
  AOI22_X1 U22526 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19546), .ZN(n20056) );
  NOR2_X2 U22527 ( .A1(n19549), .A2(n10762), .ZN(n20051) );
  INV_X1 U22528 ( .A(n20051), .ZN(n19997) );
  OAI22_X1 U22529 ( .A1(n20075), .A2(n20056), .B1(n19997), .B2(n19550), .ZN(
        n19524) );
  INV_X1 U22530 ( .A(n19524), .ZN(n19527) );
  AND2_X1 U22531 ( .A1(n20033), .A2(n19525), .ZN(n20052) );
  AOI22_X1 U22532 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19554), .B1(
        n20052), .B2(n19553), .ZN(n19526) );
  OAI211_X1 U22533 ( .C1(n20001), .C2(n19576), .A(n19527), .B(n19526), .ZN(
        P2_U3051) );
  AOI22_X2 U22534 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19546), .ZN(n20062) );
  OAI22_X2 U22535 ( .A1(n19528), .A2(n19539), .B1(n15926), .B2(n19538), .ZN(
        n20059) );
  NOR2_X2 U22536 ( .A1(n19549), .A2(n19529), .ZN(n20057) );
  AOI22_X1 U22537 ( .A1(n20059), .A2(n20082), .B1(n20057), .B2(n19542), .ZN(
        n19532) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19554), .B1(
        n20058), .B2(n19553), .ZN(n19531) );
  OAI211_X1 U22539 ( .C1(n20062), .C2(n19576), .A(n19532), .B(n19531), .ZN(
        P2_U3052) );
  AOI22_X2 U22540 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19546), .ZN(n20068) );
  OAI22_X2 U22541 ( .A1(n19533), .A2(n19539), .B1(n15917), .B2(n19538), .ZN(
        n20065) );
  NOR2_X2 U22542 ( .A1(n19549), .A2(n19534), .ZN(n20063) );
  AOI22_X1 U22543 ( .A1(n20065), .A2(n20082), .B1(n20063), .B2(n19542), .ZN(
        n19537) );
  AND2_X1 U22544 ( .A1(n20033), .A2(n19535), .ZN(n20064) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19554), .B1(
        n20064), .B2(n19553), .ZN(n19536) );
  OAI211_X1 U22546 ( .C1(n20068), .C2(n19576), .A(n19537), .B(n19536), .ZN(
        P2_U3053) );
  AOI22_X2 U22547 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19546), .ZN(n20076) );
  OAI22_X2 U22548 ( .A1(n19540), .A2(n19539), .B1(n12431), .B2(n19538), .ZN(
        n20071) );
  NOR2_X2 U22549 ( .A1(n19549), .A2(n19541), .ZN(n20069) );
  AOI22_X1 U22550 ( .A1(n20071), .A2(n20082), .B1(n20069), .B2(n19542), .ZN(
        n19545) );
  AND2_X1 U22551 ( .A1(n20033), .A2(n19543), .ZN(n20070) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19554), .B1(
        n20070), .B2(n19553), .ZN(n19544) );
  OAI211_X1 U22553 ( .C1(n20076), .C2(n19576), .A(n19545), .B(n19544), .ZN(
        P2_U3054) );
  AOI22_X2 U22554 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19546), .ZN(n20015) );
  AOI22_X1 U22555 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19547), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19546), .ZN(n20087) );
  NOR2_X2 U22556 ( .A1(n19549), .A2(n19548), .ZN(n20077) );
  INV_X1 U22557 ( .A(n20077), .ZN(n20014) );
  OAI22_X1 U22558 ( .A1(n20075), .A2(n20087), .B1(n20014), .B2(n19550), .ZN(
        n19551) );
  INV_X1 U22559 ( .A(n19551), .ZN(n19556) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19554), .B1(
        n20079), .B2(n19553), .ZN(n19555) );
  OAI211_X1 U22561 ( .C1(n20015), .C2(n19576), .A(n19556), .B(n19555), .ZN(
        P2_U3055) );
  NOR2_X1 U22562 ( .A1(n19805), .A2(n19619), .ZN(n19581) );
  INV_X1 U22563 ( .A(n19581), .ZN(n19562) );
  AND2_X1 U22564 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19562), .ZN(n19558) );
  NAND2_X1 U22565 ( .A1(n19559), .A2(n19558), .ZN(n19564) );
  OAI21_X1 U22566 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19561), .A(n20207), 
        .ZN(n19560) );
  AOI22_X1 U22567 ( .A1(n19582), .A2(n20026), .B1(n20025), .B2(n19581), .ZN(
        n19567) );
  INV_X1 U22568 ( .A(n19748), .ZN(n19618) );
  OAI21_X1 U22569 ( .B1(n19618), .B2(n19808), .A(n19561), .ZN(n19565) );
  NAND2_X1 U22570 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19562), .ZN(n19563) );
  NAND4_X1 U22571 ( .A1(n19565), .A2(n20033), .A3(n19564), .A4(n19563), .ZN(
        n19584) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19584), .B1(
        n19583), .B2(n20035), .ZN(n19566) );
  OAI211_X1 U22573 ( .C1(n20038), .C2(n19587), .A(n19567), .B(n19566), .ZN(
        P2_U3056) );
  AOI22_X1 U22574 ( .A1(n19582), .A2(n20040), .B1(n20039), .B2(n19581), .ZN(
        n19569) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19584), .B1(
        n19583), .B2(n20041), .ZN(n19568) );
  OAI211_X1 U22576 ( .C1(n20044), .C2(n19587), .A(n19569), .B(n19568), .ZN(
        P2_U3057) );
  AOI22_X1 U22577 ( .A1(n19582), .A2(n20046), .B1(n20045), .B2(n19581), .ZN(
        n19571) );
  INV_X1 U22578 ( .A(n19996), .ZN(n20047) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19584), .B1(
        n19614), .B2(n20047), .ZN(n19570) );
  OAI211_X1 U22580 ( .C1(n20050), .C2(n19576), .A(n19571), .B(n19570), .ZN(
        P2_U3058) );
  AOI22_X1 U22581 ( .A1(n19582), .A2(n20052), .B1(n20051), .B2(n19581), .ZN(
        n19573) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19584), .B1(
        n19583), .B2(n19928), .ZN(n19572) );
  OAI211_X1 U22583 ( .C1(n20001), .C2(n19587), .A(n19573), .B(n19572), .ZN(
        P2_U3059) );
  INV_X1 U22584 ( .A(n20059), .ZN(n19832) );
  AOI22_X1 U22585 ( .A1(n19582), .A2(n20058), .B1(n20057), .B2(n19581), .ZN(
        n19575) );
  INV_X1 U22586 ( .A(n20062), .ZN(n19700) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19584), .B1(
        n19614), .B2(n19700), .ZN(n19574) );
  OAI211_X1 U22588 ( .C1(n19832), .C2(n19576), .A(n19575), .B(n19574), .ZN(
        P2_U3060) );
  AOI22_X1 U22589 ( .A1(n19582), .A2(n20064), .B1(n20063), .B2(n19581), .ZN(
        n19578) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19584), .B1(
        n19583), .B2(n20065), .ZN(n19577) );
  OAI211_X1 U22591 ( .C1(n20068), .C2(n19587), .A(n19578), .B(n19577), .ZN(
        P2_U3061) );
  AOI22_X1 U22592 ( .A1(n19582), .A2(n20070), .B1(n20069), .B2(n19581), .ZN(
        n19580) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19584), .B1(
        n19583), .B2(n20071), .ZN(n19579) );
  OAI211_X1 U22594 ( .C1(n20076), .C2(n19587), .A(n19580), .B(n19579), .ZN(
        P2_U3062) );
  AOI22_X1 U22595 ( .A1(n19582), .A2(n20079), .B1(n20077), .B2(n19581), .ZN(
        n19586) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19584), .B1(
        n19583), .B2(n19939), .ZN(n19585) );
  OAI211_X1 U22597 ( .C1(n20015), .C2(n19587), .A(n19586), .B(n19585), .ZN(
        P2_U3063) );
  INV_X1 U22598 ( .A(n19588), .ZN(n19593) );
  NOR2_X1 U22599 ( .A1(n19848), .A2(n19619), .ZN(n19612) );
  INV_X1 U22600 ( .A(n19612), .ZN(n19589) );
  AND2_X1 U22601 ( .A1(n19593), .A2(n19589), .ZN(n19592) );
  INV_X1 U22602 ( .A(n19850), .ZN(n19591) );
  INV_X1 U22603 ( .A(n19619), .ZN(n19590) );
  NAND2_X1 U22604 ( .A1(n19591), .A2(n19590), .ZN(n19594) );
  AOI22_X1 U22605 ( .A1(n19613), .A2(n20026), .B1(n20025), .B2(n19612), .ZN(
        n19599) );
  AOI21_X1 U22606 ( .B1(n19593), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19597) );
  OAI21_X1 U22607 ( .B1(n19614), .B2(n19641), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19595) );
  NAND3_X1 U22608 ( .A1(n19595), .A2(n20180), .A3(n19594), .ZN(n19596) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n20035), .ZN(n19598) );
  OAI211_X1 U22610 ( .C1(n20038), .C2(n19650), .A(n19599), .B(n19598), .ZN(
        P2_U3064) );
  AOI22_X1 U22611 ( .A1(n19613), .A2(n20040), .B1(n20039), .B2(n19612), .ZN(
        n19601) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n20041), .ZN(n19600) );
  OAI211_X1 U22613 ( .C1(n20044), .C2(n19650), .A(n19601), .B(n19600), .ZN(
        P2_U3065) );
  AOI22_X1 U22614 ( .A1(n19613), .A2(n20046), .B1(n20045), .B2(n19612), .ZN(
        n19603) );
  INV_X1 U22615 ( .A(n20050), .ZN(n19925) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19925), .ZN(n19602) );
  OAI211_X1 U22617 ( .C1(n19996), .C2(n19650), .A(n19603), .B(n19602), .ZN(
        P2_U3066) );
  AOI22_X1 U22618 ( .A1(n19613), .A2(n20052), .B1(n20051), .B2(n19612), .ZN(
        n19605) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19928), .ZN(n19604) );
  OAI211_X1 U22620 ( .C1(n20001), .C2(n19650), .A(n19605), .B(n19604), .ZN(
        P2_U3067) );
  AOI22_X1 U22621 ( .A1(n19613), .A2(n20058), .B1(n20057), .B2(n19612), .ZN(
        n19607) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n20059), .ZN(n19606) );
  OAI211_X1 U22623 ( .C1(n20062), .C2(n19650), .A(n19607), .B(n19606), .ZN(
        P2_U3068) );
  AOI22_X1 U22624 ( .A1(n19613), .A2(n20064), .B1(n20063), .B2(n19612), .ZN(
        n19609) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n20065), .ZN(n19608) );
  OAI211_X1 U22626 ( .C1(n20068), .C2(n19650), .A(n19609), .B(n19608), .ZN(
        P2_U3069) );
  AOI22_X1 U22627 ( .A1(n19613), .A2(n20070), .B1(n20069), .B2(n19612), .ZN(
        n19611) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n20071), .ZN(n19610) );
  OAI211_X1 U22629 ( .C1(n20076), .C2(n19650), .A(n19611), .B(n19610), .ZN(
        P2_U3070) );
  AOI22_X1 U22630 ( .A1(n19613), .A2(n20079), .B1(n20077), .B2(n19612), .ZN(
        n19617) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19615), .B1(
        n19614), .B2(n19939), .ZN(n19616) );
  OAI211_X1 U22632 ( .C1(n20015), .C2(n19650), .A(n19617), .B(n19616), .ZN(
        P2_U3071) );
  NOR2_X1 U22633 ( .A1(n19743), .A2(n19619), .ZN(n19645) );
  AOI22_X1 U22634 ( .A1(n20035), .A2(n19641), .B1(n19645), .B2(n20025), .ZN(
        n19630) );
  NOR2_X1 U22635 ( .A1(n20205), .A2(n19619), .ZN(n19624) );
  INV_X1 U22636 ( .A(n19620), .ZN(n19625) );
  OAI21_X1 U22637 ( .B1(n19625), .B2(n20207), .A(n19977), .ZN(n19622) );
  INV_X1 U22638 ( .A(n19645), .ZN(n19621) );
  AOI21_X1 U22639 ( .B1(n19622), .B2(n19621), .A(n19978), .ZN(n19623) );
  INV_X1 U22640 ( .A(n19624), .ZN(n19627) );
  OAI21_X1 U22641 ( .B1(n19625), .B2(n19645), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19626) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19647), .B1(
        n20026), .B2(n19646), .ZN(n19629) );
  OAI211_X1 U22643 ( .C1(n20038), .C2(n19644), .A(n19630), .B(n19629), .ZN(
        P2_U3072) );
  AOI22_X1 U22644 ( .A1(n19988), .A2(n19676), .B1(n19645), .B2(n20039), .ZN(
        n19632) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19647), .B1(
        n20040), .B2(n19646), .ZN(n19631) );
  OAI211_X1 U22646 ( .C1(n19991), .C2(n19650), .A(n19632), .B(n19631), .ZN(
        P2_U3073) );
  AOI22_X1 U22647 ( .A1(n19676), .A2(n20047), .B1(n19645), .B2(n20045), .ZN(
        n19634) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19647), .B1(
        n20046), .B2(n19646), .ZN(n19633) );
  OAI211_X1 U22649 ( .C1(n20050), .C2(n19650), .A(n19634), .B(n19633), .ZN(
        P2_U3074) );
  INV_X1 U22650 ( .A(n20001), .ZN(n20053) );
  AOI22_X1 U22651 ( .A1(n19676), .A2(n20053), .B1(n19645), .B2(n20051), .ZN(
        n19636) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19647), .B1(
        n20052), .B2(n19646), .ZN(n19635) );
  OAI211_X1 U22653 ( .C1(n20056), .C2(n19650), .A(n19636), .B(n19635), .ZN(
        P2_U3075) );
  AOI22_X1 U22654 ( .A1(n20059), .A2(n19641), .B1(n19645), .B2(n20057), .ZN(
        n19638) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19647), .B1(
        n20058), .B2(n19646), .ZN(n19637) );
  OAI211_X1 U22656 ( .C1(n20062), .C2(n19644), .A(n19638), .B(n19637), .ZN(
        P2_U3076) );
  AOI22_X1 U22657 ( .A1(n20065), .A2(n19641), .B1(n19645), .B2(n20063), .ZN(
        n19640) );
  AOI22_X1 U22658 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19647), .B1(
        n20064), .B2(n19646), .ZN(n19639) );
  OAI211_X1 U22659 ( .C1(n20068), .C2(n19644), .A(n19640), .B(n19639), .ZN(
        P2_U3077) );
  AOI22_X1 U22660 ( .A1(n20071), .A2(n19641), .B1(n19645), .B2(n20069), .ZN(
        n19643) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19647), .B1(
        n20070), .B2(n19646), .ZN(n19642) );
  OAI211_X1 U22662 ( .C1(n20076), .C2(n19644), .A(n19643), .B(n19642), .ZN(
        P2_U3078) );
  INV_X1 U22663 ( .A(n20015), .ZN(n20081) );
  AOI22_X1 U22664 ( .A1(n19676), .A2(n20081), .B1(n19645), .B2(n20077), .ZN(
        n19649) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19647), .B1(
        n20079), .B2(n19646), .ZN(n19648) );
  OAI211_X1 U22666 ( .C1(n20087), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P2_U3079) );
  NOR2_X1 U22667 ( .A1(n19652), .A2(n19651), .ZN(n19914) );
  NAND2_X1 U22668 ( .A1(n19914), .A2(n20188), .ZN(n19657) );
  NAND2_X1 U22669 ( .A1(n20188), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19744) );
  OR2_X1 U22670 ( .A1(n19744), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19688) );
  NOR2_X1 U22671 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19688), .ZN(
        n19674) );
  OAI21_X1 U22672 ( .B1(n19654), .B2(n19674), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19653) );
  OAI21_X1 U22673 ( .B1(n19657), .B2(n20176), .A(n19653), .ZN(n19675) );
  AOI22_X1 U22674 ( .A1(n19675), .A2(n20026), .B1(n20025), .B2(n19674), .ZN(
        n19661) );
  INV_X1 U22675 ( .A(n19654), .ZN(n19655) );
  AOI21_X1 U22676 ( .B1(n19655), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19659) );
  OAI21_X1 U22677 ( .B1(n19676), .B2(n19709), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19656) );
  NAND2_X1 U22678 ( .A1(n19657), .A2(n19656), .ZN(n19658) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19677), .B1(
        n19676), .B2(n20035), .ZN(n19660) );
  OAI211_X1 U22680 ( .C1(n20038), .C2(n19697), .A(n19661), .B(n19660), .ZN(
        P2_U3080) );
  AOI22_X1 U22681 ( .A1(n19675), .A2(n20040), .B1(n20039), .B2(n19674), .ZN(
        n19663) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19677), .B1(
        n19676), .B2(n20041), .ZN(n19662) );
  OAI211_X1 U22683 ( .C1(n20044), .C2(n19697), .A(n19663), .B(n19662), .ZN(
        P2_U3081) );
  AOI22_X1 U22684 ( .A1(n19675), .A2(n20046), .B1(n20045), .B2(n19674), .ZN(
        n19665) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19677), .B1(
        n19676), .B2(n19925), .ZN(n19664) );
  OAI211_X1 U22686 ( .C1(n19996), .C2(n19697), .A(n19665), .B(n19664), .ZN(
        P2_U3082) );
  AOI22_X1 U22687 ( .A1(n19675), .A2(n20052), .B1(n20051), .B2(n19674), .ZN(
        n19667) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19677), .B1(
        n19676), .B2(n19928), .ZN(n19666) );
  OAI211_X1 U22689 ( .C1(n20001), .C2(n19697), .A(n19667), .B(n19666), .ZN(
        P2_U3083) );
  AOI22_X1 U22690 ( .A1(n19675), .A2(n20058), .B1(n20057), .B2(n19674), .ZN(
        n19669) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19677), .B1(
        n19676), .B2(n20059), .ZN(n19668) );
  OAI211_X1 U22692 ( .C1(n20062), .C2(n19697), .A(n19669), .B(n19668), .ZN(
        P2_U3084) );
  AOI22_X1 U22693 ( .A1(n19675), .A2(n20064), .B1(n20063), .B2(n19674), .ZN(
        n19671) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19677), .B1(
        n19676), .B2(n20065), .ZN(n19670) );
  OAI211_X1 U22695 ( .C1(n20068), .C2(n19697), .A(n19671), .B(n19670), .ZN(
        P2_U3085) );
  AOI22_X1 U22696 ( .A1(n19675), .A2(n20070), .B1(n20069), .B2(n19674), .ZN(
        n19673) );
  AOI22_X1 U22697 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19677), .B1(
        n19676), .B2(n20071), .ZN(n19672) );
  OAI211_X1 U22698 ( .C1(n20076), .C2(n19697), .A(n19673), .B(n19672), .ZN(
        P2_U3086) );
  AOI22_X1 U22699 ( .A1(n19675), .A2(n20079), .B1(n20077), .B2(n19674), .ZN(
        n19679) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19677), .B1(
        n19676), .B2(n19939), .ZN(n19678) );
  OAI211_X1 U22701 ( .C1(n20015), .C2(n19697), .A(n19679), .B(n19678), .ZN(
        P2_U3087) );
  AOI21_X1 U22702 ( .B1(n19748), .B2(n19912), .A(n20176), .ZN(n19685) );
  NAND2_X1 U22703 ( .A1(n19685), .A2(n19688), .ZN(n19683) );
  NAND2_X1 U22704 ( .A1(n19686), .A2(n19977), .ZN(n19681) );
  NOR2_X1 U22705 ( .A1(n19805), .A2(n19744), .ZN(n19718) );
  NOR2_X1 U22706 ( .A1(n20180), .A2(n19718), .ZN(n19680) );
  AOI21_X1 U22707 ( .B1(n19681), .B2(n19680), .A(n19978), .ZN(n19682) );
  INV_X1 U22708 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19692) );
  INV_X1 U22709 ( .A(n20038), .ZN(n19684) );
  AOI22_X1 U22710 ( .A1(n19738), .A2(n19684), .B1(n20025), .B2(n19718), .ZN(
        n19691) );
  INV_X1 U22711 ( .A(n19685), .ZN(n19689) );
  OAI21_X1 U22712 ( .B1(n19686), .B2(n19718), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19687) );
  AOI22_X1 U22713 ( .A1(n20026), .A2(n19710), .B1(n19709), .B2(n20035), .ZN(
        n19690) );
  OAI211_X1 U22714 ( .C1(n19704), .C2(n19692), .A(n19691), .B(n19690), .ZN(
        P2_U3088) );
  AOI22_X1 U22715 ( .A1(n19709), .A2(n20041), .B1(n20039), .B2(n19718), .ZN(
        n19694) );
  AOI22_X1 U22716 ( .A1(n20040), .A2(n19710), .B1(n19738), .B2(n19988), .ZN(
        n19693) );
  OAI211_X1 U22717 ( .C1(n19704), .C2(n10877), .A(n19694), .B(n19693), .ZN(
        P2_U3089) );
  AOI22_X1 U22718 ( .A1(n19738), .A2(n20047), .B1(n20045), .B2(n19718), .ZN(
        n19696) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19711), .B1(
        n20046), .B2(n19710), .ZN(n19695) );
  OAI211_X1 U22720 ( .C1(n20050), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        P2_U3090) );
  INV_X1 U22721 ( .A(n19738), .ZN(n19714) );
  AOI22_X1 U22722 ( .A1(n19709), .A2(n19928), .B1(n19718), .B2(n20051), .ZN(
        n19699) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19711), .B1(
        n20052), .B2(n19710), .ZN(n19698) );
  OAI211_X1 U22724 ( .C1(n20001), .C2(n19714), .A(n19699), .B(n19698), .ZN(
        P2_U3091) );
  INV_X1 U22725 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19703) );
  AOI22_X1 U22726 ( .A1(n19738), .A2(n19700), .B1(n19718), .B2(n20057), .ZN(
        n19702) );
  AOI22_X1 U22727 ( .A1(n20058), .A2(n19710), .B1(n19709), .B2(n20059), .ZN(
        n19701) );
  OAI211_X1 U22728 ( .C1(n19704), .C2(n19703), .A(n19702), .B(n19701), .ZN(
        P2_U3092) );
  AOI22_X1 U22729 ( .A1(n20065), .A2(n19709), .B1(n20063), .B2(n19718), .ZN(
        n19706) );
  AOI22_X1 U22730 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19711), .B1(
        n20064), .B2(n19710), .ZN(n19705) );
  OAI211_X1 U22731 ( .C1(n20068), .C2(n19714), .A(n19706), .B(n19705), .ZN(
        P2_U3093) );
  AOI22_X1 U22732 ( .A1(n20071), .A2(n19709), .B1(n20069), .B2(n19718), .ZN(
        n19708) );
  AOI22_X1 U22733 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19711), .B1(
        n20070), .B2(n19710), .ZN(n19707) );
  OAI211_X1 U22734 ( .C1(n20076), .C2(n19714), .A(n19708), .B(n19707), .ZN(
        P2_U3094) );
  AOI22_X1 U22735 ( .A1(n19709), .A2(n19939), .B1(n20077), .B2(n19718), .ZN(
        n19713) );
  AOI22_X1 U22736 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19711), .B1(
        n20079), .B2(n19710), .ZN(n19712) );
  OAI211_X1 U22737 ( .C1(n20015), .C2(n19714), .A(n19713), .B(n19712), .ZN(
        P2_U3095) );
  INV_X1 U22738 ( .A(n20028), .ZN(n19747) );
  NOR2_X1 U22739 ( .A1(n19848), .A2(n19744), .ZN(n19736) );
  OAI21_X1 U22740 ( .B1(n19717), .B2(n19736), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19716) );
  OAI21_X1 U22741 ( .B1(n19744), .B2(n19850), .A(n19716), .ZN(n19737) );
  AOI22_X1 U22742 ( .A1(n19737), .A2(n20026), .B1(n20025), .B2(n19736), .ZN(
        n19723) );
  INV_X1 U22743 ( .A(n19717), .ZN(n19720) );
  AOI221_X1 U22744 ( .B1(n19738), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19769), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19718), .ZN(n19719) );
  AOI211_X1 U22745 ( .C1(n19720), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19719), .ZN(n19721) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19739), .B1(
        n19738), .B2(n20035), .ZN(n19722) );
  OAI211_X1 U22747 ( .C1(n20038), .C2(n19767), .A(n19723), .B(n19722), .ZN(
        P2_U3096) );
  AOI22_X1 U22748 ( .A1(n19737), .A2(n20040), .B1(n20039), .B2(n19736), .ZN(
        n19725) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19739), .B1(
        n19738), .B2(n20041), .ZN(n19724) );
  OAI211_X1 U22750 ( .C1(n20044), .C2(n19767), .A(n19725), .B(n19724), .ZN(
        P2_U3097) );
  AOI22_X1 U22751 ( .A1(n19737), .A2(n20046), .B1(n20045), .B2(n19736), .ZN(
        n19727) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19739), .B1(
        n19738), .B2(n19925), .ZN(n19726) );
  OAI211_X1 U22753 ( .C1(n19996), .C2(n19767), .A(n19727), .B(n19726), .ZN(
        P2_U3098) );
  AOI22_X1 U22754 ( .A1(n19737), .A2(n20052), .B1(n20051), .B2(n19736), .ZN(
        n19729) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19739), .B1(
        n19738), .B2(n19928), .ZN(n19728) );
  OAI211_X1 U22756 ( .C1(n20001), .C2(n19767), .A(n19729), .B(n19728), .ZN(
        P2_U3099) );
  AOI22_X1 U22757 ( .A1(n19737), .A2(n20058), .B1(n20057), .B2(n19736), .ZN(
        n19731) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19739), .B1(
        n19738), .B2(n20059), .ZN(n19730) );
  OAI211_X1 U22759 ( .C1(n20062), .C2(n19767), .A(n19731), .B(n19730), .ZN(
        P2_U3100) );
  AOI22_X1 U22760 ( .A1(n19737), .A2(n20064), .B1(n20063), .B2(n19736), .ZN(
        n19733) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19739), .B1(
        n19738), .B2(n20065), .ZN(n19732) );
  OAI211_X1 U22762 ( .C1(n20068), .C2(n19767), .A(n19733), .B(n19732), .ZN(
        P2_U3101) );
  AOI22_X1 U22763 ( .A1(n19737), .A2(n20070), .B1(n20069), .B2(n19736), .ZN(
        n19735) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19739), .B1(
        n19738), .B2(n20071), .ZN(n19734) );
  OAI211_X1 U22765 ( .C1(n20076), .C2(n19767), .A(n19735), .B(n19734), .ZN(
        P2_U3102) );
  AOI22_X1 U22766 ( .A1(n19737), .A2(n20079), .B1(n20077), .B2(n19736), .ZN(
        n19741) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19739), .B1(
        n19738), .B2(n19939), .ZN(n19740) );
  OAI211_X1 U22768 ( .C1(n20015), .C2(n19767), .A(n19741), .B(n19740), .ZN(
        P2_U3103) );
  NAND2_X1 U22769 ( .A1(n19975), .A2(n20188), .ZN(n19749) );
  INV_X1 U22770 ( .A(n19743), .ZN(n19877) );
  INV_X1 U22771 ( .A(n19744), .ZN(n19745) );
  NAND2_X1 U22772 ( .A1(n19877), .A2(n19745), .ZN(n19775) );
  INV_X1 U22773 ( .A(n19775), .ZN(n19778) );
  OAI21_X1 U22774 ( .B1(n19752), .B2(n19778), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19746) );
  OAI21_X1 U22775 ( .B1(n19749), .B2(n20176), .A(n19746), .ZN(n19768) );
  AOI22_X1 U22776 ( .A1(n19768), .A2(n20026), .B1(n19778), .B2(n20025), .ZN(
        n19754) );
  NAND2_X1 U22777 ( .A1(n19775), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19751) );
  NAND2_X1 U22778 ( .A1(n19748), .A2(n19747), .ZN(n20177) );
  AOI22_X1 U22779 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19775), .B1(n20177), 
        .B2(n19749), .ZN(n19750) );
  OAI211_X1 U22780 ( .C1(n19752), .C2(n19751), .A(n20033), .B(n19750), .ZN(
        n19770) );
  AOI22_X1 U22781 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n20035), .ZN(n19753) );
  OAI211_X1 U22782 ( .C1(n20038), .C2(n19804), .A(n19754), .B(n19753), .ZN(
        P2_U3104) );
  AOI22_X1 U22783 ( .A1(n19768), .A2(n20040), .B1(n19778), .B2(n20039), .ZN(
        n19756) );
  AOI22_X1 U22784 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19770), .B1(
        n19794), .B2(n19988), .ZN(n19755) );
  OAI211_X1 U22785 ( .C1(n19991), .C2(n19767), .A(n19756), .B(n19755), .ZN(
        P2_U3105) );
  AOI22_X1 U22786 ( .A1(n19768), .A2(n20046), .B1(n19778), .B2(n20045), .ZN(
        n19758) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19925), .ZN(n19757) );
  OAI211_X1 U22788 ( .C1(n19996), .C2(n19804), .A(n19758), .B(n19757), .ZN(
        P2_U3106) );
  AOI22_X1 U22789 ( .A1(n19768), .A2(n20052), .B1(n19778), .B2(n20051), .ZN(
        n19760) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19928), .ZN(n19759) );
  OAI211_X1 U22791 ( .C1(n20001), .C2(n19804), .A(n19760), .B(n19759), .ZN(
        P2_U3107) );
  AOI22_X1 U22792 ( .A1(n19768), .A2(n20058), .B1(n19778), .B2(n20057), .ZN(
        n19762) );
  AOI22_X1 U22793 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n20059), .ZN(n19761) );
  OAI211_X1 U22794 ( .C1(n20062), .C2(n19804), .A(n19762), .B(n19761), .ZN(
        P2_U3108) );
  INV_X1 U22795 ( .A(n20065), .ZN(n20008) );
  AOI22_X1 U22796 ( .A1(n19768), .A2(n20064), .B1(n19778), .B2(n20063), .ZN(
        n19764) );
  INV_X1 U22797 ( .A(n20068), .ZN(n19897) );
  AOI22_X1 U22798 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19770), .B1(
        n19794), .B2(n19897), .ZN(n19763) );
  OAI211_X1 U22799 ( .C1(n20008), .C2(n19767), .A(n19764), .B(n19763), .ZN(
        P2_U3109) );
  INV_X1 U22800 ( .A(n20071), .ZN(n19904) );
  AOI22_X1 U22801 ( .A1(n19768), .A2(n20070), .B1(n19778), .B2(n20069), .ZN(
        n19766) );
  INV_X1 U22802 ( .A(n20076), .ZN(n19900) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19770), .B1(
        n19794), .B2(n19900), .ZN(n19765) );
  OAI211_X1 U22804 ( .C1(n19904), .C2(n19767), .A(n19766), .B(n19765), .ZN(
        P2_U3110) );
  AOI22_X1 U22805 ( .A1(n19768), .A2(n20079), .B1(n19778), .B2(n20077), .ZN(
        n19772) );
  AOI22_X1 U22806 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19770), .B1(
        n19769), .B2(n19939), .ZN(n19771) );
  OAI211_X1 U22807 ( .C1(n20015), .C2(n19804), .A(n19772), .B(n19771), .ZN(
        P2_U3111) );
  NAND2_X1 U22808 ( .A1(n20196), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19881) );
  NOR2_X1 U22809 ( .A1(n19881), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19810) );
  INV_X1 U22810 ( .A(n19810), .ZN(n19814) );
  NOR2_X1 U22811 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19814), .ZN(
        n19797) );
  AOI22_X1 U22812 ( .A1(n20035), .A2(n19794), .B1(n19797), .B2(n20025), .ZN(
        n19783) );
  AOI21_X1 U22813 ( .B1(n19804), .B2(n19842), .A(n20227), .ZN(n19773) );
  NOR2_X1 U22814 ( .A1(n19773), .A2(n20176), .ZN(n19777) );
  OAI21_X1 U22815 ( .B1(n19779), .B2(n20207), .A(n19977), .ZN(n19774) );
  AOI21_X1 U22816 ( .B1(n19777), .B2(n19775), .A(n19774), .ZN(n19776) );
  OAI21_X1 U22817 ( .B1(n19797), .B2(n19778), .A(n19777), .ZN(n19781) );
  OAI21_X1 U22818 ( .B1(n19779), .B2(n19797), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19780) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19801), .B1(
        n20026), .B2(n19800), .ZN(n19782) );
  OAI211_X1 U22820 ( .C1(n20038), .C2(n19842), .A(n19783), .B(n19782), .ZN(
        P2_U3112) );
  INV_X1 U22821 ( .A(n19842), .ZN(n19806) );
  AOI22_X1 U22822 ( .A1(n19988), .A2(n19806), .B1(n20039), .B2(n19797), .ZN(
        n19785) );
  AOI22_X1 U22823 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19801), .B1(
        n19800), .B2(n20040), .ZN(n19784) );
  OAI211_X1 U22824 ( .C1(n19991), .C2(n19804), .A(n19785), .B(n19784), .ZN(
        P2_U3113) );
  AOI22_X1 U22825 ( .A1(n19794), .A2(n19925), .B1(n19797), .B2(n20045), .ZN(
        n19787) );
  AOI22_X1 U22826 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19801), .B1(
        n19800), .B2(n20046), .ZN(n19786) );
  OAI211_X1 U22827 ( .C1(n19996), .C2(n19842), .A(n19787), .B(n19786), .ZN(
        P2_U3114) );
  AOI22_X1 U22828 ( .A1(n19794), .A2(n19928), .B1(n19797), .B2(n20051), .ZN(
        n19789) );
  AOI22_X1 U22829 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19801), .B1(
        n19800), .B2(n20052), .ZN(n19788) );
  OAI211_X1 U22830 ( .C1(n20001), .C2(n19842), .A(n19789), .B(n19788), .ZN(
        P2_U3115) );
  AOI22_X1 U22831 ( .A1(n20059), .A2(n19794), .B1(n20057), .B2(n19797), .ZN(
        n19791) );
  AOI22_X1 U22832 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19801), .B1(
        n19800), .B2(n20058), .ZN(n19790) );
  OAI211_X1 U22833 ( .C1(n20062), .C2(n19842), .A(n19791), .B(n19790), .ZN(
        P2_U3116) );
  AOI22_X1 U22834 ( .A1(n20065), .A2(n19794), .B1(n20063), .B2(n19797), .ZN(
        n19793) );
  AOI22_X1 U22835 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19801), .B1(
        n19800), .B2(n20064), .ZN(n19792) );
  OAI211_X1 U22836 ( .C1(n20068), .C2(n19842), .A(n19793), .B(n19792), .ZN(
        P2_U3117) );
  AOI22_X1 U22837 ( .A1(n20071), .A2(n19794), .B1(n20069), .B2(n19797), .ZN(
        n19796) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19801), .B1(
        n19800), .B2(n20070), .ZN(n19795) );
  OAI211_X1 U22839 ( .C1(n20076), .C2(n19842), .A(n19796), .B(n19795), .ZN(
        P2_U3118) );
  INV_X1 U22840 ( .A(n19797), .ZN(n19798) );
  OAI22_X1 U22841 ( .A1(n19842), .A2(n20015), .B1(n19798), .B2(n20014), .ZN(
        n19799) );
  INV_X1 U22842 ( .A(n19799), .ZN(n19803) );
  AOI22_X1 U22843 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19801), .B1(
        n19800), .B2(n20079), .ZN(n19802) );
  OAI211_X1 U22844 ( .C1(n20087), .C2(n19804), .A(n19803), .B(n19802), .ZN(
        P2_U3119) );
  NOR2_X1 U22845 ( .A1(n19805), .A2(n19881), .ZN(n19852) );
  AOI22_X1 U22846 ( .A1(n20035), .A2(n19806), .B1(n19852), .B2(n20025), .ZN(
        n19817) );
  INV_X1 U22847 ( .A(n19807), .ZN(n20184) );
  OAI21_X1 U22848 ( .B1(n20029), .B2(n19808), .A(n20180), .ZN(n19815) );
  INV_X1 U22849 ( .A(n19852), .ZN(n19841) );
  OAI211_X1 U22850 ( .C1(n19811), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19841), 
        .B(n20176), .ZN(n19809) );
  INV_X1 U22851 ( .A(n19811), .ZN(n19812) );
  OAI21_X1 U22852 ( .B1(n19812), .B2(n19852), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19813) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19845), .B1(
        n20026), .B2(n19844), .ZN(n19816) );
  OAI211_X1 U22854 ( .C1(n20038), .C2(n19837), .A(n19817), .B(n19816), .ZN(
        P2_U3120) );
  OAI22_X1 U22855 ( .A1(n19842), .A2(n19991), .B1(n19841), .B2(n19818), .ZN(
        n19819) );
  INV_X1 U22856 ( .A(n19819), .ZN(n19821) );
  AOI22_X1 U22857 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19845), .B1(
        n20040), .B2(n19844), .ZN(n19820) );
  OAI211_X1 U22858 ( .C1(n20044), .C2(n19837), .A(n19821), .B(n19820), .ZN(
        P2_U3121) );
  OAI22_X1 U22859 ( .A1(n19842), .A2(n20050), .B1(n19841), .B2(n19992), .ZN(
        n19822) );
  INV_X1 U22860 ( .A(n19822), .ZN(n19824) );
  AOI22_X1 U22861 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19845), .B1(
        n20046), .B2(n19844), .ZN(n19823) );
  OAI211_X1 U22862 ( .C1(n19996), .C2(n19837), .A(n19824), .B(n19823), .ZN(
        P2_U3122) );
  OAI22_X1 U22863 ( .A1(n19842), .A2(n20056), .B1(n19841), .B2(n19997), .ZN(
        n19825) );
  INV_X1 U22864 ( .A(n19825), .ZN(n19827) );
  AOI22_X1 U22865 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19845), .B1(
        n20052), .B2(n19844), .ZN(n19826) );
  OAI211_X1 U22866 ( .C1(n20001), .C2(n19837), .A(n19827), .B(n19826), .ZN(
        P2_U3123) );
  INV_X1 U22867 ( .A(n20057), .ZN(n19828) );
  OAI22_X1 U22868 ( .A1(n19837), .A2(n20062), .B1(n19828), .B2(n19841), .ZN(
        n19829) );
  INV_X1 U22869 ( .A(n19829), .ZN(n19831) );
  AOI22_X1 U22870 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19845), .B1(
        n20058), .B2(n19844), .ZN(n19830) );
  OAI211_X1 U22871 ( .C1(n19832), .C2(n19842), .A(n19831), .B(n19830), .ZN(
        P2_U3124) );
  INV_X1 U22872 ( .A(n20063), .ZN(n20004) );
  OAI22_X1 U22873 ( .A1(n19837), .A2(n20068), .B1(n19841), .B2(n20004), .ZN(
        n19833) );
  INV_X1 U22874 ( .A(n19833), .ZN(n19835) );
  AOI22_X1 U22875 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19845), .B1(
        n20064), .B2(n19844), .ZN(n19834) );
  OAI211_X1 U22876 ( .C1(n20008), .C2(n19842), .A(n19835), .B(n19834), .ZN(
        P2_U3125) );
  INV_X1 U22877 ( .A(n20069), .ZN(n19836) );
  OAI22_X1 U22878 ( .A1(n19837), .A2(n20076), .B1(n19841), .B2(n19836), .ZN(
        n19838) );
  INV_X1 U22879 ( .A(n19838), .ZN(n19840) );
  AOI22_X1 U22880 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19845), .B1(
        n20070), .B2(n19844), .ZN(n19839) );
  OAI211_X1 U22881 ( .C1(n19904), .C2(n19842), .A(n19840), .B(n19839), .ZN(
        P2_U3126) );
  OAI22_X1 U22882 ( .A1(n19842), .A2(n20087), .B1(n19841), .B2(n20014), .ZN(
        n19843) );
  INV_X1 U22883 ( .A(n19843), .ZN(n19847) );
  AOI22_X1 U22884 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19845), .B1(
        n20079), .B2(n19844), .ZN(n19846) );
  OAI211_X1 U22885 ( .C1(n20015), .C2(n19837), .A(n19847), .B(n19846), .ZN(
        P2_U3127) );
  NOR2_X1 U22886 ( .A1(n19848), .A2(n19881), .ZN(n19870) );
  OAI21_X1 U22887 ( .B1(n19851), .B2(n19870), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19849) );
  AOI22_X1 U22888 ( .A1(n19871), .A2(n20026), .B1(n20025), .B2(n19870), .ZN(
        n19857) );
  INV_X1 U22889 ( .A(n19851), .ZN(n19854) );
  AOI221_X1 U22890 ( .B1(n19907), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19872), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19852), .ZN(n19853) );
  AOI211_X1 U22891 ( .C1(n19854), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19853), .ZN(n19855) );
  OAI21_X2 U22892 ( .B1(n19855), .B2(n19870), .A(n20033), .ZN(n19873) );
  AOI22_X1 U22893 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19873), .B1(
        n19872), .B2(n20035), .ZN(n19856) );
  OAI211_X1 U22894 ( .C1(n20038), .C2(n19903), .A(n19857), .B(n19856), .ZN(
        P2_U3128) );
  AOI22_X1 U22895 ( .A1(n19871), .A2(n20040), .B1(n20039), .B2(n19870), .ZN(
        n19859) );
  AOI22_X1 U22896 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19873), .B1(
        n19872), .B2(n20041), .ZN(n19858) );
  OAI211_X1 U22897 ( .C1(n20044), .C2(n19903), .A(n19859), .B(n19858), .ZN(
        P2_U3129) );
  AOI22_X1 U22898 ( .A1(n19871), .A2(n20046), .B1(n20045), .B2(n19870), .ZN(
        n19861) );
  AOI22_X1 U22899 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19873), .B1(
        n19872), .B2(n19925), .ZN(n19860) );
  OAI211_X1 U22900 ( .C1(n19996), .C2(n19903), .A(n19861), .B(n19860), .ZN(
        P2_U3130) );
  AOI22_X1 U22901 ( .A1(n19871), .A2(n20052), .B1(n20051), .B2(n19870), .ZN(
        n19863) );
  AOI22_X1 U22902 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19873), .B1(
        n19872), .B2(n19928), .ZN(n19862) );
  OAI211_X1 U22903 ( .C1(n20001), .C2(n19903), .A(n19863), .B(n19862), .ZN(
        P2_U3131) );
  AOI22_X1 U22904 ( .A1(n19871), .A2(n20058), .B1(n20057), .B2(n19870), .ZN(
        n19865) );
  AOI22_X1 U22905 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19873), .B1(
        n19872), .B2(n20059), .ZN(n19864) );
  OAI211_X1 U22906 ( .C1(n20062), .C2(n19903), .A(n19865), .B(n19864), .ZN(
        P2_U3132) );
  AOI22_X1 U22907 ( .A1(n19871), .A2(n20064), .B1(n20063), .B2(n19870), .ZN(
        n19867) );
  AOI22_X1 U22908 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19873), .B1(
        n19872), .B2(n20065), .ZN(n19866) );
  OAI211_X1 U22909 ( .C1(n20068), .C2(n19903), .A(n19867), .B(n19866), .ZN(
        P2_U3133) );
  AOI22_X1 U22910 ( .A1(n19871), .A2(n20070), .B1(n20069), .B2(n19870), .ZN(
        n19869) );
  AOI22_X1 U22911 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19873), .B1(
        n19872), .B2(n20071), .ZN(n19868) );
  OAI211_X1 U22912 ( .C1(n20076), .C2(n19903), .A(n19869), .B(n19868), .ZN(
        P2_U3134) );
  AOI22_X1 U22913 ( .A1(n19871), .A2(n20079), .B1(n20077), .B2(n19870), .ZN(
        n19875) );
  AOI22_X1 U22914 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19873), .B1(
        n19872), .B2(n19939), .ZN(n19874) );
  OAI211_X1 U22915 ( .C1(n20015), .C2(n19903), .A(n19875), .B(n19874), .ZN(
        P2_U3135) );
  OR2_X1 U22916 ( .A1(n20205), .A2(n19881), .ZN(n19880) );
  INV_X1 U22917 ( .A(n19884), .ZN(n19878) );
  INV_X1 U22918 ( .A(n19881), .ZN(n19876) );
  NAND2_X1 U22919 ( .A1(n19877), .A2(n19876), .ZN(n19883) );
  INV_X1 U22920 ( .A(n19883), .ZN(n19905) );
  OAI21_X1 U22921 ( .B1(n19878), .B2(n19905), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19879) );
  OAI21_X1 U22922 ( .B1(n19880), .B2(n20176), .A(n19879), .ZN(n19906) );
  AOI22_X1 U22923 ( .A1(n19906), .A2(n20026), .B1(n20025), .B2(n19905), .ZN(
        n19888) );
  OAI22_X1 U22924 ( .A1(n20029), .A2(n19882), .B1(n19881), .B2(n20205), .ZN(
        n19886) );
  OAI211_X1 U22925 ( .C1(n19884), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19883), 
        .B(n20176), .ZN(n19885) );
  NAND3_X1 U22926 ( .A1(n19886), .A2(n20033), .A3(n19885), .ZN(n19908) );
  AOI22_X1 U22927 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n20035), .ZN(n19887) );
  OAI211_X1 U22928 ( .C1(n20038), .C2(n19911), .A(n19888), .B(n19887), .ZN(
        P2_U3136) );
  AOI22_X1 U22929 ( .A1(n19906), .A2(n20040), .B1(n20039), .B2(n19905), .ZN(
        n19890) );
  AOI22_X1 U22930 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n20041), .ZN(n19889) );
  OAI211_X1 U22931 ( .C1(n20044), .C2(n19911), .A(n19890), .B(n19889), .ZN(
        P2_U3137) );
  AOI22_X1 U22932 ( .A1(n19906), .A2(n20046), .B1(n20045), .B2(n19905), .ZN(
        n19892) );
  AOI22_X1 U22933 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n19925), .ZN(n19891) );
  OAI211_X1 U22934 ( .C1(n19996), .C2(n19911), .A(n19892), .B(n19891), .ZN(
        P2_U3138) );
  AOI22_X1 U22935 ( .A1(n19906), .A2(n20052), .B1(n20051), .B2(n19905), .ZN(
        n19894) );
  AOI22_X1 U22936 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n19928), .ZN(n19893) );
  OAI211_X1 U22937 ( .C1(n20001), .C2(n19911), .A(n19894), .B(n19893), .ZN(
        P2_U3139) );
  AOI22_X1 U22938 ( .A1(n19906), .A2(n20058), .B1(n20057), .B2(n19905), .ZN(
        n19896) );
  AOI22_X1 U22939 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n20059), .ZN(n19895) );
  OAI211_X1 U22940 ( .C1(n20062), .C2(n19911), .A(n19896), .B(n19895), .ZN(
        P2_U3140) );
  AOI22_X1 U22941 ( .A1(n19906), .A2(n20064), .B1(n20063), .B2(n19905), .ZN(
        n19899) );
  AOI22_X1 U22942 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19908), .B1(
        n19940), .B2(n19897), .ZN(n19898) );
  OAI211_X1 U22943 ( .C1(n20008), .C2(n19903), .A(n19899), .B(n19898), .ZN(
        P2_U3141) );
  AOI22_X1 U22944 ( .A1(n19906), .A2(n20070), .B1(n20069), .B2(n19905), .ZN(
        n19902) );
  AOI22_X1 U22945 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19908), .B1(
        n19940), .B2(n19900), .ZN(n19901) );
  OAI211_X1 U22946 ( .C1(n19904), .C2(n19903), .A(n19902), .B(n19901), .ZN(
        P2_U3142) );
  AOI22_X1 U22947 ( .A1(n19906), .A2(n20079), .B1(n20077), .B2(n19905), .ZN(
        n19910) );
  AOI22_X1 U22948 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19908), .B1(
        n19907), .B2(n19939), .ZN(n19909) );
  OAI211_X1 U22949 ( .C1(n20015), .C2(n19911), .A(n19910), .B(n19909), .ZN(
        P2_U3143) );
  NAND2_X1 U22950 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19914), .ZN(
        n19918) );
  OR2_X1 U22951 ( .A1(n19918), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19916) );
  NAND3_X1 U22952 ( .A1(n20205), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19948) );
  NOR2_X1 U22953 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19948), .ZN(
        n19937) );
  AOI22_X1 U22954 ( .A1(n19938), .A2(n20026), .B1(n20025), .B2(n19937), .ZN(
        n19922) );
  OAI21_X1 U22955 ( .B1(n19966), .B2(n19940), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19919) );
  AOI211_X1 U22956 ( .C1(n19919), .C2(n19918), .A(n19917), .B(n19978), .ZN(
        n19920) );
  OAI21_X1 U22957 ( .B1(n19937), .B2(n19977), .A(n19920), .ZN(n19941) );
  AOI22_X1 U22958 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19941), .B1(
        n19940), .B2(n20035), .ZN(n19921) );
  OAI211_X1 U22959 ( .C1(n20038), .C2(n19973), .A(n19922), .B(n19921), .ZN(
        P2_U3144) );
  AOI22_X1 U22960 ( .A1(n19938), .A2(n20040), .B1(n20039), .B2(n19937), .ZN(
        n19924) );
  AOI22_X1 U22961 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19941), .B1(
        n19940), .B2(n20041), .ZN(n19923) );
  OAI211_X1 U22962 ( .C1(n20044), .C2(n19973), .A(n19924), .B(n19923), .ZN(
        P2_U3145) );
  AOI22_X1 U22963 ( .A1(n19938), .A2(n20046), .B1(n20045), .B2(n19937), .ZN(
        n19927) );
  AOI22_X1 U22964 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19941), .B1(
        n19940), .B2(n19925), .ZN(n19926) );
  OAI211_X1 U22965 ( .C1(n19996), .C2(n19973), .A(n19927), .B(n19926), .ZN(
        P2_U3146) );
  AOI22_X1 U22966 ( .A1(n19938), .A2(n20052), .B1(n20051), .B2(n19937), .ZN(
        n19930) );
  AOI22_X1 U22967 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19941), .B1(
        n19940), .B2(n19928), .ZN(n19929) );
  OAI211_X1 U22968 ( .C1(n20001), .C2(n19973), .A(n19930), .B(n19929), .ZN(
        P2_U3147) );
  AOI22_X1 U22969 ( .A1(n19938), .A2(n20058), .B1(n20057), .B2(n19937), .ZN(
        n19932) );
  AOI22_X1 U22970 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19941), .B1(
        n19940), .B2(n20059), .ZN(n19931) );
  OAI211_X1 U22971 ( .C1(n20062), .C2(n19973), .A(n19932), .B(n19931), .ZN(
        P2_U3148) );
  AOI22_X1 U22972 ( .A1(n19938), .A2(n20064), .B1(n20063), .B2(n19937), .ZN(
        n19934) );
  AOI22_X1 U22973 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19941), .B1(
        n19940), .B2(n20065), .ZN(n19933) );
  OAI211_X1 U22974 ( .C1(n20068), .C2(n19973), .A(n19934), .B(n19933), .ZN(
        P2_U3149) );
  AOI22_X1 U22975 ( .A1(n19938), .A2(n20070), .B1(n20069), .B2(n19937), .ZN(
        n19936) );
  AOI22_X1 U22976 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19941), .B1(
        n19940), .B2(n20071), .ZN(n19935) );
  OAI211_X1 U22977 ( .C1(n20076), .C2(n19973), .A(n19936), .B(n19935), .ZN(
        P2_U3150) );
  AOI22_X1 U22978 ( .A1(n19938), .A2(n20079), .B1(n20077), .B2(n19937), .ZN(
        n19943) );
  AOI22_X1 U22979 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19941), .B1(
        n19940), .B2(n19939), .ZN(n19942) );
  OAI211_X1 U22980 ( .C1(n20015), .C2(n19973), .A(n19943), .B(n19942), .ZN(
        P2_U3151) );
  NOR2_X1 U22981 ( .A1(n12154), .A2(n19948), .ZN(n19981) );
  INV_X1 U22982 ( .A(n19981), .ZN(n19950) );
  NAND2_X1 U22983 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19950), .ZN(n19945) );
  OR2_X1 U22984 ( .A1(n19946), .A2(n19945), .ZN(n19952) );
  OAI21_X1 U22985 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19948), .A(n20207), 
        .ZN(n19947) );
  AOI22_X1 U22986 ( .A1(n19969), .A2(n20026), .B1(n20025), .B2(n19981), .ZN(
        n19955) );
  OAI21_X1 U22987 ( .B1(n20029), .B2(n19949), .A(n19948), .ZN(n19953) );
  NAND2_X1 U22988 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19950), .ZN(n19951) );
  NAND4_X1 U22989 ( .A1(n19953), .A2(n20033), .A3(n19952), .A4(n19951), .ZN(
        n19970) );
  AOI22_X1 U22990 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19970), .B1(
        n19966), .B2(n20035), .ZN(n19954) );
  OAI211_X1 U22991 ( .C1(n20038), .C2(n20021), .A(n19955), .B(n19954), .ZN(
        P2_U3152) );
  AOI22_X1 U22992 ( .A1(n19969), .A2(n20040), .B1(n20039), .B2(n19981), .ZN(
        n19957) );
  AOI22_X1 U22993 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19970), .B1(
        n20010), .B2(n19988), .ZN(n19956) );
  OAI211_X1 U22994 ( .C1(n19991), .C2(n19973), .A(n19957), .B(n19956), .ZN(
        P2_U3153) );
  AOI22_X1 U22995 ( .A1(n19969), .A2(n20046), .B1(n20045), .B2(n19981), .ZN(
        n19959) );
  AOI22_X1 U22996 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19970), .B1(
        n20010), .B2(n20047), .ZN(n19958) );
  OAI211_X1 U22997 ( .C1(n20050), .C2(n19973), .A(n19959), .B(n19958), .ZN(
        P2_U3154) );
  AOI22_X1 U22998 ( .A1(n19969), .A2(n20052), .B1(n20051), .B2(n19981), .ZN(
        n19961) );
  AOI22_X1 U22999 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19970), .B1(
        n20010), .B2(n20053), .ZN(n19960) );
  OAI211_X1 U23000 ( .C1(n20056), .C2(n19973), .A(n19961), .B(n19960), .ZN(
        P2_U3155) );
  AOI22_X1 U23001 ( .A1(n19969), .A2(n20058), .B1(n20057), .B2(n19981), .ZN(
        n19963) );
  AOI22_X1 U23002 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19970), .B1(
        n19966), .B2(n20059), .ZN(n19962) );
  OAI211_X1 U23003 ( .C1(n20062), .C2(n20021), .A(n19963), .B(n19962), .ZN(
        P2_U3156) );
  AOI22_X1 U23004 ( .A1(n19969), .A2(n20064), .B1(n20063), .B2(n19981), .ZN(
        n19965) );
  AOI22_X1 U23005 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19970), .B1(
        n19966), .B2(n20065), .ZN(n19964) );
  OAI211_X1 U23006 ( .C1(n20068), .C2(n20021), .A(n19965), .B(n19964), .ZN(
        P2_U3157) );
  AOI22_X1 U23007 ( .A1(n19969), .A2(n20070), .B1(n20069), .B2(n19981), .ZN(
        n19968) );
  AOI22_X1 U23008 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19970), .B1(
        n19966), .B2(n20071), .ZN(n19967) );
  OAI211_X1 U23009 ( .C1(n20076), .C2(n20021), .A(n19968), .B(n19967), .ZN(
        P2_U3158) );
  AOI22_X1 U23010 ( .A1(n19969), .A2(n20079), .B1(n20077), .B2(n19981), .ZN(
        n19972) );
  AOI22_X1 U23011 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19970), .B1(
        n20010), .B2(n20081), .ZN(n19971) );
  OAI211_X1 U23012 ( .C1(n20087), .C2(n19973), .A(n19972), .B(n19971), .ZN(
        P2_U3159) );
  NAND2_X1 U23013 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19975), .ZN(
        n20027) );
  NOR2_X1 U23014 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20027), .ZN(
        n20009) );
  AOI22_X1 U23015 ( .A1(n20035), .A2(n20010), .B1(n20025), .B2(n20009), .ZN(
        n19987) );
  NOR3_X1 U23016 ( .A1(n19982), .A2(n20009), .A3(n20207), .ZN(n19980) );
  OAI21_X1 U23017 ( .B1(n20072), .B2(n20010), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19976) );
  NAND2_X1 U23018 ( .A1(n19976), .A2(n20180), .ZN(n19985) );
  AOI221_X1 U23019 ( .B1(n19977), .B2(n19985), .C1(n19977), .C2(n19981), .A(
        n20009), .ZN(n19979) );
  NOR2_X1 U23020 ( .A1(n20009), .A2(n19981), .ZN(n19984) );
  OAI21_X1 U23021 ( .B1(n19982), .B2(n20009), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19983) );
  AOI22_X1 U23022 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20018), .B1(
        n20026), .B2(n20017), .ZN(n19986) );
  OAI211_X1 U23023 ( .C1(n20038), .C2(n20086), .A(n19987), .B(n19986), .ZN(
        P2_U3160) );
  AOI22_X1 U23024 ( .A1(n19988), .A2(n20072), .B1(n20039), .B2(n20009), .ZN(
        n19990) );
  AOI22_X1 U23025 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20018), .B1(
        n20040), .B2(n20017), .ZN(n19989) );
  OAI211_X1 U23026 ( .C1(n19991), .C2(n20021), .A(n19990), .B(n19989), .ZN(
        P2_U3161) );
  INV_X1 U23027 ( .A(n20009), .ZN(n20013) );
  OAI22_X1 U23028 ( .A1(n20021), .A2(n20050), .B1(n19992), .B2(n20013), .ZN(
        n19993) );
  INV_X1 U23029 ( .A(n19993), .ZN(n19995) );
  AOI22_X1 U23030 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20018), .B1(
        n20046), .B2(n20017), .ZN(n19994) );
  OAI211_X1 U23031 ( .C1(n19996), .C2(n20086), .A(n19995), .B(n19994), .ZN(
        P2_U3162) );
  OAI22_X1 U23032 ( .A1(n20021), .A2(n20056), .B1(n19997), .B2(n20013), .ZN(
        n19998) );
  INV_X1 U23033 ( .A(n19998), .ZN(n20000) );
  AOI22_X1 U23034 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20018), .B1(
        n20052), .B2(n20017), .ZN(n19999) );
  OAI211_X1 U23035 ( .C1(n20001), .C2(n20086), .A(n20000), .B(n19999), .ZN(
        P2_U3163) );
  AOI22_X1 U23036 ( .A1(n20059), .A2(n20010), .B1(n20057), .B2(n20009), .ZN(
        n20003) );
  AOI22_X1 U23037 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20018), .B1(
        n20058), .B2(n20017), .ZN(n20002) );
  OAI211_X1 U23038 ( .C1(n20062), .C2(n20086), .A(n20003), .B(n20002), .ZN(
        P2_U3164) );
  OAI22_X1 U23039 ( .A1(n20086), .A2(n20068), .B1(n20004), .B2(n20013), .ZN(
        n20005) );
  INV_X1 U23040 ( .A(n20005), .ZN(n20007) );
  AOI22_X1 U23041 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20018), .B1(
        n20064), .B2(n20017), .ZN(n20006) );
  OAI211_X1 U23042 ( .C1(n20008), .C2(n20021), .A(n20007), .B(n20006), .ZN(
        P2_U3165) );
  AOI22_X1 U23043 ( .A1(n20071), .A2(n20010), .B1(n20069), .B2(n20009), .ZN(
        n20012) );
  AOI22_X1 U23044 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20018), .B1(
        n20070), .B2(n20017), .ZN(n20011) );
  OAI211_X1 U23045 ( .C1(n20076), .C2(n20086), .A(n20012), .B(n20011), .ZN(
        P2_U3166) );
  OAI22_X1 U23046 ( .A1(n20086), .A2(n20015), .B1(n20014), .B2(n20013), .ZN(
        n20016) );
  INV_X1 U23047 ( .A(n20016), .ZN(n20020) );
  AOI22_X1 U23048 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20018), .B1(
        n20079), .B2(n20017), .ZN(n20019) );
  OAI211_X1 U23049 ( .C1(n20087), .C2(n20021), .A(n20020), .B(n20019), .ZN(
        P2_U3167) );
  NAND2_X1 U23050 ( .A1(n20030), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20022) );
  OR2_X1 U23051 ( .A1(n20023), .A2(n20022), .ZN(n20032) );
  OAI21_X1 U23052 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20027), .A(n20207), 
        .ZN(n20024) );
  AOI22_X1 U23053 ( .A1(n20080), .A2(n20026), .B1(n20078), .B2(n20025), .ZN(
        n20037) );
  OAI21_X1 U23054 ( .B1(n20029), .B2(n20028), .A(n20027), .ZN(n20034) );
  NAND2_X1 U23055 ( .A1(n20030), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20031) );
  NAND4_X1 U23056 ( .A1(n20034), .A2(n20033), .A3(n20032), .A4(n20031), .ZN(
        n20083) );
  AOI22_X1 U23057 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20083), .B1(
        n20072), .B2(n20035), .ZN(n20036) );
  OAI211_X1 U23058 ( .C1(n20038), .C2(n20075), .A(n20037), .B(n20036), .ZN(
        P2_U3168) );
  AOI22_X1 U23059 ( .A1(n20080), .A2(n20040), .B1(n20078), .B2(n20039), .ZN(
        n20043) );
  AOI22_X1 U23060 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20083), .B1(
        n20072), .B2(n20041), .ZN(n20042) );
  OAI211_X1 U23061 ( .C1(n20044), .C2(n20075), .A(n20043), .B(n20042), .ZN(
        P2_U3169) );
  AOI22_X1 U23062 ( .A1(n20080), .A2(n20046), .B1(n20078), .B2(n20045), .ZN(
        n20049) );
  AOI22_X1 U23063 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20083), .B1(
        n20082), .B2(n20047), .ZN(n20048) );
  OAI211_X1 U23064 ( .C1(n20050), .C2(n20086), .A(n20049), .B(n20048), .ZN(
        P2_U3170) );
  AOI22_X1 U23065 ( .A1(n20080), .A2(n20052), .B1(n20078), .B2(n20051), .ZN(
        n20055) );
  AOI22_X1 U23066 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20083), .B1(
        n20082), .B2(n20053), .ZN(n20054) );
  OAI211_X1 U23067 ( .C1(n20056), .C2(n20086), .A(n20055), .B(n20054), .ZN(
        P2_U3171) );
  AOI22_X1 U23068 ( .A1(n20080), .A2(n20058), .B1(n20078), .B2(n20057), .ZN(
        n20061) );
  AOI22_X1 U23069 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20083), .B1(
        n20072), .B2(n20059), .ZN(n20060) );
  OAI211_X1 U23070 ( .C1(n20062), .C2(n20075), .A(n20061), .B(n20060), .ZN(
        P2_U3172) );
  AOI22_X1 U23071 ( .A1(n20080), .A2(n20064), .B1(n20078), .B2(n20063), .ZN(
        n20067) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20083), .B1(
        n20072), .B2(n20065), .ZN(n20066) );
  OAI211_X1 U23073 ( .C1(n20068), .C2(n20075), .A(n20067), .B(n20066), .ZN(
        P2_U3173) );
  AOI22_X1 U23074 ( .A1(n20080), .A2(n20070), .B1(n20078), .B2(n20069), .ZN(
        n20074) );
  AOI22_X1 U23075 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20083), .B1(
        n20072), .B2(n20071), .ZN(n20073) );
  OAI211_X1 U23076 ( .C1(n20076), .C2(n20075), .A(n20074), .B(n20073), .ZN(
        P2_U3174) );
  AOI22_X1 U23077 ( .A1(n20080), .A2(n20079), .B1(n20078), .B2(n20077), .ZN(
        n20085) );
  AOI22_X1 U23078 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20083), .B1(
        n20082), .B2(n20081), .ZN(n20084) );
  OAI211_X1 U23079 ( .C1(n20087), .C2(n20086), .A(n20085), .B(n20084), .ZN(
        P2_U3175) );
  AND2_X1 U23080 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20088), .ZN(
        P2_U3179) );
  AND2_X1 U23081 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20088), .ZN(
        P2_U3180) );
  AND2_X1 U23082 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20088), .ZN(
        P2_U3181) );
  NOR2_X1 U23083 ( .A1(n21431), .A2(n20175), .ZN(P2_U3182) );
  AND2_X1 U23084 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20088), .ZN(
        P2_U3183) );
  AND2_X1 U23085 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20088), .ZN(
        P2_U3184) );
  AND2_X1 U23086 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20088), .ZN(
        P2_U3185) );
  AND2_X1 U23087 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20088), .ZN(
        P2_U3186) );
  AND2_X1 U23088 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20088), .ZN(
        P2_U3187) );
  AND2_X1 U23089 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20088), .ZN(
        P2_U3188) );
  AND2_X1 U23090 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20088), .ZN(
        P2_U3189) );
  AND2_X1 U23091 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20088), .ZN(
        P2_U3190) );
  AND2_X1 U23092 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20088), .ZN(
        P2_U3191) );
  AND2_X1 U23093 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20088), .ZN(
        P2_U3192) );
  AND2_X1 U23094 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20088), .ZN(
        P2_U3193) );
  AND2_X1 U23095 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20088), .ZN(
        P2_U3194) );
  AND2_X1 U23096 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20088), .ZN(
        P2_U3195) );
  AND2_X1 U23097 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20088), .ZN(
        P2_U3196) );
  NOR2_X1 U23098 ( .A1(n21482), .A2(n20175), .ZN(P2_U3197) );
  INV_X1 U23099 ( .A(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21280) );
  NOR2_X1 U23100 ( .A1(n21280), .A2(n20175), .ZN(P2_U3198) );
  AND2_X1 U23101 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20088), .ZN(
        P2_U3199) );
  AND2_X1 U23102 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20088), .ZN(
        P2_U3200) );
  AND2_X1 U23103 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20088), .ZN(P2_U3201) );
  AND2_X1 U23104 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20088), .ZN(P2_U3202) );
  AND2_X1 U23105 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20088), .ZN(P2_U3203) );
  AND2_X1 U23106 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20088), .ZN(P2_U3204) );
  AND2_X1 U23107 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20088), .ZN(P2_U3205) );
  AND2_X1 U23108 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20088), .ZN(P2_U3206) );
  AND2_X1 U23109 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20088), .ZN(P2_U3207) );
  AND2_X1 U23110 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20088), .ZN(P2_U3208) );
  NOR2_X1 U23111 ( .A1(n20100), .A2(n20238), .ZN(n20097) );
  INV_X1 U23112 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20098) );
  NOR3_X1 U23113 ( .A1(n20097), .A2(n20098), .A3(n20089), .ZN(n20093) );
  OAI211_X1 U23114 ( .C1(HOLD), .C2(n20098), .A(n20090), .B(n20241), .ZN(
        n20092) );
  NOR3_X1 U23115 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21099), .ZN(n20105) );
  INV_X1 U23116 ( .A(n20105), .ZN(n20091) );
  OAI211_X1 U23117 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20093), .A(n20092), 
        .B(n20091), .ZN(P2_U3209) );
  AOI21_X1 U23118 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21095), .A(n21283), 
        .ZN(n20101) );
  NOR3_X1 U23119 ( .A1(n20101), .A2(n20098), .A3(n20089), .ZN(n20094) );
  NOR2_X1 U23120 ( .A1(n20094), .A2(n20097), .ZN(n20095) );
  OAI211_X1 U23121 ( .C1(n21095), .C2(n20096), .A(n20095), .B(n20228), .ZN(
        P2_U3210) );
  AOI22_X1 U23122 ( .A1(n20099), .A2(n20098), .B1(n20097), .B2(n21099), .ZN(
        n20107) );
  OAI21_X1 U23123 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20106) );
  NOR2_X1 U23124 ( .A1(n21283), .A2(n20100), .ZN(n20102) );
  AOI21_X1 U23125 ( .B1(n20103), .B2(n20102), .A(n20101), .ZN(n20104) );
  OAI22_X1 U23126 ( .A1(n20107), .A2(n20106), .B1(n20105), .B2(n20104), .ZN(
        P2_U3211) );
  NAND2_X1 U23127 ( .A1(n20158), .A2(n21283), .ZN(n20165) );
  CLKBUF_X1 U23128 ( .A(n20165), .Z(n20161) );
  OAI222_X1 U23129 ( .A1(n20161), .A2(n20110), .B1(n20109), .B2(n20158), .C1(
        n20108), .C2(n20162), .ZN(P2_U3212) );
  OAI222_X1 U23130 ( .A1(n20165), .A2(n20112), .B1(n20111), .B2(n20158), .C1(
        n20110), .C2(n20162), .ZN(P2_U3213) );
  INV_X1 U23131 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n20114) );
  OAI222_X1 U23132 ( .A1(n20165), .A2(n20114), .B1(n20113), .B2(n20158), .C1(
        n20112), .C2(n20162), .ZN(P2_U3214) );
  OAI222_X1 U23133 ( .A1(n20165), .A2(n15747), .B1(n20115), .B2(n20158), .C1(
        n20114), .C2(n20162), .ZN(P2_U3215) );
  OAI222_X1 U23134 ( .A1(n20165), .A2(n20117), .B1(n20116), .B2(n20158), .C1(
        n15747), .C2(n20162), .ZN(P2_U3216) );
  INV_X1 U23135 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20118) );
  OAI222_X1 U23136 ( .A1(n20165), .A2(n20119), .B1(n20118), .B2(n20158), .C1(
        n20117), .C2(n20162), .ZN(P2_U3217) );
  OAI222_X1 U23137 ( .A1(n20161), .A2(n20121), .B1(n20120), .B2(n20158), .C1(
        n20119), .C2(n20162), .ZN(P2_U3218) );
  OAI222_X1 U23138 ( .A1(n20161), .A2(n20123), .B1(n20122), .B2(n20158), .C1(
        n20121), .C2(n20162), .ZN(P2_U3219) );
  OAI222_X1 U23139 ( .A1(n20161), .A2(n20125), .B1(n20124), .B2(n20158), .C1(
        n20123), .C2(n20162), .ZN(P2_U3220) );
  OAI222_X1 U23140 ( .A1(n20161), .A2(n20127), .B1(n20126), .B2(n20158), .C1(
        n20125), .C2(n20162), .ZN(P2_U3221) );
  OAI222_X1 U23141 ( .A1(n20161), .A2(n20129), .B1(n20128), .B2(n20158), .C1(
        n20127), .C2(n20162), .ZN(P2_U3222) );
  OAI222_X1 U23142 ( .A1(n20161), .A2(n15665), .B1(n20130), .B2(n20158), .C1(
        n20129), .C2(n20162), .ZN(P2_U3223) );
  OAI222_X1 U23143 ( .A1(n20165), .A2(n20132), .B1(n20131), .B2(n20158), .C1(
        n15665), .C2(n20162), .ZN(P2_U3224) );
  OAI222_X1 U23144 ( .A1(n20165), .A2(n20134), .B1(n20133), .B2(n20158), .C1(
        n20132), .C2(n20162), .ZN(P2_U3225) );
  OAI222_X1 U23145 ( .A1(n20165), .A2(n20136), .B1(n20135), .B2(n20158), .C1(
        n20134), .C2(n20162), .ZN(P2_U3226) );
  INV_X1 U23146 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20138) );
  OAI222_X1 U23147 ( .A1(n20165), .A2(n20138), .B1(n20137), .B2(n20158), .C1(
        n20136), .C2(n20162), .ZN(P2_U3227) );
  INV_X1 U23148 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20140) );
  OAI222_X1 U23149 ( .A1(n20165), .A2(n20140), .B1(n20139), .B2(n20158), .C1(
        n20138), .C2(n20162), .ZN(P2_U3228) );
  OAI222_X1 U23150 ( .A1(n20165), .A2(n20141), .B1(n21316), .B2(n20158), .C1(
        n20140), .C2(n20162), .ZN(P2_U3229) );
  OAI222_X1 U23151 ( .A1(n20161), .A2(n20143), .B1(n20142), .B2(n20158), .C1(
        n20141), .C2(n20162), .ZN(P2_U3230) );
  OAI222_X1 U23152 ( .A1(n20161), .A2(n20145), .B1(n20144), .B2(n20158), .C1(
        n20143), .C2(n20162), .ZN(P2_U3231) );
  INV_X1 U23153 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20147) );
  OAI222_X1 U23154 ( .A1(n20161), .A2(n20147), .B1(n20146), .B2(n20158), .C1(
        n20145), .C2(n20162), .ZN(P2_U3232) );
  INV_X1 U23155 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n21473) );
  OAI222_X1 U23156 ( .A1(n20161), .A2(n21473), .B1(n20148), .B2(n20158), .C1(
        n20147), .C2(n20162), .ZN(P2_U3233) );
  INV_X1 U23157 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20149) );
  OAI222_X1 U23158 ( .A1(n20161), .A2(n20149), .B1(n21337), .B2(n20158), .C1(
        n21473), .C2(n20162), .ZN(P2_U3234) );
  OAI222_X1 U23159 ( .A1(n20161), .A2(n20151), .B1(n20150), .B2(n20158), .C1(
        n20149), .C2(n20162), .ZN(P2_U3235) );
  INV_X1 U23160 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20153) );
  OAI222_X1 U23161 ( .A1(n20161), .A2(n20153), .B1(n20152), .B2(n20158), .C1(
        n20151), .C2(n20162), .ZN(P2_U3236) );
  OAI222_X1 U23162 ( .A1(n20161), .A2(n20156), .B1(n20154), .B2(n20158), .C1(
        n20153), .C2(n20162), .ZN(P2_U3237) );
  OAI222_X1 U23163 ( .A1(n20162), .A2(n20156), .B1(n20155), .B2(n20158), .C1(
        n20157), .C2(n20161), .ZN(P2_U3238) );
  INV_X1 U23164 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20159) );
  OAI222_X1 U23165 ( .A1(n20161), .A2(n20159), .B1(n21240), .B2(n20158), .C1(
        n20157), .C2(n20162), .ZN(P2_U3239) );
  INV_X1 U23166 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20163) );
  OAI222_X1 U23167 ( .A1(n20161), .A2(n20163), .B1(n20160), .B2(n20158), .C1(
        n20159), .C2(n20162), .ZN(P2_U3240) );
  OAI222_X1 U23168 ( .A1(n20165), .A2(n11825), .B1(n20164), .B2(n20158), .C1(
        n20163), .C2(n20162), .ZN(P2_U3241) );
  INV_X1 U23169 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20166) );
  AOI22_X1 U23170 ( .A1(n20158), .A2(n20167), .B1(n20166), .B2(n20241), .ZN(
        P2_U3585) );
  MUX2_X1 U23171 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20158), .Z(P2_U3586) );
  INV_X1 U23172 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20168) );
  AOI22_X1 U23173 ( .A1(n20158), .A2(n20169), .B1(n20168), .B2(n20241), .ZN(
        P2_U3587) );
  INV_X1 U23174 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20170) );
  AOI22_X1 U23175 ( .A1(n20158), .A2(n20171), .B1(n20170), .B2(n20241), .ZN(
        P2_U3588) );
  OAI21_X1 U23176 ( .B1(n20175), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20173), 
        .ZN(n20172) );
  INV_X1 U23177 ( .A(n20172), .ZN(P2_U3591) );
  OAI21_X1 U23178 ( .B1(n20175), .B2(n20174), .A(n20173), .ZN(P2_U3592) );
  OR2_X1 U23179 ( .A1(n20177), .A2(n20176), .ZN(n20186) );
  NAND2_X1 U23180 ( .A1(n20178), .A2(n20201), .ZN(n20191) );
  NAND2_X1 U23181 ( .A1(n20199), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20181) );
  AOI21_X1 U23182 ( .B1(n20181), .B2(n20180), .A(n20179), .ZN(n20189) );
  NAND2_X1 U23183 ( .A1(n20191), .A2(n20189), .ZN(n20183) );
  AOI22_X1 U23184 ( .A1(n20184), .A2(n20183), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20182), .ZN(n20185) );
  AND2_X1 U23185 ( .A1(n20186), .A2(n20185), .ZN(n20187) );
  AOI22_X1 U23186 ( .A1(n20214), .A2(n20188), .B1(n20187), .B2(n20212), .ZN(
        P2_U3602) );
  NOR2_X1 U23187 ( .A1(n20190), .A2(n20189), .ZN(n20193) );
  INV_X1 U23188 ( .A(n20191), .ZN(n20192) );
  AOI211_X1 U23189 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n20194), .A(n20193), 
        .B(n20192), .ZN(n20195) );
  AOI22_X1 U23190 ( .A1(n20214), .A2(n20196), .B1(n20195), .B2(n20212), .ZN(
        P2_U3603) );
  INV_X1 U23191 ( .A(n20210), .ZN(n20198) );
  NOR2_X1 U23192 ( .A1(n20198), .A2(n20197), .ZN(n20200) );
  MUX2_X1 U23193 ( .A(n20201), .B(n20200), .S(n20199), .Z(n20202) );
  AOI21_X1 U23194 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20203), .A(n20202), 
        .ZN(n20204) );
  AOI22_X1 U23195 ( .A1(n20214), .A2(n20205), .B1(n20204), .B2(n20212), .ZN(
        P2_U3604) );
  OAI21_X1 U23196 ( .B1(n20208), .B2(n20207), .A(n20206), .ZN(n20209) );
  AOI21_X1 U23197 ( .B1(n20211), .B2(n20210), .A(n20209), .ZN(n20213) );
  AOI22_X1 U23198 ( .A1(n20214), .A2(n12154), .B1(n20213), .B2(n20212), .ZN(
        P2_U3605) );
  INV_X1 U23199 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20215) );
  AOI22_X1 U23200 ( .A1(n20158), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20215), 
        .B2(n20241), .ZN(P2_U3608) );
  INV_X1 U23201 ( .A(n20216), .ZN(n20219) );
  INV_X1 U23202 ( .A(n20217), .ZN(n20218) );
  AOI22_X1 U23203 ( .A1(n20221), .A2(n20220), .B1(n20219), .B2(n20218), .ZN(
        n20222) );
  NAND2_X1 U23204 ( .A1(n20223), .A2(n20222), .ZN(n20225) );
  MUX2_X1 U23205 ( .A(P2_MORE_REG_SCAN_IN), .B(n20225), .S(n20224), .Z(
        P2_U3609) );
  OAI21_X1 U23206 ( .B1(n20228), .B2(n20227), .A(n20226), .ZN(n20231) );
  NAND3_X1 U23207 ( .A1(n20229), .A2(n20228), .A3(n13063), .ZN(n20230) );
  AND4_X1 U23208 ( .A1(n20231), .A2(n20238), .A3(P2_STATE2_REG_2__SCAN_IN), 
        .A4(n20230), .ZN(n20233) );
  OAI21_X1 U23209 ( .B1(n20233), .B2(n11619), .A(n20232), .ZN(n20240) );
  NOR2_X1 U23210 ( .A1(n20234), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20236) );
  AOI211_X1 U23211 ( .C1(n20238), .C2(n20237), .A(n20236), .B(n20235), .ZN(
        n20239) );
  MUX2_X1 U23212 ( .A(n20240), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n20239), 
        .Z(P2_U3610) );
  INV_X1 U23213 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20242) );
  AOI22_X1 U23214 ( .A1(n20158), .A2(n20243), .B1(n20242), .B2(n20241), .ZN(
        P2_U3611) );
  INV_X1 U23215 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21110) );
  AOI21_X1 U23216 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21110), .A(n21101), 
        .ZN(n20251) );
  INV_X1 U23217 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20245) );
  INV_X1 U23218 ( .A(n21185), .ZN(n21187) );
  AOI21_X1 U23219 ( .B1(n20251), .B2(n20245), .A(n21187), .ZN(P1_U2802) );
  OAI21_X1 U23220 ( .B1(n20247), .B2(n20246), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20248) );
  OAI21_X1 U23221 ( .B1(n20249), .B2(n21091), .A(n20248), .ZN(P1_U2803) );
  NOR2_X1 U23222 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20252) );
  OAI21_X1 U23223 ( .B1(n20252), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21185), .ZN(
        n20250) );
  OAI21_X1 U23224 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21185), .A(n20250), 
        .ZN(P1_U2804) );
  INV_X1 U23225 ( .A(n21185), .ZN(n21184) );
  NOR2_X1 U23226 ( .A1(n20251), .A2(n21184), .ZN(n21175) );
  OAI21_X1 U23227 ( .B1(BS16), .B2(n20252), .A(n21175), .ZN(n21173) );
  OAI21_X1 U23228 ( .B1(n21175), .B2(n20832), .A(n21173), .ZN(P1_U2805) );
  OAI21_X1 U23229 ( .B1(n20255), .B2(n20254), .A(n20253), .ZN(P1_U2806) );
  NOR4_X1 U23230 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20259) );
  NOR4_X1 U23231 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20258) );
  NOR4_X1 U23232 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20257) );
  NOR4_X1 U23233 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20256) );
  NAND4_X1 U23234 ( .A1(n20259), .A2(n20258), .A3(n20257), .A4(n20256), .ZN(
        n20265) );
  NOR4_X1 U23235 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20263) );
  INV_X1 U23236 ( .A(P1_DATAWIDTH_REG_24__SCAN_IN), .ZN(n21237) );
  INV_X1 U23237 ( .A(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n21266) );
  NAND2_X1 U23238 ( .A1(n21237), .A2(n21266), .ZN(n21213) );
  AOI21_X1 U23239 ( .B1(P1_DATAWIDTH_REG_1__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(n21213), .ZN(n20262) );
  NOR4_X1 U23240 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20261) );
  NOR4_X1 U23241 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20260) );
  NAND4_X1 U23242 ( .A1(n20263), .A2(n20262), .A3(n20261), .A4(n20260), .ZN(
        n20264) );
  NOR2_X1 U23243 ( .A1(n20265), .A2(n20264), .ZN(n21179) );
  INV_X1 U23244 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21168) );
  NOR3_X1 U23245 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20267) );
  OAI21_X1 U23246 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20267), .A(n21179), .ZN(
        n20266) );
  OAI21_X1 U23247 ( .B1(n21179), .B2(n21168), .A(n20266), .ZN(P1_U2807) );
  INV_X1 U23248 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21174) );
  AOI21_X1 U23249 ( .B1(n13419), .B2(n21174), .A(n20267), .ZN(n20268) );
  INV_X1 U23250 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21165) );
  INV_X1 U23251 ( .A(n21179), .ZN(n21181) );
  AOI22_X1 U23252 ( .A1(n21179), .A2(n20268), .B1(n21165), .B2(n21181), .ZN(
        P1_U2808) );
  AOI22_X1 U23253 ( .A1(n20334), .A2(P1_EBX_REG_9__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20335), .ZN(n20269) );
  OAI211_X1 U23254 ( .C1(n20294), .C2(n20270), .A(n20269), .B(n20314), .ZN(
        n20271) );
  AOI221_X1 U23255 ( .B1(n20273), .B2(P1_REIP_REG_9__SCAN_IN), .C1(n20272), 
        .C2(n15214), .A(n20271), .ZN(n20278) );
  INV_X1 U23256 ( .A(n20274), .ZN(n20275) );
  AOI22_X1 U23257 ( .A1(n20276), .A2(n20298), .B1(n20275), .B2(n20344), .ZN(
        n20277) );
  NAND2_X1 U23258 ( .A1(n20278), .A2(n20277), .ZN(P1_U2831) );
  NAND2_X1 U23259 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20284) );
  NOR3_X1 U23260 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20284), .A3(n20309), .ZN(
        n20279) );
  AOI211_X1 U23261 ( .C1(n20335), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20296), .B(n20279), .ZN(n20283) );
  INV_X1 U23262 ( .A(n20280), .ZN(n20281) );
  AOI22_X1 U23263 ( .A1(n20334), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n20333), .B2(
        n20281), .ZN(n20282) );
  AND2_X1 U23264 ( .A1(n20283), .A2(n20282), .ZN(n20289) );
  INV_X1 U23265 ( .A(n20284), .ZN(n20285) );
  INV_X1 U23266 ( .A(n20302), .ZN(n20325) );
  OAI21_X1 U23267 ( .B1(n20286), .B2(n20285), .A(n20325), .ZN(n20297) );
  AOI22_X1 U23268 ( .A1(n20287), .A2(n20298), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20297), .ZN(n20288) );
  OAI211_X1 U23269 ( .C1(n20290), .C2(n20330), .A(n20289), .B(n20288), .ZN(
        P1_U2833) );
  INV_X1 U23270 ( .A(n20349), .ZN(n20293) );
  NOR2_X1 U23271 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20309), .ZN(n20291) );
  AOI22_X1 U23272 ( .A1(n20334), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n20291), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n20292) );
  OAI21_X1 U23273 ( .B1(n20294), .B2(n20293), .A(n20292), .ZN(n20295) );
  AOI211_X1 U23274 ( .C1(n20335), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20296), .B(n20295), .ZN(n20300) );
  AOI22_X1 U23275 ( .A1(n20352), .A2(n20298), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n20297), .ZN(n20299) );
  OAI211_X1 U23276 ( .C1(n20301), .C2(n20330), .A(n20300), .B(n20299), .ZN(
        P1_U2834) );
  AOI22_X1 U23277 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20335), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n20302), .ZN(n20303) );
  OAI211_X1 U23278 ( .C1(n20305), .C2(n20304), .A(n20303), .B(n20314), .ZN(
        n20306) );
  AOI21_X1 U23279 ( .B1(n20333), .B2(n20307), .A(n20306), .ZN(n20308) );
  OAI21_X1 U23280 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20309), .A(n20308), .ZN(
        n20310) );
  AOI21_X1 U23281 ( .B1(n20311), .B2(n20327), .A(n20310), .ZN(n20312) );
  OAI21_X1 U23282 ( .B1(n20313), .B2(n20330), .A(n20312), .ZN(P1_U2835) );
  NAND2_X1 U23283 ( .A1(n20335), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20315) );
  AND2_X1 U23284 ( .A1(n20315), .A2(n20314), .ZN(n20317) );
  NAND2_X1 U23285 ( .A1(n20333), .A2(n20437), .ZN(n20316) );
  OAI211_X1 U23286 ( .C1(n20319), .C2(n20318), .A(n20317), .B(n20316), .ZN(
        n20320) );
  INV_X1 U23287 ( .A(n20320), .ZN(n20329) );
  INV_X1 U23288 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21117) );
  NAND3_X1 U23289 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20321) );
  NOR3_X1 U23290 ( .A1(n20322), .A2(P1_REIP_REG_4__SCAN_IN), .A3(n20321), .ZN(
        n20323) );
  AOI21_X1 U23291 ( .B1(n20334), .B2(P1_EBX_REG_4__SCAN_IN), .A(n20323), .ZN(
        n20324) );
  OAI21_X1 U23292 ( .B1(n20325), .B2(n21117), .A(n20324), .ZN(n20326) );
  AOI21_X1 U23293 ( .B1(n20427), .B2(n20327), .A(n20326), .ZN(n20328) );
  OAI211_X1 U23294 ( .C1(n20432), .C2(n20330), .A(n20329), .B(n20328), .ZN(
        P1_U2836) );
  AOI21_X1 U23295 ( .B1(n20337), .B2(n13419), .A(n20331), .ZN(n20348) );
  INV_X1 U23296 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21113) );
  INV_X1 U23297 ( .A(n20332), .ZN(n20453) );
  AOI22_X1 U23298 ( .A1(n20334), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n20333), .B2(
        n20453), .ZN(n20347) );
  AND2_X1 U23299 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n21113), .ZN(n20336) );
  AOI22_X1 U23300 ( .A1(n20337), .A2(n20336), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20335), .ZN(n20340) );
  INV_X1 U23301 ( .A(n12949), .ZN(n20495) );
  NAND2_X1 U23302 ( .A1(n20495), .A2(n20338), .ZN(n20339) );
  OAI211_X1 U23303 ( .C1(n20342), .C2(n20341), .A(n20340), .B(n20339), .ZN(
        n20343) );
  AOI21_X1 U23304 ( .B1(n20345), .B2(n20344), .A(n20343), .ZN(n20346) );
  OAI211_X1 U23305 ( .C1(n20348), .C2(n21113), .A(n20347), .B(n20346), .ZN(
        P1_U2838) );
  AOI22_X1 U23306 ( .A1(n20352), .A2(n20351), .B1(n20350), .B2(n20349), .ZN(
        n20353) );
  OAI21_X1 U23307 ( .B1(n20355), .B2(n20354), .A(n20353), .ZN(P1_U2866) );
  AOI22_X1 U23308 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20356) );
  OAI21_X1 U23309 ( .B1(n21259), .B2(n20384), .A(n20356), .ZN(P1_U2921) );
  AOI22_X1 U23310 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20357) );
  OAI21_X1 U23311 ( .B1(n20358), .B2(n20384), .A(n20357), .ZN(P1_U2922) );
  AOI22_X1 U23312 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20359) );
  OAI21_X1 U23313 ( .B1(n14995), .B2(n20384), .A(n20359), .ZN(P1_U2923) );
  AOI22_X1 U23314 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20360) );
  OAI21_X1 U23315 ( .B1(n14997), .B2(n20384), .A(n20360), .ZN(P1_U2924) );
  INV_X1 U23316 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20362) );
  AOI22_X1 U23317 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20361) );
  OAI21_X1 U23318 ( .B1(n20362), .B2(n20384), .A(n20361), .ZN(P1_U2925) );
  AOI22_X1 U23319 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20363) );
  OAI21_X1 U23320 ( .B1(n14999), .B2(n20384), .A(n20363), .ZN(P1_U2926) );
  AOI22_X1 U23321 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20372), .B1(n20381), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20364) );
  OAI21_X1 U23322 ( .B1(n15001), .B2(n20384), .A(n20364), .ZN(P1_U2927) );
  AOI22_X1 U23323 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20372), .B1(n20381), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20365) );
  OAI21_X1 U23324 ( .B1(n15002), .B2(n20384), .A(n20365), .ZN(P1_U2928) );
  AOI22_X1 U23325 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20372), .B1(n20381), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20366) );
  OAI21_X1 U23326 ( .B1(n20367), .B2(n20384), .A(n20366), .ZN(P1_U2929) );
  AOI22_X1 U23327 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20372), .B1(n20381), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20368) );
  OAI21_X1 U23328 ( .B1(n20369), .B2(n20384), .A(n20368), .ZN(P1_U2930) );
  AOI22_X1 U23329 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20372), .B1(n20381), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20370) );
  OAI21_X1 U23330 ( .B1(n20371), .B2(n20384), .A(n20370), .ZN(P1_U2931) );
  AOI22_X1 U23331 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20372), .B1(n20381), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20373) );
  OAI21_X1 U23332 ( .B1(n20374), .B2(n20384), .A(n20373), .ZN(P1_U2932) );
  AOI22_X1 U23333 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20375) );
  OAI21_X1 U23334 ( .B1(n20376), .B2(n20384), .A(n20375), .ZN(P1_U2933) );
  AOI22_X1 U23335 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20377) );
  OAI21_X1 U23336 ( .B1(n20378), .B2(n20384), .A(n20377), .ZN(P1_U2934) );
  AOI22_X1 U23337 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20379) );
  OAI21_X1 U23338 ( .B1(n20380), .B2(n20384), .A(n20379), .ZN(P1_U2935) );
  AOI22_X1 U23339 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20382), .B1(n20381), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20383) );
  OAI21_X1 U23340 ( .B1(n20385), .B2(n20384), .A(n20383), .ZN(P1_U2936) );
  AOI22_X1 U23341 ( .A1(n20418), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20392), .ZN(n20388) );
  INV_X1 U23342 ( .A(n20386), .ZN(n20387) );
  NAND2_X1 U23343 ( .A1(n20405), .A2(n20387), .ZN(n20407) );
  NAND2_X1 U23344 ( .A1(n20388), .A2(n20407), .ZN(P1_U2945) );
  AOI22_X1 U23345 ( .A1(n20418), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20392), .ZN(n20391) );
  INV_X1 U23346 ( .A(n20389), .ZN(n20390) );
  NAND2_X1 U23347 ( .A1(n20405), .A2(n20390), .ZN(n20409) );
  NAND2_X1 U23348 ( .A1(n20391), .A2(n20409), .ZN(P1_U2946) );
  AOI22_X1 U23349 ( .A1(n20393), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20392), .ZN(n20396) );
  INV_X1 U23350 ( .A(n20394), .ZN(n20395) );
  NAND2_X1 U23351 ( .A1(n20405), .A2(n20395), .ZN(n20411) );
  NAND2_X1 U23352 ( .A1(n20396), .A2(n20411), .ZN(P1_U2947) );
  AOI22_X1 U23353 ( .A1(n20418), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20417), .ZN(n20399) );
  INV_X1 U23354 ( .A(n20397), .ZN(n20398) );
  NAND2_X1 U23355 ( .A1(n20405), .A2(n20398), .ZN(n20413) );
  NAND2_X1 U23356 ( .A1(n20399), .A2(n20413), .ZN(P1_U2948) );
  AOI22_X1 U23357 ( .A1(n20418), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20417), .ZN(n20402) );
  INV_X1 U23358 ( .A(n20400), .ZN(n20401) );
  NAND2_X1 U23359 ( .A1(n20405), .A2(n20401), .ZN(n20415) );
  NAND2_X1 U23360 ( .A1(n20402), .A2(n20415), .ZN(P1_U2949) );
  AOI22_X1 U23361 ( .A1(n20418), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20417), .ZN(n20406) );
  INV_X1 U23362 ( .A(n20403), .ZN(n20404) );
  NAND2_X1 U23363 ( .A1(n20405), .A2(n20404), .ZN(n20419) );
  NAND2_X1 U23364 ( .A1(n20406), .A2(n20419), .ZN(P1_U2950) );
  AOI22_X1 U23365 ( .A1(n20418), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20392), .ZN(n20408) );
  NAND2_X1 U23366 ( .A1(n20408), .A2(n20407), .ZN(P1_U2960) );
  AOI22_X1 U23367 ( .A1(n20418), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20417), .ZN(n20410) );
  NAND2_X1 U23368 ( .A1(n20410), .A2(n20409), .ZN(P1_U2961) );
  AOI22_X1 U23369 ( .A1(n20418), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20392), .ZN(n20412) );
  NAND2_X1 U23370 ( .A1(n20412), .A2(n20411), .ZN(P1_U2962) );
  AOI22_X1 U23371 ( .A1(n20418), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20417), .ZN(n20414) );
  NAND2_X1 U23372 ( .A1(n20414), .A2(n20413), .ZN(P1_U2963) );
  AOI22_X1 U23373 ( .A1(n20418), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20392), .ZN(n20416) );
  NAND2_X1 U23374 ( .A1(n20416), .A2(n20415), .ZN(P1_U2964) );
  AOI22_X1 U23375 ( .A1(n20418), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20417), .ZN(n20420) );
  NAND2_X1 U23376 ( .A1(n20420), .A2(n20419), .ZN(P1_U2965) );
  AOI22_X1 U23377 ( .A1(n20421), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20436), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20431) );
  AOI21_X1 U23378 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20423), .A(
        n20422), .ZN(n20426) );
  XNOR2_X1 U23379 ( .A(n20424), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20425) );
  XNOR2_X1 U23380 ( .A(n20426), .B(n20425), .ZN(n20439) );
  AOI22_X1 U23381 ( .A1(n20439), .A2(n20429), .B1(n20428), .B2(n20427), .ZN(
        n20430) );
  OAI211_X1 U23382 ( .C1(n20433), .C2(n20432), .A(n20431), .B(n20430), .ZN(
        P1_U2995) );
  INV_X1 U23383 ( .A(n20434), .ZN(n20435) );
  OAI21_X1 U23384 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20435), .ZN(n20442) );
  AOI22_X1 U23385 ( .A1(n20454), .A2(n20437), .B1(n20436), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20441) );
  OR2_X1 U23386 ( .A1(n20452), .A2(n20438), .ZN(n20466) );
  OAI211_X1 U23387 ( .C1(n20460), .C2(n20450), .A(n20459), .B(n20466), .ZN(
        n20445) );
  AOI22_X1 U23388 ( .A1(n20439), .A2(n20477), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20445), .ZN(n20440) );
  OAI211_X1 U23389 ( .C1(n20449), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        P1_U3027) );
  AOI21_X1 U23390 ( .B1(n20454), .B2(n20444), .A(n20443), .ZN(n20448) );
  AOI22_X1 U23391 ( .A1(n20446), .A2(n20477), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20445), .ZN(n20447) );
  OAI211_X1 U23392 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20449), .A(
        n20448), .B(n20447), .ZN(P1_U3028) );
  INV_X1 U23393 ( .A(n20450), .ZN(n20451) );
  OR3_X1 U23394 ( .A1(n20452), .A2(n13344), .A3(n20451), .ZN(n20456) );
  NAND2_X1 U23395 ( .A1(n20454), .A2(n20453), .ZN(n20455) );
  OAI211_X1 U23396 ( .C1(n21113), .C2(n20457), .A(n20456), .B(n20455), .ZN(
        n20458) );
  INV_X1 U23397 ( .A(n20458), .ZN(n20468) );
  OAI21_X1 U23398 ( .B1(n20460), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20459), .ZN(n20461) );
  AOI22_X1 U23399 ( .A1(n20462), .A2(n20477), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20461), .ZN(n20467) );
  NAND3_X1 U23400 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20464), .A3(
        n20463), .ZN(n20465) );
  NAND4_X1 U23401 ( .A1(n20468), .A2(n20467), .A3(n20466), .A4(n20465), .ZN(
        P1_U3029) );
  OAI21_X1 U23402 ( .B1(n20471), .B2(n20470), .A(n20469), .ZN(n20472) );
  INV_X1 U23403 ( .A(n20472), .ZN(n20480) );
  INV_X1 U23404 ( .A(n20473), .ZN(n20478) );
  AND3_X1 U23405 ( .A1(n20475), .A2(n20481), .A3(n20474), .ZN(n20476) );
  AOI21_X1 U23406 ( .B1(n20478), .B2(n20477), .A(n20476), .ZN(n20479) );
  OAI211_X1 U23407 ( .C1(n20482), .C2(n20481), .A(n20480), .B(n20479), .ZN(
        P1_U3030) );
  NOR2_X1 U23408 ( .A1(n20484), .A2(n20483), .ZN(P1_U3032) );
  NOR2_X2 U23409 ( .A1(n20488), .A2(n20487), .ZN(n20531) );
  AOI22_X1 U23410 ( .A1(DATAI_24_), .A2(n20531), .B1(BUF1_REG_24__SCAN_IN), 
        .B2(n20486), .ZN(n20964) );
  NAND2_X1 U23411 ( .A1(n20533), .A2(n12888), .ZN(n20906) );
  NAND3_X1 U23412 ( .A1(n20834), .A2(n20830), .A3(n20905), .ZN(n20543) );
  OR2_X1 U23413 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20543), .ZN(
        n20534) );
  OAI22_X1 U23414 ( .A1(n21071), .A2(n20964), .B1(n20906), .B2(n20534), .ZN(
        n20492) );
  INV_X1 U23415 ( .A(n20492), .ZN(n20505) );
  INV_X1 U23416 ( .A(n20566), .ZN(n20493) );
  OAI21_X1 U23417 ( .B1(n20493), .B2(n21084), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20494) );
  NAND2_X1 U23418 ( .A1(n20494), .A2(n20908), .ZN(n20503) );
  OR2_X1 U23419 ( .A1(n20775), .A2(n20495), .ZN(n20610) );
  NOR2_X1 U23420 ( .A1(n20610), .A2(n20988), .ZN(n20500) );
  INV_X1 U23421 ( .A(n20776), .ZN(n20496) );
  NAND2_X1 U23422 ( .A1(n20496), .A2(n20835), .ZN(n20650) );
  AOI22_X1 U23423 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20650), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20534), .ZN(n20498) );
  INV_X1 U23424 ( .A(n20501), .ZN(n20497) );
  NOR2_X1 U23425 ( .A1(n20497), .A2(n13022), .ZN(n20647) );
  NOR2_X2 U23426 ( .A1(n20653), .A2(n20499), .ZN(n21031) );
  INV_X1 U23427 ( .A(n20500), .ZN(n20502) );
  NOR2_X1 U23428 ( .A1(n20501), .A2(n13022), .ZN(n20654) );
  INV_X1 U23429 ( .A(n20654), .ZN(n20841) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20538), .B1(
        n21031), .B2(n20537), .ZN(n20504) );
  OAI211_X1 U23431 ( .C1(n21041), .C2(n20566), .A(n20505), .B(n20504), .ZN(
        P1_U3033) );
  AOI22_X1 U23432 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20486), .B1(DATAI_17_), 
        .B2(n20531), .ZN(n21001) );
  NAND2_X1 U23433 ( .A1(n20533), .A2(n20506), .ZN(n20921) );
  OAI22_X1 U23434 ( .A1(n21071), .A2(n21047), .B1(n20921), .B2(n20534), .ZN(
        n20507) );
  INV_X1 U23435 ( .A(n20507), .ZN(n20510) );
  NOR2_X2 U23436 ( .A1(n20653), .A2(n20508), .ZN(n21042) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20538), .B1(
        n21042), .B2(n20537), .ZN(n20509) );
  OAI211_X1 U23438 ( .C1(n21001), .C2(n20566), .A(n20510), .B(n20509), .ZN(
        P1_U3034) );
  AOI22_X1 U23439 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20486), .B1(DATAI_18_), 
        .B2(n20531), .ZN(n21005) );
  OAI22_X1 U23440 ( .A1(n21071), .A2(n21053), .B1(n20925), .B2(n20534), .ZN(
        n20511) );
  INV_X1 U23441 ( .A(n20511), .ZN(n20514) );
  NOR2_X2 U23442 ( .A1(n20653), .A2(n20512), .ZN(n21048) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20538), .B1(
        n21048), .B2(n20537), .ZN(n20513) );
  OAI211_X1 U23444 ( .C1(n21005), .C2(n20566), .A(n20514), .B(n20513), .ZN(
        P1_U3035) );
  AOI22_X1 U23445 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20486), .B1(DATAI_27_), 
        .B2(n20531), .ZN(n20972) );
  NAND2_X1 U23446 ( .A1(n20533), .A2(n12892), .ZN(n20929) );
  OAI22_X1 U23447 ( .A1(n21071), .A2(n20972), .B1(n20929), .B2(n20534), .ZN(
        n20515) );
  INV_X1 U23448 ( .A(n20515), .ZN(n20518) );
  NOR2_X2 U23449 ( .A1(n20653), .A2(n20516), .ZN(n21054) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20538), .B1(
        n21054), .B2(n20537), .ZN(n20517) );
  OAI211_X1 U23451 ( .C1(n21059), .C2(n20566), .A(n20518), .B(n20517), .ZN(
        P1_U3036) );
  AOI22_X1 U23452 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20486), .B1(DATAI_20_), 
        .B2(n20531), .ZN(n21011) );
  NAND2_X1 U23453 ( .A1(n20533), .A2(n12812), .ZN(n20933) );
  OAI22_X1 U23454 ( .A1(n21071), .A2(n21065), .B1(n20933), .B2(n20534), .ZN(
        n20519) );
  INV_X1 U23455 ( .A(n20519), .ZN(n20522) );
  NOR2_X2 U23456 ( .A1(n20653), .A2(n20520), .ZN(n21060) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20538), .B1(
        n21060), .B2(n20537), .ZN(n20521) );
  OAI211_X1 U23458 ( .C1(n21011), .C2(n20566), .A(n20522), .B(n20521), .ZN(
        P1_U3037) );
  AOI22_X1 U23459 ( .A1(DATAI_21_), .A2(n20531), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20486), .ZN(n21072) );
  AOI22_X1 U23460 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20486), .B1(DATAI_29_), 
        .B2(n20531), .ZN(n20977) );
  NAND2_X1 U23461 ( .A1(n20533), .A2(n12813), .ZN(n20937) );
  OAI22_X1 U23462 ( .A1(n21071), .A2(n9923), .B1(n20937), .B2(n20534), .ZN(
        n20523) );
  INV_X1 U23463 ( .A(n20523), .ZN(n20526) );
  NOR2_X2 U23464 ( .A1(n20653), .A2(n20524), .ZN(n21066) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20538), .B1(
        n21066), .B2(n20537), .ZN(n20525) );
  OAI211_X1 U23466 ( .C1(n9921), .C2(n20566), .A(n20526), .B(n20525), .ZN(
        P1_U3038) );
  AOI22_X1 U23467 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20486), .B1(DATAI_30_), 
        .B2(n20531), .ZN(n21078) );
  NAND2_X1 U23468 ( .A1(n20533), .A2(n12819), .ZN(n20941) );
  OAI22_X1 U23469 ( .A1(n21071), .A2(n9925), .B1(n20941), .B2(n20534), .ZN(
        n20527) );
  INV_X1 U23470 ( .A(n20527), .ZN(n20530) );
  NOR2_X2 U23471 ( .A1(n20653), .A2(n20528), .ZN(n21073) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20538), .B1(
        n21073), .B2(n20537), .ZN(n20529) );
  OAI211_X1 U23473 ( .C1(n21016), .C2(n20566), .A(n20530), .B(n20529), .ZN(
        P1_U3039) );
  AOI22_X1 U23474 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20486), .B1(DATAI_23_), 
        .B2(n20531), .ZN(n21024) );
  NAND2_X1 U23475 ( .A1(n20533), .A2(n20532), .ZN(n20946) );
  OAI22_X1 U23476 ( .A1(n21071), .A2(n21089), .B1(n20946), .B2(n20534), .ZN(
        n20535) );
  INV_X1 U23477 ( .A(n20535), .ZN(n20540) );
  NOR2_X2 U23478 ( .A1(n20653), .A2(n20536), .ZN(n21080) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20538), .B1(
        n21080), .B2(n20537), .ZN(n20539) );
  OAI211_X1 U23480 ( .C1(n21024), .C2(n20566), .A(n20540), .B(n20539), .ZN(
        P1_U3040) );
  NOR2_X1 U23481 ( .A1(n20953), .A2(n20543), .ZN(n20562) );
  INV_X1 U23482 ( .A(n20610), .ZN(n20542) );
  INV_X1 U23483 ( .A(n20541), .ZN(n20954) );
  AOI21_X1 U23484 ( .B1(n20542), .B2(n20954), .A(n20562), .ZN(n20544) );
  OAI22_X1 U23485 ( .A1(n20544), .A2(n21030), .B1(n20543), .B2(n13022), .ZN(
        n20561) );
  AOI22_X1 U23486 ( .A1(n21032), .A2(n20562), .B1(n21031), .B2(n20561), .ZN(
        n20548) );
  INV_X1 U23487 ( .A(n20543), .ZN(n20546) );
  INV_X1 U23488 ( .A(n20605), .ZN(n20613) );
  OAI21_X1 U23489 ( .B1(n20613), .B2(n20804), .A(n20544), .ZN(n20545) );
  INV_X1 U23490 ( .A(n21041), .ZN(n20961) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20563), .B1(
        n20570), .B2(n20961), .ZN(n20547) );
  OAI211_X1 U23492 ( .C1(n20964), .C2(n20566), .A(n20548), .B(n20547), .ZN(
        P1_U3041) );
  AOI22_X1 U23493 ( .A1(n21043), .A2(n20562), .B1(n21042), .B2(n20561), .ZN(
        n20550) );
  INV_X1 U23494 ( .A(n21001), .ZN(n21044) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20563), .B1(
        n20570), .B2(n21044), .ZN(n20549) );
  OAI211_X1 U23496 ( .C1(n21047), .C2(n20566), .A(n20550), .B(n20549), .ZN(
        P1_U3042) );
  AOI22_X1 U23497 ( .A1(n21049), .A2(n20562), .B1(n21048), .B2(n20561), .ZN(
        n20552) );
  INV_X1 U23498 ( .A(n21005), .ZN(n21050) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20563), .B1(
        n20570), .B2(n21050), .ZN(n20551) );
  OAI211_X1 U23500 ( .C1(n21053), .C2(n20566), .A(n20552), .B(n20551), .ZN(
        P1_U3043) );
  AOI22_X1 U23501 ( .A1(n21055), .A2(n20562), .B1(n21054), .B2(n20561), .ZN(
        n20554) );
  INV_X1 U23502 ( .A(n21059), .ZN(n20969) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20563), .B1(
        n20570), .B2(n20969), .ZN(n20553) );
  OAI211_X1 U23504 ( .C1(n20972), .C2(n20566), .A(n20554), .B(n20553), .ZN(
        P1_U3044) );
  AOI22_X1 U23505 ( .A1(n21061), .A2(n20562), .B1(n21060), .B2(n20561), .ZN(
        n20556) );
  INV_X1 U23506 ( .A(n21011), .ZN(n21062) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20563), .B1(
        n20570), .B2(n21062), .ZN(n20555) );
  OAI211_X1 U23508 ( .C1(n21065), .C2(n20566), .A(n20556), .B(n20555), .ZN(
        P1_U3045) );
  AOI22_X1 U23509 ( .A1(n21067), .A2(n20562), .B1(n21066), .B2(n20561), .ZN(
        n20558) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20563), .B1(
        n20570), .B2(n9920), .ZN(n20557) );
  OAI211_X1 U23511 ( .C1(n9923), .C2(n20566), .A(n20558), .B(n20557), .ZN(
        P1_U3046) );
  AOI22_X1 U23512 ( .A1(n21074), .A2(n20562), .B1(n21073), .B2(n20561), .ZN(
        n20560) );
  INV_X1 U23513 ( .A(n21016), .ZN(n21075) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20563), .B1(
        n20570), .B2(n21075), .ZN(n20559) );
  OAI211_X1 U23515 ( .C1(n9925), .C2(n20566), .A(n20560), .B(n20559), .ZN(
        P1_U3047) );
  AOI22_X1 U23516 ( .A1(n21082), .A2(n20562), .B1(n21080), .B2(n20561), .ZN(
        n20565) );
  INV_X1 U23517 ( .A(n21024), .ZN(n21083) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20563), .B1(
        n20570), .B2(n21083), .ZN(n20564) );
  OAI211_X1 U23519 ( .C1(n21089), .C2(n20566), .A(n20565), .B(n20564), .ZN(
        P1_U3048) );
  NAND3_X1 U23520 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20834), .A3(
        n20830), .ZN(n20617) );
  NOR2_X1 U23521 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20617), .ZN(
        n20572) );
  INV_X1 U23522 ( .A(n20572), .ZN(n20598) );
  OAI22_X1 U23523 ( .A1(n20604), .A2(n20964), .B1(n20598), .B2(n20906), .ZN(
        n20569) );
  INV_X1 U23524 ( .A(n20569), .ZN(n20579) );
  NOR2_X1 U23525 ( .A1(n20570), .A2(n21030), .ZN(n20571) );
  NOR2_X1 U23526 ( .A1(n21030), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20705) );
  NOR2_X1 U23527 ( .A1(n20610), .A2(n14871), .ZN(n20575) );
  OR2_X1 U23528 ( .A1(n20835), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20712) );
  NAND2_X1 U23529 ( .A1(n20712), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20707) );
  OAI211_X1 U23530 ( .C1(n20913), .C2(n20572), .A(n20707), .B(n20836), .ZN(
        n20573) );
  INV_X1 U23531 ( .A(n20573), .ZN(n20574) );
  INV_X1 U23532 ( .A(n20575), .ZN(n20576) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20601), .B1(
        n21031), .B2(n20600), .ZN(n20578) );
  OAI211_X1 U23534 ( .C1(n21041), .C2(n20646), .A(n20579), .B(n20578), .ZN(
        P1_U3049) );
  OAI22_X1 U23535 ( .A1(n20646), .A2(n21001), .B1(n20921), .B2(n20598), .ZN(
        n20580) );
  INV_X1 U23536 ( .A(n20580), .ZN(n20582) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20601), .B1(
        n21042), .B2(n20600), .ZN(n20581) );
  OAI211_X1 U23538 ( .C1(n21047), .C2(n20604), .A(n20582), .B(n20581), .ZN(
        P1_U3050) );
  OAI22_X1 U23539 ( .A1(n20604), .A2(n21053), .B1(n20598), .B2(n20925), .ZN(
        n20583) );
  INV_X1 U23540 ( .A(n20583), .ZN(n20585) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20601), .B1(
        n21048), .B2(n20600), .ZN(n20584) );
  OAI211_X1 U23542 ( .C1(n21005), .C2(n20646), .A(n20585), .B(n20584), .ZN(
        P1_U3051) );
  OAI22_X1 U23543 ( .A1(n20604), .A2(n20972), .B1(n20598), .B2(n20929), .ZN(
        n20586) );
  INV_X1 U23544 ( .A(n20586), .ZN(n20588) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20601), .B1(
        n21054), .B2(n20600), .ZN(n20587) );
  OAI211_X1 U23546 ( .C1(n21059), .C2(n20646), .A(n20588), .B(n20587), .ZN(
        P1_U3052) );
  OAI22_X1 U23547 ( .A1(n20646), .A2(n21011), .B1(n20598), .B2(n20933), .ZN(
        n20589) );
  INV_X1 U23548 ( .A(n20589), .ZN(n20591) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20601), .B1(
        n21060), .B2(n20600), .ZN(n20590) );
  OAI211_X1 U23550 ( .C1(n21065), .C2(n20604), .A(n20591), .B(n20590), .ZN(
        P1_U3053) );
  OAI22_X1 U23551 ( .A1(n20646), .A2(n9921), .B1(n20598), .B2(n20937), .ZN(
        n20592) );
  INV_X1 U23552 ( .A(n20592), .ZN(n20594) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20601), .B1(
        n21066), .B2(n20600), .ZN(n20593) );
  OAI211_X1 U23554 ( .C1(n9923), .C2(n20604), .A(n20594), .B(n20593), .ZN(
        P1_U3054) );
  OAI22_X1 U23555 ( .A1(n20604), .A2(n9925), .B1(n20598), .B2(n20941), .ZN(
        n20595) );
  INV_X1 U23556 ( .A(n20595), .ZN(n20597) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20601), .B1(
        n21073), .B2(n20600), .ZN(n20596) );
  OAI211_X1 U23558 ( .C1(n21016), .C2(n20646), .A(n20597), .B(n20596), .ZN(
        P1_U3055) );
  OAI22_X1 U23559 ( .A1(n20646), .A2(n21024), .B1(n20598), .B2(n20946), .ZN(
        n20599) );
  INV_X1 U23560 ( .A(n20599), .ZN(n20603) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20601), .B1(
        n21080), .B2(n20600), .ZN(n20602) );
  OAI211_X1 U23562 ( .C1(n21089), .C2(n20604), .A(n20603), .B(n20602), .ZN(
        P1_U3056) );
  INV_X1 U23563 ( .A(n20606), .ZN(n20874) );
  NAND2_X1 U23564 ( .A1(n20874), .A2(n20834), .ZN(n20640) );
  OAI22_X1 U23565 ( .A1(n20646), .A2(n20964), .B1(n20906), .B2(n20640), .ZN(
        n20607) );
  INV_X1 U23566 ( .A(n20607), .ZN(n20621) );
  AND2_X1 U23567 ( .A1(n13020), .A2(n10368), .ZN(n20743) );
  INV_X1 U23568 ( .A(n20743), .ZN(n20609) );
  OR2_X1 U23569 ( .A1(n20610), .A2(n20609), .ZN(n20611) );
  INV_X1 U23570 ( .A(n20619), .ZN(n20616) );
  INV_X1 U23571 ( .A(n21035), .ZN(n20614) );
  AOI21_X1 U23572 ( .B1(n21030), .B2(n20617), .A(n20614), .ZN(n20615) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20643), .B1(
        n21031), .B2(n20642), .ZN(n20620) );
  OAI211_X1 U23574 ( .C1(n21041), .C2(n20676), .A(n20621), .B(n20620), .ZN(
        P1_U3057) );
  OAI22_X1 U23575 ( .A1(n20676), .A2(n21001), .B1(n20921), .B2(n20640), .ZN(
        n20622) );
  INV_X1 U23576 ( .A(n20622), .ZN(n20624) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20643), .B1(
        n21042), .B2(n20642), .ZN(n20623) );
  OAI211_X1 U23578 ( .C1(n21047), .C2(n20646), .A(n20624), .B(n20623), .ZN(
        P1_U3058) );
  OAI22_X1 U23579 ( .A1(n20646), .A2(n21053), .B1(n20640), .B2(n20925), .ZN(
        n20625) );
  INV_X1 U23580 ( .A(n20625), .ZN(n20627) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20643), .B1(
        n21048), .B2(n20642), .ZN(n20626) );
  OAI211_X1 U23582 ( .C1(n21005), .C2(n20676), .A(n20627), .B(n20626), .ZN(
        P1_U3059) );
  OAI22_X1 U23583 ( .A1(n20676), .A2(n21059), .B1(n20640), .B2(n20929), .ZN(
        n20628) );
  INV_X1 U23584 ( .A(n20628), .ZN(n20630) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20643), .B1(
        n21054), .B2(n20642), .ZN(n20629) );
  OAI211_X1 U23586 ( .C1(n20972), .C2(n20646), .A(n20630), .B(n20629), .ZN(
        P1_U3060) );
  OAI22_X1 U23587 ( .A1(n20676), .A2(n21011), .B1(n20933), .B2(n20640), .ZN(
        n20631) );
  INV_X1 U23588 ( .A(n20631), .ZN(n20633) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20643), .B1(
        n21060), .B2(n20642), .ZN(n20632) );
  OAI211_X1 U23590 ( .C1(n21065), .C2(n20646), .A(n20633), .B(n20632), .ZN(
        P1_U3061) );
  OAI22_X1 U23591 ( .A1(n20676), .A2(n9921), .B1(n20937), .B2(n20640), .ZN(
        n20634) );
  INV_X1 U23592 ( .A(n20634), .ZN(n20636) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20643), .B1(
        n21066), .B2(n20642), .ZN(n20635) );
  OAI211_X1 U23594 ( .C1(n9923), .C2(n20646), .A(n20636), .B(n20635), .ZN(
        P1_U3062) );
  OAI22_X1 U23595 ( .A1(n20676), .A2(n21016), .B1(n20640), .B2(n20941), .ZN(
        n20637) );
  INV_X1 U23596 ( .A(n20637), .ZN(n20639) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20643), .B1(
        n21073), .B2(n20642), .ZN(n20638) );
  OAI211_X1 U23598 ( .C1(n9925), .C2(n20646), .A(n20639), .B(n20638), .ZN(
        P1_U3063) );
  OAI22_X1 U23599 ( .A1(n20676), .A2(n21024), .B1(n20946), .B2(n20640), .ZN(
        n20641) );
  INV_X1 U23600 ( .A(n20641), .ZN(n20645) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20643), .B1(
        n21080), .B2(n20642), .ZN(n20644) );
  OAI211_X1 U23602 ( .C1(n21089), .C2(n20646), .A(n20645), .B(n20644), .ZN(
        P1_U3064) );
  NAND3_X1 U23603 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20834), .A3(
        n20905), .ZN(n20677) );
  NOR2_X1 U23604 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20677), .ZN(
        n20672) );
  INV_X1 U23605 ( .A(n20647), .ZN(n20989) );
  NOR2_X1 U23606 ( .A1(n12949), .A2(n20648), .ZN(n20744) );
  NAND3_X1 U23607 ( .A1(n20744), .A2(n20908), .A3(n14871), .ZN(n20649) );
  OAI21_X1 U23608 ( .B1(n20989), .B2(n20650), .A(n20649), .ZN(n20671) );
  AOI22_X1 U23609 ( .A1(n21032), .A2(n20672), .B1(n21031), .B2(n20671), .ZN(
        n20657) );
  AOI21_X1 U23610 ( .B1(n20676), .B2(n20703), .A(n20832), .ZN(n20651) );
  AOI21_X1 U23611 ( .B1(n20744), .B2(n14871), .A(n20651), .ZN(n20652) );
  NOR2_X1 U23612 ( .A1(n20652), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20655) );
  INV_X1 U23613 ( .A(n20676), .ZN(n20668) );
  INV_X1 U23614 ( .A(n20964), .ZN(n21038) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20673), .B1(
        n20668), .B2(n21038), .ZN(n20656) );
  OAI211_X1 U23616 ( .C1(n21041), .C2(n20703), .A(n20657), .B(n20656), .ZN(
        P1_U3065) );
  AOI22_X1 U23617 ( .A1(n21043), .A2(n20672), .B1(n21042), .B2(n20671), .ZN(
        n20659) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20673), .B1(
        n20692), .B2(n21044), .ZN(n20658) );
  OAI211_X1 U23619 ( .C1(n21047), .C2(n20676), .A(n20659), .B(n20658), .ZN(
        P1_U3066) );
  AOI22_X1 U23620 ( .A1(n21049), .A2(n20672), .B1(n21048), .B2(n20671), .ZN(
        n20661) );
  INV_X1 U23621 ( .A(n21053), .ZN(n21002) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20673), .B1(
        n20668), .B2(n21002), .ZN(n20660) );
  OAI211_X1 U23623 ( .C1(n21005), .C2(n20703), .A(n20661), .B(n20660), .ZN(
        P1_U3067) );
  AOI22_X1 U23624 ( .A1(n21055), .A2(n20672), .B1(n21054), .B2(n20671), .ZN(
        n20663) );
  INV_X1 U23625 ( .A(n20972), .ZN(n21056) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20673), .B1(
        n20668), .B2(n21056), .ZN(n20662) );
  OAI211_X1 U23627 ( .C1(n21059), .C2(n20703), .A(n20663), .B(n20662), .ZN(
        P1_U3068) );
  AOI22_X1 U23628 ( .A1(n21061), .A2(n20672), .B1(n21060), .B2(n20671), .ZN(
        n20665) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20673), .B1(
        n20692), .B2(n21062), .ZN(n20664) );
  OAI211_X1 U23630 ( .C1(n21065), .C2(n20676), .A(n20665), .B(n20664), .ZN(
        P1_U3069) );
  AOI22_X1 U23631 ( .A1(n21067), .A2(n20672), .B1(n21066), .B2(n20671), .ZN(
        n20667) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20673), .B1(
        n20692), .B2(n9920), .ZN(n20666) );
  OAI211_X1 U23633 ( .C1(n9923), .C2(n20676), .A(n20667), .B(n20666), .ZN(
        P1_U3070) );
  AOI22_X1 U23634 ( .A1(n21074), .A2(n20672), .B1(n21073), .B2(n20671), .ZN(
        n20670) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20673), .B1(
        n20668), .B2(n9924), .ZN(n20669) );
  OAI211_X1 U23636 ( .C1(n21016), .C2(n20703), .A(n20670), .B(n20669), .ZN(
        P1_U3071) );
  AOI22_X1 U23637 ( .A1(n21082), .A2(n20672), .B1(n21080), .B2(n20671), .ZN(
        n20675) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20673), .B1(
        n20692), .B2(n21083), .ZN(n20674) );
  OAI211_X1 U23639 ( .C1(n21089), .C2(n20676), .A(n20675), .B(n20674), .ZN(
        P1_U3072) );
  NOR2_X1 U23640 ( .A1(n20953), .A2(n20677), .ZN(n20698) );
  AOI21_X1 U23641 ( .B1(n20744), .B2(n20954), .A(n20698), .ZN(n20678) );
  OAI22_X1 U23642 ( .A1(n20678), .A2(n21030), .B1(n20677), .B2(n13022), .ZN(
        n20697) );
  AOI22_X1 U23643 ( .A1(n21032), .A2(n20698), .B1(n21031), .B2(n20697), .ZN(
        n20683) );
  INV_X1 U23644 ( .A(n20677), .ZN(n20681) );
  INV_X1 U23645 ( .A(n20742), .ZN(n20679) );
  OAI21_X1 U23646 ( .B1(n20679), .B2(n20804), .A(n20678), .ZN(n20680) );
  OAI221_X1 U23647 ( .B1(n20908), .B2(n20681), .C1(n21030), .C2(n20680), .A(
        n21035), .ZN(n20700) );
  INV_X1 U23648 ( .A(n20741), .ZN(n20699) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n20961), .ZN(n20682) );
  OAI211_X1 U23650 ( .C1(n20964), .C2(n20703), .A(n20683), .B(n20682), .ZN(
        P1_U3073) );
  AOI22_X1 U23651 ( .A1(n21043), .A2(n20698), .B1(n21042), .B2(n20697), .ZN(
        n20685) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n21044), .ZN(n20684) );
  OAI211_X1 U23653 ( .C1(n21047), .C2(n20703), .A(n20685), .B(n20684), .ZN(
        P1_U3074) );
  AOI22_X1 U23654 ( .A1(n21049), .A2(n20698), .B1(n21048), .B2(n20697), .ZN(
        n20687) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20700), .B1(
        n20692), .B2(n21002), .ZN(n20686) );
  OAI211_X1 U23656 ( .C1(n21005), .C2(n20741), .A(n20687), .B(n20686), .ZN(
        P1_U3075) );
  AOI22_X1 U23657 ( .A1(n21055), .A2(n20698), .B1(n21054), .B2(n20697), .ZN(
        n20689) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20700), .B1(
        n20692), .B2(n21056), .ZN(n20688) );
  OAI211_X1 U23659 ( .C1(n21059), .C2(n20741), .A(n20689), .B(n20688), .ZN(
        P1_U3076) );
  AOI22_X1 U23660 ( .A1(n21061), .A2(n20698), .B1(n21060), .B2(n20697), .ZN(
        n20691) );
  INV_X1 U23661 ( .A(n21065), .ZN(n21008) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20700), .B1(
        n20692), .B2(n21008), .ZN(n20690) );
  OAI211_X1 U23663 ( .C1(n21011), .C2(n20741), .A(n20691), .B(n20690), .ZN(
        P1_U3077) );
  AOI22_X1 U23664 ( .A1(n21067), .A2(n20698), .B1(n21066), .B2(n20697), .ZN(
        n20694) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20700), .B1(
        n20692), .B2(n9922), .ZN(n20693) );
  OAI211_X1 U23666 ( .C1(n9921), .C2(n20741), .A(n20694), .B(n20693), .ZN(
        P1_U3078) );
  AOI22_X1 U23667 ( .A1(n21074), .A2(n20698), .B1(n21073), .B2(n20697), .ZN(
        n20696) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n21075), .ZN(n20695) );
  OAI211_X1 U23669 ( .C1(n9925), .C2(n20703), .A(n20696), .B(n20695), .ZN(
        P1_U3079) );
  AOI22_X1 U23670 ( .A1(n21082), .A2(n20698), .B1(n21080), .B2(n20697), .ZN(
        n20702) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20700), .B1(
        n20699), .B2(n21083), .ZN(n20701) );
  OAI211_X1 U23672 ( .C1(n21089), .C2(n20703), .A(n20702), .B(n20701), .ZN(
        P1_U3080) );
  INV_X1 U23673 ( .A(n20751), .ZN(n20746) );
  NOR2_X1 U23674 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20746), .ZN(
        n20710) );
  INV_X1 U23675 ( .A(n20710), .ZN(n20735) );
  OAI22_X1 U23676 ( .A1(n20741), .A2(n20964), .B1(n20906), .B2(n20735), .ZN(
        n20704) );
  INV_X1 U23677 ( .A(n20704), .ZN(n20716) );
  NAND3_X1 U23678 ( .A1(n20774), .A2(n20741), .A3(n20908), .ZN(n20706) );
  INV_X1 U23679 ( .A(n20705), .ZN(n20909) );
  NAND2_X1 U23680 ( .A1(n20706), .A2(n20909), .ZN(n20711) );
  NAND2_X1 U23681 ( .A1(n20744), .A2(n20988), .ZN(n20713) );
  INV_X1 U23682 ( .A(n20707), .ZN(n20708) );
  AOI21_X1 U23683 ( .B1(n20711), .B2(n20713), .A(n20708), .ZN(n20709) );
  INV_X1 U23684 ( .A(n20711), .ZN(n20714) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20738), .B1(
        n21031), .B2(n20737), .ZN(n20715) );
  OAI211_X1 U23686 ( .C1(n21041), .C2(n20774), .A(n20716), .B(n20715), .ZN(
        P1_U3081) );
  OAI22_X1 U23687 ( .A1(n20774), .A2(n21001), .B1(n20735), .B2(n20921), .ZN(
        n20717) );
  INV_X1 U23688 ( .A(n20717), .ZN(n20719) );
  AOI22_X1 U23689 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20738), .B1(
        n21042), .B2(n20737), .ZN(n20718) );
  OAI211_X1 U23690 ( .C1(n21047), .C2(n20741), .A(n20719), .B(n20718), .ZN(
        P1_U3082) );
  OAI22_X1 U23691 ( .A1(n20741), .A2(n21053), .B1(n20925), .B2(n20735), .ZN(
        n20720) );
  INV_X1 U23692 ( .A(n20720), .ZN(n20722) );
  AOI22_X1 U23693 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20738), .B1(
        n21048), .B2(n20737), .ZN(n20721) );
  OAI211_X1 U23694 ( .C1(n21005), .C2(n20774), .A(n20722), .B(n20721), .ZN(
        P1_U3083) );
  OAI22_X1 U23695 ( .A1(n20774), .A2(n21059), .B1(n20929), .B2(n20735), .ZN(
        n20723) );
  INV_X1 U23696 ( .A(n20723), .ZN(n20725) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20738), .B1(
        n21054), .B2(n20737), .ZN(n20724) );
  OAI211_X1 U23698 ( .C1(n20972), .C2(n20741), .A(n20725), .B(n20724), .ZN(
        P1_U3084) );
  OAI22_X1 U23699 ( .A1(n20741), .A2(n21065), .B1(n20933), .B2(n20735), .ZN(
        n20726) );
  INV_X1 U23700 ( .A(n20726), .ZN(n20728) );
  AOI22_X1 U23701 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20738), .B1(
        n21060), .B2(n20737), .ZN(n20727) );
  OAI211_X1 U23702 ( .C1(n21011), .C2(n20774), .A(n20728), .B(n20727), .ZN(
        P1_U3085) );
  OAI22_X1 U23703 ( .A1(n20741), .A2(n9923), .B1(n20937), .B2(n20735), .ZN(
        n20729) );
  INV_X1 U23704 ( .A(n20729), .ZN(n20731) );
  AOI22_X1 U23705 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20738), .B1(
        n21066), .B2(n20737), .ZN(n20730) );
  OAI211_X1 U23706 ( .C1(n9921), .C2(n20774), .A(n20731), .B(n20730), .ZN(
        P1_U3086) );
  OAI22_X1 U23707 ( .A1(n20741), .A2(n9925), .B1(n20941), .B2(n20735), .ZN(
        n20732) );
  INV_X1 U23708 ( .A(n20732), .ZN(n20734) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20738), .B1(
        n21073), .B2(n20737), .ZN(n20733) );
  OAI211_X1 U23710 ( .C1(n21016), .C2(n20774), .A(n20734), .B(n20733), .ZN(
        P1_U3087) );
  OAI22_X1 U23711 ( .A1(n20774), .A2(n21024), .B1(n20735), .B2(n20946), .ZN(
        n20736) );
  INV_X1 U23712 ( .A(n20736), .ZN(n20740) );
  AOI22_X1 U23713 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20738), .B1(
        n21080), .B2(n20737), .ZN(n20739) );
  OAI211_X1 U23714 ( .C1(n21089), .C2(n20741), .A(n20740), .B(n20739), .ZN(
        P1_U3088) );
  INV_X1 U23715 ( .A(n20797), .ZN(n20768) );
  INV_X1 U23716 ( .A(n20745), .ZN(n20770) );
  NAND2_X1 U23717 ( .A1(n20743), .A2(n20908), .ZN(n21026) );
  INV_X1 U23718 ( .A(n20744), .ZN(n20747) );
  OAI222_X1 U23719 ( .A1(n21026), .A2(n20747), .B1(n13022), .B2(n20746), .C1(
        n20745), .C2(n21030), .ZN(n20769) );
  AOI22_X1 U23720 ( .A1(n21032), .A2(n20770), .B1(n21031), .B2(n20769), .ZN(
        n20754) );
  NAND3_X1 U23721 ( .A1(n20749), .A2(n20908), .A3(n20748), .ZN(n21034) );
  NOR2_X1 U23722 ( .A1(n21034), .A2(n20750), .ZN(n20752) );
  INV_X1 U23723 ( .A(n20774), .ZN(n20765) );
  AOI22_X1 U23724 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n20765), .B2(n21038), .ZN(n20753) );
  OAI211_X1 U23725 ( .C1(n21041), .C2(n20768), .A(n20754), .B(n20753), .ZN(
        P1_U3089) );
  AOI22_X1 U23726 ( .A1(n21043), .A2(n20770), .B1(n21042), .B2(n20769), .ZN(
        n20756) );
  INV_X1 U23727 ( .A(n21047), .ZN(n20998) );
  AOI22_X1 U23728 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n20765), .B2(n20998), .ZN(n20755) );
  OAI211_X1 U23729 ( .C1(n21001), .C2(n20768), .A(n20756), .B(n20755), .ZN(
        P1_U3090) );
  AOI22_X1 U23730 ( .A1(n21049), .A2(n20770), .B1(n21048), .B2(n20769), .ZN(
        n20758) );
  AOI22_X1 U23731 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n20797), .B2(n21050), .ZN(n20757) );
  OAI211_X1 U23732 ( .C1(n21053), .C2(n20774), .A(n20758), .B(n20757), .ZN(
        P1_U3091) );
  AOI22_X1 U23733 ( .A1(n21055), .A2(n20770), .B1(n21054), .B2(n20769), .ZN(
        n20760) );
  AOI22_X1 U23734 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n20765), .B2(n21056), .ZN(n20759) );
  OAI211_X1 U23735 ( .C1(n21059), .C2(n20768), .A(n20760), .B(n20759), .ZN(
        P1_U3092) );
  AOI22_X1 U23736 ( .A1(n21061), .A2(n20770), .B1(n21060), .B2(n20769), .ZN(
        n20762) );
  AOI22_X1 U23737 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n20797), .B2(n21062), .ZN(n20761) );
  OAI211_X1 U23738 ( .C1(n21065), .C2(n20774), .A(n20762), .B(n20761), .ZN(
        P1_U3093) );
  AOI22_X1 U23739 ( .A1(n21067), .A2(n20770), .B1(n21066), .B2(n20769), .ZN(
        n20764) );
  AOI22_X1 U23740 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n20797), .B2(n9920), .ZN(n20763) );
  OAI211_X1 U23741 ( .C1(n9923), .C2(n20774), .A(n20764), .B(n20763), .ZN(
        P1_U3094) );
  AOI22_X1 U23742 ( .A1(n21074), .A2(n20770), .B1(n21073), .B2(n20769), .ZN(
        n20767) );
  AOI22_X1 U23743 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n20765), .B2(n9924), .ZN(n20766) );
  OAI211_X1 U23744 ( .C1(n21016), .C2(n20768), .A(n20767), .B(n20766), .ZN(
        P1_U3095) );
  AOI22_X1 U23745 ( .A1(n21082), .A2(n20770), .B1(n21080), .B2(n20769), .ZN(
        n20773) );
  AOI22_X1 U23746 ( .A1(n20771), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n20797), .B2(n21083), .ZN(n20772) );
  OAI211_X1 U23747 ( .C1(n21089), .C2(n20774), .A(n20773), .B(n20772), .ZN(
        P1_U3096) );
  INV_X1 U23748 ( .A(n20873), .ZN(n20878) );
  NAND3_X1 U23749 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20830), .A3(
        n20905), .ZN(n20802) );
  NOR2_X1 U23750 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20802), .ZN(
        n20796) );
  NAND2_X1 U23751 ( .A1(n20775), .A2(n12949), .ZN(n20876) );
  INV_X1 U23752 ( .A(n20876), .ZN(n20801) );
  AOI21_X1 U23753 ( .B1(n20801), .B2(n14871), .A(n20796), .ZN(n20778) );
  NAND2_X1 U23754 ( .A1(n20776), .A2(n20835), .ZN(n20916) );
  OAI22_X1 U23755 ( .A1(n20778), .A2(n21030), .B1(n20841), .B2(n20916), .ZN(
        n20795) );
  AOI22_X1 U23756 ( .A1(n21032), .A2(n20796), .B1(n21031), .B2(n20795), .ZN(
        n20782) );
  INV_X1 U23757 ( .A(n20828), .ZN(n20777) );
  OAI21_X1 U23758 ( .B1(n20777), .B2(n20797), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20779) );
  NAND2_X1 U23759 ( .A1(n20779), .A2(n20778), .ZN(n20780) );
  AOI22_X1 U23760 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n21038), .ZN(n20781) );
  OAI211_X1 U23761 ( .C1(n21041), .C2(n20828), .A(n20782), .B(n20781), .ZN(
        P1_U3097) );
  AOI22_X1 U23762 ( .A1(n21043), .A2(n20796), .B1(n21042), .B2(n20795), .ZN(
        n20784) );
  AOI22_X1 U23763 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n20998), .ZN(n20783) );
  OAI211_X1 U23764 ( .C1(n21001), .C2(n20828), .A(n20784), .B(n20783), .ZN(
        P1_U3098) );
  AOI22_X1 U23765 ( .A1(n21049), .A2(n20796), .B1(n21048), .B2(n20795), .ZN(
        n20786) );
  AOI22_X1 U23766 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n21002), .ZN(n20785) );
  OAI211_X1 U23767 ( .C1(n21005), .C2(n20828), .A(n20786), .B(n20785), .ZN(
        P1_U3099) );
  AOI22_X1 U23768 ( .A1(n21055), .A2(n20796), .B1(n21054), .B2(n20795), .ZN(
        n20788) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n21056), .ZN(n20787) );
  OAI211_X1 U23770 ( .C1(n21059), .C2(n20828), .A(n20788), .B(n20787), .ZN(
        P1_U3100) );
  AOI22_X1 U23771 ( .A1(n21061), .A2(n20796), .B1(n21060), .B2(n20795), .ZN(
        n20790) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n21008), .ZN(n20789) );
  OAI211_X1 U23773 ( .C1(n21011), .C2(n20828), .A(n20790), .B(n20789), .ZN(
        P1_U3101) );
  AOI22_X1 U23774 ( .A1(n21067), .A2(n20796), .B1(n21066), .B2(n20795), .ZN(
        n20792) );
  AOI22_X1 U23775 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n9922), .ZN(n20791) );
  OAI211_X1 U23776 ( .C1(n9921), .C2(n20828), .A(n20792), .B(n20791), .ZN(
        P1_U3102) );
  AOI22_X1 U23777 ( .A1(n21074), .A2(n20796), .B1(n21073), .B2(n20795), .ZN(
        n20794) );
  AOI22_X1 U23778 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n9924), .ZN(n20793) );
  OAI211_X1 U23779 ( .C1(n21016), .C2(n20828), .A(n20794), .B(n20793), .ZN(
        P1_U3103) );
  AOI22_X1 U23780 ( .A1(n21082), .A2(n20796), .B1(n21080), .B2(n20795), .ZN(
        n20800) );
  INV_X1 U23781 ( .A(n21089), .ZN(n21019) );
  AOI22_X1 U23782 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n21019), .ZN(n20799) );
  OAI211_X1 U23783 ( .C1(n21024), .C2(n20828), .A(n20800), .B(n20799), .ZN(
        P1_U3104) );
  NOR2_X1 U23784 ( .A1(n20953), .A2(n20802), .ZN(n20823) );
  AOI21_X1 U23785 ( .B1(n20801), .B2(n20954), .A(n20823), .ZN(n20803) );
  OAI22_X1 U23786 ( .A1(n20803), .A2(n21030), .B1(n20802), .B2(n13022), .ZN(
        n20822) );
  AOI22_X1 U23787 ( .A1(n21032), .A2(n20823), .B1(n21031), .B2(n20822), .ZN(
        n20809) );
  INV_X1 U23788 ( .A(n20802), .ZN(n20806) );
  OAI21_X1 U23789 ( .B1(n20873), .B2(n20804), .A(n20803), .ZN(n20805) );
  OAI221_X1 U23790 ( .B1(n20908), .B2(n20806), .C1(n21030), .C2(n20805), .A(
        n21035), .ZN(n20825) );
  AOI22_X1 U23791 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20825), .B1(
        n20824), .B2(n20961), .ZN(n20808) );
  OAI211_X1 U23792 ( .C1(n20964), .C2(n20828), .A(n20809), .B(n20808), .ZN(
        P1_U3105) );
  AOI22_X1 U23793 ( .A1(n21043), .A2(n20823), .B1(n21042), .B2(n20822), .ZN(
        n20811) );
  AOI22_X1 U23794 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20825), .B1(
        n20824), .B2(n21044), .ZN(n20810) );
  OAI211_X1 U23795 ( .C1(n21047), .C2(n20828), .A(n20811), .B(n20810), .ZN(
        P1_U3106) );
  AOI22_X1 U23796 ( .A1(n21049), .A2(n20823), .B1(n21048), .B2(n20822), .ZN(
        n20813) );
  AOI22_X1 U23797 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20825), .B1(
        n20824), .B2(n21050), .ZN(n20812) );
  OAI211_X1 U23798 ( .C1(n21053), .C2(n20828), .A(n20813), .B(n20812), .ZN(
        P1_U3107) );
  AOI22_X1 U23799 ( .A1(n21055), .A2(n20823), .B1(n21054), .B2(n20822), .ZN(
        n20815) );
  AOI22_X1 U23800 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20825), .B1(
        n20824), .B2(n20969), .ZN(n20814) );
  OAI211_X1 U23801 ( .C1(n20972), .C2(n20828), .A(n20815), .B(n20814), .ZN(
        P1_U3108) );
  AOI22_X1 U23802 ( .A1(n21061), .A2(n20823), .B1(n21060), .B2(n20822), .ZN(
        n20817) );
  AOI22_X1 U23803 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20825), .B1(
        n20824), .B2(n21062), .ZN(n20816) );
  OAI211_X1 U23804 ( .C1(n21065), .C2(n20828), .A(n20817), .B(n20816), .ZN(
        P1_U3109) );
  AOI22_X1 U23805 ( .A1(n21067), .A2(n20823), .B1(n21066), .B2(n20822), .ZN(
        n20819) );
  AOI22_X1 U23806 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20825), .B1(
        n20824), .B2(n9920), .ZN(n20818) );
  OAI211_X1 U23807 ( .C1(n9923), .C2(n20828), .A(n20819), .B(n20818), .ZN(
        P1_U3110) );
  AOI22_X1 U23808 ( .A1(n21074), .A2(n20823), .B1(n21073), .B2(n20822), .ZN(
        n20821) );
  AOI22_X1 U23809 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20825), .B1(
        n20824), .B2(n21075), .ZN(n20820) );
  OAI211_X1 U23810 ( .C1(n9925), .C2(n20828), .A(n20821), .B(n20820), .ZN(
        P1_U3111) );
  AOI22_X1 U23811 ( .A1(n21082), .A2(n20823), .B1(n21080), .B2(n20822), .ZN(
        n20827) );
  AOI22_X1 U23812 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20825), .B1(
        n20824), .B2(n21083), .ZN(n20826) );
  OAI211_X1 U23813 ( .C1(n21089), .C2(n20828), .A(n20827), .B(n20826), .ZN(
        P1_U3112) );
  INV_X1 U23814 ( .A(n20986), .ZN(n20829) );
  NAND3_X1 U23815 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20830), .ZN(n20879) );
  NOR2_X1 U23816 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20879), .ZN(
        n20837) );
  INV_X1 U23817 ( .A(n20837), .ZN(n20864) );
  OAI22_X1 U23818 ( .A1(n20865), .A2(n20964), .B1(n20906), .B2(n20864), .ZN(
        n20831) );
  INV_X1 U23819 ( .A(n20831), .ZN(n20845) );
  AOI21_X1 U23820 ( .B1(n20891), .B2(n20865), .A(n20832), .ZN(n20833) );
  NOR2_X1 U23821 ( .A1(n20833), .A2(n21030), .ZN(n20840) );
  OR2_X1 U23822 ( .A1(n20876), .A2(n14871), .ZN(n20842) );
  OR2_X1 U23823 ( .A1(n20835), .A2(n20834), .ZN(n20990) );
  NAND2_X1 U23824 ( .A1(n20990), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20993) );
  OAI211_X1 U23825 ( .C1(n20913), .C2(n20837), .A(n20993), .B(n20836), .ZN(
        n20838) );
  AOI21_X1 U23826 ( .B1(n20840), .B2(n20842), .A(n20838), .ZN(n20839) );
  INV_X1 U23827 ( .A(n20840), .ZN(n20843) );
  AOI22_X1 U23828 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20868), .B1(
        n21031), .B2(n20867), .ZN(n20844) );
  OAI211_X1 U23829 ( .C1(n21041), .C2(n20891), .A(n20845), .B(n20844), .ZN(
        P1_U3113) );
  OAI22_X1 U23830 ( .A1(n20891), .A2(n21001), .B1(n20921), .B2(n20864), .ZN(
        n20846) );
  INV_X1 U23831 ( .A(n20846), .ZN(n20848) );
  AOI22_X1 U23832 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20868), .B1(
        n21042), .B2(n20867), .ZN(n20847) );
  OAI211_X1 U23833 ( .C1(n21047), .C2(n20865), .A(n20848), .B(n20847), .ZN(
        P1_U3114) );
  OAI22_X1 U23834 ( .A1(n20865), .A2(n21053), .B1(n20925), .B2(n20864), .ZN(
        n20849) );
  INV_X1 U23835 ( .A(n20849), .ZN(n20851) );
  AOI22_X1 U23836 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20868), .B1(
        n21048), .B2(n20867), .ZN(n20850) );
  OAI211_X1 U23837 ( .C1(n21005), .C2(n20891), .A(n20851), .B(n20850), .ZN(
        P1_U3115) );
  OAI22_X1 U23838 ( .A1(n20865), .A2(n20972), .B1(n20864), .B2(n20929), .ZN(
        n20852) );
  INV_X1 U23839 ( .A(n20852), .ZN(n20854) );
  AOI22_X1 U23840 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20868), .B1(
        n21054), .B2(n20867), .ZN(n20853) );
  OAI211_X1 U23841 ( .C1(n21059), .C2(n20891), .A(n20854), .B(n20853), .ZN(
        P1_U3116) );
  OAI22_X1 U23842 ( .A1(n20865), .A2(n21065), .B1(n20933), .B2(n20864), .ZN(
        n20855) );
  INV_X1 U23843 ( .A(n20855), .ZN(n20857) );
  AOI22_X1 U23844 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20868), .B1(
        n21060), .B2(n20867), .ZN(n20856) );
  OAI211_X1 U23845 ( .C1(n21011), .C2(n20891), .A(n20857), .B(n20856), .ZN(
        P1_U3117) );
  OAI22_X1 U23846 ( .A1(n20865), .A2(n9923), .B1(n20937), .B2(n20864), .ZN(
        n20858) );
  INV_X1 U23847 ( .A(n20858), .ZN(n20860) );
  AOI22_X1 U23848 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20868), .B1(
        n21066), .B2(n20867), .ZN(n20859) );
  OAI211_X1 U23849 ( .C1(n9921), .C2(n20891), .A(n20860), .B(n20859), .ZN(
        P1_U3118) );
  OAI22_X1 U23850 ( .A1(n20891), .A2(n21016), .B1(n20864), .B2(n20941), .ZN(
        n20861) );
  INV_X1 U23851 ( .A(n20861), .ZN(n20863) );
  AOI22_X1 U23852 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20868), .B1(
        n21073), .B2(n20867), .ZN(n20862) );
  OAI211_X1 U23853 ( .C1(n9925), .C2(n20865), .A(n20863), .B(n20862), .ZN(
        P1_U3119) );
  OAI22_X1 U23854 ( .A1(n20865), .A2(n21089), .B1(n20946), .B2(n20864), .ZN(
        n20866) );
  INV_X1 U23855 ( .A(n20866), .ZN(n20870) );
  AOI22_X1 U23856 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20868), .B1(
        n21080), .B2(n20867), .ZN(n20869) );
  OAI211_X1 U23857 ( .C1(n21024), .C2(n20891), .A(n20870), .B(n20869), .ZN(
        P1_U3120) );
  INV_X1 U23858 ( .A(n20871), .ZN(n20872) );
  NAND2_X1 U23859 ( .A1(n20874), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20875) );
  INV_X1 U23860 ( .A(n20875), .ZN(n20899) );
  OAI222_X1 U23861 ( .A1(n21026), .A2(n20876), .B1(n13022), .B2(n20879), .C1(
        n21030), .C2(n20875), .ZN(n20898) );
  AOI22_X1 U23862 ( .A1(n21032), .A2(n20899), .B1(n21031), .B2(n20898), .ZN(
        n20883) );
  AND2_X1 U23863 ( .A1(n20878), .A2(n20877), .ZN(n20881) );
  INV_X1 U23864 ( .A(n20879), .ZN(n20880) );
  INV_X1 U23865 ( .A(n20891), .ZN(n20900) );
  AOI22_X1 U23866 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20901), .B1(
        n20900), .B2(n21038), .ZN(n20882) );
  OAI211_X1 U23867 ( .C1(n21041), .C2(n20952), .A(n20883), .B(n20882), .ZN(
        P1_U3121) );
  AOI22_X1 U23868 ( .A1(n21043), .A2(n20899), .B1(n21042), .B2(n20898), .ZN(
        n20885) );
  INV_X1 U23869 ( .A(n20952), .ZN(n20888) );
  AOI22_X1 U23870 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20901), .B1(
        n20888), .B2(n21044), .ZN(n20884) );
  OAI211_X1 U23871 ( .C1(n21047), .C2(n20891), .A(n20885), .B(n20884), .ZN(
        P1_U3122) );
  AOI22_X1 U23872 ( .A1(n21049), .A2(n20899), .B1(n21048), .B2(n20898), .ZN(
        n20887) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20901), .B1(
        n20888), .B2(n21050), .ZN(n20886) );
  OAI211_X1 U23874 ( .C1(n21053), .C2(n20891), .A(n20887), .B(n20886), .ZN(
        P1_U3123) );
  AOI22_X1 U23875 ( .A1(n21055), .A2(n20899), .B1(n21054), .B2(n20898), .ZN(
        n20890) );
  AOI22_X1 U23876 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20901), .B1(
        n20888), .B2(n20969), .ZN(n20889) );
  OAI211_X1 U23877 ( .C1(n20972), .C2(n20891), .A(n20890), .B(n20889), .ZN(
        P1_U3124) );
  AOI22_X1 U23878 ( .A1(n21061), .A2(n20899), .B1(n21060), .B2(n20898), .ZN(
        n20893) );
  AOI22_X1 U23879 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20901), .B1(
        n20900), .B2(n21008), .ZN(n20892) );
  OAI211_X1 U23880 ( .C1(n21011), .C2(n20952), .A(n20893), .B(n20892), .ZN(
        P1_U3125) );
  AOI22_X1 U23881 ( .A1(n21067), .A2(n20899), .B1(n21066), .B2(n20898), .ZN(
        n20895) );
  AOI22_X1 U23882 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20901), .B1(
        n20900), .B2(n9922), .ZN(n20894) );
  OAI211_X1 U23883 ( .C1(n9921), .C2(n20952), .A(n20895), .B(n20894), .ZN(
        P1_U3126) );
  AOI22_X1 U23884 ( .A1(n21074), .A2(n20899), .B1(n21073), .B2(n20898), .ZN(
        n20897) );
  AOI22_X1 U23885 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20901), .B1(
        n20900), .B2(n9924), .ZN(n20896) );
  OAI211_X1 U23886 ( .C1(n21016), .C2(n20952), .A(n20897), .B(n20896), .ZN(
        P1_U3127) );
  AOI22_X1 U23887 ( .A1(n21082), .A2(n20899), .B1(n21080), .B2(n20898), .ZN(
        n20903) );
  AOI22_X1 U23888 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20901), .B1(
        n20900), .B2(n21019), .ZN(n20902) );
  OAI211_X1 U23889 ( .C1(n21024), .C2(n20952), .A(n20903), .B(n20902), .ZN(
        P1_U3128) );
  NAND3_X1 U23890 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20905), .ZN(n20956) );
  NOR2_X1 U23891 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20956), .ZN(
        n20914) );
  INV_X1 U23892 ( .A(n20914), .ZN(n20945) );
  OAI22_X1 U23893 ( .A1(n20985), .A2(n21041), .B1(n20906), .B2(n20945), .ZN(
        n20907) );
  INV_X1 U23894 ( .A(n20907), .ZN(n20920) );
  NAND3_X1 U23895 ( .A1(n20952), .A2(n20908), .A3(n20985), .ZN(n20910) );
  NAND2_X1 U23896 ( .A1(n20910), .A2(n20909), .ZN(n20915) );
  NOR2_X1 U23897 ( .A1(n12949), .A2(n20911), .ZN(n21025) );
  NAND2_X1 U23898 ( .A1(n21025), .A2(n14871), .ZN(n20917) );
  AOI22_X1 U23899 ( .A1(n20915), .A2(n20917), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20916), .ZN(n20912) );
  INV_X1 U23900 ( .A(n20915), .ZN(n20918) );
  AOI22_X1 U23901 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20949), .B1(
        n21031), .B2(n20948), .ZN(n20919) );
  OAI211_X1 U23902 ( .C1(n20964), .C2(n20952), .A(n20920), .B(n20919), .ZN(
        P1_U3129) );
  OAI22_X1 U23903 ( .A1(n20985), .A2(n21001), .B1(n20921), .B2(n20945), .ZN(
        n20922) );
  INV_X1 U23904 ( .A(n20922), .ZN(n20924) );
  AOI22_X1 U23905 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20949), .B1(
        n21042), .B2(n20948), .ZN(n20923) );
  OAI211_X1 U23906 ( .C1(n21047), .C2(n20952), .A(n20924), .B(n20923), .ZN(
        P1_U3130) );
  OAI22_X1 U23907 ( .A1(n20985), .A2(n21005), .B1(n20925), .B2(n20945), .ZN(
        n20926) );
  INV_X1 U23908 ( .A(n20926), .ZN(n20928) );
  AOI22_X1 U23909 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20949), .B1(
        n21048), .B2(n20948), .ZN(n20927) );
  OAI211_X1 U23910 ( .C1(n21053), .C2(n20952), .A(n20928), .B(n20927), .ZN(
        P1_U3131) );
  OAI22_X1 U23911 ( .A1(n20985), .A2(n21059), .B1(n20929), .B2(n20945), .ZN(
        n20930) );
  INV_X1 U23912 ( .A(n20930), .ZN(n20932) );
  AOI22_X1 U23913 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20949), .B1(
        n21054), .B2(n20948), .ZN(n20931) );
  OAI211_X1 U23914 ( .C1(n20972), .C2(n20952), .A(n20932), .B(n20931), .ZN(
        P1_U3132) );
  OAI22_X1 U23915 ( .A1(n20985), .A2(n21011), .B1(n20933), .B2(n20945), .ZN(
        n20934) );
  INV_X1 U23916 ( .A(n20934), .ZN(n20936) );
  AOI22_X1 U23917 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20949), .B1(
        n21060), .B2(n20948), .ZN(n20935) );
  OAI211_X1 U23918 ( .C1(n21065), .C2(n20952), .A(n20936), .B(n20935), .ZN(
        P1_U3133) );
  OAI22_X1 U23919 ( .A1(n20985), .A2(n9921), .B1(n20937), .B2(n20945), .ZN(
        n20938) );
  INV_X1 U23920 ( .A(n20938), .ZN(n20940) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20949), .B1(
        n21066), .B2(n20948), .ZN(n20939) );
  OAI211_X1 U23922 ( .C1(n9923), .C2(n20952), .A(n20940), .B(n20939), .ZN(
        P1_U3134) );
  OAI22_X1 U23923 ( .A1(n20985), .A2(n21016), .B1(n20941), .B2(n20945), .ZN(
        n20942) );
  INV_X1 U23924 ( .A(n20942), .ZN(n20944) );
  AOI22_X1 U23925 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20949), .B1(
        n21073), .B2(n20948), .ZN(n20943) );
  OAI211_X1 U23926 ( .C1(n9925), .C2(n20952), .A(n20944), .B(n20943), .ZN(
        P1_U3135) );
  OAI22_X1 U23927 ( .A1(n20985), .A2(n21024), .B1(n20946), .B2(n20945), .ZN(
        n20947) );
  INV_X1 U23928 ( .A(n20947), .ZN(n20951) );
  AOI22_X1 U23929 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20949), .B1(
        n21080), .B2(n20948), .ZN(n20950) );
  OAI211_X1 U23930 ( .C1(n21089), .C2(n20952), .A(n20951), .B(n20950), .ZN(
        P1_U3136) );
  NOR2_X1 U23931 ( .A1(n20953), .A2(n20956), .ZN(n20981) );
  AOI21_X1 U23932 ( .B1(n21025), .B2(n20954), .A(n20981), .ZN(n20955) );
  OAI22_X1 U23933 ( .A1(n20955), .A2(n21030), .B1(n20956), .B2(n13022), .ZN(
        n20980) );
  AOI22_X1 U23934 ( .A1(n21032), .A2(n20981), .B1(n21031), .B2(n20980), .ZN(
        n20963) );
  INV_X1 U23935 ( .A(n20956), .ZN(n20958) );
  INV_X1 U23936 ( .A(n20987), .ZN(n20960) );
  AOI22_X1 U23937 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20982), .B1(
        n21020), .B2(n20961), .ZN(n20962) );
  OAI211_X1 U23938 ( .C1(n20964), .C2(n20985), .A(n20963), .B(n20962), .ZN(
        P1_U3137) );
  AOI22_X1 U23939 ( .A1(n21043), .A2(n20981), .B1(n21042), .B2(n20980), .ZN(
        n20966) );
  AOI22_X1 U23940 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20982), .B1(
        n21020), .B2(n21044), .ZN(n20965) );
  OAI211_X1 U23941 ( .C1(n21047), .C2(n20985), .A(n20966), .B(n20965), .ZN(
        P1_U3138) );
  AOI22_X1 U23942 ( .A1(n21049), .A2(n20981), .B1(n21048), .B2(n20980), .ZN(
        n20968) );
  AOI22_X1 U23943 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20982), .B1(
        n21020), .B2(n21050), .ZN(n20967) );
  OAI211_X1 U23944 ( .C1(n21053), .C2(n20985), .A(n20968), .B(n20967), .ZN(
        P1_U3139) );
  AOI22_X1 U23945 ( .A1(n21055), .A2(n20981), .B1(n21054), .B2(n20980), .ZN(
        n20971) );
  AOI22_X1 U23946 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20982), .B1(
        n21020), .B2(n20969), .ZN(n20970) );
  OAI211_X1 U23947 ( .C1(n20972), .C2(n20985), .A(n20971), .B(n20970), .ZN(
        P1_U3140) );
  AOI22_X1 U23948 ( .A1(n21061), .A2(n20981), .B1(n21060), .B2(n20980), .ZN(
        n20974) );
  AOI22_X1 U23949 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20982), .B1(
        n21020), .B2(n21062), .ZN(n20973) );
  OAI211_X1 U23950 ( .C1(n21065), .C2(n20985), .A(n20974), .B(n20973), .ZN(
        P1_U3141) );
  AOI22_X1 U23951 ( .A1(n21067), .A2(n20981), .B1(n21066), .B2(n20980), .ZN(
        n20976) );
  AOI22_X1 U23952 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20982), .B1(
        n21020), .B2(n9920), .ZN(n20975) );
  OAI211_X1 U23953 ( .C1(n9923), .C2(n20985), .A(n20976), .B(n20975), .ZN(
        P1_U3142) );
  AOI22_X1 U23954 ( .A1(n21074), .A2(n20981), .B1(n21073), .B2(n20980), .ZN(
        n20979) );
  AOI22_X1 U23955 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20982), .B1(
        n21020), .B2(n21075), .ZN(n20978) );
  OAI211_X1 U23956 ( .C1(n9925), .C2(n20985), .A(n20979), .B(n20978), .ZN(
        P1_U3143) );
  AOI22_X1 U23957 ( .A1(n21082), .A2(n20981), .B1(n21080), .B2(n20980), .ZN(
        n20984) );
  AOI22_X1 U23958 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20982), .B1(
        n21020), .B2(n21083), .ZN(n20983) );
  OAI211_X1 U23959 ( .C1(n21089), .C2(n20985), .A(n20984), .B(n20983), .ZN(
        P1_U3144) );
  NOR2_X1 U23960 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21028), .ZN(
        n21018) );
  NAND2_X1 U23961 ( .A1(n21025), .A2(n20988), .ZN(n20991) );
  OAI22_X1 U23962 ( .A1(n20991), .A2(n21030), .B1(n20990), .B2(n20989), .ZN(
        n21017) );
  AOI22_X1 U23963 ( .A1(n21032), .A2(n21018), .B1(n21031), .B2(n21017), .ZN(
        n20997) );
  OAI21_X1 U23964 ( .B1(n21020), .B2(n21068), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20992) );
  AOI21_X1 U23965 ( .B1(n20992), .B2(n20991), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20995) );
  AOI22_X1 U23966 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21021), .B1(
        n21020), .B2(n21038), .ZN(n20996) );
  OAI211_X1 U23967 ( .C1(n21041), .C2(n21088), .A(n20997), .B(n20996), .ZN(
        P1_U3145) );
  AOI22_X1 U23968 ( .A1(n21043), .A2(n21018), .B1(n21042), .B2(n21017), .ZN(
        n21000) );
  AOI22_X1 U23969 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21021), .B1(
        n21020), .B2(n20998), .ZN(n20999) );
  OAI211_X1 U23970 ( .C1(n21001), .C2(n21088), .A(n21000), .B(n20999), .ZN(
        P1_U3146) );
  AOI22_X1 U23971 ( .A1(n21049), .A2(n21018), .B1(n21048), .B2(n21017), .ZN(
        n21004) );
  AOI22_X1 U23972 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21021), .B1(
        n21020), .B2(n21002), .ZN(n21003) );
  OAI211_X1 U23973 ( .C1(n21005), .C2(n21088), .A(n21004), .B(n21003), .ZN(
        P1_U3147) );
  AOI22_X1 U23974 ( .A1(n21055), .A2(n21018), .B1(n21054), .B2(n21017), .ZN(
        n21007) );
  AOI22_X1 U23975 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21021), .B1(
        n21020), .B2(n21056), .ZN(n21006) );
  OAI211_X1 U23976 ( .C1(n21059), .C2(n21088), .A(n21007), .B(n21006), .ZN(
        P1_U3148) );
  AOI22_X1 U23977 ( .A1(n21061), .A2(n21018), .B1(n21060), .B2(n21017), .ZN(
        n21010) );
  AOI22_X1 U23978 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21021), .B1(
        n21020), .B2(n21008), .ZN(n21009) );
  OAI211_X1 U23979 ( .C1(n21011), .C2(n21088), .A(n21010), .B(n21009), .ZN(
        P1_U3149) );
  AOI22_X1 U23980 ( .A1(n21067), .A2(n21018), .B1(n21066), .B2(n21017), .ZN(
        n21013) );
  AOI22_X1 U23981 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21021), .B1(
        n21020), .B2(n9922), .ZN(n21012) );
  OAI211_X1 U23982 ( .C1(n9921), .C2(n21088), .A(n21013), .B(n21012), .ZN(
        P1_U3150) );
  AOI22_X1 U23983 ( .A1(n21074), .A2(n21018), .B1(n21073), .B2(n21017), .ZN(
        n21015) );
  AOI22_X1 U23984 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21021), .B1(
        n21020), .B2(n9924), .ZN(n21014) );
  OAI211_X1 U23985 ( .C1(n21016), .C2(n21088), .A(n21015), .B(n21014), .ZN(
        P1_U3151) );
  AOI22_X1 U23986 ( .A1(n21082), .A2(n21018), .B1(n21080), .B2(n21017), .ZN(
        n21023) );
  AOI22_X1 U23987 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21021), .B1(
        n21020), .B2(n21019), .ZN(n21022) );
  OAI211_X1 U23988 ( .C1(n21024), .C2(n21088), .A(n21023), .B(n21022), .ZN(
        P1_U3152) );
  INV_X1 U23989 ( .A(n21029), .ZN(n21081) );
  INV_X1 U23990 ( .A(n21025), .ZN(n21027) );
  OAI222_X1 U23991 ( .A1(n21030), .A2(n21029), .B1(n13022), .B2(n21028), .C1(
        n21027), .C2(n21026), .ZN(n21079) );
  AOI22_X1 U23992 ( .A1(n21032), .A2(n21081), .B1(n21031), .B2(n21079), .ZN(
        n21040) );
  NOR2_X1 U23993 ( .A1(n21034), .A2(n21033), .ZN(n21037) );
  OAI21_X1 U23994 ( .B1(n21037), .B2(n21036), .A(n21035), .ZN(n21085) );
  AOI22_X1 U23995 ( .A1(n21085), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n21068), .B2(n21038), .ZN(n21039) );
  OAI211_X1 U23996 ( .C1(n21041), .C2(n21071), .A(n21040), .B(n21039), .ZN(
        P1_U3153) );
  AOI22_X1 U23997 ( .A1(n21043), .A2(n21081), .B1(n21042), .B2(n21079), .ZN(
        n21046) );
  AOI22_X1 U23998 ( .A1(n21085), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n21084), .B2(n21044), .ZN(n21045) );
  OAI211_X1 U23999 ( .C1(n21047), .C2(n21088), .A(n21046), .B(n21045), .ZN(
        P1_U3154) );
  AOI22_X1 U24000 ( .A1(n21049), .A2(n21081), .B1(n21048), .B2(n21079), .ZN(
        n21052) );
  AOI22_X1 U24001 ( .A1(n21085), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n21084), .B2(n21050), .ZN(n21051) );
  OAI211_X1 U24002 ( .C1(n21053), .C2(n21088), .A(n21052), .B(n21051), .ZN(
        P1_U3155) );
  AOI22_X1 U24003 ( .A1(n21055), .A2(n21081), .B1(n21054), .B2(n21079), .ZN(
        n21058) );
  AOI22_X1 U24004 ( .A1(n21085), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n21068), .B2(n21056), .ZN(n21057) );
  OAI211_X1 U24005 ( .C1(n21059), .C2(n21071), .A(n21058), .B(n21057), .ZN(
        P1_U3156) );
  AOI22_X1 U24006 ( .A1(n21061), .A2(n21081), .B1(n21060), .B2(n21079), .ZN(
        n21064) );
  AOI22_X1 U24007 ( .A1(n21085), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n21084), .B2(n21062), .ZN(n21063) );
  OAI211_X1 U24008 ( .C1(n21065), .C2(n21088), .A(n21064), .B(n21063), .ZN(
        P1_U3157) );
  AOI22_X1 U24009 ( .A1(n21067), .A2(n21081), .B1(n21066), .B2(n21079), .ZN(
        n21070) );
  AOI22_X1 U24010 ( .A1(n21085), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n21068), .B2(n9922), .ZN(n21069) );
  OAI211_X1 U24011 ( .C1(n9921), .C2(n21071), .A(n21070), .B(n21069), .ZN(
        P1_U3158) );
  AOI22_X1 U24012 ( .A1(n21074), .A2(n21081), .B1(n21073), .B2(n21079), .ZN(
        n21077) );
  AOI22_X1 U24013 ( .A1(n21085), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n21084), .B2(n21075), .ZN(n21076) );
  OAI211_X1 U24014 ( .C1(n9925), .C2(n21088), .A(n21077), .B(n21076), .ZN(
        P1_U3159) );
  AOI22_X1 U24015 ( .A1(n21082), .A2(n21081), .B1(n21080), .B2(n21079), .ZN(
        n21087) );
  AOI22_X1 U24016 ( .A1(n21085), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n21084), .B2(n21083), .ZN(n21086) );
  OAI211_X1 U24017 ( .C1(n21089), .C2(n21088), .A(n21087), .B(n21086), .ZN(
        P1_U3160) );
  NOR2_X1 U24018 ( .A1(n21091), .A2(n21090), .ZN(n21093) );
  OAI21_X1 U24019 ( .B1(n21093), .B2(n13022), .A(n21092), .ZN(P1_U3163) );
  INV_X1 U24020 ( .A(n21175), .ZN(n21171) );
  AND2_X1 U24021 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21171), .ZN(
        P1_U3164) );
  AND2_X1 U24022 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21171), .ZN(
        P1_U3165) );
  AND2_X1 U24023 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21171), .ZN(
        P1_U3166) );
  AND2_X1 U24024 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21171), .ZN(
        P1_U3167) );
  AND2_X1 U24025 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21171), .ZN(
        P1_U3168) );
  AND2_X1 U24026 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21171), .ZN(
        P1_U3169) );
  AND2_X1 U24027 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21171), .ZN(
        P1_U3170) );
  NOR2_X1 U24028 ( .A1(n21175), .A2(n21237), .ZN(P1_U3171) );
  AND2_X1 U24029 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21171), .ZN(
        P1_U3172) );
  AND2_X1 U24030 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21171), .ZN(
        P1_U3173) );
  AND2_X1 U24031 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21171), .ZN(
        P1_U3174) );
  AND2_X1 U24032 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21171), .ZN(
        P1_U3175) );
  AND2_X1 U24033 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21171), .ZN(
        P1_U3176) );
  AND2_X1 U24034 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21171), .ZN(
        P1_U3177) );
  AND2_X1 U24035 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21171), .ZN(
        P1_U3178) );
  AND2_X1 U24036 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21171), .ZN(
        P1_U3179) );
  AND2_X1 U24037 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21171), .ZN(
        P1_U3180) );
  AND2_X1 U24038 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21171), .ZN(
        P1_U3181) );
  INV_X1 U24039 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n21243) );
  NOR2_X1 U24040 ( .A1(n21175), .A2(n21243), .ZN(P1_U3182) );
  AND2_X1 U24041 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21171), .ZN(
        P1_U3183) );
  NOR2_X1 U24042 ( .A1(n21175), .A2(n21266), .ZN(P1_U3184) );
  AND2_X1 U24043 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21171), .ZN(
        P1_U3185) );
  AND2_X1 U24044 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21171), .ZN(P1_U3186) );
  INV_X1 U24045 ( .A(P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21464) );
  NOR2_X1 U24046 ( .A1(n21175), .A2(n21464), .ZN(P1_U3187) );
  AND2_X1 U24047 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21171), .ZN(P1_U3188) );
  AND2_X1 U24048 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21171), .ZN(P1_U3189) );
  AND2_X1 U24049 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21171), .ZN(P1_U3190) );
  AND2_X1 U24050 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21171), .ZN(P1_U3191) );
  INV_X1 U24051 ( .A(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21467) );
  NOR2_X1 U24052 ( .A1(n21175), .A2(n21467), .ZN(P1_U3192) );
  AND2_X1 U24053 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21171), .ZN(P1_U3193) );
  AOI21_X1 U24054 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21094), .A(n21101), 
        .ZN(n21109) );
  NOR2_X1 U24055 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21096) );
  NOR2_X1 U24056 ( .A1(n21096), .A2(n21095), .ZN(n21097) );
  AOI211_X1 U24057 ( .C1(NA), .C2(n21101), .A(n21097), .B(n21105), .ZN(n21098)
         );
  OAI22_X1 U24058 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21109), .B1(n21187), 
        .B2(n21098), .ZN(P1_U3194) );
  OAI21_X1 U24059 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21100), .A(n21099), 
        .ZN(n21107) );
  AOI221_X1 U24060 ( .B1(NA), .B2(n21103), .C1(n21102), .C2(n21103), .A(n21101), .ZN(n21104) );
  OAI211_X1 U24061 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21105), .A(HOLD), .B(
        n21104), .ZN(n21106) );
  OAI221_X1 U24062 ( .B1(n21109), .B2(n21108), .C1(n21109), .C2(n21107), .A(
        n21106), .ZN(P1_U3196) );
  NAND2_X1 U24063 ( .A1(n21187), .A2(n21110), .ZN(n21159) );
  INV_X1 U24064 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21111) );
  AND2_X1 U24065 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21187), .ZN(n21156) );
  INV_X1 U24066 ( .A(n21156), .ZN(n21163) );
  OAI222_X1 U24067 ( .A1(n21159), .A2(n21113), .B1(n21111), .B2(n21184), .C1(
        n13419), .C2(n21163), .ZN(P1_U3197) );
  INV_X1 U24068 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21112) );
  OAI222_X1 U24069 ( .A1(n21163), .A2(n21113), .B1(n21112), .B2(n21184), .C1(
        n21115), .C2(n21159), .ZN(P1_U3198) );
  OAI222_X1 U24070 ( .A1(n21163), .A2(n21115), .B1(n21114), .B2(n21184), .C1(
        n21117), .C2(n21159), .ZN(P1_U3199) );
  INV_X1 U24071 ( .A(n21159), .ZN(n21153) );
  AOI22_X1 U24072 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n21185), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(n21153), .ZN(n21116) );
  OAI21_X1 U24073 ( .B1(n21117), .B2(n21163), .A(n21116), .ZN(P1_U3200) );
  INV_X1 U24074 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21119) );
  AOI22_X1 U24075 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n21185), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n21153), .ZN(n21118) );
  OAI21_X1 U24076 ( .B1(n21119), .B2(n21163), .A(n21118), .ZN(P1_U3201) );
  AOI22_X1 U24077 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n21185), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n21156), .ZN(n21120) );
  OAI21_X1 U24078 ( .B1(n21122), .B2(n21159), .A(n21120), .ZN(P1_U3202) );
  AOI22_X1 U24079 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n21185), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n21153), .ZN(n21121) );
  OAI21_X1 U24080 ( .B1(n21122), .B2(n21163), .A(n21121), .ZN(P1_U3203) );
  AOI22_X1 U24081 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n21185), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n21156), .ZN(n21123) );
  OAI21_X1 U24082 ( .B1(n15214), .B2(n21159), .A(n21123), .ZN(P1_U3204) );
  AOI222_X1 U24083 ( .A1(n21156), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21185), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n21153), .ZN(n21124) );
  INV_X1 U24084 ( .A(n21124), .ZN(P1_U3205) );
  AOI222_X1 U24085 ( .A1(n21156), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n21185), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n21153), .ZN(n21125) );
  INV_X1 U24086 ( .A(n21125), .ZN(P1_U3206) );
  INV_X1 U24087 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n21126) );
  OAI222_X1 U24088 ( .A1(n21163), .A2(n21127), .B1(n21126), .B2(n21184), .C1(
        n21129), .C2(n21159), .ZN(P1_U3207) );
  INV_X1 U24089 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21128) );
  OAI222_X1 U24090 ( .A1(n21163), .A2(n21129), .B1(n21128), .B2(n21184), .C1(
        n21131), .C2(n21159), .ZN(P1_U3208) );
  INV_X1 U24091 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21130) );
  OAI222_X1 U24092 ( .A1(n21163), .A2(n21131), .B1(n21130), .B2(n21184), .C1(
        n21132), .C2(n21159), .ZN(P1_U3209) );
  INV_X1 U24093 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21133) );
  OAI222_X1 U24094 ( .A1(n21159), .A2(n21135), .B1(n21133), .B2(n21184), .C1(
        n21132), .C2(n21163), .ZN(P1_U3210) );
  INV_X1 U24095 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21134) );
  OAI222_X1 U24096 ( .A1(n21163), .A2(n21135), .B1(n21134), .B2(n21184), .C1(
        n21137), .C2(n21159), .ZN(P1_U3211) );
  INV_X1 U24097 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21136) );
  OAI222_X1 U24098 ( .A1(n21163), .A2(n21137), .B1(n21136), .B2(n21184), .C1(
        n15129), .C2(n21159), .ZN(P1_U3212) );
  INV_X1 U24099 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21138) );
  OAI222_X1 U24100 ( .A1(n21159), .A2(n21140), .B1(n21138), .B2(n21184), .C1(
        n15129), .C2(n21163), .ZN(P1_U3213) );
  AOI22_X1 U24101 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21185), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21153), .ZN(n21139) );
  OAI21_X1 U24102 ( .B1(n21140), .B2(n21163), .A(n21139), .ZN(P1_U3214) );
  AOI22_X1 U24103 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21185), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21156), .ZN(n21141) );
  OAI21_X1 U24104 ( .B1(n21143), .B2(n21159), .A(n21141), .ZN(P1_U3215) );
  INV_X1 U24105 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21142) );
  OAI222_X1 U24106 ( .A1(n21163), .A2(n21143), .B1(n21142), .B2(n21184), .C1(
        n15091), .C2(n21159), .ZN(P1_U3216) );
  INV_X1 U24107 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21144) );
  OAI222_X1 U24108 ( .A1(n21159), .A2(n21146), .B1(n21144), .B2(n21184), .C1(
        n15091), .C2(n21163), .ZN(P1_U3217) );
  INV_X1 U24109 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21145) );
  OAI222_X1 U24110 ( .A1(n21163), .A2(n21146), .B1(n21145), .B2(n21184), .C1(
        n15072), .C2(n21159), .ZN(P1_U3218) );
  INV_X1 U24111 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21147) );
  OAI222_X1 U24112 ( .A1(n21163), .A2(n15072), .B1(n21147), .B2(n21184), .C1(
        n21148), .C2(n21159), .ZN(P1_U3219) );
  INV_X1 U24113 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21350) );
  OAI222_X1 U24114 ( .A1(n21163), .A2(n21148), .B1(n21350), .B2(n21184), .C1(
        n21150), .C2(n21159), .ZN(P1_U3220) );
  INV_X1 U24115 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21149) );
  OAI222_X1 U24116 ( .A1(n21163), .A2(n21150), .B1(n21149), .B2(n21184), .C1(
        n21152), .C2(n21159), .ZN(P1_U3221) );
  INV_X1 U24117 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21151) );
  OAI222_X1 U24118 ( .A1(n21163), .A2(n21152), .B1(n21151), .B2(n21184), .C1(
        n21155), .C2(n21159), .ZN(P1_U3222) );
  AOI22_X1 U24119 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21153), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21185), .ZN(n21154) );
  OAI21_X1 U24120 ( .B1(n21155), .B2(n21163), .A(n21154), .ZN(P1_U3223) );
  AOI22_X1 U24121 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n21156), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21185), .ZN(n21157) );
  OAI21_X1 U24122 ( .B1(n21158), .B2(n21159), .A(n21157), .ZN(P1_U3224) );
  INV_X1 U24123 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21498) );
  OAI222_X1 U24124 ( .A1(n21159), .A2(n21162), .B1(n21498), .B2(n21184), .C1(
        n21158), .C2(n21163), .ZN(P1_U3225) );
  INV_X1 U24125 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21161) );
  OAI222_X1 U24126 ( .A1(n21163), .A2(n21162), .B1(n21161), .B2(n21184), .C1(
        n21160), .C2(n21159), .ZN(P1_U3226) );
  INV_X1 U24127 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21164) );
  AOI22_X1 U24128 ( .A1(n21187), .A2(n21165), .B1(n21164), .B2(n21185), .ZN(
        P1_U3458) );
  INV_X1 U24129 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21177) );
  INV_X1 U24130 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21166) );
  AOI22_X1 U24131 ( .A1(n21184), .A2(n21177), .B1(n21166), .B2(n21185), .ZN(
        P1_U3459) );
  INV_X1 U24132 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21167) );
  AOI22_X1 U24133 ( .A1(n21184), .A2(n21168), .B1(n21167), .B2(n21185), .ZN(
        P1_U3460) );
  INV_X1 U24134 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21182) );
  INV_X1 U24135 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21169) );
  AOI22_X1 U24136 ( .A1(n21184), .A2(n21182), .B1(n21169), .B2(n21185), .ZN(
        P1_U3461) );
  INV_X1 U24137 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21172) );
  INV_X1 U24138 ( .A(n21173), .ZN(n21170) );
  AOI21_X1 U24139 ( .B1(n21172), .B2(n21171), .A(n21170), .ZN(P1_U3464) );
  OAI21_X1 U24140 ( .B1(n21175), .B2(n21174), .A(n21173), .ZN(P1_U3465) );
  AOI21_X1 U24141 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21176) );
  AOI22_X1 U24142 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21176), .B2(n13419), .ZN(n21178) );
  AOI22_X1 U24143 ( .A1(n21179), .A2(n21178), .B1(n21177), .B2(n21181), .ZN(
        P1_U3481) );
  NOR2_X1 U24144 ( .A1(n21181), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21180) );
  AOI22_X1 U24145 ( .A1(n21182), .A2(n21181), .B1(n13242), .B2(n21180), .ZN(
        P1_U3482) );
  INV_X1 U24146 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21183) );
  AOI22_X1 U24147 ( .A1(n21184), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21183), 
        .B2(n21185), .ZN(P1_U3483) );
  INV_X1 U24148 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21186) );
  AOI22_X1 U24149 ( .A1(n21187), .A2(n21186), .B1(n21369), .B2(n21185), .ZN(
        P1_U3486) );
  AOI22_X1 U24150 ( .A1(n21189), .A2(P3_ADDRESS_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n21188), .ZN(n21500) );
  NOR4_X1 U24151 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(
        P1_EAX_REG_14__SCAN_IN), .A3(P3_REIP_REG_22__SCAN_IN), .A4(
        P1_UWORD_REG_0__SCAN_IN), .ZN(n21190) );
  NAND3_X1 U24152 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_ADDRESS_REG_9__SCAN_IN), .A3(n21190), .ZN(n21200) );
  NAND4_X1 U24153 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(P1_LWORD_REG_0__SCAN_IN), 
        .A3(n21386), .A4(n21384), .ZN(n21191) );
  NOR3_X1 U24154 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(n21191), .ZN(n21198) );
  NAND4_X1 U24155 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n21406), .A3(
        n21396), .A4(n21399), .ZN(n21196) );
  NAND4_X1 U24156 ( .A1(BUF1_REG_23__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_DATAO_REG_4__SCAN_IN), .A4(n21412), .ZN(n21195) );
  NAND4_X1 U24157 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n21420), .ZN(n21192) );
  NOR2_X1 U24158 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21192), .ZN(
        n21193) );
  NAND4_X1 U24159 ( .A1(n21193), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A3(
        P3_REIP_REG_0__SCAN_IN), .A4(n21415), .ZN(n21194) );
  NOR3_X1 U24160 ( .A1(n21196), .A2(n21195), .A3(n21194), .ZN(n21197) );
  NAND4_X1 U24161 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21198), .A3(n21197), 
        .A4(n21468), .ZN(n21199) );
  NOR4_X1 U24162 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(n21370), .A3(n21200), .A4(
        n21199), .ZN(n21233) );
  INV_X1 U24163 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21274) );
  NAND4_X1 U24164 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(n21274), .A4(n21268), .ZN(
        n21204) );
  NAND4_X1 U24165 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .A3(P3_UWORD_REG_1__SCAN_IN), .A4(n21259), 
        .ZN(n21203) );
  NAND4_X1 U24166 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P1_UWORD_REG_5__SCAN_IN), 
        .A3(P1_DATAO_REG_4__SCAN_IN), .A4(n21290), .ZN(n21202) );
  NAND4_X1 U24167 ( .A1(n21281), .A2(n15072), .A3(n21280), .A4(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21201) );
  NOR4_X1 U24168 ( .A1(n21204), .A2(n21203), .A3(n21202), .A4(n21201), .ZN(
        n21232) );
  NAND4_X1 U24169 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_EAX_REG_25__SCAN_IN), .A3(n21235), .A4(n19079), .ZN(n21208) );
  INV_X1 U24170 ( .A(P1_UWORD_REG_3__SCAN_IN), .ZN(n21403) );
  NAND4_X1 U24171 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n13138), .A3(n21403), 
        .A4(n21402), .ZN(n21207) );
  NAND4_X1 U24172 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_2__0__SCAN_IN), .A3(P3_DATAO_REG_25__SCAN_IN), .A4(
        n21256), .ZN(n21206) );
  INV_X1 U24173 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n21250) );
  NAND4_X1 U24174 ( .A1(P3_DATAO_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(n21250), .A4(n21249), .ZN(n21205)
         );
  NOR4_X1 U24175 ( .A1(n21208), .A2(n21207), .A3(n21206), .A4(n21205), .ZN(
        n21231) );
  NOR4_X1 U24176 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(
        P1_EBX_REG_31__SCAN_IN), .A3(P2_DATAWIDTH_REG_28__SCAN_IN), .A4(n21437), .ZN(n21212) );
  INV_X1 U24177 ( .A(P2_UWORD_REG_11__SCAN_IN), .ZN(n21474) );
  NOR4_X1 U24178 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21473), .A3(
        n21477), .A4(n21474), .ZN(n21211) );
  INV_X1 U24179 ( .A(READY22_REG_SCAN_IN), .ZN(n21483) );
  NOR4_X1 U24180 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(
        P1_EBX_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(n21483), .ZN(n21210) );
  AND4_X1 U24181 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_5__0__SCAN_IN), .A3(P1_INSTQUEUE_REG_15__0__SCAN_IN), 
        .A4(n21457), .ZN(n21209) );
  NAND4_X1 U24182 ( .A1(n21212), .A2(n21211), .A3(n21210), .A4(n21209), .ZN(
        n21229) );
  NOR4_X1 U24183 ( .A1(P3_LWORD_REG_15__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .A3(n21214), .A4(n21213), .ZN(n21217) );
  INV_X1 U24184 ( .A(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21434) );
  NOR4_X1 U24185 ( .A1(BUF2_REG_9__SCAN_IN), .A2(DATAI_11_), .A3(
        P3_INSTQUEUE_REG_11__3__SCAN_IN), .A4(n21434), .ZN(n21216) );
  INV_X1 U24186 ( .A(P3_UWORD_REG_14__SCAN_IN), .ZN(n21444) );
  NOR4_X1 U24187 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_EBX_REG_11__SCAN_IN), .A3(n12854), .A4(n21444), .ZN(n21215) );
  NAND4_X1 U24188 ( .A1(P3_UWORD_REG_8__SCAN_IN), .A2(n21217), .A3(n21216), 
        .A4(n21215), .ZN(n21228) );
  INV_X1 U24189 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n21334) );
  NOR4_X1 U24190 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A4(
        n21334), .ZN(n21221) );
  INV_X1 U24191 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n21332) );
  NOR4_X1 U24192 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n21332), .ZN(n21220) );
  INV_X1 U24193 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21348) );
  NOR4_X1 U24194 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21351), .A3(
        n21348), .A4(n21350), .ZN(n21219) );
  NOR4_X1 U24195 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_EAX_REG_24__SCAN_IN), .A3(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A4(
        P3_UWORD_REG_6__SCAN_IN), .ZN(n21218) );
  NAND4_X1 U24196 ( .A1(n21221), .A2(n21220), .A3(n21219), .A4(n21218), .ZN(
        n21227) );
  INV_X1 U24197 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n21306) );
  NOR4_X1 U24198 ( .A1(READY21_REG_SCAN_IN), .A2(P3_EAX_REG_28__SCAN_IN), .A3(
        n21306), .A4(n21307), .ZN(n21225) );
  NOR4_X1 U24199 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(
        BUF1_REG_22__SCAN_IN), .A3(P3_EBX_REG_12__SCAN_IN), .A4(n21304), .ZN(
        n21224) );
  NOR4_X1 U24200 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10595), .A3(
        n21319), .A4(n21322), .ZN(n21223) );
  NOR4_X1 U24201 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_14__3__SCAN_IN), .A3(BUF1_REG_25__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21222) );
  NAND4_X1 U24202 ( .A1(n21225), .A2(n21224), .A3(n21223), .A4(n21222), .ZN(
        n21226) );
  NOR4_X1 U24203 ( .A1(n21229), .A2(n21228), .A3(n21227), .A4(n21226), .ZN(
        n21230) );
  NAND4_X1 U24204 ( .A1(n21233), .A2(n21232), .A3(n21231), .A4(n21230), .ZN(
        n21497) );
  AOI22_X1 U24205 ( .A1(n13138), .A2(keyinput72), .B1(n21235), .B2(keyinput103), .ZN(n21234) );
  OAI221_X1 U24206 ( .B1(n13138), .B2(keyinput72), .C1(n21235), .C2(
        keyinput103), .A(n21234), .ZN(n21247) );
  AOI22_X1 U24207 ( .A1(n19079), .A2(keyinput22), .B1(keyinput47), .B2(n21237), 
        .ZN(n21236) );
  OAI221_X1 U24208 ( .B1(n19079), .B2(keyinput22), .C1(n21237), .C2(keyinput47), .A(n21236), .ZN(n21246) );
  AOI22_X1 U24209 ( .A1(n21240), .A2(keyinput100), .B1(n21239), .B2(keyinput29), .ZN(n21238) );
  OAI221_X1 U24210 ( .B1(n21240), .B2(keyinput100), .C1(n21239), .C2(
        keyinput29), .A(n21238), .ZN(n21245) );
  INV_X1 U24211 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n21242) );
  AOI22_X1 U24212 ( .A1(n21243), .A2(keyinput126), .B1(n21242), .B2(keyinput67), .ZN(n21241) );
  OAI221_X1 U24213 ( .B1(n21243), .B2(keyinput126), .C1(n21242), .C2(
        keyinput67), .A(n21241), .ZN(n21244) );
  NOR4_X1 U24214 ( .A1(n21247), .A2(n21246), .A3(n21245), .A4(n21244), .ZN(
        n21298) );
  AOI22_X1 U24215 ( .A1(n21250), .A2(keyinput104), .B1(keyinput117), .B2(
        n21249), .ZN(n21248) );
  OAI221_X1 U24216 ( .B1(n21250), .B2(keyinput104), .C1(n21249), .C2(
        keyinput117), .A(n21248), .ZN(n21263) );
  INV_X1 U24217 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n21253) );
  INV_X1 U24218 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n21252) );
  AOI22_X1 U24219 ( .A1(n21253), .A2(keyinput88), .B1(n21252), .B2(keyinput97), 
        .ZN(n21251) );
  OAI221_X1 U24220 ( .B1(n21253), .B2(keyinput88), .C1(n21252), .C2(keyinput97), .A(n21251), .ZN(n21262) );
  INV_X1 U24221 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n21255) );
  AOI22_X1 U24222 ( .A1(n21256), .A2(keyinput1), .B1(keyinput77), .B2(n21255), 
        .ZN(n21254) );
  OAI221_X1 U24223 ( .B1(n21256), .B2(keyinput1), .C1(n21255), .C2(keyinput77), 
        .A(n21254), .ZN(n21261) );
  INV_X1 U24224 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n21258) );
  AOI22_X1 U24225 ( .A1(n21259), .A2(keyinput114), .B1(keyinput4), .B2(n21258), 
        .ZN(n21257) );
  OAI221_X1 U24226 ( .B1(n21259), .B2(keyinput114), .C1(n21258), .C2(keyinput4), .A(n21257), .ZN(n21260) );
  NOR4_X1 U24227 ( .A1(n21263), .A2(n21262), .A3(n21261), .A4(n21260), .ZN(
        n21297) );
  INV_X1 U24228 ( .A(P3_UWORD_REG_1__SCAN_IN), .ZN(n21265) );
  AOI22_X1 U24229 ( .A1(n21266), .A2(keyinput113), .B1(n21265), .B2(keyinput87), .ZN(n21264) );
  OAI221_X1 U24230 ( .B1(n21266), .B2(keyinput113), .C1(n21265), .C2(
        keyinput87), .A(n21264), .ZN(n21278) );
  INV_X1 U24231 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n21269) );
  AOI22_X1 U24232 ( .A1(n21269), .A2(keyinput71), .B1(keyinput2), .B2(n21268), 
        .ZN(n21267) );
  OAI221_X1 U24233 ( .B1(n21269), .B2(keyinput71), .C1(n21268), .C2(keyinput2), 
        .A(n21267), .ZN(n21277) );
  AOI22_X1 U24234 ( .A1(n21272), .A2(keyinput19), .B1(keyinput120), .B2(n21271), .ZN(n21270) );
  OAI221_X1 U24235 ( .B1(n21272), .B2(keyinput19), .C1(n21271), .C2(
        keyinput120), .A(n21270), .ZN(n21276) );
  AOI22_X1 U24236 ( .A1(n21274), .A2(keyinput12), .B1(keyinput31), .B2(n15072), 
        .ZN(n21273) );
  OAI221_X1 U24237 ( .B1(n21274), .B2(keyinput12), .C1(n15072), .C2(keyinput31), .A(n21273), .ZN(n21275) );
  NOR4_X1 U24238 ( .A1(n21278), .A2(n21277), .A3(n21276), .A4(n21275), .ZN(
        n21296) );
  AOI22_X1 U24239 ( .A1(n21281), .A2(keyinput14), .B1(keyinput91), .B2(n21280), 
        .ZN(n21279) );
  OAI221_X1 U24240 ( .B1(n21281), .B2(keyinput14), .C1(n21280), .C2(keyinput91), .A(n21279), .ZN(n21294) );
  AOI22_X1 U24241 ( .A1(n21284), .A2(keyinput80), .B1(keyinput24), .B2(n21283), 
        .ZN(n21282) );
  OAI221_X1 U24242 ( .B1(n21284), .B2(keyinput80), .C1(n21283), .C2(keyinput24), .A(n21282), .ZN(n21293) );
  INV_X1 U24243 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n21286) );
  AOI22_X1 U24244 ( .A1(n21287), .A2(keyinput32), .B1(n21286), .B2(keyinput38), 
        .ZN(n21285) );
  OAI221_X1 U24245 ( .B1(n21287), .B2(keyinput32), .C1(n21286), .C2(keyinput38), .A(n21285), .ZN(n21292) );
  INV_X1 U24246 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n21289) );
  AOI22_X1 U24247 ( .A1(n21290), .A2(keyinput34), .B1(keyinput61), .B2(n21289), 
        .ZN(n21288) );
  OAI221_X1 U24248 ( .B1(n21290), .B2(keyinput34), .C1(n21289), .C2(keyinput61), .A(n21288), .ZN(n21291) );
  NOR4_X1 U24249 ( .A1(n21294), .A2(n21293), .A3(n21292), .A4(n21291), .ZN(
        n21295) );
  NAND4_X1 U24250 ( .A1(n21298), .A2(n21297), .A3(n21296), .A4(n21295), .ZN(
        n21495) );
  INV_X1 U24251 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n21301) );
  AOI22_X1 U24252 ( .A1(n21301), .A2(keyinput21), .B1(keyinput79), .B2(n21300), 
        .ZN(n21299) );
  OAI221_X1 U24253 ( .B1(n21301), .B2(keyinput21), .C1(n21300), .C2(keyinput79), .A(n21299), .ZN(n21314) );
  INV_X1 U24254 ( .A(READY21_REG_SCAN_IN), .ZN(n21303) );
  AOI22_X1 U24255 ( .A1(n21304), .A2(keyinput3), .B1(n21303), .B2(keyinput36), 
        .ZN(n21302) );
  OAI221_X1 U24256 ( .B1(n21304), .B2(keyinput3), .C1(n21303), .C2(keyinput36), 
        .A(n21302), .ZN(n21313) );
  AOI22_X1 U24257 ( .A1(n21307), .A2(keyinput63), .B1(n21306), .B2(keyinput23), 
        .ZN(n21305) );
  OAI221_X1 U24258 ( .B1(n21307), .B2(keyinput63), .C1(n21306), .C2(keyinput23), .A(n21305), .ZN(n21312) );
  INV_X1 U24259 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n21309) );
  AOI22_X1 U24260 ( .A1(n21310), .A2(keyinput124), .B1(n21309), .B2(keyinput66), .ZN(n21308) );
  OAI221_X1 U24261 ( .B1(n21310), .B2(keyinput124), .C1(n21309), .C2(
        keyinput66), .A(n21308), .ZN(n21311) );
  NOR4_X1 U24262 ( .A1(n21314), .A2(n21313), .A3(n21312), .A4(n21311), .ZN(
        n21364) );
  AOI22_X1 U24263 ( .A1(n21317), .A2(keyinput102), .B1(n21316), .B2(keyinput58), .ZN(n21315) );
  OAI221_X1 U24264 ( .B1(n21317), .B2(keyinput102), .C1(n21316), .C2(
        keyinput58), .A(n21315), .ZN(n21329) );
  AOI22_X1 U24265 ( .A1(n21320), .A2(keyinput10), .B1(n21319), .B2(keyinput17), 
        .ZN(n21318) );
  OAI221_X1 U24266 ( .B1(n21320), .B2(keyinput10), .C1(n21319), .C2(keyinput17), .A(n21318), .ZN(n21328) );
  AOI22_X1 U24267 ( .A1(n21323), .A2(keyinput99), .B1(keyinput111), .B2(n21322), .ZN(n21321) );
  OAI221_X1 U24268 ( .B1(n21323), .B2(keyinput99), .C1(n21322), .C2(
        keyinput111), .A(n21321), .ZN(n21327) );
  INV_X1 U24269 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n21325) );
  AOI22_X1 U24270 ( .A1(n10595), .A2(keyinput40), .B1(keyinput96), .B2(n21325), 
        .ZN(n21324) );
  OAI221_X1 U24271 ( .B1(n10595), .B2(keyinput40), .C1(n21325), .C2(keyinput96), .A(n21324), .ZN(n21326) );
  NOR4_X1 U24272 ( .A1(n21329), .A2(n21328), .A3(n21327), .A4(n21326), .ZN(
        n21363) );
  AOI22_X1 U24273 ( .A1(n21332), .A2(keyinput55), .B1(keyinput56), .B2(n21331), 
        .ZN(n21330) );
  OAI221_X1 U24274 ( .B1(n21332), .B2(keyinput55), .C1(n21331), .C2(keyinput56), .A(n21330), .ZN(n21345) );
  AOI22_X1 U24275 ( .A1(n21335), .A2(keyinput93), .B1(keyinput27), .B2(n21334), 
        .ZN(n21333) );
  OAI221_X1 U24276 ( .B1(n21335), .B2(keyinput93), .C1(n21334), .C2(keyinput27), .A(n21333), .ZN(n21344) );
  INV_X1 U24277 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n21338) );
  AOI22_X1 U24278 ( .A1(n21338), .A2(keyinput119), .B1(n21337), .B2(keyinput11), .ZN(n21336) );
  OAI221_X1 U24279 ( .B1(n21338), .B2(keyinput119), .C1(n21337), .C2(
        keyinput11), .A(n21336), .ZN(n21343) );
  INV_X1 U24280 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n21341) );
  AOI22_X1 U24281 ( .A1(n21341), .A2(keyinput116), .B1(keyinput8), .B2(n21340), 
        .ZN(n21339) );
  OAI221_X1 U24282 ( .B1(n21341), .B2(keyinput116), .C1(n21340), .C2(keyinput8), .A(n21339), .ZN(n21342) );
  NOR4_X1 U24283 ( .A1(n21345), .A2(n21344), .A3(n21343), .A4(n21342), .ZN(
        n21362) );
  INV_X1 U24284 ( .A(P3_UWORD_REG_8__SCAN_IN), .ZN(n21347) );
  AOI22_X1 U24285 ( .A1(n21348), .A2(keyinput51), .B1(keyinput15), .B2(n21347), 
        .ZN(n21346) );
  OAI221_X1 U24286 ( .B1(n21348), .B2(keyinput51), .C1(n21347), .C2(keyinput15), .A(n21346), .ZN(n21360) );
  AOI22_X1 U24287 ( .A1(n21351), .A2(keyinput92), .B1(keyinput73), .B2(n21350), 
        .ZN(n21349) );
  OAI221_X1 U24288 ( .B1(n21351), .B2(keyinput92), .C1(n21350), .C2(keyinput73), .A(n21349), .ZN(n21359) );
  INV_X1 U24289 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n21354) );
  INV_X1 U24290 ( .A(P3_UWORD_REG_6__SCAN_IN), .ZN(n21353) );
  AOI22_X1 U24291 ( .A1(n21354), .A2(keyinput33), .B1(keyinput122), .B2(n21353), .ZN(n21352) );
  OAI221_X1 U24292 ( .B1(n21354), .B2(keyinput33), .C1(n21353), .C2(
        keyinput122), .A(n21352), .ZN(n21358) );
  XNOR2_X1 U24293 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B(keyinput123), 
        .ZN(n21356) );
  XNOR2_X1 U24294 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput18), 
        .ZN(n21355) );
  NAND2_X1 U24295 ( .A1(n21356), .A2(n21355), .ZN(n21357) );
  NOR4_X1 U24296 ( .A1(n21360), .A2(n21359), .A3(n21358), .A4(n21357), .ZN(
        n21361) );
  NAND4_X1 U24297 ( .A1(n21364), .A2(n21363), .A3(n21362), .A4(n21361), .ZN(
        n21494) );
  INV_X1 U24298 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21366) );
  AOI22_X1 U24299 ( .A1(n21367), .A2(keyinput75), .B1(n21366), .B2(keyinput7), 
        .ZN(n21365) );
  OAI221_X1 U24300 ( .B1(n21367), .B2(keyinput75), .C1(n21366), .C2(keyinput7), 
        .A(n21365), .ZN(n21379) );
  AOI22_X1 U24301 ( .A1(n21370), .A2(keyinput109), .B1(keyinput125), .B2(
        n21369), .ZN(n21368) );
  OAI221_X1 U24302 ( .B1(n21370), .B2(keyinput109), .C1(n21369), .C2(
        keyinput125), .A(n21368), .ZN(n21378) );
  AOI22_X1 U24303 ( .A1(n21373), .A2(keyinput85), .B1(n21372), .B2(keyinput68), 
        .ZN(n21371) );
  OAI221_X1 U24304 ( .B1(n21373), .B2(keyinput85), .C1(n21372), .C2(keyinput68), .A(n21371), .ZN(n21377) );
  XNOR2_X1 U24305 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B(keyinput39), .ZN(
        n21375) );
  XNOR2_X1 U24306 ( .A(P1_EAX_REG_14__SCAN_IN), .B(keyinput84), .ZN(n21374) );
  NAND2_X1 U24307 ( .A1(n21375), .A2(n21374), .ZN(n21376) );
  NOR4_X1 U24308 ( .A1(n21379), .A2(n21378), .A3(n21377), .A4(n21376), .ZN(
        n21429) );
  AOI22_X1 U24309 ( .A1(n10490), .A2(keyinput57), .B1(keyinput16), .B2(n21381), 
        .ZN(n21380) );
  OAI221_X1 U24310 ( .B1(n10490), .B2(keyinput57), .C1(n21381), .C2(keyinput16), .A(n21380), .ZN(n21394) );
  AOI22_X1 U24311 ( .A1(n21384), .A2(keyinput37), .B1(n21383), .B2(keyinput5), 
        .ZN(n21382) );
  OAI221_X1 U24312 ( .B1(n21384), .B2(keyinput37), .C1(n21383), .C2(keyinput5), 
        .A(n21382), .ZN(n21393) );
  INV_X1 U24313 ( .A(P1_LWORD_REG_0__SCAN_IN), .ZN(n21387) );
  AOI22_X1 U24314 ( .A1(n21387), .A2(keyinput89), .B1(n21386), .B2(keyinput30), 
        .ZN(n21385) );
  OAI221_X1 U24315 ( .B1(n21387), .B2(keyinput89), .C1(n21386), .C2(keyinput30), .A(n21385), .ZN(n21392) );
  INV_X1 U24316 ( .A(P1_UWORD_REG_0__SCAN_IN), .ZN(n21388) );
  XOR2_X1 U24317 ( .A(n21388), .B(keyinput110), .Z(n21390) );
  XNOR2_X1 U24318 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B(keyinput59), .ZN(
        n21389) );
  NAND2_X1 U24319 ( .A1(n21390), .A2(n21389), .ZN(n21391) );
  NOR4_X1 U24320 ( .A1(n21394), .A2(n21393), .A3(n21392), .A4(n21391), .ZN(
        n21428) );
  AOI22_X1 U24321 ( .A1(n21397), .A2(keyinput82), .B1(n21396), .B2(keyinput46), 
        .ZN(n21395) );
  OAI221_X1 U24322 ( .B1(n21397), .B2(keyinput82), .C1(n21396), .C2(keyinput46), .A(n21395), .ZN(n21410) );
  AOI22_X1 U24323 ( .A1(n21400), .A2(keyinput50), .B1(keyinput64), .B2(n21399), 
        .ZN(n21398) );
  OAI221_X1 U24324 ( .B1(n21400), .B2(keyinput50), .C1(n21399), .C2(keyinput64), .A(n21398), .ZN(n21409) );
  AOI22_X1 U24325 ( .A1(n21403), .A2(keyinput44), .B1(keyinput70), .B2(n21402), 
        .ZN(n21401) );
  OAI221_X1 U24326 ( .B1(n21403), .B2(keyinput44), .C1(n21402), .C2(keyinput70), .A(n21401), .ZN(n21408) );
  AOI22_X1 U24327 ( .A1(n21406), .A2(keyinput76), .B1(keyinput49), .B2(n21405), 
        .ZN(n21404) );
  OAI221_X1 U24328 ( .B1(n21406), .B2(keyinput76), .C1(n21405), .C2(keyinput49), .A(n21404), .ZN(n21407) );
  NOR4_X1 U24329 ( .A1(n21410), .A2(n21409), .A3(n21408), .A4(n21407), .ZN(
        n21427) );
  INV_X1 U24330 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n21413) );
  AOI22_X1 U24331 ( .A1(n21413), .A2(keyinput26), .B1(n21412), .B2(keyinput35), 
        .ZN(n21411) );
  OAI221_X1 U24332 ( .B1(n21413), .B2(keyinput26), .C1(n21412), .C2(keyinput35), .A(n21411), .ZN(n21425) );
  AOI22_X1 U24333 ( .A1(n21415), .A2(keyinput106), .B1(keyinput65), .B2(n9995), 
        .ZN(n21414) );
  OAI221_X1 U24334 ( .B1(n21415), .B2(keyinput106), .C1(n9995), .C2(keyinput65), .A(n21414), .ZN(n21424) );
  INV_X1 U24335 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n21418) );
  AOI22_X1 U24336 ( .A1(n21418), .A2(keyinput101), .B1(keyinput81), .B2(n21417), .ZN(n21416) );
  OAI221_X1 U24337 ( .B1(n21418), .B2(keyinput101), .C1(n21417), .C2(
        keyinput81), .A(n21416), .ZN(n21423) );
  AOI22_X1 U24338 ( .A1(n21421), .A2(keyinput13), .B1(n21420), .B2(keyinput9), 
        .ZN(n21419) );
  OAI221_X1 U24339 ( .B1(n21421), .B2(keyinput13), .C1(n21420), .C2(keyinput9), 
        .A(n21419), .ZN(n21422) );
  NOR4_X1 U24340 ( .A1(n21425), .A2(n21424), .A3(n21423), .A4(n21422), .ZN(
        n21426) );
  NAND4_X1 U24341 ( .A1(n21429), .A2(n21428), .A3(n21427), .A4(n21426), .ZN(
        n21493) );
  INV_X1 U24342 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n21432) );
  AOI22_X1 U24343 ( .A1(n21432), .A2(keyinput25), .B1(keyinput83), .B2(n21431), 
        .ZN(n21430) );
  OAI221_X1 U24344 ( .B1(n21432), .B2(keyinput25), .C1(n21431), .C2(keyinput83), .A(n21430), .ZN(n21442) );
  AOI22_X1 U24345 ( .A1(n13132), .A2(keyinput41), .B1(n21434), .B2(keyinput20), 
        .ZN(n21433) );
  OAI221_X1 U24346 ( .B1(n13132), .B2(keyinput41), .C1(n21434), .C2(keyinput20), .A(n21433), .ZN(n21441) );
  AOI22_X1 U24347 ( .A1(n14561), .A2(keyinput48), .B1(n10953), .B2(keyinput107), .ZN(n21435) );
  OAI221_X1 U24348 ( .B1(n14561), .B2(keyinput48), .C1(n10953), .C2(
        keyinput107), .A(n21435), .ZN(n21440) );
  AOI22_X1 U24349 ( .A1(n21438), .A2(keyinput121), .B1(keyinput118), .B2(
        n21437), .ZN(n21436) );
  OAI221_X1 U24350 ( .B1(n21438), .B2(keyinput121), .C1(n21437), .C2(
        keyinput118), .A(n21436), .ZN(n21439) );
  NOR4_X1 U24351 ( .A1(n21442), .A2(n21441), .A3(n21440), .A4(n21439), .ZN(
        n21491) );
  AOI22_X1 U24352 ( .A1(keyinput112), .A2(n21444), .B1(keyinput54), .B2(n21498), .ZN(n21443) );
  OAI21_X1 U24353 ( .B1(n21444), .B2(keyinput112), .A(n21443), .ZN(n21455) );
  INV_X1 U24354 ( .A(P3_LWORD_REG_15__SCAN_IN), .ZN(n21446) );
  AOI22_X1 U24355 ( .A1(n15129), .A2(keyinput62), .B1(keyinput127), .B2(n21446), .ZN(n21445) );
  OAI221_X1 U24356 ( .B1(n15129), .B2(keyinput62), .C1(n21446), .C2(
        keyinput127), .A(n21445), .ZN(n21454) );
  INV_X1 U24357 ( .A(DATAI_11_), .ZN(n21448) );
  AOI22_X1 U24358 ( .A1(n21449), .A2(keyinput53), .B1(keyinput42), .B2(n21448), 
        .ZN(n21447) );
  OAI221_X1 U24359 ( .B1(n21449), .B2(keyinput53), .C1(n21448), .C2(keyinput42), .A(n21447), .ZN(n21453) );
  AOI22_X1 U24360 ( .A1(n21451), .A2(keyinput98), .B1(n12854), .B2(keyinput115), .ZN(n21450) );
  OAI221_X1 U24361 ( .B1(n21451), .B2(keyinput98), .C1(n12854), .C2(
        keyinput115), .A(n21450), .ZN(n21452) );
  NOR4_X1 U24362 ( .A1(n21455), .A2(n21454), .A3(n21453), .A4(n21452), .ZN(
        n21490) );
  AOI22_X1 U24363 ( .A1(n21458), .A2(keyinput90), .B1(n21457), .B2(keyinput60), 
        .ZN(n21456) );
  OAI221_X1 U24364 ( .B1(n21458), .B2(keyinput90), .C1(n21457), .C2(keyinput60), .A(n21456), .ZN(n21462) );
  XOR2_X1 U24365 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B(keyinput6), .Z(
        n21461) );
  XNOR2_X1 U24366 ( .A(n21459), .B(keyinput0), .ZN(n21460) );
  OR3_X1 U24367 ( .A1(n21462), .A2(n21461), .A3(n21460), .ZN(n21471) );
  AOI22_X1 U24368 ( .A1(n21465), .A2(keyinput69), .B1(keyinput95), .B2(n21464), 
        .ZN(n21463) );
  OAI221_X1 U24369 ( .B1(n21465), .B2(keyinput69), .C1(n21464), .C2(keyinput95), .A(n21463), .ZN(n21470) );
  AOI22_X1 U24370 ( .A1(n21468), .A2(keyinput28), .B1(keyinput52), .B2(n21467), 
        .ZN(n21466) );
  OAI221_X1 U24371 ( .B1(n21468), .B2(keyinput28), .C1(n21467), .C2(keyinput52), .A(n21466), .ZN(n21469) );
  NOR3_X1 U24372 ( .A1(n21471), .A2(n21470), .A3(n21469), .ZN(n21489) );
  AOI22_X1 U24373 ( .A1(n21474), .A2(keyinput45), .B1(n21473), .B2(keyinput86), 
        .ZN(n21472) );
  OAI221_X1 U24374 ( .B1(n21474), .B2(keyinput45), .C1(n21473), .C2(keyinput86), .A(n21472), .ZN(n21487) );
  INV_X1 U24375 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n21476) );
  AOI22_X1 U24376 ( .A1(n21477), .A2(keyinput108), .B1(n21476), .B2(keyinput78), .ZN(n21475) );
  OAI221_X1 U24377 ( .B1(n21477), .B2(keyinput108), .C1(n21476), .C2(
        keyinput78), .A(n21475), .ZN(n21486) );
  INV_X1 U24378 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21479) );
  AOI22_X1 U24379 ( .A1(n21480), .A2(keyinput74), .B1(keyinput43), .B2(n21479), 
        .ZN(n21478) );
  OAI221_X1 U24380 ( .B1(n21480), .B2(keyinput74), .C1(n21479), .C2(keyinput43), .A(n21478), .ZN(n21485) );
  AOI22_X1 U24381 ( .A1(n21483), .A2(keyinput94), .B1(keyinput105), .B2(n21482), .ZN(n21481) );
  OAI221_X1 U24382 ( .B1(n21483), .B2(keyinput94), .C1(n21482), .C2(
        keyinput105), .A(n21481), .ZN(n21484) );
  NOR4_X1 U24383 ( .A1(n21487), .A2(n21486), .A3(n21485), .A4(n21484), .ZN(
        n21488) );
  NAND4_X1 U24384 ( .A1(n21491), .A2(n21490), .A3(n21489), .A4(n21488), .ZN(
        n21492) );
  NOR4_X1 U24385 ( .A1(n21495), .A2(n21494), .A3(n21493), .A4(n21492), .ZN(
        n21496) );
  OAI221_X1 U24386 ( .B1(keyinput54), .B2(n21498), .C1(keyinput54), .C2(n21497), .A(n21496), .ZN(n21499) );
  XOR2_X1 U24387 ( .A(n21500), .B(n21499), .Z(U351) );
  AND2_X1 U13231 ( .A1(n10007), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13441) );
  INV_X2 U11332 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11030) );
  INV_X1 U11314 ( .A(n12813), .ZN(n12898) );
  NAND2_X1 U11203 ( .A1(n12814), .A2(n12892), .ZN(n12887) );
  BUF_X2 U11207 ( .A(n10855), .Z(n12395) );
  CLKBUF_X1 U11261 ( .A(n17457), .Z(n9727) );
  CLKBUF_X2 U11191 ( .A(n11892), .Z(n9723) );
  INV_X1 U11167 ( .A(n17363), .ZN(n17345) );
  AND2_X2 U12921 ( .A1(n12401), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10937) );
  OAI21_X2 U11405 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19257), .A(n17005), 
        .ZN(n18289) );
  NAND2_X1 U15831 ( .A1(n18289), .A2(n18251), .ZN(n18218) );
  CLKBUF_X1 U11172 ( .A(n14475), .Z(n14228) );
  CLKBUF_X1 U11187 ( .A(n12768), .Z(n14028) );
  CLKBUF_X1 U11209 ( .A(n12924), .Z(n12929) );
  NAND2_X2 U11260 ( .A1(n19226), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11861) );
  CLKBUF_X1 U11308 ( .A(n12976), .Z(n14314) );
  CLKBUF_X1 U11310 ( .A(n10821), .Z(n10822) );
  CLKBUF_X1 U11330 ( .A(n11293), .Z(n11716) );
  OR2_X1 U11442 ( .A1(n14206), .A2(n14205), .ZN(n14324) );
  NAND2_X1 U11727 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13476) );
  INV_X1 U11728 ( .A(n13685), .ZN(n20229) );
  INV_X2 U11936 ( .A(n18640), .ZN(n12085) );
  AND2_X1 U12613 ( .A1(n10222), .A2(n12126), .ZN(n17956) );
  CLKBUF_X2 U12633 ( .A(n10823), .Z(n13436) );
  CLKBUF_X1 U12744 ( .A(n19435), .Z(n19467) );
  CLKBUF_X1 U12778 ( .A(n16137), .Z(n16455) );
  CLKBUF_X1 U13344 ( .A(n16989), .Z(n16990) );
  AND2_X1 U13523 ( .A1(n9826), .A2(n13492), .ZN(n21501) );
  CLKBUF_X1 U13571 ( .A(n17909), .Z(n17917) );
endmodule

