

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9590, n9591, n9592, n9593, n9594, n9596, n9597, n9598, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808;

  AOI211_X1 U11034 ( .C1(n14541), .C2(n19832), .A(n13973), .B(n13972), .ZN(
        n13974) );
  XNOR2_X1 U11035 ( .A(n13989), .B(n13975), .ZN(n14316) );
  NAND2_X1 U11036 ( .A1(n15017), .A2(n9676), .ZN(n15016) );
  XNOR2_X1 U11037 ( .A(n12394), .B(n12396), .ZN(n14756) );
  NAND2_X1 U11038 ( .A1(n13654), .A2(n13657), .ZN(n13658) );
  NAND2_X1 U11039 ( .A1(n12749), .A2(n12748), .ZN(n15980) );
  AOI21_X1 U11040 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15614), .A(
        n12146), .ZN(n12153) );
  NOR2_X1 U11041 ( .A1(n10310), .A2(n10321), .ZN(n10496) );
  CLKBUF_X1 U11042 ( .A(n11054), .Z(n11294) );
  OAI21_X1 U11043 ( .B1(n12202), .B2(n12209), .A(n12201), .ZN(n12204) );
  INV_X1 U11044 ( .A(n12195), .ZN(n10101) );
  INV_X1 U11045 ( .A(n13823), .ZN(n17943) );
  CLKBUF_X2 U11046 ( .A(n10272), .Z(n10273) );
  CLKBUF_X2 U11047 ( .A(n10720), .Z(n12521) );
  AND2_X1 U11048 ( .A1(n12485), .A2(n13211), .ZN(n12341) );
  AND2_X1 U11049 ( .A1(n12484), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10388) );
  AND2_X1 U11050 ( .A1(n10335), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10482) );
  AND2_X1 U11051 ( .A1(n12315), .A2(n10332), .ZN(n12332) );
  INV_X1 U11052 ( .A(n11539), .ZN(n11484) );
  CLKBUF_X2 U11054 ( .A(n11342), .Z(n9597) );
  INV_X1 U11055 ( .A(n11579), .ZN(n11478) );
  BUF_X2 U11056 ( .A(n11377), .Z(n11916) );
  CLKBUF_X2 U11057 ( .A(n10227), .Z(n19044) );
  OR2_X2 U11058 ( .A1(n11331), .A2(n11330), .ZN(n11421) );
  CLKBUF_X1 U11059 ( .A(n13824), .Z(n15432) );
  CLKBUF_X2 U11060 ( .A(n15436), .Z(n16905) );
  INV_X1 U11061 ( .A(n13827), .ZN(n16886) );
  INV_X2 U11062 ( .A(n9644), .ZN(n16635) );
  INV_X2 U11063 ( .A(n13758), .ZN(n16895) );
  AND4_X1 U11064 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11414) );
  CLKBUF_X2 U11065 ( .A(n10194), .Z(n19023) );
  NAND2_X2 U11066 ( .A1(n10163), .A2(n10162), .ZN(n11021) );
  AND2_X1 U11067 ( .A1(n11307), .A2(n11313), .ZN(n11463) );
  AND2_X1 U11068 ( .A1(n11307), .A2(n11316), .ZN(n11498) );
  AND2_X1 U11069 ( .A1(n11313), .A2(n13116), .ZN(n11342) );
  AND2_X1 U11070 ( .A1(n9936), .A2(n13115), .ZN(n11986) );
  CLKBUF_X2 U11071 ( .A(n11332), .Z(n11985) );
  CLKBUF_X2 U11072 ( .A(n10344), .Z(n12490) );
  INV_X2 U11073 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15352) );
  AND2_X1 U11074 ( .A1(n10216), .A2(n10240), .ZN(n11213) );
  CLKBUF_X3 U11075 ( .A(n11332), .Z(n12069) );
  AOI211_X1 U11076 ( .C1(n10644), .C2(P2_REIP_REG_1__SCAN_IN), .A(n10245), .B(
        n10244), .ZN(n10246) );
  NAND2_X1 U11077 ( .A1(n12838), .A2(n12837), .ZN(n12866) );
  OR2_X1 U11078 ( .A1(n14334), .A2(n9851), .ZN(n9852) );
  AND2_X2 U11079 ( .A1(n19932), .A2(n11424), .ZN(n13949) );
  NOR2_X1 U11080 ( .A1(n19954), .A2(n19949), .ZN(n13124) );
  AND2_X1 U11081 ( .A1(n12315), .A2(n10343), .ZN(n12342) );
  INV_X1 U11082 ( .A(n12197), .ZN(n10321) );
  OR2_X1 U11083 ( .A1(n16557), .A2(n13757), .ZN(n10112) );
  AND4_X1 U11084 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11413) );
  CLKBUF_X2 U11085 ( .A(n13342), .Z(n13938) );
  OR2_X1 U11086 ( .A1(n14294), .A2(n9898), .ZN(n14308) );
  INV_X1 U11087 ( .A(n19949), .ZN(n9937) );
  AND3_X1 U11088 ( .A1(n11420), .A2(n11419), .A3(n11418), .ZN(n11431) );
  INV_X1 U11089 ( .A(n10865), .ZN(n10895) );
  OR2_X2 U11090 ( .A1(n11215), .A2(n10125), .ZN(n13256) );
  NOR2_X1 U11091 ( .A1(n10310), .A2(n9592), .ZN(n19084) );
  OR2_X1 U11092 ( .A1(n10320), .A2(n10313), .ZN(n19417) );
  OR2_X1 U11093 ( .A1(n10320), .A2(n10315), .ZN(n19489) );
  NAND2_X1 U11095 ( .A1(n13045), .A2(n13044), .ZN(n13093) );
  NAND2_X1 U11096 ( .A1(n9982), .A2(n11646), .ZN(n13137) );
  OR2_X1 U11098 ( .A1(n10314), .A2(n10313), .ZN(n19137) );
  CLKBUF_X3 U11099 ( .A(n10719), .Z(n19028) );
  INV_X1 U11100 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13211) );
  INV_X1 U11101 ( .A(n19843), .ZN(n19822) );
  INV_X1 U11102 ( .A(n11438), .ZN(n14209) );
  NAND4_X2 U11103 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n19932) );
  OAI21_X1 U11104 ( .B1(n13238), .B2(n11021), .A(n10721), .ZN(n12501) );
  INV_X1 U11105 ( .A(n18676), .ZN(n9969) );
  NOR2_X2 U11106 ( .A1(n15980), .A2(n15981), .ZN(n15979) );
  OR2_X1 U11107 ( .A1(n14316), .A2(n19924), .ZN(n9897) );
  AOI211_X1 U11108 ( .C1(n15950), .C2(n15828), .A(n14904), .B(n14903), .ZN(
        n14905) );
  NAND2_X1 U11109 ( .A1(n10309), .A2(n10283), .ZN(n12202) );
  INV_X1 U11111 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19544) );
  NOR2_X2 U11112 ( .A1(n9719), .A2(n9718), .ZN(n16702) );
  INV_X1 U11113 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18385) );
  OR2_X1 U11114 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13755), .ZN(
        n9590) );
  OR2_X1 U11115 ( .A1(n18426), .A2(n17568), .ZN(n9591) );
  AND2_X1 U11116 ( .A1(n11315), .A2(n11316), .ZN(n11377) );
  AOI21_X2 U11117 ( .B1(n13256), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10224), 
        .ZN(n10225) );
  NOR2_X2 U11118 ( .A1(n16864), .A2(n16433), .ZN(n16865) );
  AND2_X4 U11120 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10341) );
  MUX2_X2 U11122 ( .A(n9667), .B(n14310), .S(n14492), .Z(n14311) );
  XNOR2_X1 U11123 ( .A(n13093), .B(n13046), .ZN(n13092) );
  NAND2_X2 U11124 ( .A1(n10012), .A2(n10010), .ZN(n10719) );
  XNOR2_X2 U11125 ( .A(n15492), .B(n15491), .ZN(n17514) );
  NAND2_X2 U11126 ( .A1(n17525), .A2(n15489), .ZN(n15492) );
  NOR2_X2 U11127 ( .A1(n10736), .A2(n10735), .ZN(n10770) );
  XNOR2_X1 U11128 ( .A(n10309), .B(n10308), .ZN(n12197) );
  NOR3_X2 U11129 ( .A1(n14375), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14324), .ZN(n14343) );
  NAND2_X2 U11130 ( .A1(n10868), .A2(n10867), .ZN(n14916) );
  XNOR2_X2 U11131 ( .A(n10759), .B(n10739), .ZN(n13621) );
  NAND2_X2 U11132 ( .A1(n10738), .A2(n18788), .ZN(n10759) );
  AND2_X1 U11133 ( .A1(n9611), .A2(n9703), .ZN(n10930) );
  NAND2_X1 U11135 ( .A1(n10839), .A2(n15281), .ZN(n14949) );
  NAND2_X1 U11136 ( .A1(n14756), .A2(n14755), .ZN(n14754) );
  AND2_X1 U11137 ( .A1(n10018), .A2(n10021), .ZN(n12394) );
  OR2_X1 U11138 ( .A1(n13602), .A2(n13688), .ZN(n9734) );
  INV_X1 U11139 ( .A(n13658), .ZN(n14492) );
  AND2_X1 U11140 ( .A1(n10302), .A2(n12845), .ZN(n13454) );
  AND2_X1 U11141 ( .A1(n10302), .A2(n10101), .ZN(n19370) );
  AND2_X1 U11142 ( .A1(n9854), .A2(n11606), .ZN(n9853) );
  CLKBUF_X2 U11143 ( .A(n12210), .Z(n18983) );
  AND2_X1 U11144 ( .A1(n12714), .A2(n12713), .ZN(n11043) );
  AND2_X1 U11145 ( .A1(n10237), .A2(n10236), .ZN(n10971) );
  NAND3_X1 U11146 ( .A1(n9939), .A2(n12904), .A3(n9938), .ZN(n12156) );
  AND2_X1 U11147 ( .A1(n12501), .A2(n10233), .ZN(n10237) );
  BUF_X1 U11148 ( .A(n11436), .Z(n13073) );
  NOR2_X1 U11149 ( .A1(n10721), .A2(n18596), .ZN(n10241) );
  AND2_X1 U11150 ( .A1(n13238), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12601) );
  INV_X1 U11151 ( .A(n11021), .ZN(n11023) );
  NAND2_X1 U11152 ( .A1(n10227), .A2(n19016), .ZN(n10214) );
  CLKBUF_X2 U11153 ( .A(n10205), .Z(n19033) );
  NAND2_X2 U11154 ( .A1(n13238), .A2(n11021), .ZN(n10721) );
  INV_X2 U11155 ( .A(n9590), .ZN(n9608) );
  CLKBUF_X2 U11156 ( .A(n15436), .Z(n16810) );
  CLKBUF_X2 U11157 ( .A(n11463), .Z(n12071) );
  CLKBUF_X2 U11158 ( .A(n12046), .Z(n12079) );
  BUF_X2 U11159 ( .A(n11468), .Z(n12082) );
  CLKBUF_X2 U11160 ( .A(n9604), .Z(n9606) );
  BUF_X2 U11161 ( .A(n11986), .Z(n12073) );
  AND2_X1 U11162 ( .A1(n10041), .A2(n10039), .ZN(n11304) );
  AOI21_X1 U11163 ( .B1(n11302), .B2(n18977), .A(n10040), .ZN(n10039) );
  XNOR2_X1 U11164 ( .A(n14876), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14873) );
  XNOR2_X1 U11165 ( .A(n10006), .B(n12100), .ZN(n13885) );
  NAND2_X1 U11166 ( .A1(n9850), .A2(n14308), .ZN(n14318) );
  AOI21_X1 U11167 ( .B1(n14561), .B2(n15692), .A(n14331), .ZN(n14332) );
  NAND2_X1 U11168 ( .A1(n14308), .A2(n9799), .ZN(n14295) );
  CLKBUF_X1 U11169 ( .A(n15008), .Z(n15220) );
  NOR2_X2 U11170 ( .A1(n14037), .A2(n14039), .ZN(n14027) );
  NAND2_X1 U11171 ( .A1(n17250), .A2(n17253), .ZN(n17249) );
  XNOR2_X1 U11172 ( .A(n12419), .B(n9697), .ZN(n14751) );
  NAND2_X1 U11173 ( .A1(n14754), .A2(n12398), .ZN(n12419) );
  AOI21_X1 U11174 ( .B1(n9919), .B2(n9613), .A(n9627), .ZN(n9773) );
  NOR2_X1 U11175 ( .A1(n15795), .A2(n15794), .ZN(n15793) );
  NAND3_X1 U11176 ( .A1(n10495), .A2(n10107), .A3(n10449), .ZN(n13619) );
  AND2_X1 U11177 ( .A1(n9957), .A2(n9956), .ZN(n15795) );
  INV_X1 U11178 ( .A(n13616), .ZN(n10495) );
  AND2_X1 U11179 ( .A1(n9775), .A2(n9777), .ZN(n9776) );
  OR2_X1 U11180 ( .A1(n13587), .A2(n11746), .ZN(n13736) );
  AOI21_X1 U11181 ( .B1(n12352), .B2(n10020), .A(n9696), .ZN(n10021) );
  OR2_X1 U11182 ( .A1(n14844), .A2(n10019), .ZN(n10018) );
  AOI21_X1 U11183 ( .B1(n14431), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14492), .ZN(n9856) );
  NAND2_X1 U11184 ( .A1(n14896), .A2(n14907), .ZN(n9772) );
  AND2_X1 U11185 ( .A1(n9780), .A2(n11745), .ZN(n9775) );
  NOR2_X1 U11186 ( .A1(n15687), .A2(n9962), .ZN(n9961) );
  NAND2_X1 U11187 ( .A1(n10416), .A2(n10417), .ZN(n10108) );
  NOR2_X1 U11188 ( .A1(n9955), .A2(n9953), .ZN(n9952) );
  AOI21_X1 U11189 ( .B1(n14444), .B2(n14430), .A(n14446), .ZN(n14431) );
  OR2_X1 U11190 ( .A1(n13653), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15688) );
  OR2_X1 U11191 ( .A1(n14286), .A2(n14464), .ZN(n14444) );
  NAND2_X1 U11192 ( .A1(n14443), .A2(n14454), .ZN(n9955) );
  AND2_X1 U11193 ( .A1(n11654), .A2(n11653), .ZN(n9793) );
  OR2_X1 U11194 ( .A1(n13658), .A2(n14668), .ZN(n14454) );
  NAND2_X1 U11195 ( .A1(n9810), .A2(n13157), .ZN(n13333) );
  INV_X4 U11196 ( .A(n14492), .ZN(n9593) );
  OAI21_X1 U11197 ( .B1(n17389), .B2(n10115), .A(n17483), .ZN(n15500) );
  AND2_X1 U11198 ( .A1(n13654), .A2(n11672), .ZN(n13476) );
  INV_X1 U11199 ( .A(n9591), .ZN(n9610) );
  NAND2_X1 U11200 ( .A1(n9811), .A2(n13094), .ZN(n13154) );
  NAND2_X1 U11201 ( .A1(n11669), .A2(n11668), .ZN(n13654) );
  AND4_X1 U11202 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10369) );
  NOR2_X2 U11203 ( .A1(n17068), .A2(n17577), .ZN(n17484) );
  NOR4_X2 U11204 ( .A1(n17028), .A2(n17119), .A3(n17121), .A4(n16952), .ZN(
        n16993) );
  CLKBUF_X1 U11205 ( .A(n12185), .Z(n14268) );
  INV_X1 U11206 ( .A(n19417), .ZN(n19414) );
  NAND2_X1 U11207 ( .A1(n11578), .A2(n9853), .ZN(n11671) );
  AND2_X1 U11208 ( .A1(n11635), .A2(n13075), .ZN(n9789) );
  NAND2_X1 U11209 ( .A1(n9884), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17481) );
  OR2_X1 U11210 ( .A1(n10314), .A2(n10315), .ZN(n19211) );
  NAND2_X2 U11211 ( .A1(n14270), .A2(n13074), .ZN(n14279) );
  AND2_X1 U11212 ( .A1(n10298), .A2(n12845), .ZN(n13490) );
  AND2_X1 U11213 ( .A1(n10301), .A2(n12845), .ZN(n19240) );
  AND2_X1 U11214 ( .A1(n12729), .A2(n10299), .ZN(n10302) );
  AND2_X1 U11215 ( .A1(n12729), .A2(n10300), .ZN(n10298) );
  AND2_X1 U11216 ( .A1(n18983), .A2(n10299), .ZN(n10301) );
  XNOR2_X1 U11217 ( .A(n11555), .B(n11554), .ZN(n11613) );
  CLKBUF_X1 U11218 ( .A(n13138), .Z(n20010) );
  NAND2_X1 U11219 ( .A1(n9784), .A2(n9657), .ZN(n11555) );
  NAND2_X1 U11220 ( .A1(n12885), .A2(n12884), .ZN(n13042) );
  XNOR2_X1 U11221 ( .A(n10279), .B(n10278), .ZN(n12210) );
  XNOR2_X1 U11222 ( .A(n11622), .B(n11522), .ZN(n13138) );
  NAND2_X1 U11223 ( .A1(n9787), .A2(n9786), .ZN(n9785) );
  NAND2_X1 U11224 ( .A1(n9905), .A2(n9660), .ZN(n20009) );
  NAND2_X1 U11225 ( .A1(n9880), .A2(n9757), .ZN(n17503) );
  NOR2_X1 U11226 ( .A1(n19007), .A2(n19046), .ZN(n19504) );
  NOR2_X1 U11227 ( .A1(n19047), .A2(n19046), .ZN(n19536) );
  NOR2_X1 U11228 ( .A1(n19034), .A2(n19046), .ZN(n19529) );
  NOR2_X1 U11229 ( .A1(n19029), .A2(n19046), .ZN(n19525) );
  NOR2_X1 U11230 ( .A1(n19017), .A2(n19046), .ZN(n19515) );
  NOR2_X1 U11231 ( .A1(n19011), .A2(n19046), .ZN(n19509) );
  NAND2_X1 U11232 ( .A1(n10821), .A2(n10794), .ZN(n10812) );
  NOR2_X1 U11233 ( .A1(n13444), .A2(n13443), .ZN(n9910) );
  INV_X2 U11234 ( .A(n18851), .ZN(n18843) );
  NAND2_X4 U11235 ( .A1(n20399), .A2(n11533), .ZN(n13879) );
  NOR2_X2 U11236 ( .A1(n10819), .A2(n10814), .ZN(n10821) );
  AOI221_X1 U11237 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15632), .C1(n19729), .C2(
        n15632), .A(n19553), .ZN(n19721) );
  OAI21_X1 U11238 ( .B1(n11631), .B2(n9942), .A(n9940), .ZN(n11497) );
  NAND2_X1 U11239 ( .A1(n11562), .A2(n11561), .ZN(n20087) );
  OAI211_X1 U11240 ( .C1(n15611), .C2(n20220), .A(n11536), .B(n11535), .ZN(
        n11537) );
  XNOR2_X1 U11241 ( .A(n10608), .B(n10607), .ZN(n10606) );
  OR2_X1 U11242 ( .A1(n10782), .A2(n12521), .ZN(n10874) );
  OR2_X1 U11243 ( .A1(n11534), .A2(n13112), .ZN(n11536) );
  NAND2_X1 U11244 ( .A1(n12595), .A2(n19617), .ZN(n18961) );
  NAND2_X1 U11245 ( .A1(n10261), .A2(n10260), .ZN(n10282) );
  INV_X2 U11246 ( .A(n17166), .ZN(n17196) );
  AOI21_X1 U11247 ( .B1(n9878), .B2(n15486), .A(n9877), .ZN(n9876) );
  NAND2_X1 U11248 ( .A1(n10295), .A2(n10294), .ZN(n10608) );
  NAND2_X1 U11249 ( .A1(n11516), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11529) );
  NAND2_X1 U11250 ( .A1(n15360), .A2(n15361), .ZN(n15633) );
  AND4_X1 U11251 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10261) );
  NAND2_X1 U11252 ( .A1(n11493), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11628) );
  CLKBUF_X1 U11253 ( .A(n11215), .Z(n13233) );
  NAND2_X1 U11254 ( .A1(n10218), .A2(n10217), .ZN(n12504) );
  NAND2_X1 U11255 ( .A1(n11428), .A2(n11427), .ZN(n12911) );
  AND2_X1 U11256 ( .A1(n11440), .A2(n11455), .ZN(n12779) );
  NOR2_X1 U11257 ( .A1(n18357), .A2(n9714), .ZN(n15358) );
  NAND2_X1 U11258 ( .A1(n17950), .A2(n13823), .ZN(n9714) );
  AND3_X1 U11259 ( .A1(n9937), .A2(n19954), .A3(n19932), .ZN(n12904) );
  AND2_X2 U11260 ( .A1(n11007), .A2(n12418), .ZN(n11180) );
  NAND3_X1 U11261 ( .A1(n10223), .A2(n10221), .A3(n10222), .ZN(n10240) );
  AND2_X1 U11262 ( .A1(n10987), .A2(n12601), .ZN(n10248) );
  NOR2_X1 U11263 ( .A1(n11434), .A2(n19949), .ZN(n12881) );
  NAND3_X1 U11264 ( .A1(n13794), .A2(n13793), .A3(n13792), .ZN(n17102) );
  OR2_X1 U11265 ( .A1(n11476), .A2(n11475), .ZN(n13660) );
  AND2_X1 U11266 ( .A1(n10413), .A2(n10412), .ZN(n11048) );
  NOR2_X2 U11267 ( .A1(n13822), .A2(n13821), .ZN(n17927) );
  AND2_X1 U11268 ( .A1(n10205), .A2(n10719), .ZN(n10228) );
  NOR2_X1 U11269 ( .A1(n11021), .A2(n19010), .ZN(n10972) );
  INV_X1 U11270 ( .A(n10194), .ZN(n10977) );
  NAND2_X2 U11271 ( .A1(n9824), .A2(n9823), .ZN(n19010) );
  NOR2_X1 U11272 ( .A1(n11367), .A2(n11366), .ZN(n11372) );
  OR2_X2 U11273 ( .A1(n11361), .A2(n11360), .ZN(n19954) );
  AND2_X1 U11274 ( .A1(n11341), .A2(n10133), .ZN(n11630) );
  NAND2_X1 U11275 ( .A1(n9727), .A2(n9722), .ZN(n19016) );
  AND4_X1 U11276 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11393) );
  AND4_X1 U11277 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11412) );
  AND4_X1 U11278 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n11341) );
  AND4_X1 U11279 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11392) );
  NAND2_X1 U11280 ( .A1(n10204), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9823) );
  AND4_X1 U11281 ( .A1(n11311), .A2(n11310), .A3(n11309), .A4(n11308), .ZN(
        n11321) );
  NAND2_X1 U11282 ( .A1(n10199), .A2(n13211), .ZN(n9824) );
  AND4_X1 U11283 ( .A1(n11410), .A2(n11409), .A3(n11408), .A4(n11407), .ZN(
        n11411) );
  NOR2_X2 U11284 ( .A1(n19925), .A2(n19924), .ZN(n19926) );
  INV_X2 U11285 ( .A(n9590), .ZN(n9609) );
  INV_X2 U11286 ( .A(n14848), .ZN(n14847) );
  BUF_X4 U11287 ( .A(n15468), .Z(n9598) );
  AND4_X1 U11288 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11391) );
  INV_X1 U11289 ( .A(n16907), .ZN(n15473) );
  AND4_X1 U11290 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11390) );
  AND2_X1 U11291 ( .A1(n10164), .A2(n13211), .ZN(n9771) );
  AND2_X1 U11292 ( .A1(n10169), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9769) );
  INV_X1 U11293 ( .A(n16895), .ZN(n9594) );
  CLKBUF_X2 U11294 ( .A(n13825), .Z(n16894) );
  CLKBUF_X3 U11295 ( .A(n13826), .Z(n16909) );
  NAND2_X1 U11297 ( .A1(n9754), .A2(n9753), .ZN(n16907) );
  BUF_X2 U11298 ( .A(n15418), .Z(n16610) );
  INV_X2 U11299 ( .A(n16163), .ZN(U215) );
  INV_X1 U11300 ( .A(n16845), .ZN(n9596) );
  BUF_X2 U11301 ( .A(n11332), .Z(n11921) );
  BUF_X2 U11302 ( .A(n12072), .Z(n12051) );
  BUF_X2 U11303 ( .A(n11470), .Z(n11901) );
  INV_X2 U11304 ( .A(n16166), .ZN(n16168) );
  BUF_X2 U11305 ( .A(n13824), .Z(n16658) );
  AND2_X2 U11306 ( .A1(n10335), .A2(n13211), .ZN(n13224) );
  CLKBUF_X3 U11307 ( .A(n10328), .Z(n12486) );
  CLKBUF_X2 U11308 ( .A(n9603), .Z(n9605) );
  BUF_X2 U11309 ( .A(n12479), .Z(n12489) );
  INV_X2 U11310 ( .A(n19735), .ZN(n19672) );
  AND2_X1 U11311 ( .A1(n11306), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11314) );
  NAND2_X1 U11312 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18528), .ZN(
        n13750) );
  AND2_X1 U11313 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13115) );
  CLKBUF_X1 U11314 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n12789) );
  INV_X2 U11315 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18528) );
  INV_X2 U11316 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18549) );
  INV_X2 U11317 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18535) );
  NOR2_X2 U11318 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10343) );
  NOR2_X2 U11319 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13205) );
  AND2_X1 U11320 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10581) );
  NOR3_X2 U11321 ( .A1(n15378), .A2(n16837), .A3(n16835), .ZN(n16822) );
  INV_X2 U11322 ( .A(n9639), .ZN(n15468) );
  INV_X4 U11324 ( .A(n16907), .ZN(n16889) );
  BUF_X4 U11325 ( .A(n15418), .Z(n16888) );
  INV_X1 U11327 ( .A(n18576), .ZN(n17922) );
  NOR2_X2 U11328 ( .A1(n13837), .A2(n13836), .ZN(n18576) );
  BUF_X1 U11329 ( .A(n10272), .Z(n9601) );
  AOI21_X2 U11330 ( .B1(n10239), .B2(n13202), .A(n18596), .ZN(n10272) );
  AND2_X2 U11331 ( .A1(n14027), .A2(n9791), .ZN(n9612) );
  OAI21_X2 U11332 ( .B1(n14423), .B2(n14292), .A(n9954), .ZN(n14381) );
  AND2_X4 U11333 ( .A1(n10343), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9602) );
  OAI21_X2 U11334 ( .B1(n14916), .B2(n10869), .A(n10870), .ZN(n9896) );
  NOR2_X4 U11335 ( .A1(n9638), .A2(n13991), .ZN(n13993) );
  OR3_X4 U11336 ( .A1(n14077), .A2(n9931), .A3(n14003), .ZN(n9638) );
  NOR4_X1 U11337 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n18549), .A4(n18528), .ZN(
        n9603) );
  NOR4_X1 U11338 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n18549), .A4(n18528), .ZN(
        n9604) );
  NOR3_X2 U11339 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n16557), .ZN(n15418) );
  NAND2_X2 U11340 ( .A1(n18542), .A2(n18549), .ZN(n16557) );
  NOR2_X4 U11341 ( .A1(n15008), .A2(n10559), .ZN(n14994) );
  NAND2_X2 U11342 ( .A1(n15032), .A2(n15222), .ZN(n15008) );
  NOR2_X1 U11343 ( .A1(n13823), .A2(n16953), .ZN(n13838) );
  NOR2_X2 U11344 ( .A1(n13804), .A2(n13803), .ZN(n16953) );
  XNOR2_X1 U11345 ( .A(n11525), .B(n11523), .ZN(n11621) );
  INV_X1 U11346 ( .A(n10937), .ZN(n10223) );
  NOR2_X1 U11347 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12315) );
  NAND2_X1 U11348 ( .A1(n9838), .A2(n9837), .ZN(n9924) );
  NOR2_X1 U11349 ( .A1(n14916), .A2(n10869), .ZN(n9837) );
  XNOR2_X1 U11350 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n16008), .ZN(
        n16478) );
  CLKBUF_X1 U11351 ( .A(n11402), .Z(n12083) );
  OAI21_X1 U11352 ( .B1(n12156), .B2(n12696), .A(n12911), .ZN(n11429) );
  NAND2_X1 U11353 ( .A1(n11497), .A2(n11496), .ZN(n11525) );
  INV_X1 U11354 ( .A(n11628), .ZN(n9942) );
  AOI21_X1 U11355 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20276), .A(
        n12132), .ZN(n12147) );
  AND2_X1 U11356 ( .A1(n9893), .A2(n10493), .ZN(n10127) );
  INV_X1 U11357 ( .A(n10228), .ZN(n10938) );
  NAND2_X1 U11358 ( .A1(n13473), .A2(n13555), .ZN(n10003) );
  AND2_X1 U11359 ( .A1(n11671), .A2(n11608), .ZN(n13322) );
  NAND2_X1 U11360 ( .A1(n11578), .A2(n9854), .ZN(n11607) );
  NOR2_X2 U11361 ( .A1(n19968), .A2(n11609), .ZN(n11800) );
  NAND2_X1 U11362 ( .A1(n11424), .A2(n11421), .ZN(n13655) );
  NOR2_X1 U11363 ( .A1(n12936), .A2(n12751), .ZN(n12891) );
  NAND2_X1 U11364 ( .A1(n10156), .A2(n13211), .ZN(n10163) );
  NAND2_X1 U11365 ( .A1(n12397), .A2(n12396), .ZN(n12398) );
  AND2_X1 U11366 ( .A1(n12710), .A2(n19006), .ZN(n12854) );
  INV_X1 U11367 ( .A(n10205), .ZN(n12509) );
  INV_X1 U11368 ( .A(n10719), .ZN(n10720) );
  AOI21_X1 U11369 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10277), .ZN(n10286) );
  OR2_X1 U11370 ( .A1(n10557), .A2(n10773), .ZN(n10558) );
  INV_X1 U11371 ( .A(n11294), .ZN(n11210) );
  NAND2_X1 U11372 ( .A1(n10445), .A2(n9766), .ZN(n10447) );
  OAI21_X1 U11373 ( .B1(n10240), .B2(n10939), .A(n10231), .ZN(n10232) );
  INV_X1 U11374 ( .A(n12854), .ZN(n12413) );
  NOR3_X1 U11375 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n13756), .ZN(n13825) );
  NOR3_X1 U11376 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18371), .ZN(n13824) );
  NOR2_X1 U11377 ( .A1(n16557), .A2(n13750), .ZN(n16625) );
  NAND2_X1 U11378 ( .A1(n17488), .A2(n15499), .ZN(n9884) );
  NAND2_X1 U11379 ( .A1(n17553), .A2(n15482), .ZN(n15485) );
  OR2_X1 U11380 ( .A1(n17879), .A2(n15481), .ZN(n15482) );
  NAND2_X1 U11381 ( .A1(n13845), .A2(n15518), .ZN(n13868) );
  OR2_X1 U11382 ( .A1(n20611), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12938) );
  AND2_X1 U11383 ( .A1(n11609), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12097) );
  NOR2_X1 U11384 ( .A1(n12156), .A2(n19741), .ZN(n12157) );
  NAND2_X1 U11385 ( .A1(n9963), .A2(n9961), .ZN(n9964) );
  INV_X1 U11386 ( .A(n13644), .ZN(n9962) );
  INV_X1 U11387 ( .A(n19986), .ZN(n20097) );
  AND2_X1 U11388 ( .A1(n20010), .A2(n19929), .ZN(n20326) );
  NOR2_X1 U11389 ( .A1(n15852), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15837) );
  AND2_X1 U11390 ( .A1(n10024), .A2(n12227), .ZN(n9735) );
  NAND2_X1 U11391 ( .A1(n12476), .A2(n9744), .ZN(n9743) );
  AOI21_X1 U11392 ( .B1(n14740), .B2(n9745), .A(n12471), .ZN(n14730) );
  XNOR2_X1 U11393 ( .A(n12351), .B(n12374), .ZN(n14844) );
  NAND2_X1 U11394 ( .A1(n10054), .A2(n10053), .ZN(n10052) );
  NOR2_X1 U11395 ( .A1(n14746), .A2(n14727), .ZN(n10053) );
  NAND2_X1 U11396 ( .A1(n9838), .A2(n9926), .ZN(n9925) );
  INV_X1 U11397 ( .A(n9927), .ZN(n9926) );
  AOI21_X1 U11398 ( .B1(n10912), .B2(n10881), .A(n9839), .ZN(n9927) );
  AND4_X1 U11399 ( .A1(n10540), .A2(n10539), .A3(n10538), .A4(n10537), .ZN(
        n10552) );
  NOR3_X1 U11400 ( .A1(n14855), .A2(n10075), .A3(n14856), .ZN(n15176) );
  NAND2_X1 U11401 ( .A1(n10959), .A2(n12613), .ZN(n11218) );
  NAND2_X1 U11402 ( .A1(n12191), .A2(n19544), .ZN(n12215) );
  NAND2_X1 U11403 ( .A1(n10931), .A2(n10710), .ZN(n13237) );
  NAND2_X1 U11404 ( .A1(n10709), .A2(n12601), .ZN(n10710) );
  INV_X1 U11405 ( .A(n16003), .ZN(n12613) );
  NOR2_X2 U11406 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19688) );
  AND2_X1 U11407 ( .A1(n19277), .A2(n19715), .ZN(n19207) );
  NOR2_X1 U11408 ( .A1(n17943), .A2(n13868), .ZN(n13848) );
  OAI21_X1 U11409 ( .B1(n13866), .B2(n15523), .A(n13873), .ZN(n18403) );
  AND2_X1 U11410 ( .A1(n9875), .A2(n16478), .ZN(n16219) );
  OR2_X1 U11411 ( .A1(n16229), .A2(n16230), .ZN(n9875) );
  INV_X1 U11412 ( .A(n17248), .ZN(n9868) );
  AND2_X1 U11413 ( .A1(n17244), .A2(n9628), .ZN(n16039) );
  NOR2_X1 U11414 ( .A1(n9882), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9760) );
  OR2_X1 U11415 ( .A1(n17312), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9882) );
  NAND2_X1 U11416 ( .A1(n15485), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15486) );
  INV_X1 U11417 ( .A(n19922), .ZN(n13153) );
  XNOR2_X1 U11418 ( .A(n9637), .B(n10968), .ZN(n14871) );
  INV_X1 U11419 ( .A(n15939), .ZN(n15947) );
  INV_X1 U11420 ( .A(n18986), .ZN(n15982) );
  NAND2_X1 U11421 ( .A1(n20220), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12104) );
  INV_X1 U11422 ( .A(n13159), .ZN(n13323) );
  NOR2_X1 U11423 ( .A1(n11549), .A2(n11548), .ZN(n13051) );
  NAND2_X1 U11424 ( .A1(n10105), .A2(n10555), .ZN(n10104) );
  INV_X1 U11425 ( .A(n10553), .ZN(n10105) );
  AND4_X1 U11426 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10508) );
  AND2_X1 U11427 ( .A1(n10397), .A2(n9829), .ZN(n10727) );
  NOR3_X1 U11428 ( .A1(n10396), .A2(n9654), .A3(n9830), .ZN(n9829) );
  INV_X1 U11429 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n9716) );
  NOR2_X1 U11430 ( .A1(n9930), .A2(n13896), .ZN(n9929) );
  INV_X1 U11431 ( .A(n13889), .ZN(n9930) );
  NOR2_X1 U11432 ( .A1(n11437), .A2(n11421), .ZN(n12168) );
  NOR2_X1 U11433 ( .A1(n13990), .A2(n10005), .ZN(n10004) );
  INV_X1 U11434 ( .A(n14002), .ZN(n10005) );
  NOR2_X1 U11435 ( .A1(n9672), .A2(n9988), .ZN(n9987) );
  INV_X1 U11436 ( .A(n14073), .ZN(n9988) );
  INV_X1 U11437 ( .A(n9992), .ZN(n9788) );
  NOR2_X2 U11438 ( .A1(n11818), .A2(n15614), .ZN(n12092) );
  NOR2_X1 U11439 ( .A1(n9997), .A2(n14190), .ZN(n9994) );
  NOR2_X1 U11440 ( .A1(n10003), .A2(n10002), .ZN(n10001) );
  INV_X1 U11441 ( .A(n13588), .ZN(n10002) );
  INV_X1 U11442 ( .A(n12864), .ZN(n11635) );
  INV_X1 U11443 ( .A(n12643), .ZN(n11448) );
  NAND2_X1 U11444 ( .A1(n9932), .A2(n13942), .ZN(n9931) );
  INV_X1 U11445 ( .A(n9933), .ZN(n9932) );
  INV_X1 U11446 ( .A(n9806), .ZN(n14293) );
  NAND2_X1 U11447 ( .A1(n9809), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9808) );
  NAND2_X1 U11448 ( .A1(n9593), .A2(n14291), .ZN(n9809) );
  OR2_X1 U11449 ( .A1(n11490), .A2(n11489), .ZN(n13048) );
  INV_X1 U11450 ( .A(n19932), .ZN(n13280) );
  NAND2_X1 U11451 ( .A1(n11527), .A2(n11526), .ZN(n11614) );
  INV_X1 U11452 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13112) );
  AND2_X1 U11453 ( .A1(n11431), .A2(n11422), .ZN(n12752) );
  OR2_X1 U11454 ( .A1(n11534), .A2(n11305), .ZN(n11562) );
  NAND2_X1 U11455 ( .A1(n9832), .A2(n13070), .ZN(n9831) );
  INV_X1 U11456 ( .A(n9833), .ZN(n9832) );
  AND2_X1 U11457 ( .A1(n10730), .A2(n10753), .ZN(n10758) );
  AND2_X1 U11458 ( .A1(n14779), .A2(n15870), .ZN(n10025) );
  NOR2_X1 U11459 ( .A1(n12228), .A2(n10009), .ZN(n10008) );
  INV_X1 U11460 ( .A(n18838), .ZN(n10009) );
  OR2_X1 U11461 ( .A1(n10523), .A2(n10522), .ZN(n11069) );
  NAND2_X1 U11462 ( .A1(n9974), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9973) );
  NAND2_X1 U11463 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U11464 ( .A1(n14785), .A2(n11212), .ZN(n10058) );
  INV_X1 U11465 ( .A(n10887), .ZN(n9838) );
  AND2_X1 U11466 ( .A1(n10908), .A2(n14906), .ZN(n10909) );
  INV_X1 U11467 ( .A(n15173), .ZN(n10075) );
  AOI21_X1 U11468 ( .B1(n14954), .B2(n10080), .A(n14953), .ZN(n10079) );
  INV_X1 U11469 ( .A(n15259), .ZN(n10080) );
  INV_X1 U11470 ( .A(n14954), .ZN(n10082) );
  OR2_X1 U11471 ( .A1(n15053), .A2(n14952), .ZN(n10084) );
  NOR2_X1 U11472 ( .A1(n12970), .A2(n10047), .ZN(n10046) );
  INV_X1 U11473 ( .A(n12858), .ZN(n10047) );
  NAND2_X1 U11474 ( .A1(n10536), .A2(n10535), .ZN(n10557) );
  NAND2_X1 U11475 ( .A1(n10289), .A2(n10288), .ZN(n9818) );
  NAND2_X1 U11476 ( .A1(n9600), .A2(n11055), .ZN(n10351) );
  INV_X1 U11477 ( .A(n9916), .ZN(n9914) );
  NOR2_X1 U11478 ( .A1(n13575), .A2(n13402), .ZN(n9916) );
  NOR2_X1 U11479 ( .A1(n10895), .A2(n13402), .ZN(n9917) );
  AND2_X1 U11480 ( .A1(n18983), .A2(n10300), .ZN(n10076) );
  NAND2_X1 U11481 ( .A1(n9767), .A2(n12729), .ZN(n10322) );
  NAND2_X1 U11482 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n9731) );
  AOI22_X1 U11483 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U11484 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n9729) );
  NAND2_X1 U11485 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n9724) );
  NAND2_X1 U11486 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n9726) );
  NOR2_X1 U11487 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12587) );
  OAI21_X1 U11488 ( .B1(n16176), .B2(n15514), .A(n18413), .ZN(n13867) );
  NOR4_X1 U11489 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n18549), .ZN(n15424) );
  NOR4_X1 U11490 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n18549), .A4(n18528), .ZN(
        n15423) );
  AOI21_X1 U11491 ( .B1(n16810), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n15422), .ZN(n15430) );
  NOR2_X1 U11492 ( .A1(n17075), .A2(n15490), .ZN(n15466) );
  NAND2_X1 U11493 ( .A1(n15517), .A2(n13874), .ZN(n15360) );
  AND2_X1 U11494 ( .A1(n19954), .A2(n11424), .ZN(n12643) );
  OR2_X1 U11495 ( .A1(n20628), .A2(n13280), .ZN(n13300) );
  AND2_X1 U11496 ( .A1(n13304), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13308) );
  INV_X1 U11497 ( .A(n11424), .ZN(n12979) );
  NOR2_X1 U11498 ( .A1(n9993), .A2(n9999), .ZN(n9992) );
  INV_X1 U11499 ( .A(n14146), .ZN(n9999) );
  INV_X1 U11500 ( .A(n9994), .ZN(n9993) );
  CLKBUF_X1 U11501 ( .A(n14122), .Z(n14123) );
  OR2_X1 U11502 ( .A1(n13387), .A2(n9781), .ZN(n9777) );
  NAND2_X1 U11503 ( .A1(n13387), .A2(n9779), .ZN(n9778) );
  AND2_X1 U11504 ( .A1(n9782), .A2(n9781), .ZN(n9779) );
  AOI21_X1 U11505 ( .B1(n13322), .B2(n11800), .A(n11612), .ZN(n13361) );
  INV_X1 U11506 ( .A(n19741), .ZN(n12937) );
  INV_X1 U11507 ( .A(n13949), .ZN(n13945) );
  OR2_X1 U11508 ( .A1(n14327), .A2(n14325), .ZN(n9813) );
  INV_X1 U11509 ( .A(n14375), .ZN(n14353) );
  NAND2_X1 U11510 ( .A1(n9964), .A2(n9901), .ZN(n9904) );
  INV_X1 U11511 ( .A(n15688), .ZN(n9902) );
  NAND2_X1 U11512 ( .A1(n9648), .A2(n13512), .ZN(n13562) );
  AOI21_X1 U11513 ( .B1(n13480), .B2(n9796), .A(n9664), .ZN(n9795) );
  INV_X1 U11514 ( .A(n13480), .ZN(n9797) );
  AND2_X1 U11515 ( .A1(n14679), .A2(n19914), .ZN(n15740) );
  NAND2_X1 U11516 ( .A1(n13333), .A2(n13332), .ZN(n9798) );
  NAND2_X1 U11517 ( .A1(n9801), .A2(n11447), .ZN(n11518) );
  INV_X1 U11518 ( .A(n11446), .ZN(n11447) );
  INV_X1 U11519 ( .A(n11818), .ZN(n14710) );
  AND2_X1 U11520 ( .A1(n12752), .A2(n13289), .ZN(n14712) );
  INV_X1 U11521 ( .A(n11637), .ZN(n20197) );
  AND2_X1 U11522 ( .A1(n20428), .A2(n20097), .ZN(n20278) );
  INV_X1 U11523 ( .A(n20323), .ZN(n20327) );
  INV_X1 U11524 ( .A(n20127), .ZN(n20396) );
  NOR2_X1 U11525 ( .A1(n20010), .A2(n19929), .ZN(n20350) );
  AND2_X1 U11526 ( .A1(n20281), .A2(n20097), .ZN(n20435) );
  INV_X1 U11527 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20467) );
  INV_X1 U11528 ( .A(n20149), .ZN(n20425) );
  AND2_X1 U11529 ( .A1(n9816), .A2(n20197), .ZN(n20426) );
  OR2_X1 U11530 ( .A1(n12153), .A2(n12165), .ZN(n12154) );
  AND2_X1 U11531 ( .A1(n12936), .A2(n12935), .ZN(n15597) );
  OR2_X1 U11532 ( .A1(n15820), .A2(n9959), .ZN(n9957) );
  NAND2_X1 U11533 ( .A1(n11223), .A2(n9960), .ZN(n9959) );
  INV_X1 U11534 ( .A(n15819), .ZN(n9960) );
  NAND2_X1 U11535 ( .A1(n18764), .A2(n11223), .ZN(n9958) );
  NOR2_X1 U11536 ( .A1(n18764), .A2(n15829), .ZN(n15820) );
  NAND2_X1 U11537 ( .A1(n10854), .A2(n9631), .ZN(n15852) );
  NOR2_X1 U11538 ( .A1(n10831), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10805) );
  OR2_X1 U11539 ( .A1(n18631), .A2(n18632), .ZN(n9971) );
  INV_X1 U11540 ( .A(n13565), .ZN(n12228) );
  AND2_X1 U11541 ( .A1(n9625), .A2(n9685), .ZN(n10024) );
  NAND2_X1 U11542 ( .A1(n9736), .A2(n9659), .ZN(n12855) );
  INV_X1 U11543 ( .A(n13424), .ZN(n9736) );
  OAI22_X1 U11544 ( .A1(n14751), .A2(n9748), .B1(n9751), .B2(n12438), .ZN(
        n14734) );
  NAND2_X1 U11545 ( .A1(n9750), .A2(n9749), .ZN(n9748) );
  INV_X1 U11546 ( .A(n14750), .ZN(n9749) );
  NAND2_X1 U11547 ( .A1(n9690), .A2(n9733), .ZN(n9732) );
  INV_X1 U11548 ( .A(n15866), .ZN(n9733) );
  AND3_X1 U11549 ( .A1(n11123), .A2(n11122), .A3(n11121), .ZN(n15303) );
  INV_X1 U11550 ( .A(n13427), .ZN(n10064) );
  OAI22_X1 U11551 ( .A1(n12844), .A2(n12843), .B1(n12509), .B2(n12220), .ZN(
        n13424) );
  AND2_X1 U11552 ( .A1(n12503), .A2(n12502), .ZN(n12607) );
  NAND2_X1 U11553 ( .A1(n10975), .A2(n19016), .ZN(n10218) );
  NOR2_X1 U11554 ( .A1(n12580), .A2(n9600), .ZN(n12595) );
  INV_X1 U11555 ( .A(n10054), .ZN(n10051) );
  NAND2_X1 U11556 ( .A1(n9984), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9983) );
  NOR2_X1 U11557 ( .A1(n11229), .A2(n14900), .ZN(n9984) );
  INV_X1 U11558 ( .A(n11252), .ZN(n9972) );
  NOR3_X1 U11559 ( .A1(n9636), .A2(n10059), .A3(n10061), .ZN(n11211) );
  NOR2_X1 U11560 ( .A1(n9636), .A2(n10059), .ZN(n14796) );
  OR2_X1 U11561 ( .A1(n15816), .A2(n10865), .ZN(n10912) );
  AND2_X1 U11562 ( .A1(n10908), .A2(n10907), .ZN(n14896) );
  NOR2_X1 U11563 ( .A1(n9658), .A2(n9886), .ZN(n9885) );
  INV_X1 U11564 ( .A(n14934), .ZN(n9886) );
  INV_X1 U11565 ( .A(n14935), .ZN(n9889) );
  OR3_X1 U11566 ( .A1(n15575), .A2(n10865), .A3(n20668), .ZN(n14934) );
  AND2_X1 U11567 ( .A1(n14949), .A2(n10840), .ZN(n9888) );
  INV_X1 U11568 ( .A(n14975), .ZN(n10090) );
  NAND2_X1 U11569 ( .A1(n10093), .A2(n10090), .ZN(n10089) );
  NOR2_X1 U11570 ( .A1(n10095), .A2(n10094), .ZN(n10093) );
  INV_X1 U11571 ( .A(n14990), .ZN(n10094) );
  INV_X1 U11572 ( .A(n14960), .ZN(n10092) );
  AND2_X1 U11573 ( .A1(n11190), .A2(n11189), .ZN(n14856) );
  NAND2_X1 U11574 ( .A1(n9848), .A2(n10895), .ZN(n9847) );
  INV_X1 U11575 ( .A(n14957), .ZN(n9848) );
  INV_X1 U11576 ( .A(n15315), .ZN(n10097) );
  INV_X1 U11577 ( .A(n9919), .ZN(n9918) );
  AOI21_X1 U11578 ( .B1(n15057), .B2(n10553), .A(n10106), .ZN(n10102) );
  NAND2_X1 U11579 ( .A1(n13533), .A2(n20652), .ZN(n10107) );
  NAND2_X1 U11580 ( .A1(n13391), .A2(n10756), .ZN(n13535) );
  XNOR2_X1 U11581 ( .A(n10446), .B(n10447), .ZN(n13533) );
  CLKBUF_X1 U11582 ( .A(n10341), .Z(n10342) );
  NAND2_X1 U11583 ( .A1(n12548), .A2(n12207), .ZN(n12725) );
  OR2_X1 U11584 ( .A1(n12413), .A2(n12208), .ZN(n12723) );
  NAND2_X1 U11585 ( .A1(n12217), .A2(n12216), .ZN(n12726) );
  NAND2_X1 U11586 ( .A1(n9737), .A2(n13457), .ZN(n12614) );
  OR2_X1 U11587 ( .A1(n19139), .A2(n19709), .ZN(n19445) );
  NOR2_X1 U11588 ( .A1(n15995), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10713) );
  NAND2_X1 U11589 ( .A1(n9706), .A2(n17938), .ZN(n13839) );
  INV_X1 U11590 ( .A(n13838), .ZN(n9706) );
  NOR2_X1 U11591 ( .A1(n16272), .A2(n16529), .ZN(n9866) );
  NOR2_X1 U11592 ( .A1(n9868), .A2(n16529), .ZN(n9867) );
  INV_X1 U11593 ( .A(n17294), .ZN(n9862) );
  NAND2_X1 U11594 ( .A1(n16317), .A2(n9863), .ZN(n9861) );
  NOR2_X1 U11595 ( .A1(n17294), .A2(n9865), .ZN(n9863) );
  INV_X1 U11596 ( .A(n17306), .ZN(n9865) );
  INV_X1 U11597 ( .A(n13875), .ZN(n15635) );
  NAND2_X1 U11598 ( .A1(n15500), .A2(n9759), .ZN(n17362) );
  AND2_X1 U11599 ( .A1(n10034), .A2(n9679), .ZN(n9759) );
  OR2_X1 U11600 ( .A1(n17710), .A2(n17704), .ZN(n10034) );
  AOI21_X1 U11601 ( .B1(n15494), .B2(n17840), .A(n9881), .ZN(n9880) );
  NAND2_X1 U11602 ( .A1(n9758), .A2(n15494), .ZN(n9757) );
  INV_X1 U11603 ( .A(n17505), .ZN(n9881) );
  NAND2_X1 U11604 ( .A1(n17514), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17513) );
  INV_X1 U11605 ( .A(n15486), .ZN(n9879) );
  INV_X1 U11606 ( .A(n17543), .ZN(n9878) );
  NAND2_X1 U11607 ( .A1(n17544), .A2(n17543), .ZN(n17542) );
  INV_X1 U11608 ( .A(n18403), .ZN(n16171) );
  INV_X1 U11609 ( .A(n13750), .ZN(n9717) );
  NOR2_X1 U11610 ( .A1(n12976), .A2(n12642), .ZN(n20628) );
  NAND2_X1 U11611 ( .A1(n14270), .A2(n12184), .ZN(n14263) );
  INV_X1 U11612 ( .A(n14270), .ZN(n14275) );
  NAND2_X1 U11613 ( .A1(n9906), .A2(n11628), .ZN(n9905) );
  NAND2_X1 U11614 ( .A1(n11627), .A2(n11629), .ZN(n9906) );
  NAND2_X1 U11615 ( .A1(n9785), .A2(n12767), .ZN(n13102) );
  AND2_X1 U11616 ( .A1(n9816), .A2(n11637), .ZN(n20199) );
  INV_X1 U11617 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20276) );
  AOI21_X1 U11618 ( .B1(n13136), .B2(n13135), .A(n20097), .ZN(n19922) );
  OR2_X1 U11619 ( .A1(n20049), .A2(n20047), .ZN(n20094) );
  NOR3_X1 U11620 ( .A1(n10782), .A2(n10780), .A3(P2_EBX_REG_9__SCAN_IN), .ZN(
        n10784) );
  AND2_X1 U11621 ( .A1(n18851), .A2(n19044), .ZN(n18848) );
  AND2_X1 U11622 ( .A1(n12534), .A2(n12613), .ZN(n18851) );
  OAI211_X1 U11623 ( .C1(n14730), .C2(n9743), .A(n9740), .B(n9738), .ZN(n12535) );
  INV_X1 U11624 ( .A(n9739), .ZN(n9738) );
  OAI22_X1 U11625 ( .A1(n14729), .A2(n9743), .B1(n12476), .B2(n9744), .ZN(
        n9739) );
  INV_X1 U11626 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14900) );
  NAND2_X1 U11627 ( .A1(n12586), .A2(n10591), .ZN(n15953) );
  AND2_X1 U11628 ( .A1(n15953), .A2(n12672), .ZN(n15944) );
  NAND3_X1 U11629 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19688), .A3(n19553), 
        .ZN(n15063) );
  AND2_X1 U11630 ( .A1(n10590), .A2(n12418), .ZN(n15939) );
  INV_X1 U11631 ( .A(n11219), .ZN(n10057) );
  XNOR2_X1 U11632 ( .A(n10966), .B(n10965), .ZN(n14875) );
  INV_X1 U11633 ( .A(n15330), .ZN(n18982) );
  INV_X1 U11634 ( .A(n15978), .ZN(n18977) );
  OR2_X1 U11635 ( .A1(n11218), .A2(n11217), .ZN(n18986) );
  INV_X1 U11636 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19720) );
  OR2_X1 U11637 ( .A1(n12204), .A2(n12711), .ZN(n19715) );
  INV_X1 U11638 ( .A(n18573), .ZN(n18589) );
  AOI21_X1 U11639 ( .B1(n16225), .B2(n16578), .A(n16214), .ZN(n9874) );
  NAND2_X1 U11640 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16473), .ZN(n16549) );
  INV_X1 U11641 ( .A(n17036), .ZN(n17959) );
  NOR2_X2 U11642 ( .A1(n15397), .A2(n15396), .ZN(n17068) );
  NAND2_X1 U11643 ( .A1(n16062), .A2(n17565), .ZN(n10028) );
  NAND2_X1 U11644 ( .A1(n10032), .A2(n10030), .ZN(n16061) );
  NAND2_X1 U11645 ( .A1(n16016), .A2(n10031), .ZN(n10030) );
  NAND2_X1 U11646 ( .A1(n16021), .A2(n16022), .ZN(n10032) );
  INV_X1 U11647 ( .A(n16022), .ZN(n10031) );
  OR2_X1 U11648 ( .A1(n11602), .A2(n11601), .ZN(n13325) );
  OR2_X1 U11649 ( .A1(n11508), .A2(n11507), .ZN(n13049) );
  AOI21_X1 U11650 ( .B1(n11628), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9941), 
        .ZN(n9940) );
  INV_X1 U11651 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10135) );
  AND2_X1 U11652 ( .A1(n12104), .A2(n12103), .ZN(n12107) );
  AND2_X1 U11653 ( .A1(n12106), .A2(n12104), .ZN(n12133) );
  XNOR2_X1 U11654 ( .A(n11305), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12134) );
  OR2_X1 U11655 ( .A1(n12119), .A2(n12120), .ZN(n12121) );
  INV_X1 U11656 ( .A(n11645), .ZN(n9855) );
  INV_X1 U11657 ( .A(n11636), .ZN(n11578) );
  INV_X1 U11658 ( .A(n19954), .ZN(n11434) );
  OR2_X1 U11659 ( .A1(n11664), .A2(n11663), .ZN(n13648) );
  INV_X1 U11660 ( .A(n13325), .ZN(n13327) );
  OR2_X1 U11661 ( .A1(n11590), .A2(n11589), .ZN(n13159) );
  NOR2_X1 U11662 ( .A1(n11512), .A2(n9803), .ZN(n9804) );
  CLKBUF_X1 U11663 ( .A(n12353), .Z(n12483) );
  OR2_X1 U11664 ( .A1(n14764), .A2(n14843), .ZN(n10019) );
  NAND2_X1 U11665 ( .A1(n10077), .A2(n10127), .ZN(n10534) );
  AND2_X1 U11666 ( .A1(n12587), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10224) );
  NOR2_X1 U11667 ( .A1(n19044), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11020) );
  INV_X1 U11668 ( .A(n19010), .ZN(n10943) );
  OR2_X1 U11669 ( .A1(n13860), .A2(n13861), .ZN(n13856) );
  NAND2_X1 U11670 ( .A1(n18549), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13756) );
  NAND2_X1 U11671 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U11672 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18535), .ZN(
        n13757) );
  INV_X1 U11673 ( .A(n13757), .ZN(n9753) );
  NOR2_X1 U11674 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12105), .ZN(
        n12164) );
  INV_X1 U11675 ( .A(n9990), .ZN(n9989) );
  AND2_X1 U11676 ( .A1(n9991), .A2(n14098), .ZN(n9990) );
  INV_X1 U11677 ( .A(n14108), .ZN(n9991) );
  NOR2_X1 U11678 ( .A1(n9593), .A2(n14290), .ZN(n9953) );
  NOR2_X1 U11679 ( .A1(n11779), .A2(n11775), .ZN(n11805) );
  INV_X1 U11680 ( .A(n14159), .ZN(n9998) );
  INV_X1 U11681 ( .A(n11746), .ZN(n9781) );
  XNOR2_X1 U11682 ( .A(n13654), .B(n11683), .ZN(n13646) );
  NAND2_X1 U11683 ( .A1(n14573), .A2(n14562), .ZN(n9851) );
  NAND2_X1 U11684 ( .A1(n13933), .A2(n9934), .ZN(n9933) );
  INV_X1 U11685 ( .A(n14065), .ZN(n9934) );
  INV_X1 U11686 ( .A(n13927), .ZN(n13937) );
  NAND2_X1 U11687 ( .A1(n13977), .A2(n13949), .ZN(n13927) );
  INV_X1 U11688 ( .A(n13660), .ZN(n11681) );
  NAND2_X1 U11689 ( .A1(n11437), .A2(n19932), .ZN(n12757) );
  NOR2_X1 U11690 ( .A1(n12794), .A2(n9803), .ZN(n9802) );
  INV_X1 U11691 ( .A(n11621), .ZN(n11622) );
  OR2_X1 U11692 ( .A1(n12757), .A2(n15614), .ZN(n12145) );
  NAND2_X1 U11693 ( .A1(n12757), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12118) );
  OR2_X1 U11694 ( .A1(n11574), .A2(n11573), .ZN(n13089) );
  INV_X1 U11695 ( .A(n9936), .ZN(n13103) );
  OAI21_X1 U11696 ( .B1(n13134), .B2(n15781), .A(n20609), .ZN(n19930) );
  AND2_X1 U11697 ( .A1(n10732), .A2(n10722), .ZN(n10704) );
  NOR2_X1 U11698 ( .A1(n10889), .A2(n10888), .ZN(n10892) );
  INV_X1 U11699 ( .A(n10861), .ZN(n9835) );
  INV_X1 U11700 ( .A(n18632), .ZN(n9968) );
  NAND2_X1 U11701 ( .A1(n12959), .A2(n9834), .ZN(n9833) );
  NAND2_X1 U11702 ( .A1(n9828), .A2(n9827), .ZN(n10750) );
  NAND2_X1 U11703 ( .A1(n12521), .A2(n10728), .ZN(n9827) );
  NAND2_X1 U11704 ( .A1(n10727), .A2(n19028), .ZN(n9828) );
  NAND2_X1 U11705 ( .A1(n10007), .A2(n9626), .ZN(n13602) );
  NOR2_X1 U11706 ( .A1(n11236), .A2(n10598), .ZN(n11232) );
  NOR2_X1 U11707 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  INV_X1 U11708 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U11709 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9976) );
  NOR2_X1 U11710 ( .A1(n10056), .A2(n10055), .ZN(n10054) );
  INV_X1 U11711 ( .A(n10919), .ZN(n10055) );
  NAND2_X1 U11712 ( .A1(n10907), .A2(n9840), .ZN(n9839) );
  NOR2_X1 U11713 ( .A1(n14895), .A2(n9841), .ZN(n9840) );
  INV_X1 U11714 ( .A(n10870), .ZN(n9841) );
  NAND2_X1 U11715 ( .A1(n14794), .A2(n10060), .ZN(n10059) );
  INV_X1 U11716 ( .A(n14805), .ZN(n10060) );
  OR2_X1 U11717 ( .A1(n10885), .A2(n10884), .ZN(n10908) );
  NOR2_X1 U11718 ( .A1(n15118), .A2(n10994), .ZN(n10110) );
  OAI21_X1 U11719 ( .B1(n10839), .B2(n9891), .A(n9761), .ZN(n9764) );
  NOR2_X1 U11720 ( .A1(n9765), .A2(n9662), .ZN(n9761) );
  INV_X1 U11721 ( .A(n15281), .ZN(n9762) );
  INV_X1 U11722 ( .A(n9885), .ZN(n9765) );
  NAND2_X1 U11723 ( .A1(n10072), .A2(n10071), .ZN(n10070) );
  INV_X1 U11724 ( .A(n10073), .ZN(n10072) );
  NOR2_X1 U11725 ( .A1(n10075), .A2(n15147), .ZN(n10071) );
  NAND2_X1 U11726 ( .A1(n12565), .A2(n10074), .ZN(n10073) );
  INV_X1 U11727 ( .A(n14856), .ZN(n10074) );
  OR2_X1 U11728 ( .A1(n18635), .A2(n10865), .ZN(n10843) );
  OR2_X1 U11729 ( .A1(n18654), .A2(n10865), .ZN(n10848) );
  AND2_X1 U11730 ( .A1(n15048), .A2(n15162), .ZN(n15032) );
  NAND2_X1 U11731 ( .A1(n10767), .A2(n9629), .ZN(n9919) );
  OR2_X1 U11732 ( .A1(n10557), .A2(n10865), .ZN(n10556) );
  AND2_X1 U11733 ( .A1(n10526), .A2(n10525), .ZN(n10535) );
  NAND2_X1 U11734 ( .A1(n10718), .A2(n10865), .ZN(n10738) );
  NAND2_X1 U11735 ( .A1(n13397), .A2(n10427), .ZN(n10446) );
  OR2_X1 U11736 ( .A1(n10350), .A2(n10349), .ZN(n11055) );
  XNOR2_X1 U11737 ( .A(n10262), .B(n10263), .ZN(n10284) );
  OR2_X1 U11738 ( .A1(n10381), .A2(n10380), .ZN(n11032) );
  NAND2_X1 U11739 ( .A1(n10255), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10256) );
  AND2_X1 U11740 ( .A1(n19028), .A2(n19544), .ZN(n11007) );
  CLKBUF_X1 U11741 ( .A(n10971), .Z(n13248) );
  OR2_X1 U11742 ( .A1(n12413), .A2(n12203), .ZN(n12205) );
  AND2_X1 U11743 ( .A1(n12854), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12196) );
  OAI21_X1 U11744 ( .B1(n12195), .B2(n12209), .A(n12194), .ZN(n12221) );
  NAND2_X1 U11745 ( .A1(n10101), .A2(n12202), .ZN(n10320) );
  NAND2_X1 U11746 ( .A1(n10017), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10016) );
  NAND2_X1 U11747 ( .A1(n9770), .A2(n9768), .ZN(n10194) );
  NOR2_X1 U11748 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18549), .ZN(
        n13869) );
  OAI22_X1 U11749 ( .A1(n18535), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13860) );
  NAND3_X1 U11750 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18542), .ZN(n13755) );
  NOR2_X1 U11751 ( .A1(n13750), .A2(n13756), .ZN(n13826) );
  NOR2_X1 U11752 ( .A1(n13749), .A2(n16557), .ZN(n15436) );
  AOI21_X1 U11753 ( .B1(n16887), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(n9755), .ZN(n15439) );
  AND3_X1 U11754 ( .A1(n9754), .A2(n9753), .A3(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n9755) );
  AOI21_X1 U11755 ( .B1(n16635), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(n9715), .ZN(n15433) );
  NOR2_X1 U11756 ( .A1(n13827), .A2(n9716), .ZN(n9715) );
  NOR2_X1 U11757 ( .A1(n17219), .A2(n9858), .ZN(n9857) );
  NAND2_X1 U11758 ( .A1(n17244), .A2(n9620), .ZN(n16040) );
  NAND2_X1 U11759 ( .A1(n16015), .A2(n17483), .ZN(n16018) );
  OR2_X1 U11760 ( .A1(n17312), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10036) );
  NAND2_X1 U11761 ( .A1(n17503), .A2(n15496), .ZN(n15497) );
  INV_X1 U11762 ( .A(n17514), .ZN(n9758) );
  XNOR2_X1 U11763 ( .A(n15546), .B(n17092), .ZN(n15481) );
  OR2_X1 U11764 ( .A1(n18528), .A2(n13755), .ZN(n10126) );
  NOR2_X1 U11765 ( .A1(n9708), .A2(n9707), .ZN(n13823) );
  NAND2_X1 U11766 ( .A1(n20628), .A2(n13287), .ZN(n13304) );
  OR2_X1 U11767 ( .A1(n13300), .A2(n13299), .ZN(n19790) );
  OR2_X1 U11768 ( .A1(n14088), .A2(n14075), .ZN(n14077) );
  AND2_X1 U11769 ( .A1(n13915), .A2(n13914), .ZN(n14100) );
  NOR2_X1 U11770 ( .A1(n14113), .A2(n14100), .ZN(n14099) );
  NAND2_X1 U11771 ( .A1(n14200), .A2(n13889), .ZN(n14204) );
  OAI211_X1 U11772 ( .C1(n15680), .C2(n12065), .A(n11731), .B(n11730), .ZN(
        n13588) );
  INV_X1 U11773 ( .A(n10003), .ZN(n10000) );
  AOI21_X1 U11774 ( .B1(n13476), .B2(n11800), .A(n11680), .ZN(n13386) );
  XNOR2_X1 U11775 ( .A(n13283), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14302) );
  OR2_X1 U11776 ( .A1(n13282), .A2(n13281), .ZN(n13283) );
  AOI22_X1 U11777 ( .A1(n13980), .A2(n12096), .B1(n12095), .B2(n12094), .ZN(
        n13975) );
  AOI22_X1 U11778 ( .A1(n14328), .A2(n12096), .B1(n12039), .B2(n12038), .ZN(
        n14002) );
  AND2_X1 U11779 ( .A1(n12003), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12004) );
  NAND2_X1 U11780 ( .A1(n12004), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12040) );
  NOR2_X1 U11781 ( .A1(n14014), .A2(n9792), .ZN(n9791) );
  INV_X1 U11782 ( .A(n14028), .ZN(n9792) );
  NAND2_X1 U11783 ( .A1(n11960), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12002) );
  CLKBUF_X1 U11784 ( .A(n14037), .Z(n14038) );
  NOR2_X1 U11785 ( .A1(n11914), .A2(n14386), .ZN(n11915) );
  NAND2_X1 U11786 ( .A1(n11915), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11958) );
  CLKBUF_X1 U11787 ( .A(n14060), .Z(n14061) );
  OR2_X1 U11788 ( .A1(n11883), .A2(n11882), .ZN(n11885) );
  OR2_X1 U11789 ( .A1(n11885), .A2(n11884), .ZN(n11914) );
  NAND2_X1 U11790 ( .A1(n11853), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11883) );
  NAND2_X1 U11791 ( .A1(n11838), .A2(n11837), .ZN(n11839) );
  AND2_X1 U11792 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11837) );
  NOR2_X1 U11793 ( .A1(n11808), .A2(n15643), .ZN(n11838) );
  NAND2_X1 U11794 ( .A1(n14447), .A2(n14457), .ZN(n14446) );
  NAND2_X1 U11795 ( .A1(n11805), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U11796 ( .A1(n11776), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11779) );
  NOR2_X1 U11797 ( .A1(n11758), .A2(n11757), .ZN(n11776) );
  NAND2_X1 U11798 ( .A1(n11732), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11758) );
  INV_X1 U11799 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U11800 ( .A1(n9783), .A2(n11746), .ZN(n9780) );
  NOR2_X1 U11801 ( .A1(n11718), .A2(n19767), .ZN(n11732) );
  NAND2_X1 U11802 ( .A1(n11714), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11718) );
  CLKBUF_X1 U11803 ( .A(n13387), .Z(n13388) );
  NAND2_X1 U11804 ( .A1(n11674), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11684) );
  INV_X1 U11805 ( .A(n13361), .ZN(n11654) );
  INV_X1 U11806 ( .A(n11615), .ZN(n11638) );
  NAND2_X1 U11807 ( .A1(n11638), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11649) );
  NAND2_X1 U11808 ( .A1(n11620), .A2(n11619), .ZN(n9790) );
  OAI21_X1 U11809 ( .B1(n20009), .B2(n13655), .A(n12879), .ZN(n12943) );
  OAI21_X1 U11810 ( .B1(n14334), .B2(n9702), .A(n9616), .ZN(n9799) );
  INV_X1 U11811 ( .A(n14295), .ZN(n14296) );
  NAND2_X1 U11812 ( .A1(n9899), .A2(n14528), .ZN(n9898) );
  NOR2_X1 U11813 ( .A1(n14077), .A2(n9933), .ZN(n14041) );
  NOR2_X1 U11814 ( .A1(n14077), .A2(n14065), .ZN(n14064) );
  AND2_X1 U11815 ( .A1(n14531), .A2(n14530), .ZN(n14583) );
  OR2_X1 U11816 ( .A1(n9808), .A2(n9593), .ZN(n9807) );
  OR2_X1 U11817 ( .A1(n14127), .A2(n14111), .ZN(n14113) );
  INV_X1 U11818 ( .A(n14138), .ZN(n9928) );
  NAND2_X1 U11819 ( .A1(n14200), .A2(n9622), .ZN(n14148) );
  AND2_X1 U11820 ( .A1(n13726), .A2(n13725), .ZN(n14200) );
  AND2_X1 U11821 ( .A1(n13743), .A2(n13742), .ZN(n14202) );
  AND2_X1 U11822 ( .A1(n14280), .A2(n9655), .ZN(n9903) );
  NOR2_X1 U11823 ( .A1(n13597), .A2(n13596), .ZN(n13726) );
  NAND2_X1 U11824 ( .A1(n9908), .A2(n9907), .ZN(n13597) );
  INV_X1 U11825 ( .A(n13563), .ZN(n9907) );
  INV_X1 U11826 ( .A(n13562), .ZN(n9908) );
  INV_X1 U11827 ( .A(n15761), .ZN(n9909) );
  AND2_X1 U11828 ( .A1(n13442), .A2(n13441), .ZN(n13443) );
  INV_X1 U11829 ( .A(n9910), .ZN(n15760) );
  OR2_X1 U11830 ( .A1(n13347), .A2(n13346), .ZN(n13444) );
  NAND2_X1 U11831 ( .A1(n13169), .A2(n13168), .ZN(n13347) );
  NOR2_X1 U11832 ( .A1(n13084), .A2(n13083), .ZN(n13169) );
  NAND2_X1 U11833 ( .A1(n9922), .A2(n9921), .ZN(n13084) );
  INV_X1 U11834 ( .A(n12872), .ZN(n9921) );
  INV_X1 U11835 ( .A(n12873), .ZN(n9922) );
  NAND2_X1 U11836 ( .A1(n13047), .A2(n13645), .ZN(n13056) );
  AND2_X1 U11837 ( .A1(n15740), .A2(n19915), .ZN(n14660) );
  INV_X1 U11838 ( .A(n11437), .ZN(n12901) );
  INV_X1 U11839 ( .A(n12786), .ZN(n11428) );
  INV_X1 U11840 ( .A(n9816), .ZN(n19927) );
  AND2_X1 U11841 ( .A1(n12828), .A2(n12765), .ZN(n15585) );
  NOR2_X2 U11842 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20398) );
  AND2_X1 U11843 ( .A1(n19931), .A2(n19930), .ZN(n19974) );
  NAND2_X1 U11844 ( .A1(n11636), .A2(n11637), .ZN(n9982) );
  AOI21_X1 U11845 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20397), .A(n19986), 
        .ZN(n20476) );
  NAND2_X1 U11846 ( .A1(n15614), .A2(n19930), .ZN(n19986) );
  INV_X1 U11847 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15606) );
  AND2_X1 U11848 ( .A1(n10577), .A2(n10576), .ZN(n19726) );
  OR2_X1 U11849 ( .A1(n10575), .A2(n10574), .ZN(n10577) );
  NOR2_X1 U11850 ( .A1(n15820), .A2(n15819), .ZN(n15818) );
  NAND2_X1 U11851 ( .A1(n10854), .A2(n9630), .ZN(n10871) );
  NAND2_X1 U11852 ( .A1(n10854), .A2(n10855), .ZN(n10862) );
  NAND2_X1 U11853 ( .A1(n10805), .A2(n10803), .ZN(n10857) );
  NAND2_X1 U11854 ( .A1(n9836), .A2(n9695), .ZN(n10831) );
  NAND2_X1 U11855 ( .A1(n10836), .A2(n10791), .ZN(n10819) );
  NOR3_X1 U11856 ( .A1(n10782), .A2(n10780), .A3(n9833), .ZN(n10835) );
  OR2_X1 U11857 ( .A1(n12289), .A2(n12288), .ZN(n15870) );
  NAND2_X1 U11858 ( .A1(n15027), .A2(n10043), .ZN(n10042) );
  NOR2_X1 U11859 ( .A1(n13566), .A2(n13691), .ZN(n10043) );
  OR2_X1 U11860 ( .A1(n11135), .A2(n11134), .ZN(n13065) );
  INV_X1 U11861 ( .A(n12499), .ZN(n9744) );
  NOR2_X1 U11862 ( .A1(n9742), .A2(n9744), .ZN(n9741) );
  INV_X1 U11863 ( .A(n14729), .ZN(n9742) );
  NAND2_X1 U11864 ( .A1(n9747), .A2(n9752), .ZN(n9746) );
  OR2_X1 U11865 ( .A1(n14751), .A2(n14750), .ZN(n9752) );
  AND2_X1 U11866 ( .A1(n11201), .A2(n11200), .ZN(n14811) );
  AND2_X1 U11867 ( .A1(n13687), .A2(n14779), .ZN(n15871) );
  NAND2_X1 U11868 ( .A1(n12221), .A2(n12196), .ZN(n13421) );
  INV_X1 U11869 ( .A(n12519), .ZN(n14848) );
  OAI21_X1 U11870 ( .B1(n12518), .B2(n12517), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12519) );
  INV_X1 U11871 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14890) );
  INV_X1 U11872 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U11873 ( .A1(n11232), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11234) );
  NAND2_X1 U11874 ( .A1(n14780), .A2(n9677), .ZN(n14941) );
  INV_X1 U11875 ( .A(n14938), .ZN(n10049) );
  NOR2_X2 U11876 ( .A1(n14941), .A2(n12573), .ZN(n14769) );
  NAND2_X1 U11877 ( .A1(n14780), .A2(n9619), .ZN(n14983) );
  NAND2_X1 U11878 ( .A1(n14780), .A2(n9623), .ZN(n14939) );
  AND2_X1 U11879 ( .A1(n14780), .A2(n14781), .ZN(n14981) );
  AND2_X1 U11880 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10595) );
  NOR2_X1 U11881 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  INV_X1 U11882 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9950) );
  AND2_X1 U11883 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10593) );
  INV_X1 U11884 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13547) );
  AND2_X1 U11885 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11263) );
  INV_X1 U11886 ( .A(n10286), .ZN(n10278) );
  INV_X1 U11887 ( .A(n14880), .ZN(n9923) );
  INV_X1 U11888 ( .A(n10912), .ZN(n10910) );
  AND2_X1 U11889 ( .A1(n11198), .A2(n11197), .ZN(n14832) );
  NAND2_X1 U11890 ( .A1(n14994), .A2(n9633), .ZN(n14966) );
  NAND2_X1 U11891 ( .A1(n10096), .A2(n14958), .ZN(n10095) );
  INV_X1 U11892 ( .A(n15001), .ZN(n10096) );
  NOR2_X1 U11893 ( .A1(n15234), .A2(n15233), .ZN(n15235) );
  NAND2_X1 U11894 ( .A1(n15955), .A2(n13438), .ZN(n15234) );
  CLKBUF_X1 U11895 ( .A(n15032), .Z(n15033) );
  NOR2_X1 U11896 ( .A1(n10083), .A2(n10082), .ZN(n10081) );
  INV_X1 U11897 ( .A(n10079), .ZN(n10078) );
  INV_X1 U11898 ( .A(n10084), .ZN(n10083) );
  NOR2_X1 U11899 ( .A1(n15957), .A2(n15956), .ZN(n15955) );
  NAND2_X1 U11900 ( .A1(n13180), .A2(n13179), .ZN(n15957) );
  NAND2_X1 U11901 ( .A1(n10085), .A2(n10084), .ZN(n15258) );
  AND2_X2 U11902 ( .A1(n15979), .A2(n10066), .ZN(n13180) );
  AND2_X1 U11903 ( .A1(n10067), .A2(n9621), .ZN(n10066) );
  INV_X1 U11904 ( .A(n13150), .ZN(n10067) );
  NOR2_X1 U11905 ( .A1(n10069), .A2(n15303), .ZN(n10068) );
  INV_X1 U11906 ( .A(n12825), .ZN(n10069) );
  NAND2_X1 U11907 ( .A1(n15979), .A2(n9621), .ZN(n15283) );
  NOR2_X1 U11908 ( .A1(n15049), .A2(n15318), .ZN(n15293) );
  NAND2_X1 U11909 ( .A1(n15979), .A2(n12825), .ZN(n15304) );
  INV_X1 U11910 ( .A(n12962), .ZN(n10048) );
  NAND2_X1 U11911 ( .A1(n10768), .A2(n10767), .ZN(n9920) );
  XNOR2_X1 U11912 ( .A(n10557), .B(n10865), .ZN(n15058) );
  NAND2_X1 U11913 ( .A1(n10533), .A2(n10532), .ZN(n15057) );
  NAND2_X1 U11914 ( .A1(n10062), .A2(n10065), .ZN(n13426) );
  AND2_X1 U11915 ( .A1(n9912), .A2(n9683), .ZN(n9911) );
  NAND2_X1 U11916 ( .A1(n9915), .A2(n9846), .ZN(n13391) );
  AND2_X1 U11917 ( .A1(n13575), .A2(n13402), .ZN(n9846) );
  NOR2_X1 U11918 ( .A1(n11218), .A2(n13236), .ZN(n18973) );
  OAI22_X1 U11919 ( .A1(n10265), .A2(n10248), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10663), .ZN(n10251) );
  NOR2_X1 U11920 ( .A1(n19033), .A2(n18596), .ZN(n12710) );
  AOI21_X1 U11921 ( .B1(n10321), .B2(n12200), .A(n12199), .ZN(n12547) );
  CLKBUF_X1 U11922 ( .A(n10329), .Z(n10330) );
  OAI21_X1 U11923 ( .B1(n12219), .B2(n12726), .A(n12218), .ZN(n12843) );
  NOR2_X1 U11924 ( .A1(n12725), .A2(n12723), .ZN(n12219) );
  CLKBUF_X1 U11925 ( .A(n10581), .Z(n13216) );
  AND2_X1 U11926 ( .A1(n12212), .A2(n19278), .ZN(n19213) );
  AND2_X1 U11927 ( .A1(n19277), .A2(n19276), .ZN(n19238) );
  AND2_X1 U11928 ( .A1(n19139), .A2(n18992), .ZN(n19308) );
  AND2_X1 U11929 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19368) );
  AND2_X1 U11930 ( .A1(n19139), .A2(n19709), .ZN(n19375) );
  INV_X1 U11931 ( .A(n19485), .ZN(n19411) );
  INV_X1 U11932 ( .A(n19445), .ZN(n19450) );
  OAI21_X1 U11933 ( .B1(n9728), .B2(n9720), .A(n13211), .ZN(n9727) );
  OAI21_X1 U11934 ( .B1(n9723), .B2(n9721), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9722) );
  INV_X1 U11935 ( .A(n19022), .ZN(n19043) );
  INV_X1 U11936 ( .A(n19553), .ZN(n19046) );
  INV_X1 U11937 ( .A(n19041), .ZN(n19037) );
  INV_X1 U11938 ( .A(n19042), .ZN(n19039) );
  NOR2_X2 U11939 ( .A1(n14847), .A2(n15063), .ZN(n19042) );
  OR2_X1 U11940 ( .A1(n19277), .A2(n19715), .ZN(n19446) );
  OR2_X1 U11941 ( .A1(n19277), .A2(n19276), .ZN(n19485) );
  OR2_X1 U11942 ( .A1(n19139), .A2(n18992), .ZN(n19484) );
  INV_X1 U11943 ( .A(n19484), .ZN(n19548) );
  NOR2_X1 U11944 ( .A1(n17916), .A2(n17922), .ZN(n15516) );
  NAND2_X1 U11945 ( .A1(n16865), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n15378) );
  NAND2_X1 U11946 ( .A1(n16925), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n16902) );
  NOR2_X1 U11947 ( .A1(n18576), .A2(n17916), .ZN(n15362) );
  AND3_X1 U11948 ( .A1(n10038), .A2(n15429), .A3(n9653), .ZN(n15536) );
  AND2_X1 U11949 ( .A1(n15430), .A2(n15431), .ZN(n10038) );
  NOR2_X1 U11950 ( .A1(n13823), .A2(n17950), .ZN(n18379) );
  AOI221_X1 U11951 ( .B1(n18571), .B2(n18413), .C1(n17165), .C2(n18413), .A(
        n17164), .ZN(n17166) );
  NAND2_X1 U11952 ( .A1(n17244), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17218) );
  NOR2_X1 U11953 ( .A1(n17258), .A2(n17259), .ZN(n17244) );
  NOR2_X1 U11954 ( .A1(n17301), .A2(n17302), .ZN(n17281) );
  INV_X1 U11955 ( .A(n16337), .ZN(n17292) );
  NAND2_X1 U11956 ( .A1(n17321), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17301) );
  NOR2_X1 U11957 ( .A1(n17333), .A2(n17335), .ZN(n17321) );
  NAND2_X1 U11958 ( .A1(n17358), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17333) );
  NOR2_X1 U11959 ( .A1(n17397), .A2(n9872), .ZN(n9871) );
  AND2_X1 U11960 ( .A1(n9871), .A2(n17509), .ZN(n17415) );
  INV_X1 U11961 ( .A(n17481), .ZN(n17771) );
  NAND2_X1 U11962 ( .A1(n17509), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17473) );
  NOR2_X1 U11963 ( .A1(n17516), .A2(n17515), .ZN(n17509) );
  AND2_X1 U11964 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17535) );
  NOR2_X1 U11965 ( .A1(n17232), .A2(n15511), .ZN(n15616) );
  NAND2_X1 U11966 ( .A1(n15466), .A2(n15538), .ZN(n16072) );
  NOR2_X1 U11967 ( .A1(n17601), .A2(n17636), .ZN(n17264) );
  NOR2_X1 U11968 ( .A1(n17638), .A2(n17601), .ZN(n17255) );
  NOR2_X1 U11969 ( .A1(n17327), .A2(n15505), .ZN(n17275) );
  INV_X1 U11970 ( .A(n15504), .ZN(n15505) );
  NOR2_X1 U11971 ( .A1(n17712), .A2(n17718), .ZN(n17370) );
  NAND2_X1 U11972 ( .A1(n15563), .A2(n17470), .ZN(n17768) );
  NOR2_X1 U11973 ( .A1(n17425), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17404) );
  NOR2_X1 U11974 ( .A1(n17731), .A2(n17481), .ZN(n17396) );
  OR2_X1 U11975 ( .A1(n17480), .A2(n10035), .ZN(n17425) );
  OR2_X1 U11976 ( .A1(n10036), .A2(n10037), .ZN(n10035) );
  NAND2_X1 U11977 ( .A1(n17442), .A2(n17782), .ZN(n10037) );
  NAND2_X1 U11978 ( .A1(n18380), .A2(n18374), .ZN(n17780) );
  OR2_X1 U11979 ( .A1(n17480), .A2(n10036), .ZN(n17446) );
  NAND2_X1 U11980 ( .A1(n9756), .A2(n17811), .ZN(n17480) );
  INV_X1 U11981 ( .A(n9884), .ZN(n9756) );
  INV_X1 U11982 ( .A(n17703), .ZN(n17808) );
  XNOR2_X1 U11983 ( .A(n15497), .B(n10033), .ZN(n17489) );
  INV_X1 U11984 ( .A(n15498), .ZN(n10033) );
  NAND2_X1 U11985 ( .A1(n17489), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17488) );
  XNOR2_X1 U11986 ( .A(n15481), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17555) );
  NAND2_X1 U11987 ( .A1(n17555), .A2(n17554), .ZN(n17553) );
  NAND2_X1 U11988 ( .A1(n18576), .A2(n17703), .ZN(n17769) );
  XNOR2_X1 U11989 ( .A(n15536), .B(n15467), .ZN(n17563) );
  NAND2_X1 U11990 ( .A1(n18401), .A2(n13850), .ZN(n18370) );
  NOR2_X1 U11991 ( .A1(n18359), .A2(n15519), .ZN(n15513) );
  INV_X1 U11992 ( .A(n18370), .ZN(n18368) );
  NAND2_X1 U11993 ( .A1(n18588), .A2(n15517), .ZN(n18374) );
  NOR2_X1 U11994 ( .A1(n15530), .A2(n13877), .ZN(n18388) );
  INV_X1 U11995 ( .A(n18374), .ZN(n18404) );
  NAND2_X1 U11996 ( .A1(n15513), .A2(n18368), .ZN(n18400) );
  INV_X1 U11997 ( .A(n17102), .ZN(n17916) );
  INV_X1 U11998 ( .A(n16953), .ZN(n17950) );
  INV_X1 U11999 ( .A(n18561), .ZN(n18405) );
  NAND2_X1 U12000 ( .A1(n15516), .A2(n13848), .ZN(n18413) );
  NOR2_X1 U12001 ( .A1(n18428), .A2(n18415), .ZN(n18569) );
  NAND2_X1 U12002 ( .A1(n15611), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19741) );
  OR2_X1 U12003 ( .A1(n13300), .A2(n13292), .ZN(n19791) );
  NAND2_X1 U12004 ( .A1(n14302), .A2(n13308), .ZN(n19771) );
  INV_X1 U12005 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19781) );
  INV_X1 U12006 ( .A(n19771), .ZN(n19796) );
  AND2_X1 U12007 ( .A1(n13304), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19830) );
  INV_X1 U12008 ( .A(n19790), .ZN(n19834) );
  INV_X1 U12009 ( .A(n19791), .ZN(n19832) );
  AND2_X1 U12010 ( .A1(n13304), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19837) );
  INV_X1 U12011 ( .A(n19801), .ZN(n19777) );
  INV_X1 U12012 ( .A(n14196), .ZN(n19846) );
  NAND2_X1 U12013 ( .A1(n19850), .A2(n14209), .ZN(n14206) );
  AND2_X1 U12014 ( .A1(n12829), .A2(n12937), .ZN(n19850) );
  INV_X1 U12015 ( .A(n19846), .ZN(n14208) );
  INV_X1 U12016 ( .A(n14263), .ZN(n14257) );
  INV_X1 U12017 ( .A(n14272), .ZN(n14277) );
  NAND2_X1 U12018 ( .A1(n12172), .A2(n12171), .ZN(n14270) );
  OR2_X1 U12019 ( .A1(n14275), .A2(n13074), .ZN(n14272) );
  AND2_X1 U12020 ( .A1(n12797), .A2(n15603), .ZN(n19860) );
  OAI21_X1 U12021 ( .B1(n14421), .B2(n14291), .A(n9593), .ZN(n14382) );
  INV_X1 U12022 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20756) );
  NAND2_X1 U12023 ( .A1(n9995), .A2(n9992), .ZN(n14134) );
  INV_X1 U12024 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13433) );
  AND2_X2 U12025 ( .A1(n19748), .A2(n12940), .ZN(n15686) );
  INV_X1 U12026 ( .A(n15696), .ZN(n15681) );
  INV_X1 U12027 ( .A(n15686), .ZN(n14459) );
  NAND2_X2 U12028 ( .A1(n15597), .A2(n12937), .ZN(n19748) );
  NAND2_X1 U12029 ( .A1(n12934), .A2(n20398), .ZN(n19924) );
  XNOR2_X1 U12030 ( .A(n9812), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14561) );
  INV_X1 U12031 ( .A(n14326), .ZN(n9814) );
  NAND2_X1 U12032 ( .A1(n14327), .A2(n14573), .ZN(n9815) );
  NOR2_X1 U12033 ( .A1(n14294), .A2(n14585), .ZN(n14336) );
  OR2_X1 U12034 ( .A1(n14674), .A2(n14514), .ZN(n14508) );
  OR2_X1 U12035 ( .A1(n15730), .A2(n14657), .ZN(n14509) );
  AND2_X1 U12036 ( .A1(n9904), .A2(n9655), .ZN(n14281) );
  NAND2_X1 U12037 ( .A1(n9964), .A2(n15688), .ZN(n13709) );
  NAND2_X1 U12038 ( .A1(n9963), .A2(n13644), .ZN(n15691) );
  NOR2_X1 U12039 ( .A1(n15737), .A2(n13667), .ZN(n15771) );
  NAND2_X1 U12040 ( .A1(n9798), .A2(n13335), .ZN(n13481) );
  AND2_X1 U12041 ( .A1(n14679), .A2(n14715), .ZN(n13061) );
  INV_X1 U12042 ( .A(n15736), .ZN(n19915) );
  INV_X1 U12043 ( .A(n14704), .ZN(n19913) );
  INV_X1 U12044 ( .A(n11517), .ZN(n11461) );
  NAND2_X1 U12045 ( .A1(n9817), .A2(n19927), .ZN(n20323) );
  INV_X1 U12046 ( .A(n12789), .ZN(n12794) );
  INV_X1 U12047 ( .A(n20041), .ZN(n20012) );
  OAI22_X1 U12048 ( .A1(n20019), .A2(n20018), .B1(n20158), .B2(n20281), .ZN(
        n20043) );
  OAI221_X1 U12049 ( .B1(n20117), .B2(n20357), .C1(n20117), .C2(n20098), .A(
        n20435), .ZN(n20119) );
  OAI211_X1 U12050 ( .C1(n10124), .C2(n20357), .A(n20278), .B(n20226), .ZN(
        n20242) );
  AND2_X1 U12051 ( .A1(n20199), .A2(n20326), .ZN(n20644) );
  OAI211_X1 U12052 ( .C1(n20390), .C2(n20357), .A(n20435), .B(n20356), .ZN(
        n20392) );
  OAI211_X1 U12053 ( .C1(n20457), .C2(n20436), .A(n20435), .B(n20434), .ZN(
        n20460) );
  INV_X1 U12054 ( .A(n20271), .ZN(n20474) );
  INV_X1 U12055 ( .A(n20286), .ZN(n20484) );
  INV_X1 U12056 ( .A(n20293), .ZN(n20496) );
  INV_X1 U12057 ( .A(n20297), .ZN(n20641) );
  INV_X1 U12058 ( .A(n20380), .ZN(n20504) );
  INV_X1 U12059 ( .A(n20304), .ZN(n20510) );
  NAND2_X1 U12060 ( .A1(n20426), .A2(n20425), .ZN(n20526) );
  INV_X1 U12061 ( .A(n20309), .ZN(n20520) );
  NAND2_X1 U12062 ( .A1(n12936), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20609) );
  INV_X1 U12063 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20357) );
  OR2_X1 U12064 ( .A1(n13272), .A2(n12550), .ZN(n12580) );
  NOR2_X1 U12065 ( .A1(n12585), .A2(n16003), .ZN(n18598) );
  AND2_X1 U12066 ( .A1(n9958), .A2(n9969), .ZN(n9956) );
  AND2_X1 U12067 ( .A1(n10875), .A2(n10900), .ZN(n15826) );
  NAND2_X1 U12068 ( .A1(n18764), .A2(n14919), .ZN(n9977) );
  NOR2_X1 U12069 ( .A1(n14926), .A2(n15851), .ZN(n9979) );
  NOR2_X1 U12070 ( .A1(n15571), .A2(n18676), .ZN(n12571) );
  NOR2_X1 U12071 ( .A1(n12571), .A2(n14926), .ZN(n12570) );
  AND2_X1 U12072 ( .A1(n9970), .A2(n9969), .ZN(n12561) );
  AND2_X1 U12073 ( .A1(n9971), .A2(n9969), .ZN(n18623) );
  AND2_X1 U12074 ( .A1(n12595), .A2(n11281), .ZN(n18775) );
  NOR2_X1 U12075 ( .A1(n18676), .A2(n18641), .ZN(n18631) );
  AOI21_X1 U12076 ( .B1(n18651), .B2(n18661), .A(n18676), .ZN(n18650) );
  NOR2_X1 U12077 ( .A1(n18642), .A2(n18650), .ZN(n18641) );
  INV_X1 U12078 ( .A(n18825), .ZN(n18807) );
  AND2_X1 U12079 ( .A1(n12595), .A2(n11277), .ZN(n18831) );
  AND2_X1 U12080 ( .A1(n14747), .A2(n14743), .ZN(n10920) );
  NOR2_X1 U12081 ( .A1(n13375), .A2(n12228), .ZN(n18839) );
  OR2_X1 U12082 ( .A1(n11165), .A2(n11164), .ZN(n13377) );
  OR2_X1 U12083 ( .A1(n11120), .A2(n11119), .ZN(n12951) );
  OR2_X1 U12084 ( .A1(n11106), .A2(n11105), .ZN(n12948) );
  INV_X1 U12085 ( .A(n19709), .ZN(n18992) );
  INV_X1 U12086 ( .A(n18848), .ZN(n18844) );
  INV_X1 U12087 ( .A(n15786), .ZN(n18853) );
  NOR2_X1 U12088 ( .A1(n14765), .A2(n14764), .ZN(n14763) );
  AND2_X1 U12089 ( .A1(n10023), .A2(n10022), .ZN(n14765) );
  INV_X1 U12090 ( .A(n10023), .ZN(n14842) );
  AND2_X1 U12091 ( .A1(n12520), .A2(n14847), .ZN(n18858) );
  AND2_X1 U12092 ( .A1(n12520), .A2(n14848), .ZN(n18859) );
  INV_X1 U12093 ( .A(n14859), .ZN(n18857) );
  NOR2_X1 U12094 ( .A1(n12921), .A2(n10063), .ZN(n13624) );
  NAND2_X1 U12095 ( .A1(n10065), .A2(n10064), .ZN(n10063) );
  AND2_X1 U12096 ( .A1(n18861), .A2(n18862), .ZN(n18890) );
  INV_X1 U12097 ( .A(n18862), .ZN(n18852) );
  NAND2_X1 U12098 ( .A1(n12607), .A2(n12506), .ZN(n12507) );
  INV_X1 U12099 ( .A(n13439), .ZN(n18883) );
  INV_X1 U12100 ( .A(n19715), .ZN(n19276) );
  INV_X1 U12101 ( .A(n18861), .ZN(n18884) );
  NOR2_X1 U12102 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12610), .ZN(n12636) );
  AND2_X1 U12103 ( .A1(n12600), .A2(n19623), .ZN(n18894) );
  OR2_X1 U12104 ( .A1(n18894), .A2(n18924), .ZN(n18911) );
  INV_X2 U12105 ( .A(n18911), .ZN(n18923) );
  INV_X2 U12106 ( .A(n12666), .ZN(n18958) );
  NAND2_X1 U12107 ( .A1(n9947), .A2(n10599), .ZN(n9943) );
  AND2_X1 U12108 ( .A1(n13567), .A2(n13381), .ZN(n18692) );
  INV_X1 U12109 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15914) );
  INV_X1 U12110 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15954) );
  INV_X1 U12111 ( .A(n15944), .ZN(n15922) );
  INV_X1 U12112 ( .A(n15953), .ZN(n15915) );
  XNOR2_X1 U12113 ( .A(n10691), .B(n10690), .ZN(n15862) );
  NOR2_X1 U12114 ( .A1(n9637), .A2(n10968), .ZN(n10691) );
  OAI21_X1 U12115 ( .B1(n15786), .B2(n18986), .A(n10114), .ZN(n10040) );
  NAND2_X1 U12116 ( .A1(n9924), .A2(n9925), .ZN(n14882) );
  OR2_X1 U12117 ( .A1(n11211), .A2(n14786), .ZN(n15803) );
  NAND2_X1 U12118 ( .A1(n9763), .A2(n9885), .ZN(n14924) );
  NAND2_X1 U12119 ( .A1(n9887), .A2(n10853), .ZN(n14937) );
  NAND2_X1 U12120 ( .A1(n9892), .A2(n9888), .ZN(n9887) );
  AOI21_X1 U12121 ( .B1(n10092), .B2(n10090), .A(n10088), .ZN(n10087) );
  NOR2_X1 U12122 ( .A1(n14855), .A2(n14856), .ZN(n15174) );
  AND2_X1 U12123 ( .A1(n15264), .A2(n15897), .ZN(n15905) );
  AND2_X1 U12124 ( .A1(n10098), .A2(n9650), .ZN(n15295) );
  NAND2_X1 U12125 ( .A1(n10098), .A2(n10779), .ZN(n15317) );
  NOR2_X1 U12126 ( .A1(n10992), .A2(n13701), .ZN(n15987) );
  NAND2_X1 U12127 ( .A1(n10107), .A2(n10449), .ZN(n13615) );
  NOR2_X1 U12128 ( .A1(n12921), .A2(n11053), .ZN(n13181) );
  CLKBUF_X1 U12129 ( .A(n13397), .Z(n13398) );
  OR2_X1 U12130 ( .A1(n11218), .A2(n10970), .ZN(n15330) );
  INV_X1 U12131 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20684) );
  NAND2_X1 U12132 ( .A1(n13237), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15995) );
  INV_X1 U12133 ( .A(n19150), .ZN(n19167) );
  NOR2_X1 U12134 ( .A1(n19140), .A2(n19445), .ZN(n19202) );
  NAND2_X1 U12135 ( .A1(n19411), .A2(n19308), .ZN(n19324) );
  INV_X1 U12136 ( .A(n19324), .ZN(n19333) );
  NOR2_X1 U12137 ( .A1(n19446), .A2(n19309), .ZN(n19363) );
  INV_X1 U12138 ( .A(n19565), .ZN(n19503) );
  AND2_X1 U12139 ( .A1(n19006), .A2(n19043), .ZN(n19502) );
  AND2_X1 U12140 ( .A1(n19010), .A2(n19043), .ZN(n19507) );
  AND2_X1 U12141 ( .A1(n19016), .A2(n19043), .ZN(n19513) );
  OAI22_X1 U12142 ( .A1(n19021), .A2(n19039), .B1(n19020), .B2(n19037), .ZN(
        n19518) );
  AND2_X1 U12143 ( .A1(n19028), .A2(n19043), .ZN(n19522) );
  NOR2_X1 U12144 ( .A1(n19446), .A2(n19445), .ZN(n19523) );
  AND2_X1 U12145 ( .A1(n19033), .A2(n19043), .ZN(n19528) );
  OAI21_X1 U12146 ( .B1(n19498), .B2(n19497), .A(n19496), .ZN(n19535) );
  AND2_X1 U12147 ( .A1(n19044), .A2(n19043), .ZN(n19533) );
  INV_X1 U12148 ( .A(n19396), .ZN(n19584) );
  INV_X1 U12149 ( .A(n19518), .ZN(n19587) );
  NOR2_X2 U12150 ( .A1(n19446), .A2(n19484), .ZN(n19599) );
  INV_X1 U12151 ( .A(n19541), .ZN(n19609) );
  NOR2_X2 U12152 ( .A1(n19485), .A2(n19484), .ZN(n19610) );
  INV_X1 U12153 ( .A(n19534), .ZN(n19615) );
  NAND2_X1 U12154 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19617) );
  OR2_X1 U12155 ( .A1(n11283), .A2(n13409), .ZN(n16003) );
  CLKBUF_X1 U12156 ( .A(n11284), .Z(n18819) );
  AOI21_X1 U12157 ( .B1(n13848), .B2(n13847), .A(n13854), .ZN(n16176) );
  NAND2_X1 U12158 ( .A1(n18569), .A2(n16171), .ZN(n17164) );
  AOI21_X1 U12159 ( .B1(n18401), .B2(n18400), .A(n17164), .ZN(n18573) );
  NAND2_X1 U12160 ( .A1(n18569), .A2(n16007), .ZN(n16177) );
  OAI22_X1 U12161 ( .A1(n18560), .A2(n18405), .B1(n18562), .B2(n17769), .ZN(
        n16007) );
  INV_X1 U12162 ( .A(n9875), .ZN(n16228) );
  AOI21_X1 U12163 ( .B1(n16272), .B2(n9868), .A(n16529), .ZN(n16251) );
  NOR2_X1 U12164 ( .A1(n16272), .A2(n16529), .ZN(n16265) );
  NOR2_X1 U12165 ( .A1(n16265), .A2(n17248), .ZN(n16264) );
  INV_X1 U12166 ( .A(n16561), .ZN(n16517) );
  NOR2_X1 U12167 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16322), .ZN(n16306) );
  AND2_X1 U12168 ( .A1(n9861), .A2(n16478), .ZN(n16296) );
  NOR2_X1 U12169 ( .A1(n16319), .A2(n16529), .ZN(n16305) );
  NAND2_X1 U12170 ( .A1(n9861), .A2(n9860), .ZN(n16304) );
  NAND2_X1 U12171 ( .A1(n16529), .A2(n9862), .ZN(n9860) );
  NOR2_X1 U12172 ( .A1(n9865), .A2(n9864), .ZN(n16319) );
  INV_X1 U12173 ( .A(n16317), .ZN(n9864) );
  NOR2_X1 U12174 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16432), .ZN(n16415) );
  NOR2_X1 U12175 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16453), .ZN(n16445) );
  NAND2_X1 U12176 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18435), .ZN(n16531) );
  INV_X1 U12177 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16508) );
  INV_X1 U12178 ( .A(n16549), .ZN(n16564) );
  NOR2_X1 U12179 ( .A1(n18414), .A2(n16197), .ZN(n16561) );
  NOR2_X1 U12180 ( .A1(n16927), .A2(n9709), .ZN(n16693) );
  INV_X1 U12181 ( .A(n16708), .ZN(n9719) );
  AND2_X1 U12182 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16712), .ZN(n16707) );
  NOR2_X1 U12183 ( .A1(n16725), .A2(n16680), .ZN(n16708) );
  AND2_X1 U12184 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16708), .ZN(n16712) );
  NAND2_X1 U12185 ( .A1(n16738), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n16725) );
  NOR2_X1 U12186 ( .A1(n16736), .A2(n17959), .ZN(n16738) );
  NOR2_X1 U12187 ( .A1(n16750), .A2(n16792), .ZN(n16780) );
  NOR2_X1 U12188 ( .A1(n16807), .A2(n16821), .ZN(n16793) );
  NAND2_X1 U12189 ( .A1(n16822), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n16821) );
  INV_X1 U12190 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16835) );
  NOR2_X1 U12191 ( .A1(n16462), .A2(n16902), .ZN(n16884) );
  NAND2_X1 U12192 ( .A1(n16926), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n16922) );
  NOR2_X1 U12193 ( .A1(n16922), .A2(n16486), .ZN(n16925) );
  NOR2_X2 U12194 ( .A1(n13784), .A2(n13783), .ZN(n17036) );
  NOR2_X1 U12195 ( .A1(n16930), .A2(n16508), .ZN(n16926) );
  NAND3_X1 U12196 ( .A1(n15362), .A2(n18569), .A3(n15633), .ZN(n16948) );
  NAND2_X1 U12197 ( .A1(n16962), .A2(n17086), .ZN(n16960) );
  AND2_X1 U12198 ( .A1(n16974), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n16963) );
  NAND2_X1 U12199 ( .A1(n16963), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n16962) );
  INV_X1 U12200 ( .A(n16963), .ZN(n16969) );
  NOR2_X1 U12201 ( .A1(n17109), .A2(n16978), .ZN(n16974) );
  NAND2_X1 U12202 ( .A1(n16982), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n16978) );
  NOR2_X1 U12203 ( .A1(n16987), .A2(n17113), .ZN(n16982) );
  NOR2_X1 U12204 ( .A1(n16992), .A2(n17959), .ZN(n16988) );
  NAND2_X1 U12205 ( .A1(n16988), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n16987) );
  NOR3_X1 U12206 ( .A1(n17959), .A2(n17028), .A3(n17169), .ZN(n17020) );
  NAND2_X1 U12207 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17032), .ZN(n17028) );
  NOR2_X1 U12208 ( .A1(n17214), .A2(n17039), .ZN(n17032) );
  NOR2_X1 U12209 ( .A1(n17096), .A2(n9704), .ZN(n17062) );
  INV_X1 U12210 ( .A(n17067), .ZN(n9705) );
  NOR2_X1 U12211 ( .A1(n15417), .A2(n15416), .ZN(n17082) );
  NAND2_X1 U12212 ( .A1(n18379), .A2(n16950), .ZN(n17088) );
  INV_X1 U12213 ( .A(n17094), .ZN(n17091) );
  NAND2_X1 U12214 ( .A1(n16950), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17096) );
  NOR2_X1 U12215 ( .A1(n18379), .A2(n17086), .ZN(n17094) );
  INV_X1 U12216 ( .A(n17088), .ZN(n17093) );
  NOR2_X1 U12217 ( .A1(n17922), .A2(n17196), .ZN(n17179) );
  INV_X1 U12218 ( .A(n17213), .ZN(n17205) );
  INV_X1 U12219 ( .A(n17179), .ZN(n17213) );
  INV_X1 U12220 ( .A(n17710), .ZN(n17636) );
  AND3_X1 U12221 ( .A1(n9871), .A2(n9647), .A3(n9869), .ZN(n17358) );
  AND2_X1 U12222 ( .A1(n17509), .A2(n9870), .ZN(n9869) );
  INV_X1 U12223 ( .A(n17376), .ZN(n9870) );
  NOR2_X1 U12224 ( .A1(n17469), .A2(n17689), .ZN(n17382) );
  NAND2_X1 U12225 ( .A1(n17370), .A2(n17768), .ZN(n17638) );
  NOR2_X1 U12226 ( .A1(n17492), .A2(n17475), .ZN(n17477) );
  INV_X1 U12227 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17475) );
  INV_X1 U12228 ( .A(n17421), .ZN(n17485) );
  INV_X1 U12229 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17492) );
  NAND2_X1 U12230 ( .A1(n18264), .A2(n18118), .ZN(n17958) );
  INV_X1 U12231 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17560) );
  INV_X1 U12232 ( .A(n17567), .ZN(n17557) );
  INV_X1 U12233 ( .A(n17958), .ZN(n18299) );
  NAND2_X1 U12234 ( .A1(n17573), .A2(n17534), .ZN(n17568) );
  NAND2_X1 U12235 ( .A1(n17359), .A2(n9591), .ZN(n17567) );
  OAI21_X1 U12236 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18568), .A(n16177), 
        .ZN(n17573) );
  INV_X1 U12237 ( .A(n17565), .ZN(n17578) );
  NAND2_X1 U12238 ( .A1(n17249), .A2(n15510), .ZN(n16066) );
  INV_X1 U12239 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18415) );
  INV_X1 U12240 ( .A(n9883), .ZN(n17361) );
  INV_X1 U12241 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17704) );
  NOR2_X1 U12242 ( .A1(n17780), .A2(n18378), .ZN(n17703) );
  INV_X1 U12243 ( .A(n17814), .ZN(n17788) );
  NAND2_X1 U12244 ( .A1(n17513), .A2(n15494), .ZN(n17504) );
  NOR2_X1 U12245 ( .A1(n18405), .A2(n17886), .ZN(n17834) );
  NAND2_X1 U12246 ( .A1(n17542), .A2(n15486), .ZN(n17526) );
  INV_X1 U12247 ( .A(n17880), .ZN(n17888) );
  NOR2_X1 U12248 ( .A1(n17769), .A2(n17886), .ZN(n17885) );
  NOR2_X2 U12249 ( .A1(n15513), .A2(n18370), .ZN(n18380) );
  INV_X1 U12250 ( .A(n17885), .ZN(n17900) );
  INV_X1 U12251 ( .A(n17886), .ZN(n17892) );
  INV_X1 U12252 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18390) );
  INV_X1 U12253 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18399) );
  INV_X2 U12254 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18542) );
  AND2_X2 U12255 ( .A1(n12183), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19925)
         );
  XNOR2_X1 U12257 ( .A(n9816), .B(n20194), .ZN(n13152) );
  NAND2_X1 U12258 ( .A1(n12535), .A2(n18848), .ZN(n12539) );
  OAI21_X1 U12259 ( .B1(n14871), .B2(n18843), .A(n12536), .ZN(n12537) );
  AOI21_X1 U12260 ( .B1(n14873), .B2(n15939), .A(n14872), .ZN(n14874) );
  OAI21_X1 U12261 ( .B1(n14875), .B2(n15309), .A(n9663), .ZN(P2_U3016) );
  AND2_X1 U12262 ( .A1(n9665), .A2(n10057), .ZN(n9935) );
  OR2_X1 U12263 ( .A1(n15135), .A2(n15309), .ZN(n9819) );
  INV_X1 U12264 ( .A(n9873), .ZN(n16215) );
  INV_X1 U12265 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16540) );
  NOR2_X1 U12266 ( .A1(n9712), .A2(n9711), .ZN(n9710) );
  NAND2_X1 U12267 ( .A1(n10029), .A2(n9615), .ZN(P3_U2799) );
  NAND2_X1 U12268 ( .A1(n16061), .A2(n17484), .ZN(n10029) );
  INV_X2 U12269 ( .A(n11226), .ZN(n18676) );
  AND2_X2 U12270 ( .A1(n14994), .A2(n9614), .ZN(n9611) );
  CLKBUF_X3 U12271 ( .A(n13826), .Z(n16870) );
  AND2_X1 U12272 ( .A1(n15297), .A2(n9650), .ZN(n9613) );
  NAND2_X1 U12273 ( .A1(n9986), .A2(n9990), .ZN(n14084) );
  AND2_X2 U12274 ( .A1(n10552), .A2(n10551), .ZN(n10865) );
  AND2_X1 U12275 ( .A1(n9634), .A2(n9825), .ZN(n9614) );
  AND2_X2 U12276 ( .A1(n10248), .A2(n10243), .ZN(n10663) );
  AND3_X1 U12277 ( .A1(n11024), .A2(n12418), .A3(n19044), .ZN(n11054) );
  INV_X1 U12278 ( .A(n13734), .ZN(n9995) );
  INV_X1 U12279 ( .A(n9593), .ZN(n9954) );
  NAND2_X1 U12280 ( .A1(n9948), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11257) );
  NAND2_X1 U12281 ( .A1(n14027), .A2(n14028), .ZN(n14013) );
  NAND2_X1 U12282 ( .A1(n9995), .A2(n9996), .ZN(n14158) );
  INV_X1 U12283 ( .A(n11629), .ZN(n9941) );
  NOR2_X1 U12284 ( .A1(n14107), .A2(n9672), .ZN(n14072) );
  AND2_X1 U12285 ( .A1(n11313), .A2(n11315), .ZN(n11468) );
  AND3_X1 U12286 ( .A1(n16023), .A2(n9680), .A3(n10028), .ZN(n9615) );
  INV_X1 U12287 ( .A(n14734), .ZN(n9745) );
  INV_X1 U12288 ( .A(n16695), .ZN(n9709) );
  NAND2_X1 U12289 ( .A1(n14994), .A2(n9701), .ZN(n14909) );
  OR2_X1 U12290 ( .A1(n9954), .A2(n9700), .ZN(n9616) );
  AND2_X1 U12291 ( .A1(n10065), .A2(n9661), .ZN(n9617) );
  AND2_X1 U12292 ( .A1(n10228), .A2(n19023), .ZN(n9618) );
  AND2_X2 U12293 ( .A1(n11313), .A2(n13115), .ZN(n11584) );
  OR2_X1 U12294 ( .A1(n9938), .A2(n11609), .ZN(n10121) );
  NAND2_X1 U12295 ( .A1(n9972), .A2(n9974), .ZN(n11245) );
  AND2_X1 U12296 ( .A1(n14980), .A2(n14781), .ZN(n9619) );
  AND2_X1 U12297 ( .A1(n9857), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9620) );
  AND2_X1 U12298 ( .A1(n10068), .A2(n15284), .ZN(n9621) );
  NAND2_X1 U12299 ( .A1(n13687), .A2(n9690), .ZN(n14771) );
  AND2_X1 U12300 ( .A1(n9929), .A2(n14149), .ZN(n9622) );
  AND2_X1 U12301 ( .A1(n9619), .A2(n10050), .ZN(n9623) );
  OR3_X1 U12302 ( .A1(n13567), .A2(n10044), .A3(n13566), .ZN(n9624) );
  AND2_X1 U12303 ( .A1(n12225), .A2(n10128), .ZN(n9625) );
  AND2_X1 U12304 ( .A1(n10008), .A2(n12253), .ZN(n9626) );
  NAND2_X1 U12305 ( .A1(n15296), .A2(n15294), .ZN(n9627) );
  AND2_X1 U12306 ( .A1(n9620), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9628) );
  AND2_X1 U12307 ( .A1(n10100), .A2(n10099), .ZN(n9629) );
  NAND2_X1 U12308 ( .A1(n12856), .A2(n12858), .ZN(n12857) );
  AND2_X1 U12309 ( .A1(n10855), .A2(n9835), .ZN(n9630) );
  AND2_X1 U12310 ( .A1(n9630), .A2(n15853), .ZN(n9631) );
  AND4_X1 U12311 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n9632) );
  AND2_X1 U12312 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n9633) );
  AND2_X1 U12313 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n9633), .ZN(
        n9634) );
  AND2_X1 U12314 ( .A1(n10110), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9635) );
  CLKBUF_X3 U12315 ( .A(n11351), .Z(n12070) );
  OR2_X1 U12316 ( .A1(n14825), .A2(n14811), .ZN(n9636) );
  OR2_X1 U12317 ( .A1(n14760), .A2(n10052), .ZN(n9637) );
  AND2_X1 U12318 ( .A1(n10208), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10383) );
  OR2_X1 U12319 ( .A1(n13749), .A2(n13756), .ZN(n9639) );
  OR3_X1 U12320 ( .A1(n9636), .A2(n10059), .A3(n10058), .ZN(n9640) );
  OR2_X1 U12321 ( .A1(n11234), .A2(n9983), .ZN(n9641) );
  AND2_X1 U12322 ( .A1(n14994), .A2(n9634), .ZN(n9642) );
  OR2_X1 U12323 ( .A1(n14844), .A2(n14843), .ZN(n10023) );
  AND2_X1 U12324 ( .A1(n9995), .A2(n9994), .ZN(n9643) );
  OR2_X1 U12325 ( .A1(n18371), .A2(n13749), .ZN(n9644) );
  NAND2_X1 U12326 ( .A1(n14994), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14978) );
  NAND2_X1 U12327 ( .A1(n10131), .A2(n10132), .ZN(n11438) );
  INV_X1 U12328 ( .A(n14209), .ZN(n9938) );
  OR2_X1 U12329 ( .A1(n14855), .A2(n10070), .ZN(n9645) );
  NOR2_X1 U12330 ( .A1(n14060), .A2(n14062), .ZN(n14050) );
  NOR2_X1 U12331 ( .A1(n13734), .A2(n14199), .ZN(n14157) );
  NOR2_X1 U12332 ( .A1(n14107), .A2(n14108), .ZN(n14097) );
  NAND2_X1 U12333 ( .A1(n14730), .A2(n14729), .ZN(n14731) );
  AND4_X1 U12334 ( .A1(n11320), .A2(n11319), .A3(n11318), .A4(n11317), .ZN(
        n9646) );
  AND2_X1 U12335 ( .A1(n17413), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9647) );
  AND2_X1 U12336 ( .A1(n9910), .A2(n9909), .ZN(n9648) );
  INV_X1 U12337 ( .A(n19016), .ZN(n10238) );
  AOI21_X1 U12338 ( .B1(n15040), .B2(n15038), .A(n14955), .ZN(n15025) );
  OR3_X1 U12339 ( .A1(n10782), .A2(n10780), .A3(n9831), .ZN(n9649) );
  AND2_X1 U12340 ( .A1(n10097), .A2(n10779), .ZN(n9650) );
  INV_X1 U12341 ( .A(n10102), .ZN(n15930) );
  XOR2_X1 U12342 ( .A(n10901), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(
        n9651) );
  AND2_X1 U12343 ( .A1(n11314), .A2(n11315), .ZN(n12072) );
  NAND2_X2 U12344 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18371) );
  INV_X1 U12345 ( .A(n18371), .ZN(n9754) );
  NOR2_X1 U12346 ( .A1(n13764), .A2(n13763), .ZN(n15359) );
  INV_X1 U12347 ( .A(n15359), .ZN(n17938) );
  OR2_X1 U12348 ( .A1(n10782), .A2(n10780), .ZN(n9652) );
  AND4_X1 U12349 ( .A1(n15428), .A2(n15427), .A3(n15426), .A4(n15425), .ZN(
        n9653) );
  AND2_X1 U12350 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n9654) );
  AND2_X1 U12351 ( .A1(n10104), .A2(n15931), .ZN(n10103) );
  NAND2_X1 U12352 ( .A1(n13707), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9655) );
  OR2_X1 U12353 ( .A1(n14077), .A2(n9931), .ZN(n9656) );
  NAND2_X1 U12354 ( .A1(n11372), .A2(n10130), .ZN(n19949) );
  OR2_X1 U12355 ( .A1(n13051), .A2(n11550), .ZN(n9657) );
  NOR2_X1 U12356 ( .A1(n10853), .A2(n9889), .ZN(n9658) );
  NAND2_X1 U12358 ( .A1(n12221), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9659) );
  OR2_X1 U12359 ( .A1(n11628), .A2(n9941), .ZN(n9660) );
  AND2_X1 U12360 ( .A1(n10064), .A2(n13625), .ZN(n9661) );
  INV_X1 U12361 ( .A(n9836), .ZN(n10827) );
  NOR2_X1 U12362 ( .A1(n10812), .A2(n10796), .ZN(n9836) );
  BUF_X1 U12363 ( .A(n10284), .Z(n10308) );
  NAND2_X1 U12364 ( .A1(n9774), .A2(n9773), .ZN(n15279) );
  AND2_X1 U12365 ( .A1(n9890), .A2(n9762), .ZN(n9662) );
  AND2_X1 U12366 ( .A1(n11220), .A2(n9935), .ZN(n9663) );
  AND2_X1 U12367 ( .A1(n13482), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9664) );
  INV_X1 U12368 ( .A(n9891), .ZN(n9890) );
  NAND2_X1 U12369 ( .A1(n10840), .A2(n14935), .ZN(n9891) );
  NAND2_X1 U12370 ( .A1(n15258), .A2(n15259), .ZN(n15257) );
  OR2_X1 U12371 ( .A1(n11275), .A2(n18986), .ZN(n9665) );
  INV_X1 U12372 ( .A(n9783), .ZN(n9782) );
  AND3_X1 U12373 ( .A1(n13812), .A2(n13810), .A3(n13808), .ZN(n9666) );
  INV_X1 U12374 ( .A(n10027), .ZN(n17266) );
  NAND2_X1 U12375 ( .A1(n11613), .A2(n11556), .ZN(n11636) );
  OR3_X1 U12376 ( .A1(n14294), .A2(n9898), .A3(n9900), .ZN(n9667) );
  AND2_X1 U12377 ( .A1(n10046), .A2(n10048), .ZN(n9668) );
  NOR2_X1 U12378 ( .A1(n15818), .A2(n18764), .ZN(n9669) );
  INV_X1 U12379 ( .A(n10555), .ZN(n10106) );
  AND2_X1 U12380 ( .A1(n10227), .A2(n19010), .ZN(n9670) );
  AND2_X1 U12381 ( .A1(n14949), .A2(n9890), .ZN(n9671) );
  INV_X1 U12382 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U12383 ( .A1(n14122), .A2(n14124), .ZN(n14107) );
  NAND2_X1 U12384 ( .A1(n9794), .A2(n11653), .ZN(n13191) );
  NOR2_X1 U12385 ( .A1(n11252), .A2(n18685), .ZN(n11248) );
  INV_X1 U12386 ( .A(n9734), .ZN(n13687) );
  NOR2_X1 U12387 ( .A1(n11255), .A2(n15914), .ZN(n11253) );
  NOR2_X1 U12388 ( .A1(n11259), .A2(n15954), .ZN(n11260) );
  NOR2_X1 U12389 ( .A1(n11252), .A2(n9976), .ZN(n11249) );
  NOR2_X1 U12390 ( .A1(n11256), .A2(n9951), .ZN(n11254) );
  NAND2_X1 U12391 ( .A1(n13687), .A2(n10025), .ZN(n14772) );
  OR2_X1 U12392 ( .A1(n9989), .A2(n14085), .ZN(n9672) );
  AND3_X1 U12393 ( .A1(n13387), .A2(n13472), .A3(n13473), .ZN(n9673) );
  AND2_X1 U12394 ( .A1(n11253), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11251) );
  NOR2_X2 U12395 ( .A1(n17068), .A2(n16072), .ZN(n17312) );
  INV_X1 U12396 ( .A(n17312), .ZN(n17483) );
  AND2_X1 U12397 ( .A1(n14200), .A2(n9929), .ZN(n9674) );
  OR3_X1 U12398 ( .A1(n14855), .A2(n10073), .A3(n10075), .ZN(n9675) );
  INV_X1 U12399 ( .A(n14974), .ZN(n10088) );
  AND2_X1 U12400 ( .A1(n14958), .A2(n15018), .ZN(n9676) );
  INV_X1 U12401 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n15614) );
  AND2_X1 U12402 ( .A1(n9623), .A2(n10049), .ZN(n9677) );
  NOR2_X1 U12403 ( .A1(n13567), .A2(n10042), .ZN(n10045) );
  INV_X1 U12404 ( .A(n9997), .ZN(n9996) );
  OR2_X1 U12405 ( .A1(n14199), .A2(n9998), .ZN(n9997) );
  OR2_X1 U12406 ( .A1(n9788), .A2(n14135), .ZN(n9678) );
  INV_X1 U12407 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18596) );
  INV_X1 U12408 ( .A(n12418), .ZN(n19006) );
  INV_X1 U12409 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18685) );
  INV_X1 U12410 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18741) );
  OR2_X1 U12411 ( .A1(n17483), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9679) );
  OR2_X1 U12412 ( .A1(n16065), .A2(n17421), .ZN(n9680) );
  AND2_X1 U12413 ( .A1(n13975), .A2(n10004), .ZN(n9681) );
  NOR2_X1 U12414 ( .A1(n17480), .A2(n17312), .ZN(n9682) );
  OR2_X1 U12415 ( .A1(n9917), .A2(n9916), .ZN(n9683) );
  AND3_X1 U12416 ( .A1(n13387), .A2(n13472), .A3(n10000), .ZN(n9684) );
  AND2_X1 U12417 ( .A1(n13065), .A2(n12226), .ZN(n9685) );
  AND2_X1 U12418 ( .A1(n9777), .A2(n9780), .ZN(n9686) );
  AND2_X1 U12419 ( .A1(n9622), .A2(n9928), .ZN(n9687) );
  OR2_X1 U12420 ( .A1(n9867), .A2(n16252), .ZN(n9688) );
  AND2_X1 U12421 ( .A1(n10108), .A2(n10444), .ZN(n9689) );
  OR2_X1 U12422 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n12065) );
  NAND2_X1 U12423 ( .A1(n12855), .A2(n12225), .ZN(n12848) );
  AND2_X1 U12424 ( .A1(n12855), .A2(n10024), .ZN(n13142) );
  NAND2_X1 U12425 ( .A1(n12855), .A2(n9625), .ZN(n12950) );
  INV_X1 U12426 ( .A(n10335), .ZN(n10336) );
  NOR2_X1 U12427 ( .A1(n9641), .A2(n14890), .ZN(n10923) );
  NOR2_X1 U12428 ( .A1(n11240), .A2(n10597), .ZN(n11238) );
  NAND2_X1 U12429 ( .A1(n12855), .A2(n9735), .ZN(n13375) );
  INV_X1 U12430 ( .A(n13375), .ZN(n10007) );
  NAND2_X1 U12431 ( .A1(n10007), .A2(n10008), .ZN(n13603) );
  NOR2_X1 U12432 ( .A1(n11252), .A2(n9973), .ZN(n11242) );
  AND2_X1 U12433 ( .A1(n10025), .A2(n12302), .ZN(n9690) );
  AND2_X1 U12434 ( .A1(n13539), .A2(n13538), .ZN(n12856) );
  NAND2_X1 U12435 ( .A1(n12856), .A2(n10046), .ZN(n12961) );
  INV_X1 U12436 ( .A(n12563), .ZN(n10050) );
  OR3_X1 U12437 ( .A1(n16529), .A2(n16220), .A3(n16531), .ZN(n9691) );
  AND2_X1 U12438 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9692) );
  INV_X1 U12439 ( .A(n14926), .ZN(n9981) );
  INV_X1 U12440 ( .A(n13137), .ZN(n9817) );
  AND2_X1 U12441 ( .A1(n15979), .A2(n10068), .ZN(n9693) );
  OR3_X1 U12442 ( .A1(n11234), .A2(n9985), .A3(n11229), .ZN(n9694) );
  NAND2_X1 U12443 ( .A1(n9790), .A2(n13075), .ZN(n12863) );
  OR2_X1 U12444 ( .A1(n19028), .A2(n10801), .ZN(n9695) );
  INV_X1 U12445 ( .A(n12438), .ZN(n9750) );
  INV_X1 U12446 ( .A(n13078), .ZN(n9794) );
  NAND2_X1 U12447 ( .A1(n12168), .A2(n11630), .ZN(n12892) );
  INV_X1 U12448 ( .A(n12892), .ZN(n9939) );
  AND2_X1 U12449 ( .A1(n12374), .A2(n12373), .ZN(n9696) );
  INV_X1 U12450 ( .A(n9947), .ZN(n9946) );
  NAND2_X1 U12451 ( .A1(n9692), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9947) );
  AND2_X1 U12452 ( .A1(n12415), .A2(n12435), .ZN(n9697) );
  INV_X1 U12453 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17800) );
  AND2_X1 U12454 ( .A1(n10923), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10922) );
  AND2_X1 U12455 ( .A1(n9946), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9698) );
  INV_X1 U12456 ( .A(n11060), .ZN(n10443) );
  OR2_X1 U12457 ( .A1(n10442), .A2(n10441), .ZN(n11060) );
  AND2_X1 U12458 ( .A1(n10923), .A2(n9692), .ZN(n11270) );
  AND4_X1 U12459 ( .A1(n11059), .A2(n11058), .A3(n11057), .A4(n11056), .ZN(
        n9699) );
  INV_X1 U12460 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17811) );
  AND2_X1 U12461 ( .A1(n18767), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15932) );
  INV_X1 U12462 ( .A(n15932), .ZN(n10099) );
  NAND2_X1 U12463 ( .A1(n17244), .A2(n9857), .ZN(n9859) );
  INV_X1 U12464 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17163) );
  NOR2_X1 U12465 ( .A1(n12938), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19819) );
  INV_X1 U12466 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n9834) );
  INV_X1 U12467 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9858) );
  INV_X1 U12468 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9872) );
  OR2_X1 U12469 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9700) );
  INV_X1 U12470 ( .A(n14585), .ZN(n9899) );
  INV_X1 U12471 ( .A(n11298), .ZN(n10109) );
  AND2_X1 U12472 ( .A1(n9614), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9701) );
  OR2_X1 U12473 ( .A1(n9700), .A2(n9851), .ZN(n9702) );
  AND2_X1 U12474 ( .A1(n9635), .A2(n10109), .ZN(n9703) );
  INV_X1 U12475 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9900) );
  INV_X1 U12476 ( .A(n15137), .ZN(n9825) );
  OR2_X1 U12477 ( .A1(n10713), .A2(n10712), .ZN(n19553) );
  AOI22_X2 U12478 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19973), .B1(DATAI_21_), 
        .B2(n19926), .ZN(n20508) );
  AOI22_X2 U12479 ( .A1(DATAI_17_), .A2(n19926), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n19973), .ZN(n20443) );
  AOI22_X2 U12480 ( .A1(DATAI_24_), .A2(n19926), .B1(BUF1_REG_24__SCAN_IN), 
        .B2(n19973), .ZN(n20364) );
  AOI22_X2 U12481 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19973), .B1(DATAI_27_), 
        .B2(n19926), .ZN(n20376) );
  AOI22_X2 U12482 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19973), .B1(DATAI_30_), 
        .B2(n19926), .ZN(n20389) );
  AOI22_X2 U12483 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19973), .B1(DATAI_31_), 
        .B2(n19926), .ZN(n20527) );
  AOI22_X2 U12484 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19041), .ZN(n19558) );
  NOR2_X2 U12485 ( .A1(n14848), .A2(n15063), .ZN(n19041) );
  AOI22_X2 U12486 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19973), .B1(DATAI_18_), 
        .B2(n19926), .ZN(n20494) );
  NAND3_X1 U12487 ( .A1(n9632), .A2(P3_EAX_REG_0__SCAN_IN), .A3(n9705), .ZN(
        n9704) );
  AOI21_X2 U12488 ( .B1(n15635), .B2(n15634), .A(n18422), .ZN(n16950) );
  NAND3_X1 U12489 ( .A1(n13809), .A2(n13805), .A3(n13811), .ZN(n9707) );
  NAND3_X1 U12490 ( .A1(n13807), .A2(n13806), .A3(n9666), .ZN(n9708) );
  NOR2_X2 U12491 ( .A1(n13867), .A2(n13849), .ZN(n18401) );
  NOR2_X2 U12492 ( .A1(n16693), .A2(n9713), .ZN(n16689) );
  OAI21_X1 U12493 ( .B1(n16691), .B2(P3_EBX_REG_28__SCAN_IN), .A(n9710), .ZN(
        P3_U2675) );
  INV_X1 U12494 ( .A(n16688), .ZN(n9711) );
  NOR2_X1 U12495 ( .A1(n16689), .A2(n16690), .ZN(n9712) );
  AND2_X1 U12496 ( .A1(n16947), .A2(n16681), .ZN(n9713) );
  NAND3_X1 U12497 ( .A1(n18358), .A2(n17927), .A3(n9714), .ZN(n13841) );
  NAND3_X1 U12498 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .ZN(n9718) );
  NOR2_X2 U12499 ( .A1(n13868), .A2(n18358), .ZN(n15517) );
  XNOR2_X2 U12500 ( .A(n9818), .B(n10606), .ZN(n12195) );
  AOI22_X1 U12501 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U12502 ( .A1(n10207), .A2(n10206), .ZN(n9720) );
  NAND2_X1 U12503 ( .A1(n10210), .A2(n10209), .ZN(n9721) );
  NAND3_X1 U12504 ( .A1(n9726), .A2(n9725), .A3(n9724), .ZN(n9723) );
  NAND3_X1 U12505 ( .A1(n9731), .A2(n9730), .A3(n9729), .ZN(n9728) );
  NOR2_X2 U12506 ( .A1(n9734), .A2(n9732), .ZN(n12351) );
  NAND4_X1 U12507 ( .A1(n10228), .A2(n10238), .A3(n19023), .A4(n9670), .ZN(
        n10220) );
  INV_X1 U12508 ( .A(n10220), .ZN(n9737) );
  NAND2_X1 U12509 ( .A1(n14730), .A2(n9741), .ZN(n9740) );
  INV_X1 U12510 ( .A(n12420), .ZN(n9751) );
  AND2_X2 U12511 ( .A1(n9746), .A2(n9745), .ZN(n14742) );
  NOR2_X1 U12512 ( .A1(n12420), .A2(n9750), .ZN(n9747) );
  INV_X1 U12513 ( .A(n9752), .ZN(n14749) );
  AND2_X2 U12514 ( .A1(n9883), .A2(n17483), .ZN(n17327) );
  OR2_X2 U12515 ( .A1(n17362), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9883) );
  NAND2_X1 U12516 ( .A1(n16066), .A2(n17588), .ZN(n16069) );
  AND2_X1 U12517 ( .A1(n16066), .A2(n9760), .ZN(n15617) );
  NAND2_X1 U12518 ( .A1(n9671), .A2(n9892), .ZN(n9763) );
  OAI211_X1 U12519 ( .C1(n9892), .C2(n9765), .A(n9764), .B(n14923), .ZN(n10868) );
  OR2_X2 U12520 ( .A1(n14948), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9892) );
  XNOR2_X2 U12521 ( .A(n9766), .B(n10127), .ZN(n10718) );
  INV_X2 U12522 ( .A(n10077), .ZN(n9766) );
  AND3_X2 U12523 ( .A1(n10418), .A2(n10419), .A3(n11060), .ZN(n10077) );
  INV_X1 U12524 ( .A(n10320), .ZN(n9767) );
  NAND4_X1 U12525 ( .A1(n10170), .A2(n9769), .A3(n10168), .A4(n10171), .ZN(
        n9768) );
  NAND4_X1 U12526 ( .A1(n10165), .A2(n9771), .A3(n10167), .A4(n10166), .ZN(
        n9770) );
  XNOR2_X2 U12527 ( .A(n10911), .B(n10910), .ZN(n14887) );
  OAI21_X2 U12528 ( .B1(n9896), .B2(n9772), .A(n10909), .ZN(n10911) );
  NAND3_X1 U12529 ( .A1(n13703), .A2(n9613), .A3(n13704), .ZN(n9774) );
  XNOR2_X1 U12530 ( .A(n10766), .B(n10992), .ZN(n13704) );
  NAND2_X1 U12531 ( .A1(n13387), .A2(n9782), .ZN(n13587) );
  NAND2_X1 U12532 ( .A1(n9778), .A2(n9686), .ZN(n13719) );
  NAND2_X1 U12533 ( .A1(n9778), .A2(n9776), .ZN(n13716) );
  NAND2_X1 U12534 ( .A1(n13472), .A2(n10001), .ZN(n9783) );
  NAND3_X1 U12535 ( .A1(n9785), .A2(n12767), .A3(n9803), .ZN(n9784) );
  INV_X1 U12536 ( .A(n11537), .ZN(n9786) );
  INV_X1 U12537 ( .A(n11538), .ZN(n9787) );
  NOR2_X2 U12538 ( .A1(n13734), .A2(n9678), .ZN(n14122) );
  NAND2_X1 U12539 ( .A1(n9790), .A2(n9789), .ZN(n12862) );
  NAND2_X1 U12540 ( .A1(n9612), .A2(n14002), .ZN(n14001) );
  NAND2_X1 U12541 ( .A1(n9794), .A2(n9793), .ZN(n13359) );
  INV_X1 U12542 ( .A(n13335), .ZN(n9796) );
  OAI21_X2 U12543 ( .B1(n9798), .B2(n9797), .A(n9795), .ZN(n13642) );
  NAND3_X1 U12544 ( .A1(n11613), .A2(n11556), .A3(n20197), .ZN(n11646) );
  NAND2_X2 U12545 ( .A1(n14343), .A2(n14294), .ZN(n14334) );
  OAI211_X2 U12546 ( .C1(n9808), .C2(n14421), .A(n14381), .B(n9807), .ZN(
        n14375) );
  NAND2_X2 U12547 ( .A1(n14423), .A2(n14422), .ZN(n14421) );
  OAI21_X2 U12548 ( .B1(n14688), .B2(n9856), .A(n9952), .ZN(n14423) );
  NAND2_X1 U12549 ( .A1(n9849), .A2(n9804), .ZN(n9800) );
  NAND2_X1 U12550 ( .A1(n9800), .A2(n11514), .ZN(n9805) );
  NAND2_X1 U12551 ( .A1(n9849), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11534) );
  NAND2_X1 U12552 ( .A1(n9849), .A2(n9802), .ZN(n9801) );
  INV_X1 U12553 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U12554 ( .A1(n20050), .A2(n11519), .ZN(n11533) );
  AND2_X1 U12555 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  XNOR2_X2 U12556 ( .A(n9805), .B(n11529), .ZN(n20050) );
  AOI21_X2 U12557 ( .B1(n14421), .B2(n9593), .A(n9808), .ZN(n9806) );
  NAND2_X1 U12558 ( .A1(n13154), .A2(n13155), .ZN(n9810) );
  NAND2_X1 U12559 ( .A1(n13091), .A2(n13092), .ZN(n9811) );
  NAND3_X1 U12560 ( .A1(n9815), .A2(n9814), .A3(n9813), .ZN(n9812) );
  CLKBUF_X1 U12561 ( .A(n13047), .Z(n9816) );
  NAND3_X1 U12562 ( .A1(n9816), .A2(n20398), .A3(n20194), .ZN(n20475) );
  NAND2_X2 U12563 ( .A1(n14687), .A2(n14283), .ZN(n14688) );
  NAND2_X2 U12564 ( .A1(n9904), .A2(n9903), .ZN(n14687) );
  AOI21_X1 U12565 ( .B1(n9818), .B2(n10610), .A(n10609), .ZN(n13539) );
  NAND2_X1 U12566 ( .A1(n15134), .A2(n9819), .ZN(P2_U3022) );
  NAND3_X1 U12567 ( .A1(n9822), .A2(n9820), .A3(n10558), .ZN(n15048) );
  NAND2_X1 U12568 ( .A1(n13695), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10533) );
  NAND2_X1 U12569 ( .A1(n10103), .A2(n9821), .ZN(n9820) );
  NAND2_X1 U12570 ( .A1(n10532), .A2(n10555), .ZN(n9821) );
  NAND3_X1 U12571 ( .A1(n10103), .A2(n13695), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n9822) );
  NOR2_X2 U12572 ( .A1(n19016), .A2(n19010), .ZN(n10987) );
  NAND2_X1 U12573 ( .A1(n9826), .A2(n11304), .ZN(P2_U3015) );
  NAND2_X1 U12574 ( .A1(n10904), .A2(n11303), .ZN(n9826) );
  XNOR2_X1 U12575 ( .A(n10902), .B(n9651), .ZN(n10904) );
  AND2_X4 U12576 ( .A1(n10341), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10335) );
  NAND3_X1 U12577 ( .A1(n10393), .A2(n10394), .A3(n10395), .ZN(n9830) );
  INV_X1 U12578 ( .A(n10871), .ZN(n15854) );
  NAND3_X1 U12579 ( .A1(n9925), .A2(n9924), .A3(n9923), .ZN(n10961) );
  NAND2_X2 U12580 ( .A1(n10259), .A2(n10219), .ZN(n10265) );
  AND2_X2 U12581 ( .A1(n9845), .A2(n9842), .ZN(n10259) );
  NAND2_X1 U12582 ( .A1(n9843), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U12583 ( .A1(n10980), .A2(n9844), .ZN(n9843) );
  NAND2_X1 U12584 ( .A1(n10983), .A2(n13457), .ZN(n9844) );
  NAND2_X1 U12585 ( .A1(n11213), .A2(n12601), .ZN(n9845) );
  NAND2_X1 U12586 ( .A1(n10768), .A2(n9918), .ZN(n10098) );
  NAND2_X1 U12587 ( .A1(n13703), .A2(n13704), .ZN(n10768) );
  AOI21_X2 U12588 ( .B1(n15016), .B2(n10086), .A(n15000), .ZN(n14992) );
  OAI21_X2 U12589 ( .B1(n15025), .B2(n15026), .A(n9847), .ZN(n15017) );
  NAND2_X1 U12590 ( .A1(n11445), .A2(n11515), .ZN(n9849) );
  NAND2_X1 U12591 ( .A1(n9852), .A2(n9954), .ZN(n9850) );
  INV_X1 U12592 ( .A(n9852), .ZN(n14309) );
  NOR2_X2 U12593 ( .A1(n11637), .A2(n9855), .ZN(n9854) );
  INV_X1 U12594 ( .A(n9859), .ZN(n16038) );
  NOR2_X1 U12595 ( .A1(n9866), .A2(n9688), .ZN(n16250) );
  NAND3_X1 U12596 ( .A1(n9871), .A2(n9647), .A3(n17509), .ZN(n17372) );
  OAI21_X1 U12597 ( .B1(n16219), .B2(n9691), .A(n9874), .ZN(n9873) );
  INV_X2 U12598 ( .A(n15536), .ZN(n17092) );
  NAND2_X1 U12599 ( .A1(n15443), .A2(n15444), .ZN(n15546) );
  OAI21_X1 U12600 ( .B1(n9879), .B2(n17544), .A(n9876), .ZN(n17525) );
  INV_X1 U12601 ( .A(n17527), .ZN(n9877) );
  XNOR2_X1 U12602 ( .A(n15485), .B(n15483), .ZN(n17544) );
  NOR2_X2 U12603 ( .A1(n17481), .A2(n17689), .ZN(n17710) );
  NAND2_X1 U12604 ( .A1(n15279), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10839) );
  AND2_X2 U12605 ( .A1(n10415), .A2(n10414), .ZN(n10418) );
  NAND2_X2 U12606 ( .A1(n10352), .A2(n10351), .ZN(n10419) );
  NAND2_X1 U12607 ( .A1(n9895), .A2(n9894), .ZN(n9893) );
  NOR2_X1 U12608 ( .A1(n10479), .A2(n10478), .ZN(n9894) );
  INV_X1 U12609 ( .A(n10477), .ZN(n9895) );
  NAND2_X1 U12610 ( .A1(n14315), .A2(n9897), .ZN(P1_U2969) );
  NOR2_X1 U12611 ( .A1(n9902), .A2(n13708), .ZN(n9901) );
  AOI21_X2 U12612 ( .B1(n20221), .B2(n15614), .A(n11577), .ZN(n11637) );
  XNOR2_X2 U12613 ( .A(n12767), .B(n20087), .ZN(n20221) );
  NAND2_X2 U12614 ( .A1(n11538), .A2(n11537), .ZN(n12767) );
  NAND2_X1 U12615 ( .A1(n10418), .A2(n10419), .ZN(n10444) );
  NAND2_X1 U12616 ( .A1(n9913), .A2(n9911), .ZN(n13390) );
  NAND3_X1 U12617 ( .A1(n10418), .A2(n10419), .A3(n9914), .ZN(n9912) );
  NAND3_X1 U12618 ( .A1(n10416), .A2(n10417), .A3(n9914), .ZN(n9913) );
  NAND3_X1 U12619 ( .A1(n10108), .A2(n10444), .A3(n10865), .ZN(n9915) );
  AOI21_X1 U12620 ( .B1(n9920), .B2(n15933), .A(n15932), .ZN(n15938) );
  XNOR2_X1 U12621 ( .A(n9920), .B(n15060), .ZN(n15333) );
  NAND2_X1 U12622 ( .A1(n12867), .A2(n12866), .ZN(n12873) );
  NAND2_X1 U12623 ( .A1(n14200), .A2(n9687), .ZN(n14136) );
  AND2_X2 U12624 ( .A1(n11315), .A2(n9936), .ZN(n11351) );
  AND2_X2 U12625 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U12626 ( .A1(n9936), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13122) );
  AND2_X2 U12627 ( .A1(n9936), .A2(n13116), .ZN(n11402) );
  AND2_X1 U12628 ( .A1(n11307), .A2(n9936), .ZN(n11563) );
  NOR2_X1 U12629 ( .A1(n11316), .A2(n9936), .ZN(n14711) );
  XNOR2_X2 U12630 ( .A(n11518), .B(n11461), .ZN(n11631) );
  NAND2_X1 U12631 ( .A1(n11631), .A2(n15614), .ZN(n11627) );
  OR2_X1 U12632 ( .A1(n10923), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9945) );
  NAND2_X1 U12633 ( .A1(n10923), .A2(n9698), .ZN(n9944) );
  NAND3_X1 U12634 ( .A1(n9945), .A2(n9944), .A3(n9943), .ZN(n11222) );
  INV_X1 U12635 ( .A(n11256), .ZN(n9948) );
  NAND2_X1 U12636 ( .A1(n9948), .A2(n9949), .ZN(n11255) );
  NAND2_X1 U12637 ( .A1(n9957), .A2(n9958), .ZN(n15808) );
  NAND2_X1 U12638 ( .A1(n13642), .A2(n13641), .ZN(n9963) );
  NAND2_X1 U12639 ( .A1(n9967), .A2(n9965), .ZN(n9970) );
  NOR2_X1 U12640 ( .A1(n9966), .A2(n18624), .ZN(n9965) );
  NOR2_X1 U12641 ( .A1(n18764), .A2(n9968), .ZN(n9966) );
  NAND2_X1 U12642 ( .A1(n18631), .A2(n9969), .ZN(n9967) );
  INV_X1 U12643 ( .A(n9971), .ZN(n18630) );
  INV_X1 U12644 ( .A(n9970), .ZN(n18622) );
  AOI21_X1 U12645 ( .B1(n15571), .B2(n9981), .A(n18676), .ZN(n9980) );
  NAND2_X1 U12646 ( .A1(n9978), .A2(n9977), .ZN(n15850) );
  NAND2_X1 U12647 ( .A1(n15571), .A2(n9979), .ZN(n9978) );
  NAND3_X1 U12648 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11261) );
  OAI21_X2 U12649 ( .B1(n13137), .B2(n13655), .A(n13090), .ZN(n13156) );
  NOR2_X1 U12650 ( .A1(n11234), .A2(n11229), .ZN(n11228) );
  INV_X1 U12651 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n9985) );
  NAND3_X1 U12652 ( .A1(n11431), .A2(n11422), .A3(n12979), .ZN(n12766) );
  INV_X1 U12653 ( .A(n14107), .ZN(n9986) );
  NAND2_X1 U12654 ( .A1(n9986), .A2(n9987), .ZN(n14060) );
  AND2_X1 U12655 ( .A1(n9612), .A2(n10004), .ZN(n13989) );
  NAND2_X1 U12656 ( .A1(n9612), .A2(n9681), .ZN(n10006) );
  NAND2_X1 U12657 ( .A1(n10011), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10010) );
  NAND4_X1 U12658 ( .A1(n10143), .A2(n10142), .A3(n10141), .A4(n10140), .ZN(
        n10011) );
  NAND2_X1 U12659 ( .A1(n10013), .A2(n13211), .ZN(n10012) );
  NAND4_X1 U12660 ( .A1(n10139), .A2(n10138), .A3(n10136), .A4(n10137), .ZN(
        n10013) );
  NAND2_X2 U12661 ( .A1(n10016), .A2(n10014), .ZN(n10205) );
  NAND2_X1 U12662 ( .A1(n10015), .A2(n13211), .ZN(n10014) );
  NAND4_X1 U12663 ( .A1(n10145), .A2(n10146), .A3(n10147), .A4(n10144), .ZN(
        n10015) );
  NAND4_X1 U12664 ( .A1(n10151), .A2(n10150), .A3(n10149), .A4(n10148), .ZN(
        n10017) );
  INV_X1 U12665 ( .A(n12352), .ZN(n10022) );
  INV_X1 U12666 ( .A(n14764), .ZN(n10020) );
  NAND3_X1 U12667 ( .A1(n17278), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n10027), .ZN(n15509) );
  NAND2_X1 U12668 ( .A1(n17275), .A2(n17620), .ZN(n10027) );
  OR2_X1 U12669 ( .A1(n17266), .A2(n10026), .ZN(n17623) );
  NOR2_X1 U12670 ( .A1(n17275), .A2(n17620), .ZN(n10026) );
  NOR2_X2 U12671 ( .A1(n16066), .A2(n17588), .ZN(n16071) );
  AND2_X2 U12672 ( .A1(n15508), .A2(n15507), .ZN(n17250) );
  OR2_X1 U12673 ( .A1(n15330), .A2(n15862), .ZN(n10041) );
  NOR2_X1 U12674 ( .A1(n13567), .A2(n13566), .ZN(n15028) );
  INV_X1 U12675 ( .A(n15027), .ZN(n10044) );
  INV_X1 U12676 ( .A(n10045), .ZN(n15004) );
  NAND2_X1 U12677 ( .A1(n12856), .A2(n9668), .ZN(n13008) );
  NOR2_X1 U12678 ( .A1(n14760), .A2(n14746), .ZN(n14747) );
  OR3_X1 U12679 ( .A1(n14760), .A2(n10051), .A3(n14746), .ZN(n10918) );
  INV_X1 U12680 ( .A(n14743), .ZN(n10056) );
  NAND2_X1 U12681 ( .A1(n15235), .A2(n13606), .ZN(n13681) );
  NOR2_X1 U12682 ( .A1(n9636), .A2(n14805), .ZN(n14795) );
  INV_X1 U12683 ( .A(n14785), .ZN(n10061) );
  INV_X1 U12684 ( .A(n12921), .ZN(n10062) );
  NAND2_X1 U12685 ( .A1(n10062), .A2(n9617), .ZN(n11071) );
  NOR2_X2 U12686 ( .A1(n11053), .A2(n9699), .ZN(n10065) );
  OR2_X2 U12687 ( .A1(n10205), .A2(n10719), .ZN(n10937) );
  AND2_X2 U12688 ( .A1(n10101), .A2(n10076), .ZN(n10354) );
  AND2_X2 U12689 ( .A1(n12845), .A2(n10076), .ZN(n19179) );
  AOI21_X2 U12690 ( .B1(n10085), .B2(n10081), .A(n10078), .ZN(n15040) );
  NAND2_X1 U12691 ( .A1(n14949), .A2(n14948), .ZN(n15054) );
  NAND3_X1 U12692 ( .A1(n14949), .A2(n14948), .A3(n14951), .ZN(n10085) );
  INV_X1 U12693 ( .A(n10095), .ZN(n10086) );
  NAND2_X1 U12694 ( .A1(n15016), .A2(n14958), .ZN(n15015) );
  AOI21_X1 U12695 ( .B1(n15016), .B2(n10093), .A(n10092), .ZN(n14977) );
  OAI21_X1 U12696 ( .B1(n10091), .B2(n10089), .A(n10087), .ZN(n14965) );
  INV_X1 U12697 ( .A(n15016), .ZN(n10091) );
  INV_X1 U12698 ( .A(n15935), .ZN(n10100) );
  AND2_X1 U12699 ( .A1(n10298), .A2(n10101), .ZN(n19314) );
  AND2_X1 U12700 ( .A1(n10301), .A2(n10101), .ZN(n10353) );
  NAND3_X1 U12701 ( .A1(n10108), .A2(n10444), .A3(n13396), .ZN(n13397) );
  NAND2_X1 U12702 ( .A1(n9611), .A2(n9635), .ZN(n14902) );
  AND2_X1 U12703 ( .A1(n9611), .A2(n10110), .ZN(n14901) );
  NOR2_X1 U12704 ( .A1(n15793), .A2(n18676), .ZN(n11273) );
  NAND2_X1 U12705 ( .A1(n14050), .A2(n14051), .ZN(n14037) );
  INV_X1 U12706 ( .A(n10227), .ZN(n12508) );
  NAND2_X1 U12707 ( .A1(n13716), .A2(n13736), .ZN(n11763) );
  NAND2_X1 U12708 ( .A1(n14873), .A2(n18977), .ZN(n11220) );
  NAND2_X1 U12709 ( .A1(n11763), .A2(n13735), .ZN(n13734) );
  OAI211_X1 U12710 ( .C1(n10961), .C2(n10964), .A(n10962), .B(n14878), .ZN(
        n10902) );
  OAI22_X2 U12711 ( .A1(n14887), .A2(n15097), .B1(n10913), .B2(n10912), .ZN(
        n10916) );
  AOI21_X1 U12712 ( .B1(n15089), .B2(n18977), .A(n15088), .ZN(n15090) );
  AND2_X1 U12713 ( .A1(n12351), .A2(n12374), .ZN(n12352) );
  NAND2_X1 U12714 ( .A1(n10904), .A2(n10903), .ZN(n10905) );
  NAND2_X1 U12715 ( .A1(n10988), .A2(n10238), .ZN(n10217) );
  AND2_X1 U12716 ( .A1(n10977), .A2(n19044), .ZN(n10233) );
  NOR2_X1 U12717 ( .A1(n10977), .A2(n19010), .ZN(n10221) );
  INV_X1 U12718 ( .A(n10240), .ZN(n10242) );
  NAND2_X1 U12719 ( .A1(n10226), .A2(n10225), .ZN(n10262) );
  XNOR2_X1 U12720 ( .A(n11050), .B(n11049), .ZN(n12920) );
  NAND2_X1 U12721 ( .A1(n10272), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10260) );
  AOI211_X2 U12722 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15085), .A(
        n15084), .B(n15083), .ZN(n15086) );
  XNOR2_X1 U12723 ( .A(n12844), .B(n12843), .ZN(n19277) );
  OAI21_X1 U12724 ( .B1(n12221), .B2(n12196), .A(n13421), .ZN(n12844) );
  NAND2_X4 U12725 ( .A1(n10193), .A2(n10192), .ZN(n13238) );
  BUF_X4 U12726 ( .A(n11470), .Z(n12081) );
  OR2_X1 U12727 ( .A1(n11275), .A2(n18862), .ZN(n12530) );
  NOR2_X1 U12728 ( .A1(n18823), .A2(n11275), .ZN(n11291) );
  INV_X1 U12729 ( .A(n10685), .ZN(n10644) );
  INV_X1 U12730 ( .A(n10234), .ZN(n11041) );
  NAND2_X1 U12731 ( .A1(n12732), .A2(n10234), .ZN(n13439) );
  OR2_X1 U12732 ( .A1(n18881), .A2(n10234), .ZN(n18861) );
  NOR2_X1 U12733 ( .A1(n15005), .A2(n14780), .ZN(n10111) );
  INV_X1 U12734 ( .A(n11232), .ZN(n11233) );
  CLKBUF_X3 U12735 ( .A(n13825), .Z(n16872) );
  NOR2_X1 U12737 ( .A1(n13757), .A2(n13756), .ZN(n15435) );
  INV_X1 U12738 ( .A(n18759), .ZN(n18823) );
  OR4_X1 U12739 ( .A1(n15070), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n11299), .A4(n11298), .ZN(n10113) );
  AND3_X1 U12740 ( .A1(n11301), .A2(n11300), .A3(n10113), .ZN(n10114) );
  INV_X1 U12741 ( .A(n15309), .ZN(n11303) );
  NAND2_X1 U12742 ( .A1(n17758), .A2(n17718), .ZN(n10115) );
  INV_X1 U12743 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18756) );
  INV_X1 U12744 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15483) );
  INV_X1 U12745 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17718) );
  NOR2_X1 U12746 ( .A1(n12110), .A2(n11425), .ZN(n10116) );
  INV_X1 U12747 ( .A(n11426), .ZN(n11427) );
  OR2_X1 U12748 ( .A1(n9600), .A2(n15336), .ZN(n10117) );
  AND4_X1 U12749 ( .A1(n10972), .A2(n13457), .A3(n10720), .A4(n19033), .ZN(
        n10118) );
  INV_X1 U12750 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12211) );
  OR2_X1 U12751 ( .A1(n17483), .A2(n17579), .ZN(n10119) );
  AND2_X1 U12752 ( .A1(n10238), .A2(n19044), .ZN(n10120) );
  INV_X1 U12753 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14928) );
  INV_X1 U12754 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10596) );
  INV_X1 U12755 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15031) );
  INV_X1 U12756 ( .A(n19170), .ZN(n19212) );
  AND2_X1 U12757 ( .A1(n10744), .A2(n10586), .ZN(n10122) );
  NAND2_X1 U12758 ( .A1(n16009), .A2(n17573), .ZN(n17359) );
  NAND2_X1 U12759 ( .A1(n18596), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12209) );
  NOR2_X2 U12760 ( .A1(n18807), .A2(n19544), .ZN(n18802) );
  AND2_X1 U12761 ( .A1(n12530), .A2(n12529), .ZN(n10123) );
  NOR2_X1 U12762 ( .A1(n20351), .A2(n20316), .ZN(n10124) );
  INV_X1 U12763 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12771) );
  AND2_X1 U12764 ( .A1(n10118), .A2(n10120), .ZN(n10125) );
  INV_X1 U12765 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17758) );
  INV_X1 U12766 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15336) );
  AND2_X1 U12767 ( .A1(n12948), .A2(n12951), .ZN(n10128) );
  OR2_X1 U12768 ( .A1(n12586), .A2(n9600), .ZN(n15946) );
  AND2_X1 U12769 ( .A1(n13227), .A2(n13226), .ZN(n15355) );
  INV_X1 U12770 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13264) );
  INV_X2 U12771 ( .A(n16927), .ZN(n16941) );
  INV_X1 U12772 ( .A(n11020), .ZN(n11186) );
  OR2_X1 U12773 ( .A1(n15805), .A2(n15063), .ZN(n10129) );
  OR2_X1 U12774 ( .A1(n18595), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15891) );
  INV_X1 U12775 ( .A(n18791), .ZN(n18970) );
  INV_X1 U12776 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10711) );
  AND4_X1 U12778 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n10130) );
  AND4_X1 U12779 ( .A1(n11346), .A2(n11345), .A3(n11344), .A4(n11343), .ZN(
        n10131) );
  AND4_X1 U12780 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n10132) );
  INV_X1 U12781 ( .A(n11522), .ZN(n12880) );
  AND4_X1 U12782 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n10133) );
  INV_X1 U12783 ( .A(n12145), .ZN(n12138) );
  OR2_X1 U12784 ( .A1(n13656), .A2(n15614), .ZN(n11496) );
  OR2_X1 U12785 ( .A1(n12127), .A2(n12979), .ZN(n12140) );
  INV_X1 U12786 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10562) );
  AND2_X1 U12787 ( .A1(n11511), .A2(n11510), .ZN(n11523) );
  INV_X1 U12788 ( .A(n10342), .ZN(n13200) );
  NAND2_X1 U12789 ( .A1(n11438), .A2(n11437), .ZN(n11417) );
  INV_X1 U12790 ( .A(n13718), .ZN(n11745) );
  OR2_X1 U12791 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  INV_X1 U12792 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10597) );
  AND2_X1 U12793 ( .A1(n10663), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U12794 ( .A1(n19720), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10578) );
  NOR2_X1 U12795 ( .A1(n12133), .A2(n12134), .ZN(n12132) );
  INV_X1 U12796 ( .A(n13193), .ZN(n11653) );
  INV_X1 U12797 ( .A(n11421), .ZN(n12116) );
  AND4_X1 U12798 ( .A1(n11458), .A2(n11457), .A3(n12903), .A4(n12758), .ZN(
        n11459) );
  NOR2_X1 U12799 ( .A1(n12145), .A2(n13655), .ZN(n12150) );
  NAND2_X1 U12800 ( .A1(n10566), .A2(n10565), .ZN(n10570) );
  NAND2_X1 U12801 ( .A1(n10297), .A2(n10296), .ZN(n10607) );
  INV_X1 U12802 ( .A(n12395), .ZN(n12396) );
  NOR2_X1 U12803 ( .A1(n13614), .A2(n10535), .ZN(n10527) );
  NAND2_X1 U12804 ( .A1(n10977), .A2(n10234), .ZN(n10944) );
  AND2_X1 U12805 ( .A1(n18832), .A2(n10285), .ZN(n10299) );
  OR2_X1 U12806 ( .A1(n11952), .A2(n11951), .ZN(n11975) );
  NAND2_X1 U12807 ( .A1(n19968), .A2(n11438), .ZN(n11426) );
  AND2_X1 U12808 ( .A1(n12041), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12042) );
  AND2_X1 U12809 ( .A1(n11959), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11960) );
  INV_X1 U12810 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11884) );
  INV_X1 U12811 ( .A(n12097), .ZN(n11804) );
  NAND2_X1 U12812 ( .A1(n12901), .A2(n11421), .ZN(n11432) );
  INV_X1 U12813 ( .A(n12938), .ZN(n11560) );
  NAND2_X1 U12814 ( .A1(n11460), .A2(n11459), .ZN(n11517) );
  AOI21_X1 U12815 ( .B1(n10570), .B2(n10568), .A(n10567), .ZN(n10575) );
  INV_X1 U12816 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11262) );
  AND2_X1 U12817 ( .A1(n12419), .A2(n9697), .ZN(n12420) );
  OR2_X1 U12818 ( .A1(n12349), .A2(n12348), .ZN(n12368) );
  OR2_X1 U12819 ( .A1(n12240), .A2(n12239), .ZN(n18838) );
  OR2_X1 U12820 ( .A1(n15104), .A2(n11002), .ZN(n15070) );
  INV_X1 U12821 ( .A(n10762), .ZN(n10530) );
  NAND3_X1 U12822 ( .A1(n10234), .A2(n11023), .A3(n10988), .ZN(n10983) );
  INV_X1 U12823 ( .A(n12198), .ZN(n12199) );
  OAI21_X1 U12824 ( .B1(n17369), .B2(n17614), .A(n15503), .ZN(n15504) );
  AOI21_X1 U12825 ( .B1(n18385), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13855), .ZN(n13861) );
  NOR2_X1 U12826 ( .A1(n17036), .A2(n17933), .ZN(n15518) );
  AND2_X1 U12827 ( .A1(n13595), .A2(n13594), .ZN(n13596) );
  NAND2_X1 U12828 ( .A1(n12979), .A2(n19932), .ZN(n12756) );
  NAND2_X1 U12829 ( .A1(n12042), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13282) );
  AND2_X1 U12830 ( .A1(n12915), .A2(n13105), .ZN(n15736) );
  NAND2_X1 U12831 ( .A1(n12901), .A2(n13660), .ZN(n13656) );
  INV_X1 U12832 ( .A(n20274), .ZN(n20319) );
  OR2_X1 U12833 ( .A1(n11149), .A2(n11148), .ZN(n12226) );
  OR2_X1 U12834 ( .A1(n11091), .A2(n11090), .ZN(n12223) );
  AND2_X1 U12835 ( .A1(n12330), .A2(n12329), .ZN(n12371) );
  AND2_X1 U12836 ( .A1(n11184), .A2(n11183), .ZN(n15233) );
  OR2_X1 U12837 ( .A1(n18672), .A2(n10865), .ZN(n10850) );
  INV_X1 U12838 ( .A(n10718), .ZN(n10494) );
  OR2_X1 U12839 ( .A1(n13490), .A2(n13489), .ZN(n13498) );
  INV_X1 U12840 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n13409) );
  NOR3_X1 U12841 ( .A1(n17353), .A2(n15506), .A3(n17357), .ZN(n17278) );
  OAI211_X1 U12842 ( .C1(n13861), .C2(n13860), .A(n13870), .B(n13859), .ZN(
        n15523) );
  INV_X1 U12843 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15643) );
  INV_X1 U12844 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19767) );
  AND2_X1 U12845 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n11673), .ZN(
        n11674) );
  INV_X1 U12846 ( .A(n19830), .ZN(n19782) );
  INV_X1 U12847 ( .A(n11425), .ZN(n13309) );
  OR2_X1 U12848 ( .A1(n12826), .A2(n13945), .ZN(n12827) );
  INV_X1 U12849 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14386) );
  NOR2_X1 U12850 ( .A1(n11839), .A2(n20756), .ZN(n11853) );
  OR2_X1 U12851 ( .A1(n14618), .A2(n14525), .ZN(n14595) );
  AND2_X1 U12852 ( .A1(n13906), .A2(n13905), .ZN(n14125) );
  OR2_X1 U12853 ( .A1(n15740), .A2(n13061), .ZN(n15730) );
  AND2_X1 U12854 ( .A1(n12910), .A2(n12909), .ZN(n14520) );
  AND2_X1 U12855 ( .A1(n20052), .A2(n20080), .ZN(n20059) );
  INV_X1 U12856 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20397) );
  INV_X1 U12857 ( .A(n20009), .ZN(n19929) );
  AND2_X2 U12858 ( .A1(n12155), .A2(n12154), .ZN(n12936) );
  INV_X1 U12859 ( .A(n13232), .ZN(n11282) );
  OAI22_X1 U12860 ( .A1(n11222), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n18596), 
        .B2(n11221), .ZN(n11226) );
  INV_X1 U12861 ( .A(n10273), .ZN(n10689) );
  OR2_X1 U12862 ( .A1(n11019), .A2(n11018), .ZN(n13376) );
  AND2_X1 U12863 ( .A1(n11203), .A2(n11202), .ZN(n14805) );
  AND3_X1 U12864 ( .A1(n11063), .A2(n11062), .A3(n11061), .ZN(n13427) );
  AND2_X1 U12865 ( .A1(n11194), .A2(n11193), .ZN(n15147) );
  OR2_X1 U12866 ( .A1(n10850), .A2(n15250), .ZN(n15039) );
  XNOR2_X1 U12867 ( .A(n10556), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15931) );
  OR2_X1 U12868 ( .A1(n15203), .A2(n18963), .ZN(n15267) );
  OR2_X1 U12869 ( .A1(n10584), .A2(n19717), .ZN(n15631) );
  OR2_X1 U12870 ( .A1(n12547), .A2(n12546), .ZN(n12549) );
  OR2_X1 U12871 ( .A1(n19240), .A2(n19239), .ZN(n19248) );
  INV_X1 U12872 ( .A(n19308), .ZN(n19309) );
  OR2_X1 U12873 ( .A1(n19376), .A2(n19373), .ZN(n19404) );
  NAND2_X1 U12874 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19553), .ZN(n19022) );
  OR2_X1 U12875 ( .A1(n19550), .A2(n19545), .ZN(n19607) );
  NOR2_X1 U12876 ( .A1(n17808), .A2(n15525), .ZN(n18561) );
  NOR2_X1 U12877 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16361), .ZN(n16348) );
  NOR2_X1 U12878 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16485), .ZN(n16467) );
  INV_X1 U12879 ( .A(n16562), .ZN(n16569) );
  NAND2_X1 U12880 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16884), .ZN(n16864) );
  NAND2_X1 U12881 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17281), .ZN(
        n17258) );
  NOR2_X1 U12882 ( .A1(n17428), .A2(n17418), .ZN(n17413) );
  INV_X1 U12883 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17418) );
  AND2_X1 U12884 ( .A1(n17265), .A2(n10119), .ZN(n15510) );
  OR2_X1 U12885 ( .A1(n17614), .A2(n17620), .ZN(n17601) );
  INV_X1 U12886 ( .A(n17866), .ZN(n17849) );
  INV_X1 U12887 ( .A(n17370), .ZN(n17689) );
  INV_X1 U12888 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15467) );
  INV_X1 U12889 ( .A(n18189), .ZN(n18165) );
  NOR2_X1 U12890 ( .A1(n13774), .A2(n13773), .ZN(n17933) );
  INV_X1 U12891 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18395) );
  AND2_X1 U12892 ( .A1(n12887), .A2(n12752), .ZN(n19739) );
  AND2_X1 U12893 ( .A1(n14069), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14058) );
  NAND2_X1 U12894 ( .A1(n13958), .A2(n13304), .ZN(n19801) );
  NOR2_X1 U12895 ( .A1(n19817), .A2(n13517), .ZN(n13720) );
  NOR2_X1 U12896 ( .A1(n11649), .A2(n13433), .ZN(n11673) );
  INV_X1 U12897 ( .A(n19850), .ZN(n14197) );
  INV_X1 U12898 ( .A(n14206), .ZN(n19845) );
  NAND2_X1 U12899 ( .A1(n12976), .A2(n12158), .ZN(n12172) );
  INV_X2 U12900 ( .A(n13006), .ZN(n19904) );
  AND2_X1 U12901 ( .A1(n12936), .A2(n12157), .ZN(n12976) );
  INV_X1 U12902 ( .A(n19748), .ZN(n15692) );
  NOR2_X1 U12903 ( .A1(n11684), .A2(n19781), .ZN(n11714) );
  AND2_X1 U12904 ( .A1(n12862), .A2(n12865), .ZN(n13356) );
  AND2_X1 U12905 ( .A1(n14587), .A2(n14533), .ZN(n14575) );
  OR2_X1 U12906 ( .A1(n14615), .A2(n14524), .ZN(n14606) );
  NOR2_X1 U12907 ( .A1(n14650), .A2(n14519), .ZN(n14635) );
  INV_X1 U12908 ( .A(n14520), .ZN(n15735) );
  NAND2_X1 U12909 ( .A1(n12897), .A2(n12896), .ZN(n12915) );
  AND2_X1 U12910 ( .A1(n12915), .A2(n12912), .ZN(n19911) );
  OAI22_X1 U12911 ( .A1(n19942), .A2(n19941), .B1(n20281), .B2(n20088), .ZN(
        n19979) );
  OR2_X1 U12912 ( .A1(n20010), .A2(n20009), .ZN(n20127) );
  NAND2_X1 U12913 ( .A1(n19927), .A2(n13137), .ZN(n20049) );
  INV_X1 U12914 ( .A(n20094), .ZN(n20118) );
  INV_X1 U12915 ( .A(n20187), .ZN(n20144) );
  INV_X1 U12916 ( .A(n20310), .ZN(n20266) );
  OAI22_X1 U12917 ( .A1(n20283), .A2(n20282), .B1(n20281), .B2(n20427), .ZN(
        n20312) );
  OAI22_X1 U12918 ( .A1(n20361), .A2(n20360), .B1(n20428), .B2(n20359), .ZN(
        n20391) );
  AND2_X1 U12919 ( .A1(n20426), .A2(n20350), .ZN(n20421) );
  INV_X1 U12920 ( .A(n20437), .ZN(n20459) );
  INV_X1 U12921 ( .A(n20515), .ZN(n20522) );
  AND2_X1 U12922 ( .A1(n15606), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15611) );
  INV_X1 U12923 ( .A(n20623), .ZN(n20631) );
  INV_X1 U12924 ( .A(n20598), .ZN(n20592) );
  OAI21_X1 U12925 ( .B1(n14871), .B2(n18796), .A(n11289), .ZN(n11290) );
  INV_X1 U12926 ( .A(n18775), .ZN(n18822) );
  AND2_X1 U12927 ( .A1(n18958), .A2(n11276), .ZN(n18759) );
  OR3_X1 U12928 ( .A1(n18598), .A2(n16001), .A3(n11285), .ZN(n18825) );
  OR2_X1 U12929 ( .A1(n11179), .A2(n11178), .ZN(n13565) );
  NAND2_X2 U12930 ( .A1(n12507), .A2(n12613), .ZN(n18881) );
  INV_X1 U12931 ( .A(n18961), .ZN(n18955) );
  INV_X1 U12932 ( .A(n15946), .ZN(n10903) );
  INV_X1 U12933 ( .A(n15063), .ZN(n15950) );
  INV_X1 U12934 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12684) );
  INV_X1 U12935 ( .A(n12743), .ZN(n18963) );
  OR2_X1 U12936 ( .A1(n18973), .A2(n18964), .ZN(n15203) );
  NAND2_X1 U12937 ( .A1(n12549), .A2(n12548), .ZN(n19709) );
  OAI21_X1 U12938 ( .B1(n19003), .B2(n19002), .A(n19001), .ZN(n19048) );
  INV_X1 U12939 ( .A(n19074), .ZN(n19078) );
  INV_X1 U12940 ( .A(n19069), .ZN(n19108) );
  AND2_X1 U12941 ( .A1(n19207), .A2(n19375), .ZN(n19131) );
  AND2_X1 U12942 ( .A1(n19238), .A2(n19375), .ZN(n19166) );
  AND2_X1 U12943 ( .A1(n19238), .A2(n19450), .ZN(n19234) );
  INV_X1 U12944 ( .A(n19275), .ZN(n19267) );
  INV_X1 U12945 ( .A(n19307), .ZN(n19299) );
  INV_X1 U12946 ( .A(n19395), .ZN(n19406) );
  INV_X1 U12947 ( .A(n19483), .ZN(n19471) );
  INV_X1 U12948 ( .A(n19572), .ZN(n19508) );
  OAI22_X1 U12949 ( .A1(n19040), .A2(n19039), .B1(n19038), .B2(n19037), .ZN(
        n19534) );
  INV_X1 U12950 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19639) );
  NOR2_X1 U12951 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16277), .ZN(n16263) );
  NOR2_X1 U12952 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16299), .ZN(n16286) );
  NOR2_X1 U12953 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16340), .ZN(n16327) );
  NOR2_X1 U12954 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16387), .ZN(n16374) );
  NOR2_X1 U12955 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16409), .ZN(n16391) );
  INV_X1 U12956 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16433) );
  NOR2_X1 U12957 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16507), .ZN(n16489) );
  OAI211_X1 U12958 ( .C1(n18428), .C2(n18419), .A(n16523), .B(n18589), .ZN(
        n16473) );
  NAND2_X1 U12959 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16793), .ZN(n16792) );
  NOR2_X1 U12960 ( .A1(n17125), .A2(n17016), .ZN(n17011) );
  INV_X1 U12961 ( .A(n17086), .ZN(n17063) );
  INV_X1 U12962 ( .A(n16009), .ZN(n17574) );
  NOR2_X1 U12963 ( .A1(n17164), .A2(n17101), .ZN(n17132) );
  INV_X1 U12964 ( .A(n17207), .ZN(n17211) );
  INV_X1 U12965 ( .A(n17573), .ZN(n17559) );
  NOR2_X1 U12966 ( .A1(n18576), .A2(n16177), .ZN(n16014) );
  OAI21_X2 U12967 ( .B1(n18357), .B2(n18370), .A(n18356), .ZN(n18378) );
  NOR2_X1 U12968 ( .A1(n17635), .A2(n17634), .ZN(n17672) );
  NAND2_X1 U12969 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17396), .ZN(
        n17395) );
  NOR2_X2 U12970 ( .A1(n17068), .A2(n17898), .ZN(n17814) );
  INV_X1 U12971 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20762) );
  NAND2_X1 U12972 ( .A1(n17563), .A2(n17571), .ZN(n17562) );
  NOR3_X1 U12973 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18575), .ZN(n18118) );
  INV_X1 U12974 ( .A(n18530), .ZN(n18545) );
  NOR2_X1 U12975 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17914), .ZN(n18264) );
  INV_X1 U12976 ( .A(n17992), .ZN(n18024) );
  INV_X1 U12977 ( .A(n18057), .ZN(n18067) );
  INV_X1 U12978 ( .A(n18082), .ZN(n18090) );
  INV_X1 U12979 ( .A(n18131), .ZN(n18141) );
  INV_X1 U12980 ( .A(n18128), .ZN(n18161) );
  INV_X1 U12981 ( .A(n18303), .ZN(n18259) );
  INV_X1 U12982 ( .A(n18419), .ZN(n18429) );
  INV_X1 U12983 ( .A(n18577), .ZN(n18571) );
  INV_X1 U12984 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18452) );
  INV_X1 U12985 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18441) );
  AND2_X1 U12986 ( .A1(n19739), .A2(n12937), .ZN(n12642) );
  INV_X1 U12987 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20429) );
  OR3_X1 U12988 ( .A1(n14009), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n13996), .ZN(
        n13998) );
  OR2_X1 U12989 ( .A1(n14103), .A2(n20577), .ZN(n14096) );
  NAND2_X1 U12990 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13720), .ZN(n19776) );
  NAND2_X1 U12991 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n13316), .ZN(n19817) );
  OR2_X1 U12992 ( .A1(n14302), .A2(n13288), .ZN(n19843) );
  NAND2_X1 U12993 ( .A1(n19850), .A2(n9938), .ZN(n14196) );
  NAND2_X1 U12994 ( .A1(n19860), .A2(n19932), .ZN(n19851) );
  INV_X1 U12995 ( .A(n19860), .ZN(n19885) );
  AND2_X1 U12996 ( .A1(n12976), .A2(n12975), .ZN(n13006) );
  INV_X1 U12997 ( .A(n19905), .ZN(n13017) );
  OR2_X1 U12998 ( .A1(n15686), .A2(n13351), .ZN(n15696) );
  AND2_X1 U12999 ( .A1(n14414), .A2(n14413), .ZN(n14653) );
  INV_X1 U13000 ( .A(n19911), .ZN(n15775) );
  NAND2_X1 U13001 ( .A1(n12915), .A2(n12902), .ZN(n14704) );
  INV_X1 U13002 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20220) );
  NOR2_X1 U13003 ( .A1(n12769), .A2(n19931), .ZN(n20613) );
  NAND2_X1 U13004 ( .A1(n19928), .A2(n20350), .ZN(n20008) );
  OR2_X1 U13005 ( .A1(n20049), .A2(n20127), .ZN(n20041) );
  OR2_X1 U13006 ( .A1(n20049), .A2(n20149), .ZN(n20081) );
  NAND2_X1 U13007 ( .A1(n20199), .A2(n20350), .ZN(n20148) );
  NAND2_X1 U13008 ( .A1(n20199), .A2(n20396), .ZN(n20187) );
  NAND2_X1 U13009 ( .A1(n20199), .A2(n20425), .ZN(n20646) );
  NAND2_X1 U13010 ( .A1(n20327), .A2(n20350), .ZN(n20270) );
  NAND2_X1 U13011 ( .A1(n20327), .A2(n20396), .ZN(n20310) );
  NAND2_X1 U13012 ( .A1(n20327), .A2(n20425), .ZN(n20343) );
  NAND2_X1 U13013 ( .A1(n20327), .A2(n20326), .ZN(n20395) );
  NAND2_X1 U13014 ( .A1(n20426), .A2(n20396), .ZN(n20437) );
  NAND2_X1 U13015 ( .A1(n20426), .A2(n20326), .ZN(n20515) );
  NOR2_X1 U13016 ( .A1(n11609), .A2(n15606), .ZN(n15781) );
  INV_X1 U13017 ( .A(n20606), .ZN(n20530) );
  INV_X1 U13018 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20532) );
  NAND2_X1 U13019 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20637), .ZN(n20594) );
  NAND2_X1 U13020 ( .A1(n20637), .A2(n20545), .ZN(n20598) );
  NAND2_X1 U13021 ( .A1(n10589), .A2(n12613), .ZN(n12586) );
  NOR2_X1 U13022 ( .A1(n11291), .A2(n11290), .ZN(n11292) );
  INV_X1 U13023 ( .A(n18831), .ZN(n18796) );
  INV_X1 U13024 ( .A(n18802), .ZN(n18833) );
  INV_X1 U13025 ( .A(n11284), .ZN(n18811) );
  INV_X1 U13026 ( .A(n12537), .ZN(n12538) );
  XNOR2_X1 U13027 ( .A(n12727), .B(n12726), .ZN(n19139) );
  INV_X1 U13028 ( .A(n18881), .ZN(n14858) );
  OR2_X1 U13029 ( .A1(n18881), .A2(n19044), .ZN(n18862) );
  INV_X1 U13030 ( .A(n12636), .ZN(n18909) );
  INV_X1 U13031 ( .A(n18894), .ZN(n18926) );
  OR2_X1 U13032 ( .A1(n18955), .A2(n18958), .ZN(n12650) );
  OR2_X1 U13033 ( .A1(n12580), .A2(n19006), .ZN(n12666) );
  INV_X1 U13034 ( .A(n12210), .ZN(n12729) );
  OR2_X1 U13035 ( .A1(n11218), .A2(n19724), .ZN(n15978) );
  OR2_X1 U13036 ( .A1(n11218), .A2(n10967), .ZN(n15309) );
  NAND2_X1 U13037 ( .A1(n19308), .A2(n19207), .ZN(n19074) );
  INV_X1 U13038 ( .A(n19131), .ZN(n19112) );
  INV_X1 U13039 ( .A(n19133), .ZN(n19125) );
  AND2_X1 U13040 ( .A1(n19144), .A2(n19143), .ZN(n19150) );
  INV_X1 U13041 ( .A(n19202), .ZN(n19196) );
  INV_X1 U13042 ( .A(n19234), .ZN(n19215) );
  NAND2_X1 U13043 ( .A1(n19548), .A2(n19207), .ZN(n19275) );
  NAND2_X1 U13044 ( .A1(n19238), .A2(n19548), .ZN(n19307) );
  INV_X1 U13045 ( .A(n19363), .ZN(n19338) );
  NAND2_X1 U13046 ( .A1(n19411), .A2(n19375), .ZN(n19395) );
  NAND2_X1 U13047 ( .A1(n19411), .A2(n19450), .ZN(n19483) );
  AND2_X1 U13048 ( .A1(n19492), .A2(n19491), .ZN(n19524) );
  INV_X1 U13049 ( .A(n19687), .ZN(n19616) );
  NAND2_X1 U13050 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19621), .ZN(n19735) );
  INV_X1 U13051 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18575) );
  INV_X1 U13052 ( .A(n16559), .ZN(n16570) );
  INV_X1 U13053 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17515) );
  NOR2_X2 U13054 ( .A1(n17036), .A2(n16948), .ZN(n16927) );
  NOR2_X1 U13055 ( .A1(n15407), .A2(n15406), .ZN(n17075) );
  OR2_X1 U13056 ( .A1(n18426), .A2(n17574), .ZN(n18570) );
  INV_X1 U13057 ( .A(n17132), .ZN(n17162) );
  INV_X1 U13058 ( .A(n17484), .ZN(n17458) );
  INV_X1 U13059 ( .A(n16014), .ZN(n17577) );
  OAI21_X2 U13060 ( .B1(n15530), .B2(n15529), .A(n18569), .ZN(n17886) );
  INV_X1 U13061 ( .A(n17834), .ZN(n17898) );
  INV_X1 U13062 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18166) );
  INV_X1 U13063 ( .A(n18113), .ZN(n18105) );
  INV_X1 U13064 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n20659) );
  INV_X1 U13065 ( .A(n18185), .ZN(n18177) );
  INV_X1 U13066 ( .A(n18210), .ZN(n18202) );
  INV_X1 U13067 ( .A(n18318), .ZN(n18281) );
  INV_X1 U13068 ( .A(n18347), .ZN(n18315) );
  INV_X1 U13069 ( .A(n18569), .ZN(n18422) );
  INV_X1 U13070 ( .A(n16531), .ZN(n18432) );
  INV_X1 U13071 ( .A(n18517), .ZN(n18436) );
  OAI211_X1 U13072 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18449), .B(n18513), .ZN(n18574) );
  INV_X2 U13073 ( .A(n18585), .ZN(n18584) );
  NOR2_X1 U13074 ( .A1(n14847), .A2(n12544), .ZN(n16085) );
  NOR2_X1 U13075 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12544), .ZN(n16156)
         );
  INV_X1 U13076 ( .A(n16126), .ZN(n16131) );
  INV_X1 U13077 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19643) );
  OR4_X1 U13078 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        P2_U2854) );
  AND2_X4 U13079 ( .A1(n13205), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12353) );
  AND2_X4 U13080 ( .A1(n10341), .A2(n15352), .ZN(n12461) );
  AOI22_X1 U13081 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10139) );
  NOR2_X2 U13082 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10134) );
  AND2_X2 U13083 ( .A1(n10134), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10344) );
  BUF_X4 U13084 ( .A(n10344), .Z(n10208) );
  AND3_X4 U13085 ( .A1(n10329), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12485) );
  AOI22_X1 U13086 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10138) );
  AND2_X4 U13087 ( .A1(n10581), .A2(n10135), .ZN(n12479) );
  AOI22_X1 U13088 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10137) );
  AND2_X4 U13089 ( .A1(n10343), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12484) );
  AND2_X4 U13090 ( .A1(n13205), .A2(n10135), .ZN(n10328) );
  AOI22_X1 U13091 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U13092 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U13093 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10142) );
  AOI22_X1 U13094 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U13095 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U13096 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U13097 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13098 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U13099 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10144) );
  AOI22_X1 U13100 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13101 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U13102 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13103 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10148) );
  NAND2_X2 U13104 ( .A1(n10719), .A2(n12509), .ZN(n10234) );
  AOI22_X1 U13105 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12353), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U13106 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13107 ( .A1(n10328), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U13108 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10152) );
  NAND4_X1 U13109 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10156) );
  AOI22_X1 U13110 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13111 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13112 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13113 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10157) );
  NAND4_X1 U13114 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(
        n10161) );
  NAND2_X1 U13115 ( .A1(n10161), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10162) );
  AOI22_X1 U13116 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U13117 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U13118 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13119 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U13120 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U13121 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13122 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13123 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U13124 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13125 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U13126 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U13127 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10172) );
  NAND4_X1 U13128 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10181) );
  AOI22_X1 U13129 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13130 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10178) );
  AOI22_X1 U13131 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U13132 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10176) );
  NAND4_X1 U13133 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10180) );
  MUX2_X2 U13134 ( .A(n10181), .B(n10180), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10227) );
  NAND4_X2 U13135 ( .A1(n10720), .A2(n19023), .A3(n12508), .A4(n19033), .ZN(
        n10988) );
  AOI22_X1 U13136 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13137 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13138 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U13139 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10182) );
  NAND4_X1 U13140 ( .A1(n10185), .A2(n10184), .A3(n10183), .A4(n10182), .ZN(
        n10186) );
  NAND2_X1 U13141 ( .A1(n10186), .A2(n13211), .ZN(n10193) );
  AOI22_X1 U13142 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13143 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U13144 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13145 ( .A1(n10208), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10187) );
  NAND4_X1 U13146 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10191) );
  NAND2_X1 U13147 ( .A1(n10191), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10192) );
  INV_X2 U13148 ( .A(n13238), .ZN(n13457) );
  MUX2_X1 U13149 ( .A(n19033), .B(n10227), .S(n10977), .Z(n10212) );
  AOI22_X1 U13150 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U13151 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13152 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13153 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10195) );
  NAND4_X1 U13154 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10199) );
  AOI22_X1 U13155 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U13156 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13157 ( .A1(n12353), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13158 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10200) );
  NAND4_X1 U13159 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10204) );
  AOI22_X1 U13160 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13161 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10206) );
  AOI22_X1 U13162 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10328), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U13163 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10209) );
  NAND2_X1 U13164 ( .A1(n10234), .A2(n19016), .ZN(n10211) );
  NAND4_X1 U13165 ( .A1(n10212), .A2(n10943), .A3(n10938), .A4(n10211), .ZN(
        n10213) );
  NAND3_X1 U13166 ( .A1(n10213), .A2(n13457), .A3(n10220), .ZN(n10980) );
  INV_X1 U13167 ( .A(n10214), .ZN(n10222) );
  NOR2_X1 U13168 ( .A1(n10214), .A2(n19010), .ZN(n10215) );
  NAND2_X1 U13169 ( .A1(n9618), .A2(n10215), .ZN(n10585) );
  NAND3_X1 U13170 ( .A1(n10585), .A2(n10943), .A3(n11021), .ZN(n10216) );
  NAND3_X1 U13171 ( .A1(n10937), .A2(n19023), .A3(n10938), .ZN(n10934) );
  NAND3_X1 U13172 ( .A1(n10934), .A2(n10944), .A3(n19044), .ZN(n10975) );
  NAND2_X1 U13173 ( .A1(n12504), .A2(n10241), .ZN(n10219) );
  NAND2_X1 U13174 ( .A1(n10265), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10226) );
  AND3_X1 U13175 ( .A1(n10223), .A2(n10222), .A3(n10221), .ZN(n10932) );
  NAND2_X1 U13176 ( .A1(n10932), .A2(n13238), .ZN(n13272) );
  NAND2_X1 U13177 ( .A1(n12614), .A2(n13272), .ZN(n11215) );
  NAND2_X1 U13178 ( .A1(n11023), .A2(n13238), .ZN(n10939) );
  AND2_X1 U13179 ( .A1(n19023), .A2(n19044), .ZN(n10230) );
  NOR2_X1 U13180 ( .A1(n10943), .A2(n13238), .ZN(n10229) );
  NAND4_X1 U13181 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10238), .ZN(
        n10231) );
  NOR2_X1 U13182 ( .A1(n10125), .A2(n10232), .ZN(n10239) );
  NOR2_X1 U13183 ( .A1(n10937), .A2(n11021), .ZN(n10235) );
  MUX2_X1 U13184 ( .A(n10235), .B(n11041), .S(n19016), .Z(n10236) );
  NAND2_X2 U13185 ( .A1(n10971), .A2(n10987), .ZN(n13202) );
  NAND2_X1 U13186 ( .A1(n10272), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10247) );
  NAND2_X4 U13187 ( .A1(n10242), .A2(n10241), .ZN(n10685) );
  NOR2_X1 U13188 ( .A1(n10988), .A2(n11023), .ZN(n10243) );
  AND2_X1 U13189 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10244) );
  NAND2_X1 U13190 ( .A1(n10247), .A2(n10246), .ZN(n10263) );
  INV_X1 U13191 ( .A(n13202), .ZN(n10249) );
  AOI22_X1 U13192 ( .A1(n10249), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12587), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U13193 ( .A1(n10251), .A2(n10250), .ZN(n10281) );
  NAND3_X1 U13194 ( .A1(n12504), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10983), 
        .ZN(n10258) );
  INV_X1 U13195 ( .A(n12587), .ZN(n10253) );
  NAND2_X1 U13196 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10252) );
  NAND2_X1 U13197 ( .A1(n10253), .A2(n10252), .ZN(n10254) );
  AOI21_X1 U13198 ( .B1(n10663), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10254), .ZN(
        n10257) );
  INV_X1 U13199 ( .A(n10685), .ZN(n10255) );
  AND2_X2 U13200 ( .A1(n10281), .A2(n10282), .ZN(n10280) );
  OR2_X1 U13201 ( .A1(n10263), .A2(n10262), .ZN(n10264) );
  OAI21_X2 U13202 ( .B1(n10284), .B2(n10280), .A(n10264), .ZN(n10271) );
  INV_X1 U13203 ( .A(n10271), .ZN(n10268) );
  NAND2_X1 U13204 ( .A1(n10265), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10267) );
  AOI21_X1 U13205 ( .B1(n18596), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U13206 ( .A1(n10267), .A2(n10266), .ZN(n10269) );
  NAND2_X1 U13207 ( .A1(n10268), .A2(n10269), .ZN(n10287) );
  INV_X1 U13208 ( .A(n10269), .ZN(n10270) );
  NAND2_X1 U13209 ( .A1(n10271), .A2(n10270), .ZN(n10288) );
  NAND2_X1 U13210 ( .A1(n10287), .A2(n10288), .ZN(n10279) );
  INV_X1 U13211 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10276) );
  CLKBUF_X3 U13212 ( .A(n10663), .Z(n10679) );
  NAND2_X1 U13213 ( .A1(n10679), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U13214 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10274) );
  OAI211_X1 U13215 ( .C1(n10685), .C2(n10276), .A(n10275), .B(n10274), .ZN(
        n10277) );
  INV_X1 U13216 ( .A(n10280), .ZN(n10309) );
  OR2_X1 U13217 ( .A1(n10282), .A2(n10281), .ZN(n10283) );
  INV_X1 U13218 ( .A(n12202), .ZN(n18832) );
  INV_X1 U13219 ( .A(n10308), .ZN(n10285) );
  NAND2_X1 U13220 ( .A1(n10287), .A2(n10286), .ZN(n10289) );
  NAND2_X1 U13221 ( .A1(n9601), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10295) );
  INV_X1 U13222 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10292) );
  NAND2_X1 U13223 ( .A1(n10679), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U13224 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10290) );
  OAI211_X1 U13225 ( .C1(n10685), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        n10293) );
  INV_X1 U13226 ( .A(n10293), .ZN(n10294) );
  NAND2_X1 U13227 ( .A1(n10265), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U13228 ( .A1(n12587), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10296) );
  AND2_X1 U13229 ( .A1(n10308), .A2(n18832), .ZN(n10300) );
  AOI22_X1 U13230 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19370), .B1(
        n19314), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13232 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n13490), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13233 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19179), .B1(
        n19240), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13234 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13454), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10303) );
  AND4_X1 U13235 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10326) );
  NAND2_X1 U13236 ( .A1(n12195), .A2(n12202), .ZN(n10314) );
  INV_X1 U13237 ( .A(n10314), .ZN(n10307) );
  NAND2_X1 U13238 ( .A1(n10307), .A2(n12729), .ZN(n10310) );
  AOI22_X1 U13239 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19084), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10325) );
  INV_X1 U13240 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10312) );
  NAND2_X1 U13241 ( .A1(n18983), .A2(n10321), .ZN(n10315) );
  NAND2_X1 U13242 ( .A1(n18983), .A2(n9592), .ZN(n10313) );
  INV_X1 U13243 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10311) );
  OAI22_X1 U13244 ( .A1(n10312), .A2(n19211), .B1(n19417), .B2(n10311), .ZN(
        n10319) );
  INV_X1 U13245 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10317) );
  INV_X1 U13246 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10316) );
  OAI22_X1 U13247 ( .A1(n10317), .A2(n19137), .B1(n19489), .B2(n10316), .ZN(
        n10318) );
  NOR2_X1 U13248 ( .A1(n10319), .A2(n10318), .ZN(n10324) );
  NOR2_X2 U13249 ( .A1(n10322), .A2(n9592), .ZN(n19339) );
  NOR2_X2 U13250 ( .A1(n10322), .A2(n10321), .ZN(n10473) );
  AOI22_X1 U13251 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19339), .B1(
        n10473), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10323) );
  NAND4_X1 U13252 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10327) );
  NAND2_X1 U13253 ( .A1(n10327), .A2(n19006), .ZN(n10352) );
  AND2_X2 U13254 ( .A1(n12486), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10428) );
  AOI22_X1 U13255 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10340) );
  AND2_X1 U13256 ( .A1(n10330), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10331) );
  AND2_X2 U13257 ( .A1(n12315), .A2(n10331), .ZN(n12333) );
  NOR2_X1 U13258 ( .A1(n10330), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10332) );
  AOI22_X1 U13259 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10334) );
  AND2_X2 U13260 ( .A1(n12484), .A2(n13211), .ZN(n12331) );
  NAND2_X1 U13261 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10333) );
  AND2_X1 U13262 ( .A1(n10334), .A2(n10333), .ZN(n10339) );
  AND2_X2 U13263 ( .A1(n12353), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10511) );
  AOI22_X1 U13265 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13266 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10337) );
  NAND4_X1 U13267 ( .A1(n10340), .A2(n10339), .A3(n10338), .A4(n10337), .ZN(
        n10350) );
  AND2_X2 U13268 ( .A1(n12489), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10382) );
  AND2_X2 U13269 ( .A1(n12489), .A2(n13211), .ZN(n12340) );
  AOI22_X1 U13270 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10348) );
  AND2_X2 U13271 ( .A1(n12485), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10436) );
  AOI22_X1 U13272 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10347) );
  AND2_X2 U13273 ( .A1(n12315), .A2(n10342), .ZN(n12343) );
  AOI22_X1 U13274 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10346) );
  NAND2_X1 U13275 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10345) );
  NAND4_X1 U13276 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10349) );
  INV_X1 U13277 ( .A(n10419), .ZN(n10417) );
  AOI22_X1 U13278 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19179), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13279 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n13490), .B1(
        n19314), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13280 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19240), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U13281 ( .A1(n19414), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10355) );
  INV_X1 U13282 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10361) );
  AOI21_X1 U13283 ( .B1(n19370), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n9600), .ZN(n10360) );
  NAND2_X1 U13284 ( .A1(n13454), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10359) );
  OAI211_X1 U13285 ( .C1(n19137), .C2(n10361), .A(n10360), .B(n10359), .ZN(
        n10362) );
  AOI21_X1 U13286 ( .B1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n19339), .A(
        n10362), .ZN(n10368) );
  AOI22_X1 U13287 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10496), .B1(
        n10473), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10367) );
  INV_X1 U13288 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10364) );
  INV_X1 U13289 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10363) );
  OAI22_X1 U13290 ( .A1(n10364), .A2(n19211), .B1(n19489), .B2(n10363), .ZN(
        n10365) );
  AOI21_X1 U13291 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n19084), .A(
        n10365), .ZN(n10366) );
  NAND4_X1 U13292 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10415) );
  AOI22_X1 U13293 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n10388), .B1(
        n10428), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U13294 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n12333), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10371) );
  NAND2_X1 U13295 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10370) );
  AND2_X1 U13296 ( .A1(n10371), .A2(n10370), .ZN(n10374) );
  AOI22_X1 U13297 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13298 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10482), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10372) );
  NAND4_X1 U13299 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        n10381) );
  AOI22_X1 U13300 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12340), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10379) );
  INV_X1 U13301 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19501) );
  AOI22_X1 U13302 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12341), .B1(
        n10436), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13303 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12343), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10377) );
  NAND2_X1 U13304 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10376) );
  NAND4_X1 U13305 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10380) );
  AND2_X1 U13306 ( .A1(n12418), .A2(n11032), .ZN(n10421) );
  AOI22_X1 U13307 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12340), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13308 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12341), .B1(
        n10436), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13309 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12343), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U13310 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10384) );
  AND4_X1 U13311 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n10397) );
  AOI22_X1 U13312 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12333), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U13313 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10391) );
  NAND2_X1 U13314 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10390) );
  NAND2_X1 U13315 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10389) );
  NAND4_X1 U13316 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10396) );
  NAND2_X1 U13317 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10395) );
  NAND2_X1 U13318 ( .A1(n10431), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10394) );
  NAND2_X1 U13319 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10393) );
  INV_X1 U13320 ( .A(n10727), .ZN(n11037) );
  NAND2_X1 U13321 ( .A1(n10421), .A2(n11037), .ZN(n10420) );
  AOI22_X1 U13322 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10382), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13323 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10383), .B1(
        n10436), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13324 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12343), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U13325 ( .A1(n12341), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10398) );
  AND4_X1 U13326 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10413) );
  AOI22_X1 U13327 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12333), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U13328 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13329 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U13330 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10402) );
  NAND4_X1 U13331 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10411) );
  NAND2_X1 U13332 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10409) );
  NAND2_X1 U13333 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10408) );
  NAND2_X1 U13334 ( .A1(n10431), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10407) );
  NAND2_X1 U13335 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10406) );
  NAND4_X1 U13336 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10410) );
  NOR2_X1 U13337 ( .A1(n10411), .A2(n10410), .ZN(n10412) );
  NAND2_X1 U13338 ( .A1(n10420), .A2(n11048), .ZN(n10414) );
  INV_X1 U13339 ( .A(n10418), .ZN(n10416) );
  XOR2_X1 U13340 ( .A(n11048), .B(n10420), .Z(n12690) );
  INV_X1 U13341 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18990) );
  OR2_X1 U13342 ( .A1(n10421), .A2(n15336), .ZN(n12667) );
  XOR2_X1 U13343 ( .A(n11032), .B(n10727), .Z(n10422) );
  NOR2_X1 U13344 ( .A1(n12667), .A2(n10422), .ZN(n10423) );
  INV_X1 U13345 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15340) );
  XNOR2_X1 U13346 ( .A(n12667), .B(n10422), .ZN(n12676) );
  NOR2_X1 U13347 ( .A1(n15340), .A2(n12676), .ZN(n12675) );
  NOR2_X1 U13348 ( .A1(n10423), .A2(n12675), .ZN(n10424) );
  XNOR2_X1 U13349 ( .A(n18990), .B(n10424), .ZN(n12689) );
  NOR2_X1 U13350 ( .A1(n12690), .A2(n12689), .ZN(n12688) );
  NOR2_X1 U13351 ( .A1(n10424), .A2(n18990), .ZN(n10425) );
  OR2_X1 U13352 ( .A1(n12688), .A2(n10425), .ZN(n10426) );
  INV_X1 U13353 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13402) );
  XNOR2_X1 U13354 ( .A(n10426), .B(n13402), .ZN(n13396) );
  NAND2_X1 U13355 ( .A1(n10426), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10427) );
  AOI22_X1 U13356 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13357 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U13358 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10429) );
  AND2_X1 U13359 ( .A1(n10430), .A2(n10429), .ZN(n10434) );
  AOI22_X1 U13360 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13361 ( .A1(n10431), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10432) );
  NAND4_X1 U13362 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10442) );
  AOI22_X1 U13363 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10440) );
  AOI22_X1 U13364 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13365 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U13366 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10437) );
  NAND4_X1 U13367 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10441) );
  NAND2_X1 U13368 ( .A1(n10444), .A2(n10443), .ZN(n10445) );
  INV_X1 U13369 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20652) );
  INV_X1 U13370 ( .A(n10446), .ZN(n10448) );
  NAND2_X1 U13371 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  INV_X1 U13372 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10453) );
  INV_X1 U13373 ( .A(n19370), .ZN(n10452) );
  INV_X1 U13374 ( .A(n10353), .ZN(n10451) );
  INV_X1 U13375 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10450) );
  OAI22_X1 U13376 ( .A1(n10453), .A2(n10452), .B1(n10451), .B2(n10450), .ZN(
        n10459) );
  INV_X1 U13377 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10457) );
  INV_X1 U13378 ( .A(n13454), .ZN(n10456) );
  INV_X1 U13379 ( .A(n13490), .ZN(n10455) );
  INV_X1 U13380 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10454) );
  OAI22_X1 U13381 ( .A1(n10457), .A2(n10456), .B1(n10455), .B2(n10454), .ZN(
        n10458) );
  NOR2_X1 U13382 ( .A1(n10459), .A2(n10458), .ZN(n10471) );
  INV_X1 U13383 ( .A(n19211), .ZN(n19209) );
  AOI22_X1 U13384 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19209), .B1(
        n19414), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10470) );
  INV_X1 U13385 ( .A(n19137), .ZN(n19145) );
  INV_X1 U13386 ( .A(n19489), .ZN(n19495) );
  AOI22_X1 U13387 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19145), .B1(
        n19495), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10469) );
  INV_X1 U13388 ( .A(n10354), .ZN(n10461) );
  INV_X1 U13389 ( .A(n19314), .ZN(n19311) );
  INV_X1 U13390 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10460) );
  OAI22_X1 U13391 ( .A1(n20661), .A2(n10461), .B1(n19311), .B2(n10460), .ZN(
        n10467) );
  INV_X1 U13392 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10465) );
  INV_X1 U13393 ( .A(n19179), .ZN(n10464) );
  INV_X1 U13394 ( .A(n19240), .ZN(n10463) );
  INV_X1 U13395 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10462) );
  OAI22_X1 U13396 ( .A1(n10465), .A2(n10464), .B1(n10463), .B2(n10462), .ZN(
        n10466) );
  NOR2_X1 U13397 ( .A1(n10467), .A2(n10466), .ZN(n10468) );
  NAND4_X1 U13398 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n10479) );
  INV_X1 U13399 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10472) );
  INV_X1 U13400 ( .A(n19084), .ZN(n19087) );
  INV_X1 U13401 ( .A(n10496), .ZN(n18998) );
  INV_X1 U13402 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12967) );
  OAI22_X1 U13403 ( .A1(n10472), .A2(n19087), .B1(n18998), .B2(n12967), .ZN(
        n10478) );
  INV_X1 U13404 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10476) );
  INV_X1 U13405 ( .A(n19339), .ZN(n19343) );
  INV_X1 U13406 ( .A(n10473), .ZN(n10475) );
  INV_X1 U13407 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10474) );
  OAI22_X1 U13408 ( .A1(n10476), .A2(n19343), .B1(n10475), .B2(n10474), .ZN(
        n10477) );
  AOI22_X1 U13409 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13410 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U13411 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10480) );
  AND2_X1 U13412 ( .A1(n10481), .A2(n10480), .ZN(n10485) );
  AOI22_X1 U13413 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13414 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10483) );
  NAND4_X1 U13415 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10492) );
  AOI22_X1 U13416 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13417 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13418 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U13419 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10487) );
  NAND4_X1 U13420 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10491) );
  NOR2_X1 U13421 ( .A1(n10492), .A2(n10491), .ZN(n11064) );
  NAND2_X1 U13422 ( .A1(n11064), .A2(n12418), .ZN(n10493) );
  INV_X1 U13423 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10739) );
  AND2_X1 U13424 ( .A1(n10494), .A2(n10739), .ZN(n13616) );
  NAND2_X1 U13425 ( .A1(n10718), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13614) );
  NAND2_X1 U13426 ( .A1(n13619), .A2(n13614), .ZN(n10531) );
  AOI22_X1 U13427 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19084), .B1(
        n10496), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13428 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19339), .B1(
        n10473), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13429 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19370), .B1(
        n19314), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13430 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n13490), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13431 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19179), .B1(
        n19240), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13432 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13454), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10497) );
  INV_X1 U13433 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10502) );
  INV_X1 U13434 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10501) );
  OAI22_X1 U13435 ( .A1(n10502), .A2(n19211), .B1(n19417), .B2(n10501), .ZN(
        n10506) );
  INV_X1 U13436 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10504) );
  INV_X1 U13437 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10503) );
  OAI22_X1 U13438 ( .A1(n10504), .A2(n19137), .B1(n19489), .B2(n10503), .ZN(
        n10505) );
  NOR2_X1 U13439 ( .A1(n10506), .A2(n10505), .ZN(n10507) );
  NAND4_X1 U13440 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10526) );
  AOI22_X1 U13441 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12331), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13442 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10513) );
  NAND2_X1 U13443 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10512) );
  AND2_X1 U13444 ( .A1(n10513), .A2(n10512), .ZN(n10516) );
  AOI22_X1 U13445 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13446 ( .A1(n10431), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10514) );
  NAND4_X1 U13447 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10523) );
  AOI22_X1 U13448 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13449 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13450 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10519) );
  NAND2_X1 U13451 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10518) );
  NAND4_X1 U13452 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10522) );
  INV_X1 U13453 ( .A(n11069), .ZN(n10524) );
  NAND2_X1 U13454 ( .A1(n10524), .A2(n9600), .ZN(n10525) );
  XNOR2_X1 U13455 ( .A(n10534), .B(n10535), .ZN(n10762) );
  INV_X1 U13456 ( .A(n13619), .ZN(n10528) );
  AOI21_X1 U13457 ( .B1(n10528), .B2(n10530), .A(n10527), .ZN(n10529) );
  OAI21_X2 U13458 ( .B1(n10531), .B2(n10530), .A(n10529), .ZN(n13695) );
  NAND2_X1 U13459 ( .A1(n10531), .A2(n10762), .ZN(n10532) );
  INV_X1 U13460 ( .A(n10534), .ZN(n10536) );
  AOI22_X1 U13461 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13462 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13463 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U13464 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10537) );
  AOI22_X1 U13465 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U13466 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10543) );
  NAND2_X1 U13467 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10542) );
  NAND2_X1 U13468 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10541) );
  NAND4_X1 U13469 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10550) );
  NAND2_X1 U13470 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10548) );
  NAND2_X1 U13471 ( .A1(n10431), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10547) );
  NAND2_X1 U13472 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10546) );
  NAND2_X1 U13473 ( .A1(n13224), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10545) );
  NAND4_X1 U13474 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n10549) );
  NOR2_X1 U13475 ( .A1(n10550), .A2(n10549), .ZN(n10551) );
  INV_X1 U13476 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15328) );
  NAND2_X1 U13477 ( .A1(n15058), .A2(n15328), .ZN(n10553) );
  INV_X1 U13478 ( .A(n15058), .ZN(n10554) );
  NAND2_X1 U13479 ( .A1(n10554), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10555) );
  INV_X1 U13480 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11079) );
  OR2_X1 U13481 ( .A1(n10865), .A2(n11079), .ZN(n10773) );
  INV_X1 U13482 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15972) );
  INV_X1 U13483 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15280) );
  NOR2_X1 U13484 ( .A1(n10786), .A2(n15280), .ZN(n15266) );
  NAND2_X1 U13485 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15266), .ZN(
        n15269) );
  NOR2_X1 U13486 ( .A1(n15972), .A2(n15269), .ZN(n15050) );
  NAND2_X1 U13487 ( .A1(n15050), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15958) );
  INV_X1 U13488 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15898) );
  NOR2_X1 U13489 ( .A1(n15958), .A2(n15898), .ZN(n15162) );
  AND2_X1 U13490 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15222) );
  NAND2_X1 U13491 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10559) );
  INV_X1 U13492 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15183) );
  INV_X1 U13493 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14967) );
  NAND2_X1 U13494 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15137) );
  INV_X1 U13495 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15118) );
  AND2_X1 U13496 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15072) );
  NAND2_X1 U13497 ( .A1(n15072), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11298) );
  NAND2_X1 U13498 ( .A1(n10930), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10560) );
  XNOR2_X1 U13499 ( .A(n10560), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11302) );
  OAI21_X1 U13500 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19720), .A(
        n10578), .ZN(n10697) );
  INV_X1 U13501 ( .A(n10697), .ZN(n10744) );
  MUX2_X1 U13502 ( .A(n10562), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10586) );
  INV_X1 U13503 ( .A(n10578), .ZN(n10561) );
  NAND2_X1 U13504 ( .A1(n10586), .A2(n10561), .ZN(n10564) );
  NAND2_X1 U13505 ( .A1(n10562), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10563) );
  NAND2_X1 U13506 ( .A1(n10564), .A2(n10563), .ZN(n10573) );
  MUX2_X1 U13507 ( .A(n12211), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10571) );
  NAND2_X1 U13508 ( .A1(n10573), .A2(n10571), .ZN(n10566) );
  NAND2_X1 U13509 ( .A1(n12211), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10565) );
  MUX2_X1 U13510 ( .A(n13264), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10568) );
  NOR2_X1 U13511 ( .A1(n13211), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10567) );
  NOR2_X1 U13512 ( .A1(n20684), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10574) );
  NAND2_X1 U13513 ( .A1(n10575), .A2(n10574), .ZN(n10732) );
  INV_X1 U13514 ( .A(n10568), .ZN(n10569) );
  XNOR2_X1 U13515 ( .A(n10570), .B(n10569), .ZN(n10722) );
  INV_X1 U13516 ( .A(n10571), .ZN(n10572) );
  XNOR2_X1 U13517 ( .A(n10573), .B(n10572), .ZN(n10692) );
  AND2_X1 U13518 ( .A1(n10704), .A2(n10692), .ZN(n10580) );
  NAND2_X1 U13519 ( .A1(n20684), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10576) );
  XNOR2_X1 U13520 ( .A(n10586), .B(n10578), .ZN(n10695) );
  NAND2_X1 U13521 ( .A1(n10695), .A2(n10580), .ZN(n10579) );
  NAND2_X1 U13522 ( .A1(n19726), .A2(n10579), .ZN(n13232) );
  AOI211_X1 U13523 ( .C1(n10744), .C2(n10580), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n13232), .ZN(n10584) );
  NAND2_X1 U13524 ( .A1(n13216), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10582) );
  NAND2_X1 U13525 ( .A1(n10582), .A2(n12220), .ZN(n13240) );
  INV_X1 U13526 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12611) );
  OAI21_X1 U13527 ( .B1(n10436), .B2(n13240), .A(n12611), .ZN(n10583) );
  AND2_X1 U13528 ( .A1(n10583), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19717) );
  NOR2_X1 U13529 ( .A1(n10585), .A2(n10721), .ZN(n19728) );
  NAND2_X1 U13530 ( .A1(n15631), .A2(n19728), .ZN(n10588) );
  NOR2_X1 U13531 ( .A1(n10585), .A2(n10939), .ZN(n10960) );
  NAND2_X1 U13532 ( .A1(n10721), .A2(n10692), .ZN(n10693) );
  OAI21_X1 U13533 ( .B1(n10721), .B2(n11048), .A(n10693), .ZN(n10729) );
  OR2_X1 U13534 ( .A1(n10729), .A2(n10122), .ZN(n10587) );
  NAND2_X1 U13535 ( .A1(n10587), .A2(n10704), .ZN(n19725) );
  NAND3_X1 U13536 ( .A1(n10960), .A2(n19726), .A3(n19725), .ZN(n10953) );
  NAND2_X1 U13537 ( .A1(n10588), .A2(n10953), .ZN(n10589) );
  NAND2_X1 U13538 ( .A1(n10711), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11283) );
  INV_X1 U13539 ( .A(n12586), .ZN(n10590) );
  NOR2_X1 U13540 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15342) );
  OR2_X1 U13541 ( .A1(n19688), .A2(n15342), .ZN(n19713) );
  NAND2_X1 U13542 ( .A1(n19713), .A2(n18596), .ZN(n10591) );
  INV_X1 U13543 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n18993) );
  NAND2_X1 U13544 ( .A1(n18993), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U13545 ( .A1(n12209), .A2(n10592), .ZN(n12672) );
  INV_X1 U13546 ( .A(n11261), .ZN(n10594) );
  NAND2_X1 U13547 ( .A1(n10594), .A2(n10593), .ZN(n11259) );
  NAND2_X1 U13548 ( .A1(n11260), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11256) );
  NAND2_X1 U13549 ( .A1(n11251), .A2(n10595), .ZN(n11252) );
  NAND2_X1 U13550 ( .A1(n11242), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11240) );
  NAND2_X1 U13551 ( .A1(n11238), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11236) );
  INV_X1 U13552 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10598) );
  INV_X1 U13553 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U13554 ( .A1(n10273), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10605) );
  INV_X1 U13555 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U13556 ( .A1(n10679), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13557 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10600) );
  OAI211_X1 U13558 ( .C1(n10685), .C2(n10602), .A(n10601), .B(n10600), .ZN(
        n10603) );
  INV_X1 U13559 ( .A(n10603), .ZN(n10604) );
  NAND2_X1 U13560 ( .A1(n10605), .A2(n10604), .ZN(n13195) );
  INV_X1 U13561 ( .A(n10606), .ZN(n10610) );
  NOR2_X1 U13562 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  INV_X1 U13563 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10613) );
  NAND2_X1 U13564 ( .A1(n10273), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10612) );
  AOI22_X1 U13565 ( .A1(n10679), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10611) );
  OAI211_X1 U13566 ( .C1(n10685), .C2(n10613), .A(n10612), .B(n10611), .ZN(
        n13538) );
  INV_X1 U13567 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13626) );
  NAND2_X1 U13568 ( .A1(n10273), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10615) );
  AOI22_X1 U13569 ( .A1(n10663), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10614) );
  OAI211_X1 U13570 ( .C1(n10685), .C2(n13626), .A(n10615), .B(n10614), .ZN(
        n12858) );
  INV_X1 U13571 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10618) );
  NAND2_X1 U13572 ( .A1(n10679), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13573 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10616) );
  OAI211_X1 U13574 ( .C1(n10685), .C2(n10618), .A(n10617), .B(n10616), .ZN(
        n10619) );
  AOI21_X1 U13575 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10619), .ZN(n12970) );
  INV_X1 U13576 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10622) );
  NAND2_X1 U13577 ( .A1(n10679), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U13578 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10620) );
  OAI211_X1 U13579 ( .C1(n10685), .C2(n10622), .A(n10621), .B(n10620), .ZN(
        n10623) );
  AOI21_X1 U13580 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10623), .ZN(n12962) );
  INV_X1 U13581 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11092) );
  NAND2_X1 U13582 ( .A1(n10679), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U13583 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10624) );
  OAI211_X1 U13584 ( .C1(n10685), .C2(n11092), .A(n10625), .B(n10624), .ZN(
        n10626) );
  AOI21_X1 U13585 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10626), .ZN(n13007) );
  NOR2_X2 U13586 ( .A1(n13008), .A2(n13007), .ZN(n13009) );
  INV_X1 U13587 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15320) );
  NAND2_X1 U13588 ( .A1(n10273), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10628) );
  AOI22_X1 U13589 ( .A1(n10679), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10627) );
  OAI211_X1 U13590 ( .C1(n10685), .C2(n15320), .A(n10628), .B(n10627), .ZN(
        n12849) );
  NAND2_X1 U13591 ( .A1(n13009), .A2(n12849), .ZN(n12953) );
  INV_X1 U13592 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10631) );
  NAND2_X1 U13593 ( .A1(n10679), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10630) );
  NAND2_X1 U13594 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10629) );
  OAI211_X1 U13595 ( .C1(n10685), .C2(n10631), .A(n10630), .B(n10629), .ZN(
        n10632) );
  AOI21_X1 U13596 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10632), .ZN(n12954) );
  NOR2_X2 U13597 ( .A1(n12953), .A2(n12954), .ZN(n13066) );
  INV_X1 U13598 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U13599 ( .A1(n10273), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10634) );
  AOI22_X1 U13600 ( .A1(n10663), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10633) );
  OAI211_X1 U13601 ( .C1(n10685), .C2(n10635), .A(n10634), .B(n10633), .ZN(
        n13067) );
  NAND2_X1 U13602 ( .A1(n13066), .A2(n13067), .ZN(n13068) );
  INV_X1 U13603 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11151) );
  AOI22_X1 U13604 ( .A1(n10679), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10636) );
  OAI21_X1 U13605 ( .B1(n10685), .B2(n11151), .A(n10636), .ZN(n10637) );
  AOI21_X1 U13606 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10637), .ZN(n13141) );
  NOR2_X2 U13607 ( .A1(n13068), .A2(n13141), .ZN(n13194) );
  NAND2_X1 U13608 ( .A1(n13195), .A2(n13194), .ZN(n13380) );
  INV_X1 U13609 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U13610 ( .A1(n10679), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10639) );
  NAND2_X1 U13611 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10638) );
  OAI211_X1 U13612 ( .C1(n10685), .C2(n11025), .A(n10639), .B(n10638), .ZN(
        n10640) );
  AOI21_X1 U13613 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10640), .ZN(n13379) );
  OR2_X2 U13614 ( .A1(n13380), .A2(n13379), .ZN(n13567) );
  INV_X1 U13615 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15042) );
  NAND2_X1 U13616 ( .A1(n10679), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13617 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10641) );
  OAI211_X1 U13618 ( .C1(n10685), .C2(n15042), .A(n10642), .B(n10641), .ZN(
        n10643) );
  AOI21_X1 U13619 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10643), .ZN(n13566) );
  INV_X1 U13620 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13621 ( .A1(n10679), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10646) );
  NAND2_X1 U13622 ( .A1(n10644), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10645) );
  OAI211_X1 U13623 ( .C1(n10689), .C2(n10842), .A(n10646), .B(n10645), .ZN(
        n15027) );
  INV_X1 U13624 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19656) );
  NAND2_X1 U13625 ( .A1(n10663), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10648) );
  NAND2_X1 U13626 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10647) );
  OAI211_X1 U13627 ( .C1(n10685), .C2(n19656), .A(n10648), .B(n10647), .ZN(
        n10649) );
  AOI21_X1 U13628 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10649), .ZN(n13691) );
  INV_X1 U13629 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19658) );
  NAND2_X1 U13630 ( .A1(n10679), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10651) );
  NAND2_X1 U13631 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10650) );
  OAI211_X1 U13632 ( .C1(n10685), .C2(n19658), .A(n10651), .B(n10650), .ZN(
        n10652) );
  AOI21_X1 U13633 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10652), .ZN(n15003) );
  NOR2_X2 U13634 ( .A1(n15004), .A2(n15003), .ZN(n14780) );
  INV_X1 U13635 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U13636 ( .A1(n10679), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10654) );
  INV_X1 U13637 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19660) );
  OR2_X1 U13638 ( .A1(n10685), .A2(n19660), .ZN(n10653) );
  OAI211_X1 U13639 ( .C1(n10689), .C2(n15195), .A(n10654), .B(n10653), .ZN(
        n14781) );
  AOI22_X1 U13640 ( .A1(n10679), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10656) );
  INV_X1 U13641 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19661) );
  OR2_X1 U13642 ( .A1(n10685), .A2(n19661), .ZN(n10655) );
  OAI211_X1 U13643 ( .C1(n10689), .C2(n15183), .A(n10656), .B(n10655), .ZN(
        n14980) );
  INV_X1 U13644 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20723) );
  NAND2_X1 U13645 ( .A1(n10679), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U13646 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10657) );
  OAI211_X1 U13647 ( .C1(n10685), .C2(n20723), .A(n10658), .B(n10657), .ZN(
        n10659) );
  AOI21_X1 U13648 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10659), .ZN(n12563) );
  INV_X1 U13649 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n14942) );
  NAND2_X1 U13650 ( .A1(n10679), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10661) );
  NAND2_X1 U13651 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10660) );
  OAI211_X1 U13652 ( .C1(n10685), .C2(n14942), .A(n10661), .B(n10660), .ZN(
        n10662) );
  AOI21_X1 U13653 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10662), .ZN(n14938) );
  INV_X1 U13654 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19665) );
  NAND2_X1 U13655 ( .A1(n10663), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13656 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10664) );
  OAI211_X1 U13657 ( .C1(n10685), .C2(n19665), .A(n10665), .B(n10664), .ZN(
        n10666) );
  AOI21_X1 U13658 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10666), .ZN(n12573) );
  INV_X1 U13659 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U13660 ( .A1(n10679), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10668) );
  INV_X1 U13661 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19667) );
  OR2_X1 U13662 ( .A1(n10685), .A2(n19667), .ZN(n10667) );
  OAI211_X1 U13663 ( .C1(n10689), .C2(n10994), .A(n10668), .B(n10667), .ZN(
        n14768) );
  NAND2_X1 U13664 ( .A1(n14769), .A2(n14768), .ZN(n14757) );
  INV_X1 U13665 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19669) );
  NAND2_X1 U13666 ( .A1(n10679), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U13667 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10669) );
  OAI211_X1 U13668 ( .C1(n10685), .C2(n19669), .A(n10670), .B(n10669), .ZN(
        n10671) );
  AOI21_X1 U13669 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10671), .ZN(n14758) );
  OR2_X2 U13670 ( .A1(n14757), .A2(n14758), .ZN(n14760) );
  INV_X1 U13671 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n14898) );
  NAND2_X1 U13672 ( .A1(n10679), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10673) );
  NAND2_X1 U13673 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10672) );
  OAI211_X1 U13674 ( .C1(n10685), .C2(n14898), .A(n10673), .B(n10672), .ZN(
        n10674) );
  AOI21_X1 U13675 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10674), .ZN(n14746) );
  INV_X1 U13676 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15097) );
  AOI22_X1 U13677 ( .A1(n10679), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10676) );
  INV_X1 U13678 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19674) );
  OR2_X1 U13679 ( .A1(n10685), .A2(n19674), .ZN(n10675) );
  OAI211_X1 U13680 ( .C1(n10689), .C2(n15097), .A(n10676), .B(n10675), .ZN(
        n14743) );
  INV_X1 U13681 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n20769) );
  AOI22_X1 U13682 ( .A1(n10679), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10678) );
  NAND2_X1 U13683 ( .A1(n10255), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10677) );
  OAI211_X1 U13684 ( .C1(n10689), .C2(n20769), .A(n10678), .B(n10677), .ZN(
        n10919) );
  INV_X1 U13685 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20752) );
  NAND2_X1 U13686 ( .A1(n10679), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10681) );
  NAND2_X1 U13687 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10680) );
  OAI211_X1 U13688 ( .C1(n10685), .C2(n20752), .A(n10681), .B(n10680), .ZN(
        n10682) );
  AOI21_X1 U13689 ( .B1(n10273), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n10682), .ZN(n14727) );
  INV_X1 U13690 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U13691 ( .A1(n10679), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10684) );
  NAND2_X1 U13692 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10683) );
  OAI211_X1 U13693 ( .C1(n10685), .C2(n11209), .A(n10684), .B(n10683), .ZN(
        n10686) );
  AOI21_X1 U13694 ( .B1(n9601), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10686), .ZN(n10968) );
  INV_X1 U13695 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U13696 ( .A1(n10679), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10688) );
  NAND2_X1 U13697 ( .A1(n10644), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n10687) );
  OAI211_X1 U13698 ( .C1(n10689), .C2(n11221), .A(n10688), .B(n10687), .ZN(
        n10690) );
  INV_X1 U13699 ( .A(n10692), .ZN(n10698) );
  OAI21_X1 U13700 ( .B1(n12601), .B2(n12418), .A(n10698), .ZN(n10694) );
  NAND2_X1 U13701 ( .A1(n10694), .A2(n10693), .ZN(n10703) );
  INV_X1 U13702 ( .A(n10695), .ZN(n10696) );
  OAI21_X1 U13703 ( .B1(n19006), .B2(n10698), .A(n10696), .ZN(n10700) );
  NAND2_X1 U13704 ( .A1(n10698), .A2(n10697), .ZN(n10699) );
  NAND3_X1 U13705 ( .A1(n10700), .A2(n13457), .A3(n10699), .ZN(n10701) );
  OAI21_X1 U13706 ( .B1(n10122), .B2(n10721), .A(n10701), .ZN(n10702) );
  NAND3_X1 U13707 ( .A1(n10703), .A2(n10704), .A3(n10702), .ZN(n10707) );
  OAI21_X1 U13708 ( .B1(n10704), .B2(n10721), .A(n19726), .ZN(n10705) );
  INV_X1 U13709 ( .A(n10705), .ZN(n10706) );
  NAND2_X1 U13710 ( .A1(n10707), .A2(n10706), .ZN(n10708) );
  MUX2_X1 U13711 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10708), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n10931) );
  INV_X1 U13712 ( .A(n19726), .ZN(n10709) );
  AOI21_X1 U13713 ( .B1(n13409), .B2(n10711), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n15994) );
  NAND2_X1 U13714 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12610) );
  AND2_X1 U13715 ( .A1(n15994), .A2(n12610), .ZN(n10712) );
  OR2_X1 U13716 ( .A1(n15862), .A2(n15063), .ZN(n10716) );
  NAND2_X1 U13717 ( .A1(n19688), .A2(n10711), .ZN(n18595) );
  INV_X2 U13718 ( .A(n15891), .ZN(n18791) );
  INV_X1 U13719 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n10714) );
  NOR2_X1 U13720 ( .A1(n18970), .A2(n10714), .ZN(n11297) );
  AOI21_X1 U13721 ( .B1(n15915), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n11297), .ZN(n10715) );
  OAI211_X1 U13722 ( .C1(n15922), .C2(n11222), .A(n10716), .B(n10715), .ZN(
        n10717) );
  AOI21_X1 U13723 ( .B1(n11302), .B2(n15939), .A(n10717), .ZN(n10906) );
  INV_X1 U13724 ( .A(n10721), .ZN(n10986) );
  NAND2_X1 U13725 ( .A1(n10986), .A2(n19028), .ZN(n10748) );
  NAND2_X1 U13726 ( .A1(n12521), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10725) );
  AND2_X1 U13727 ( .A1(n10721), .A2(n19028), .ZN(n10745) );
  INV_X1 U13728 ( .A(n10722), .ZN(n10723) );
  NAND2_X1 U13729 ( .A1(n10745), .A2(n10723), .ZN(n10724) );
  OAI211_X1 U13730 ( .C1(n10748), .C2(n11055), .A(n10725), .B(n10724), .ZN(
        n10740) );
  INV_X1 U13731 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10726) );
  INV_X1 U13732 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n18827) );
  NAND2_X1 U13733 ( .A1(n10726), .A2(n18827), .ZN(n10728) );
  NOR2_X1 U13734 ( .A1(n10740), .A2(n10750), .ZN(n10730) );
  INV_X1 U13735 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12728) );
  MUX2_X1 U13736 ( .A(n10729), .B(n12728), .S(n12521), .Z(n10753) );
  INV_X1 U13737 ( .A(n10748), .ZN(n10731) );
  NAND2_X1 U13738 ( .A1(n10731), .A2(n11060), .ZN(n10734) );
  NAND2_X1 U13739 ( .A1(n10745), .A2(n10732), .ZN(n10733) );
  OAI211_X1 U13740 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n19028), .A(n10734), .B(
        n10733), .ZN(n10757) );
  NAND2_X1 U13741 ( .A1(n10758), .A2(n10757), .ZN(n10736) );
  MUX2_X1 U13742 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n11064), .S(n19028), .Z(
        n10735) );
  AND2_X1 U13743 ( .A1(n10736), .A2(n10735), .ZN(n10737) );
  OR2_X1 U13744 ( .A1(n10737), .A2(n10770), .ZN(n18788) );
  INV_X1 U13745 ( .A(n10758), .ZN(n10743) );
  INV_X1 U13746 ( .A(n10750), .ZN(n10752) );
  NAND2_X1 U13747 ( .A1(n10753), .A2(n10752), .ZN(n10741) );
  NAND2_X1 U13748 ( .A1(n10741), .A2(n10740), .ZN(n10742) );
  NAND2_X1 U13749 ( .A1(n10743), .A2(n10742), .ZN(n13575) );
  INV_X1 U13750 ( .A(n11032), .ZN(n12668) );
  NAND2_X1 U13751 ( .A1(n12521), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10747) );
  NAND2_X1 U13752 ( .A1(n10745), .A2(n10744), .ZN(n10746) );
  OAI211_X1 U13753 ( .C1(n10748), .C2(n12668), .A(n10747), .B(n10746), .ZN(
        n18820) );
  NAND2_X1 U13754 ( .A1(n18820), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12678) );
  NAND3_X1 U13755 ( .A1(n12521), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10749) );
  NAND2_X1 U13756 ( .A1(n10750), .A2(n10749), .ZN(n12679) );
  NOR2_X1 U13757 ( .A1(n12678), .A2(n12679), .ZN(n10751) );
  NAND2_X1 U13758 ( .A1(n12678), .A2(n12679), .ZN(n12677) );
  OAI21_X1 U13759 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10751), .A(
        n12677), .ZN(n12687) );
  XNOR2_X1 U13760 ( .A(n10753), .B(n10752), .ZN(n13523) );
  XNOR2_X1 U13761 ( .A(n13523), .B(n18990), .ZN(n12686) );
  OR2_X1 U13762 ( .A1(n12687), .A2(n12686), .ZN(n18975) );
  INV_X1 U13763 ( .A(n13523), .ZN(n10754) );
  NAND2_X1 U13764 ( .A1(n10754), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10755) );
  AND2_X1 U13765 ( .A1(n18975), .A2(n10755), .ZN(n13392) );
  NAND2_X1 U13766 ( .A1(n13390), .A2(n13392), .ZN(n10756) );
  XNOR2_X1 U13767 ( .A(n10758), .B(n10757), .ZN(n18805) );
  XNOR2_X1 U13768 ( .A(n18805), .B(n20652), .ZN(n13534) );
  OAI22_X1 U13769 ( .A1(n13535), .A2(n13534), .B1(n18805), .B2(n20652), .ZN(
        n13620) );
  NAND2_X1 U13770 ( .A1(n13621), .A2(n13620), .ZN(n10761) );
  NAND2_X1 U13771 ( .A1(n10759), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10760) );
  NAND2_X1 U13772 ( .A1(n10761), .A2(n10760), .ZN(n13703) );
  NAND2_X1 U13773 ( .A1(n10762), .A2(n10865), .ZN(n10765) );
  INV_X1 U13774 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12974) );
  MUX2_X1 U13775 ( .A(n12974), .B(n11069), .S(n19028), .Z(n10769) );
  INV_X1 U13776 ( .A(n10769), .ZN(n10763) );
  XNOR2_X1 U13777 ( .A(n10770), .B(n10763), .ZN(n18776) );
  INV_X1 U13778 ( .A(n18776), .ZN(n10764) );
  NAND2_X1 U13779 ( .A1(n10765), .A2(n10764), .ZN(n10766) );
  INV_X1 U13780 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U13781 ( .A1(n10766), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10767) );
  NAND2_X1 U13782 ( .A1(n10770), .A2(n10769), .ZN(n10777) );
  MUX2_X1 U13783 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n10865), .S(n19028), .Z(
        n10775) );
  OR2_X2 U13784 ( .A1(n10777), .A2(n10775), .ZN(n10782) );
  INV_X1 U13785 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10771) );
  NOR2_X1 U13786 ( .A1(n19028), .A2(n10771), .ZN(n10780) );
  INV_X1 U13787 ( .A(n10780), .ZN(n10772) );
  XNOR2_X1 U13788 ( .A(n10782), .B(n10772), .ZN(n18754) );
  INV_X1 U13789 ( .A(n10773), .ZN(n10774) );
  AND2_X1 U13790 ( .A1(n18754), .A2(n10774), .ZN(n15935) );
  INV_X1 U13791 ( .A(n10775), .ZN(n10776) );
  XNOR2_X1 U13792 ( .A(n10777), .B(n10776), .ZN(n18767) );
  NAND2_X1 U13793 ( .A1(n18754), .A2(n10895), .ZN(n10778) );
  NAND2_X1 U13794 ( .A1(n10778), .A2(n11079), .ZN(n15934) );
  OR2_X1 U13795 ( .A1(n18767), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15933) );
  AND2_X1 U13796 ( .A1(n15934), .A2(n15933), .ZN(n10779) );
  NAND2_X1 U13797 ( .A1(n12521), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10781) );
  XNOR2_X1 U13798 ( .A(n9652), .B(n10781), .ZN(n18739) );
  AOI21_X1 U13799 ( .B1(n18739), .B2(n10895), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15315) );
  INV_X1 U13800 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12959) );
  NAND2_X1 U13801 ( .A1(n12521), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10783) );
  OAI21_X1 U13802 ( .B1(n10784), .B2(n10783), .A(n10874), .ZN(n10785) );
  OR2_X1 U13803 ( .A1(n10835), .A2(n10785), .ZN(n18730) );
  INV_X1 U13804 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10786) );
  OAI21_X1 U13805 ( .B1(n18730), .B2(n10865), .A(n10786), .ZN(n15297) );
  INV_X1 U13806 ( .A(n18730), .ZN(n10788) );
  NOR2_X1 U13807 ( .A1(n10865), .A2(n10786), .ZN(n10787) );
  NAND2_X1 U13808 ( .A1(n10788), .A2(n10787), .ZN(n15296) );
  INV_X1 U13809 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15318) );
  NOR2_X1 U13810 ( .A1(n10865), .A2(n15318), .ZN(n10789) );
  NAND2_X1 U13811 ( .A1(n18739), .A2(n10789), .ZN(n15294) );
  INV_X1 U13812 ( .A(n15279), .ZN(n10790) );
  NAND2_X1 U13813 ( .A1(n10790), .A2(n15280), .ZN(n14948) );
  NAND2_X1 U13814 ( .A1(n12521), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10797) );
  INV_X1 U13815 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13070) );
  NAND2_X1 U13816 ( .A1(n10874), .A2(n9649), .ZN(n10836) );
  NAND2_X1 U13817 ( .A1(n12521), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10791) );
  INV_X1 U13818 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10792) );
  NOR2_X1 U13819 ( .A1(n19028), .A2(n10792), .ZN(n10814) );
  INV_X1 U13820 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13384) );
  INV_X1 U13821 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n18673) );
  NAND2_X1 U13822 ( .A1(n13384), .A2(n18673), .ZN(n10793) );
  NAND2_X1 U13823 ( .A1(n12521), .A2(n10793), .ZN(n10794) );
  NOR2_X1 U13824 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n10795) );
  NOR2_X1 U13825 ( .A1(n19028), .A2(n10795), .ZN(n10796) );
  MUX2_X1 U13826 ( .A(n12521), .B(n10797), .S(n10827), .Z(n10798) );
  INV_X1 U13827 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15879) );
  NAND2_X1 U13828 ( .A1(n9836), .A2(n15879), .ZN(n10799) );
  NAND2_X1 U13829 ( .A1(n10798), .A2(n10799), .ZN(n18645) );
  INV_X1 U13830 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15209) );
  OAI21_X1 U13831 ( .B1(n18645), .B2(n10865), .A(n15209), .ZN(n14991) );
  NAND3_X1 U13832 ( .A1(n10799), .A2(n12521), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n10802) );
  INV_X1 U13833 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10800) );
  AND2_X1 U13834 ( .A1(n15879), .A2(n10800), .ZN(n10801) );
  NAND2_X1 U13835 ( .A1(n10802), .A2(n10831), .ZN(n18635) );
  NAND2_X1 U13836 ( .A1(n10843), .A2(n15195), .ZN(n14989) );
  AND2_X1 U13837 ( .A1(n14991), .A2(n14989), .ZN(n14960) );
  NAND2_X1 U13838 ( .A1(n12521), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10804) );
  INV_X1 U13839 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10803) );
  OAI211_X1 U13840 ( .C1(n10805), .C2(n10804), .A(n10874), .B(n10857), .ZN(
        n12562) );
  OR2_X1 U13841 ( .A1(n12562), .A2(n10865), .ZN(n10806) );
  NAND2_X1 U13842 ( .A1(n10806), .A2(n14967), .ZN(n14962) );
  INV_X1 U13843 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10807) );
  NOR2_X1 U13844 ( .A1(n19028), .A2(n10807), .ZN(n10809) );
  INV_X1 U13845 ( .A(n10874), .ZN(n10808) );
  AOI21_X1 U13846 ( .B1(n10812), .B2(n10809), .A(n10808), .ZN(n10810) );
  OR2_X1 U13847 ( .A1(n10812), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13848 ( .A1(n10810), .A2(n10826), .ZN(n18666) );
  OR2_X1 U13849 ( .A1(n18666), .A2(n10865), .ZN(n10811) );
  XNOR2_X1 U13850 ( .A(n10811), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14956) );
  NAND2_X1 U13851 ( .A1(n10821), .A2(n13384), .ZN(n10823) );
  NAND3_X1 U13852 ( .A1(n10823), .A2(n12521), .A3(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n10813) );
  NAND2_X1 U13853 ( .A1(n10813), .A2(n10812), .ZN(n18672) );
  INV_X1 U13854 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15250) );
  NAND2_X1 U13855 ( .A1(n10850), .A2(n15250), .ZN(n15038) );
  AND2_X1 U13856 ( .A1(n10819), .A2(n10814), .ZN(n10815) );
  OR2_X1 U13857 ( .A1(n10815), .A2(n10821), .ZN(n18696) );
  INV_X1 U13858 ( .A(n18696), .ZN(n10816) );
  NAND2_X1 U13859 ( .A1(n10816), .A2(n10895), .ZN(n10846) );
  INV_X1 U13860 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10817) );
  NAND2_X1 U13861 ( .A1(n10846), .A2(n10817), .ZN(n15259) );
  NAND3_X1 U13862 ( .A1(n12521), .A2(n9649), .A3(P2_EBX_REG_12__SCAN_IN), .ZN(
        n10818) );
  AND2_X1 U13863 ( .A1(n10819), .A2(n10818), .ZN(n18711) );
  NAND2_X1 U13864 ( .A1(n18711), .A2(n10895), .ZN(n14950) );
  NAND2_X1 U13865 ( .A1(n14950), .A2(n15972), .ZN(n14951) );
  AND3_X1 U13866 ( .A1(n15038), .A2(n15259), .A3(n14951), .ZN(n10829) );
  NOR2_X1 U13867 ( .A1(n10821), .A2(n13384), .ZN(n10820) );
  MUX2_X1 U13868 ( .A(n10821), .B(n10820), .S(n12521), .Z(n10822) );
  INV_X1 U13869 ( .A(n10822), .ZN(n10824) );
  NAND2_X1 U13870 ( .A1(n10824), .A2(n10823), .ZN(n18690) );
  OR2_X1 U13871 ( .A1(n18690), .A2(n10865), .ZN(n10825) );
  NAND2_X1 U13872 ( .A1(n10825), .A2(n15898), .ZN(n15894) );
  NAND3_X1 U13873 ( .A1(n10826), .A2(n12521), .A3(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n10828) );
  NAND2_X1 U13874 ( .A1(n10828), .A2(n10827), .ZN(n18654) );
  INV_X1 U13875 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15009) );
  NAND2_X1 U13876 ( .A1(n10848), .A2(n15009), .ZN(n15018) );
  AND4_X1 U13877 ( .A1(n14956), .A2(n10829), .A3(n15894), .A4(n15018), .ZN(
        n10833) );
  NAND2_X1 U13878 ( .A1(n12521), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10830) );
  XNOR2_X1 U13879 ( .A(n10831), .B(n10830), .ZN(n18618) );
  NAND2_X1 U13880 ( .A1(n18618), .A2(n10895), .ZN(n10832) );
  NAND2_X1 U13881 ( .A1(n10832), .A2(n15183), .ZN(n14974) );
  AND4_X1 U13882 ( .A1(n14960), .A2(n14962), .A3(n10833), .A4(n14974), .ZN(
        n10840) );
  NAND2_X1 U13883 ( .A1(n12521), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10834) );
  OR2_X1 U13884 ( .A1(n10835), .A2(n10834), .ZN(n10838) );
  INV_X1 U13885 ( .A(n10836), .ZN(n10837) );
  AND2_X1 U13886 ( .A1(n10838), .A2(n10837), .ZN(n18722) );
  NAND2_X1 U13887 ( .A1(n18722), .A2(n10895), .ZN(n15281) );
  OR2_X1 U13888 ( .A1(n12562), .A2(n14967), .ZN(n14963) );
  INV_X1 U13889 ( .A(n18645), .ZN(n10841) );
  NAND2_X1 U13890 ( .A1(n10841), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14959) );
  OR2_X1 U13891 ( .A1(n18666), .A2(n10842), .ZN(n14957) );
  NAND2_X1 U13892 ( .A1(n18618), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14961) );
  NAND4_X1 U13893 ( .A1(n14963), .A2(n14959), .A3(n14957), .A4(n14961), .ZN(
        n10852) );
  INV_X1 U13894 ( .A(n10843), .ZN(n10844) );
  NAND2_X1 U13895 ( .A1(n10844), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14990) );
  OR2_X1 U13896 ( .A1(n10865), .A2(n15898), .ZN(n10845) );
  OR2_X1 U13897 ( .A1(n18690), .A2(n10845), .ZN(n15893) );
  INV_X1 U13898 ( .A(n10846), .ZN(n10847) );
  NAND2_X1 U13899 ( .A1(n10847), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15892) );
  AND2_X1 U13900 ( .A1(n15893), .A2(n15892), .ZN(n14954) );
  INV_X1 U13901 ( .A(n10848), .ZN(n10849) );
  NAND2_X1 U13902 ( .A1(n10849), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14958) );
  NAND4_X1 U13903 ( .A1(n14990), .A2(n14954), .A3(n14958), .A4(n15039), .ZN(
        n10851) );
  AOI21_X1 U13904 ( .B1(n10895), .B2(n10852), .A(n10851), .ZN(n10853) );
  NAND2_X1 U13905 ( .A1(n10857), .A2(n10874), .ZN(n10854) );
  NAND2_X1 U13906 ( .A1(n12521), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10855) );
  INV_X1 U13907 ( .A(n10855), .ZN(n10856) );
  NAND2_X1 U13908 ( .A1(n10857), .A2(n10856), .ZN(n10858) );
  NAND2_X1 U13909 ( .A1(n10862), .A2(n10858), .ZN(n15575) );
  OR2_X1 U13910 ( .A1(n15575), .A2(n10865), .ZN(n10859) );
  INV_X1 U13911 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20668) );
  NAND2_X1 U13912 ( .A1(n10859), .A2(n20668), .ZN(n14935) );
  INV_X1 U13913 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10860) );
  NOR2_X1 U13914 ( .A1(n19028), .A2(n10860), .ZN(n10861) );
  NAND2_X1 U13915 ( .A1(n10862), .A2(n10861), .ZN(n10863) );
  NAND2_X1 U13916 ( .A1(n10871), .A2(n10863), .ZN(n12572) );
  OR2_X1 U13917 ( .A1(n12572), .A2(n10865), .ZN(n10864) );
  XNOR2_X1 U13918 ( .A(n10864), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14923) );
  INV_X1 U13919 ( .A(n12572), .ZN(n10866) );
  NAND3_X1 U13920 ( .A1(n10866), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n10895), .ZN(n10867) );
  NAND2_X1 U13921 ( .A1(n10874), .A2(n10895), .ZN(n14914) );
  NOR2_X1 U13922 ( .A1(n14914), .A2(n10994), .ZN(n10869) );
  NAND2_X1 U13923 ( .A1(n14914), .A2(n10994), .ZN(n10870) );
  INV_X1 U13924 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15853) );
  NAND2_X1 U13925 ( .A1(n12521), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10872) );
  OR2_X1 U13926 ( .A1(n15837), .A2(n10872), .ZN(n10875) );
  INV_X1 U13927 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10873) );
  NAND2_X1 U13928 ( .A1(n15837), .A2(n10873), .ZN(n10878) );
  NAND2_X1 U13929 ( .A1(n10874), .A2(n10878), .ZN(n10876) );
  INV_X1 U13930 ( .A(n10876), .ZN(n10900) );
  NAND2_X1 U13931 ( .A1(n15826), .A2(n10895), .ZN(n10885) );
  INV_X1 U13932 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10884) );
  NAND2_X1 U13933 ( .A1(n10885), .A2(n10884), .ZN(n10907) );
  NAND2_X1 U13934 ( .A1(n12521), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U13935 ( .A1(n10876), .A2(n10877), .ZN(n10889) );
  INV_X1 U13936 ( .A(n10877), .ZN(n10879) );
  NAND2_X1 U13937 ( .A1(n10879), .A2(n10878), .ZN(n10880) );
  NAND2_X1 U13938 ( .A1(n10889), .A2(n10880), .ZN(n15816) );
  INV_X1 U13939 ( .A(n15072), .ZN(n10881) );
  AND2_X1 U13940 ( .A1(n14914), .A2(n15118), .ZN(n14895) );
  NOR2_X1 U13941 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10886) );
  INV_X1 U13942 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10882) );
  NOR2_X1 U13943 ( .A1(n19028), .A2(n10882), .ZN(n10888) );
  INV_X1 U13944 ( .A(n10888), .ZN(n10883) );
  XNOR2_X1 U13945 ( .A(n10889), .B(n10883), .ZN(n15804) );
  NAND2_X1 U13946 ( .A1(n15804), .A2(n10895), .ZN(n10914) );
  OR2_X1 U13947 ( .A1(n14914), .A2(n15118), .ZN(n14906) );
  OAI21_X1 U13948 ( .B1(n10886), .B2(n10914), .A(n10909), .ZN(n10887) );
  NAND2_X1 U13949 ( .A1(n12521), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10891) );
  INV_X1 U13950 ( .A(n10891), .ZN(n10890) );
  XNOR2_X1 U13951 ( .A(n10892), .B(n10890), .ZN(n15796) );
  AOI21_X1 U13952 ( .B1(n15796), .B2(n10895), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14880) );
  NAND2_X1 U13953 ( .A1(n10892), .A2(n10891), .ZN(n10898) );
  INV_X1 U13954 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10893) );
  NOR2_X1 U13955 ( .A1(n19028), .A2(n10893), .ZN(n10894) );
  XNOR2_X1 U13956 ( .A(n10898), .B(n10894), .ZN(n11287) );
  INV_X1 U13957 ( .A(n11287), .ZN(n10896) );
  AOI21_X1 U13958 ( .B1(n10896), .B2(n10895), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10964) );
  INV_X1 U13959 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11299) );
  OR3_X1 U13960 ( .A1(n11287), .A2(n10865), .A3(n11299), .ZN(n10962) );
  INV_X1 U13961 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15071) );
  NOR2_X1 U13962 ( .A1(n10865), .A2(n15071), .ZN(n10897) );
  NAND2_X1 U13963 ( .A1(n15796), .A2(n10897), .ZN(n14878) );
  NOR2_X1 U13964 ( .A1(n10898), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10899) );
  MUX2_X1 U13965 ( .A(n10900), .B(n10899), .S(n12521), .Z(n15784) );
  NAND2_X1 U13966 ( .A1(n15784), .A2(n10895), .ZN(n10901) );
  NAND2_X1 U13967 ( .A1(n10906), .A2(n10905), .ZN(P2_U2983) );
  INV_X1 U13968 ( .A(n14895), .ZN(n14907) );
  INV_X1 U13969 ( .A(n10911), .ZN(n10913) );
  XNOR2_X1 U13970 ( .A(n10914), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10915) );
  XNOR2_X1 U13971 ( .A(n10916), .B(n10915), .ZN(n15091) );
  INV_X1 U13972 ( .A(n14902), .ZN(n10917) );
  NAND2_X1 U13973 ( .A1(n10917), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14888) );
  XNOR2_X1 U13974 ( .A(n14888), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15089) );
  OR2_X1 U13975 ( .A1(n10920), .A2(n10919), .ZN(n10921) );
  NAND2_X2 U13976 ( .A1(n10918), .A2(n10921), .ZN(n15805) );
  NOR2_X1 U13977 ( .A1(n10923), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10924) );
  OR2_X1 U13978 ( .A1(n10922), .A2(n10924), .ZN(n11223) );
  NAND2_X1 U13979 ( .A1(n18791), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15082) );
  NAND2_X1 U13980 ( .A1(n15915), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10925) );
  OAI211_X1 U13981 ( .C1(n15922), .C2(n11223), .A(n15082), .B(n10925), .ZN(
        n10926) );
  INV_X1 U13982 ( .A(n10926), .ZN(n10927) );
  NAND2_X1 U13983 ( .A1(n10129), .A2(n10927), .ZN(n10928) );
  AOI21_X1 U13984 ( .B1(n15089), .B2(n15939), .A(n10928), .ZN(n10929) );
  OAI21_X1 U13985 ( .B1(n15091), .B2(n15946), .A(n10929), .ZN(P2_U2986) );
  INV_X1 U13986 ( .A(n10930), .ZN(n14876) );
  INV_X1 U13987 ( .A(n10585), .ZN(n13239) );
  NAND3_X1 U13988 ( .A1(n15631), .A2(n13239), .A3(n19006), .ZN(n10958) );
  AOI21_X1 U13989 ( .B1(n10931), .B2(n13457), .A(n19023), .ZN(n10955) );
  NAND2_X1 U13990 ( .A1(n13237), .A2(n19006), .ZN(n12599) );
  INV_X1 U13991 ( .A(n10932), .ZN(n10949) );
  NOR2_X1 U13992 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19630) );
  AOI211_X1 U13993 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19630), .ZN(n19623) );
  NAND2_X1 U13994 ( .A1(n19623), .A2(n19617), .ZN(n12603) );
  NOR2_X1 U13995 ( .A1(n10949), .A2(n12603), .ZN(n10936) );
  INV_X1 U13996 ( .A(n10987), .ZN(n10933) );
  NAND2_X1 U13997 ( .A1(n10934), .A2(n10933), .ZN(n10935) );
  AOI21_X1 U13998 ( .B1(n10936), .B2(n11282), .A(n10935), .ZN(n10948) );
  NAND2_X1 U13999 ( .A1(n10938), .A2(n10937), .ZN(n10940) );
  AOI21_X1 U14000 ( .B1(n10940), .B2(n19044), .A(n10939), .ZN(n10974) );
  OAI21_X1 U14001 ( .B1(n19023), .B2(n19006), .A(n13457), .ZN(n10941) );
  AOI21_X1 U14002 ( .B1(n10941), .B2(n19044), .A(n19010), .ZN(n10942) );
  NOR2_X1 U14003 ( .A1(n10974), .A2(n10942), .ZN(n10947) );
  NAND2_X1 U14004 ( .A1(n10944), .A2(n10943), .ZN(n10945) );
  NAND2_X1 U14005 ( .A1(n12614), .A2(n10945), .ZN(n10946) );
  AND3_X1 U14006 ( .A1(n10948), .A2(n10947), .A3(n10946), .ZN(n12608) );
  NAND2_X1 U14007 ( .A1(n10949), .A2(n19006), .ZN(n10951) );
  INV_X1 U14008 ( .A(n10972), .ZN(n10950) );
  NAND4_X1 U14009 ( .A1(n10951), .A2(n11282), .A3(n19617), .A4(n10950), .ZN(
        n10952) );
  NAND3_X1 U14010 ( .A1(n12608), .A2(n10953), .A3(n10952), .ZN(n10954) );
  AOI21_X1 U14011 ( .B1(n10955), .B2(n12599), .A(n10954), .ZN(n10957) );
  INV_X1 U14012 ( .A(n12599), .ZN(n12605) );
  INV_X1 U14013 ( .A(n12603), .ZN(n12584) );
  NAND3_X1 U14014 ( .A1(n12605), .A2(n12584), .A3(n19010), .ZN(n10956) );
  NAND3_X1 U14015 ( .A1(n10958), .A2(n10957), .A3(n10956), .ZN(n10959) );
  INV_X1 U14016 ( .A(n10960), .ZN(n19724) );
  NAND2_X1 U14017 ( .A1(n10961), .A2(n14878), .ZN(n10966) );
  INV_X1 U14018 ( .A(n10962), .ZN(n10963) );
  NOR2_X1 U14019 ( .A1(n10964), .A2(n10963), .ZN(n10965) );
  INV_X1 U14020 ( .A(n19728), .ZN(n10967) );
  NAND2_X1 U14021 ( .A1(n13256), .A2(n12418), .ZN(n10969) );
  AND2_X1 U14022 ( .A1(n10969), .A2(n13202), .ZN(n10970) );
  NAND2_X1 U14023 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15986) );
  INV_X1 U14024 ( .A(n15986), .ZN(n10993) );
  NAND2_X1 U14025 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13622) );
  INV_X1 U14026 ( .A(n13622), .ZN(n10997) );
  AND2_X1 U14027 ( .A1(n10972), .A2(n19028), .ZN(n10973) );
  NAND2_X1 U14028 ( .A1(n13248), .A2(n10973), .ZN(n13236) );
  NAND2_X1 U14029 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18965) );
  NOR2_X1 U14030 ( .A1(n18990), .A2(n18965), .ZN(n18972) );
  NAND2_X1 U14031 ( .A1(n18990), .A2(n18965), .ZN(n10991) );
  INV_X1 U14032 ( .A(n10974), .ZN(n10976) );
  NAND2_X1 U14033 ( .A1(n10975), .A2(n19006), .ZN(n13249) );
  NAND2_X1 U14034 ( .A1(n10976), .A2(n13249), .ZN(n10982) );
  NAND2_X1 U14035 ( .A1(n13238), .A2(n19010), .ZN(n10979) );
  INV_X1 U14036 ( .A(n12501), .ZN(n12591) );
  OAI21_X1 U14037 ( .B1(n10987), .B2(n10977), .A(n12591), .ZN(n10978) );
  NAND3_X1 U14038 ( .A1(n10980), .A2(n10979), .A3(n10978), .ZN(n10981) );
  AOI21_X1 U14039 ( .B1(n10982), .B2(n19016), .A(n10981), .ZN(n10985) );
  OAI211_X1 U14040 ( .C1(n12504), .C2(n10118), .A(n10987), .B(n10983), .ZN(
        n10984) );
  NAND2_X1 U14041 ( .A1(n10985), .A2(n10984), .ZN(n13252) );
  NAND2_X1 U14042 ( .A1(n10987), .A2(n10986), .ZN(n10989) );
  NOR2_X1 U14043 ( .A1(n10989), .A2(n10988), .ZN(n12533) );
  NOR2_X1 U14044 ( .A1(n13252), .A2(n12533), .ZN(n10990) );
  NOR2_X1 U14045 ( .A1(n11218), .A2(n10990), .ZN(n18964) );
  OAI211_X1 U14046 ( .C1(n18973), .C2(n18972), .A(n10991), .B(n15203), .ZN(
        n13401) );
  NOR2_X1 U14047 ( .A1(n13402), .A2(n13401), .ZN(n13623) );
  NAND2_X1 U14048 ( .A1(n10997), .A2(n13623), .ZN(n13701) );
  NAND2_X1 U14049 ( .A1(n10993), .A2(n15987), .ZN(n15959) );
  NAND2_X1 U14050 ( .A1(n15222), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15204) );
  NOR2_X1 U14051 ( .A1(n15204), .A2(n15209), .ZN(n15163) );
  NAND2_X1 U14052 ( .A1(n15162), .A2(n15163), .ZN(n15177) );
  NAND2_X1 U14053 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15178) );
  NOR2_X1 U14054 ( .A1(n15177), .A2(n15178), .ZN(n15159) );
  NAND2_X1 U14055 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15159), .ZN(
        n10998) );
  NOR2_X1 U14056 ( .A1(n15959), .A2(n10998), .ZN(n15148) );
  NOR2_X1 U14057 ( .A1(n15137), .A2(n10994), .ZN(n10995) );
  NAND2_X1 U14058 ( .A1(n15148), .A2(n10995), .ZN(n15104) );
  NAND2_X1 U14059 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11002) );
  NOR2_X1 U14060 ( .A1(n15070), .A2(n11298), .ZN(n11005) );
  NAND2_X1 U14061 ( .A1(n11218), .A2(n15891), .ZN(n12743) );
  INV_X1 U14062 ( .A(n15267), .ZN(n13537) );
  INV_X1 U14063 ( .A(n18972), .ZN(n10996) );
  AND2_X1 U14064 ( .A1(n18964), .A2(n10996), .ZN(n18967) );
  AND3_X1 U14065 ( .A1(n18990), .A2(n18965), .A3(n18973), .ZN(n18968) );
  NOR4_X1 U14066 ( .A1(n18967), .A2(n18963), .A3(n18968), .A4(n13402), .ZN(
        n13536) );
  NAND3_X1 U14067 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13536), .A3(
        n10997), .ZN(n13696) );
  OR2_X1 U14068 ( .A1(n13696), .A2(n15986), .ZN(n15268) );
  NAND2_X1 U14069 ( .A1(n15268), .A2(n15267), .ZN(n15319) );
  NAND2_X1 U14070 ( .A1(n15267), .A2(n10998), .ZN(n10999) );
  NAND2_X1 U14071 ( .A1(n15319), .A2(n10999), .ZN(n15150) );
  NAND2_X1 U14072 ( .A1(n15267), .A2(n15137), .ZN(n11000) );
  NAND2_X1 U14073 ( .A1(n11000), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11001) );
  NOR2_X1 U14074 ( .A1(n15150), .A2(n11001), .ZN(n15130) );
  INV_X1 U14075 ( .A(n11002), .ZN(n11003) );
  NAND2_X1 U14076 ( .A1(n15130), .A2(n11003), .ZN(n11004) );
  NAND2_X1 U14077 ( .A1(n11004), .A2(n15267), .ZN(n15098) );
  OAI211_X1 U14078 ( .C1(n13537), .C2(n10109), .A(n15098), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11296) );
  OAI21_X1 U14079 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n11005), .A(
        n11296), .ZN(n11006) );
  OR2_X1 U14080 ( .A1(n15891), .A2(n11209), .ZN(n14866) );
  OAI211_X1 U14081 ( .C1(n14871), .C2(n15330), .A(n11006), .B(n14866), .ZN(
        n11219) );
  AOI22_X1 U14082 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10428), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14083 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U14084 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11008) );
  AND2_X1 U14085 ( .A1(n11009), .A2(n11008), .ZN(n11012) );
  AOI22_X1 U14086 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U14087 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11010) );
  NAND4_X1 U14088 ( .A1(n11013), .A2(n11012), .A3(n11011), .A4(n11010), .ZN(
        n11019) );
  AOI22_X1 U14089 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U14090 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10436), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U14091 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11015) );
  NAND2_X1 U14092 ( .A1(n12341), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11014) );
  NAND4_X1 U14093 ( .A1(n11017), .A2(n11016), .A3(n11015), .A4(n11014), .ZN(
        n11018) );
  INV_X1 U14094 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n11022) );
  AND2_X2 U14095 ( .A1(n11021), .A2(n19544), .ZN(n11076) );
  INV_X1 U14096 ( .A(n11076), .ZN(n11185) );
  OAI22_X1 U14097 ( .A1(n11186), .A2(n11022), .B1(n11185), .B2(n15898), .ZN(
        n11027) );
  NOR2_X1 U14098 ( .A1(n19028), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11024) );
  NOR2_X1 U14099 ( .A1(n11210), .A2(n11025), .ZN(n11026) );
  AOI211_X1 U14100 ( .C1(n11180), .C2(n13376), .A(n11027), .B(n11026), .ZN(
        n15956) );
  NAND2_X1 U14101 ( .A1(n11054), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11031) );
  INV_X1 U14102 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11028) );
  OAI211_X1 U14103 ( .C1(n19044), .C2(n11028), .A(n10117), .B(n19544), .ZN(
        n11029) );
  INV_X1 U14104 ( .A(n11029), .ZN(n11030) );
  NAND2_X1 U14105 ( .A1(n11031), .A2(n11030), .ZN(n12714) );
  NAND2_X1 U14106 ( .A1(n11180), .A2(n11032), .ZN(n11034) );
  NAND2_X1 U14107 ( .A1(n11041), .A2(n11076), .ZN(n11046) );
  NAND2_X1 U14108 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11033) );
  NAND4_X1 U14109 ( .A1(n11034), .A2(n11186), .A3(n11046), .A4(n11033), .ZN(
        n12713) );
  AOI22_X1 U14110 ( .A1(n11020), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11076), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U14111 ( .A1(n11054), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11035) );
  NAND2_X1 U14112 ( .A1(n11036), .A2(n11035), .ZN(n11042) );
  XNOR2_X1 U14113 ( .A(n11043), .B(n11042), .ZN(n12553) );
  NAND2_X1 U14114 ( .A1(n19044), .A2(n19544), .ZN(n11040) );
  NAND2_X1 U14115 ( .A1(n11180), .A2(n11037), .ZN(n11039) );
  NAND2_X1 U14116 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11038) );
  OAI211_X1 U14117 ( .C1(n11041), .C2(n11040), .A(n11039), .B(n11038), .ZN(
        n12552) );
  NOR2_X1 U14118 ( .A1(n12553), .A2(n12552), .ZN(n11045) );
  NOR2_X1 U14119 ( .A1(n11043), .A2(n11042), .ZN(n11044) );
  NOR2_X2 U14120 ( .A1(n11045), .A2(n11044), .ZN(n11050) );
  INV_X1 U14121 ( .A(n11180), .ZN(n11150) );
  NAND2_X1 U14122 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11047) );
  OAI211_X1 U14123 ( .C1(n11150), .C2(n11048), .A(n11047), .B(n11046), .ZN(
        n11049) );
  NOR2_X1 U14124 ( .A1(n11050), .A2(n11049), .ZN(n11053) );
  INV_X2 U14125 ( .A(n11186), .ZN(n11207) );
  AOI22_X1 U14126 ( .A1(n11207), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11076), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11052) );
  NAND2_X1 U14127 ( .A1(n11294), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11051) );
  NAND2_X1 U14128 ( .A1(n11052), .A2(n11051), .ZN(n12919) );
  NOR2_X1 U14129 ( .A1(n12920), .A2(n12919), .ZN(n12921) );
  NAND2_X1 U14130 ( .A1(n11294), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14131 ( .A1(n11076), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11058) );
  NAND2_X1 U14132 ( .A1(n11180), .A2(n11055), .ZN(n11057) );
  NAND2_X1 U14133 ( .A1(n11207), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11056) );
  NAND2_X1 U14134 ( .A1(n11294), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14135 ( .A1(n11207), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11076), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U14136 ( .A1(n11180), .A2(n11060), .ZN(n11061) );
  AOI22_X1 U14137 ( .A1(n11294), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11207), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11068) );
  NOR2_X1 U14138 ( .A1(n11064), .A2(n12521), .ZN(n11065) );
  MUX2_X1 U14139 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11065), .S(n9600), .Z(n11066) );
  NAND2_X1 U14140 ( .A1(n11066), .A2(n19544), .ZN(n11067) );
  NAND2_X1 U14141 ( .A1(n11068), .A2(n11067), .ZN(n13625) );
  NAND2_X1 U14142 ( .A1(n11180), .A2(n11069), .ZN(n11070) );
  NAND2_X1 U14143 ( .A1(n11071), .A2(n11070), .ZN(n12734) );
  AOI22_X1 U14144 ( .A1(n11207), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11076), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11073) );
  NAND2_X1 U14145 ( .A1(n11294), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11072) );
  NAND2_X1 U14146 ( .A1(n11073), .A2(n11072), .ZN(n12733) );
  NAND2_X1 U14147 ( .A1(n12734), .A2(n12733), .ZN(n11075) );
  NAND2_X1 U14148 ( .A1(n11180), .A2(n10895), .ZN(n11074) );
  NAND2_X1 U14149 ( .A1(n11075), .A2(n11074), .ZN(n12749) );
  AOI22_X1 U14150 ( .A1(n11207), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11076), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U14151 ( .A1(n11294), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11077) );
  NAND2_X1 U14152 ( .A1(n11078), .A2(n11077), .ZN(n12748) );
  NOR2_X1 U14153 ( .A1(n11185), .A2(n11079), .ZN(n11094) );
  AOI22_X1 U14154 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n10511), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14155 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12332), .B1(
        n12333), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U14156 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11080) );
  AND2_X1 U14157 ( .A1(n11081), .A2(n11080), .ZN(n11084) );
  AOI22_X1 U14158 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U14159 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n10431), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11082) );
  NAND4_X1 U14160 ( .A1(n11085), .A2(n11084), .A3(n11083), .A4(n11082), .ZN(
        n11091) );
  AOI22_X1 U14161 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n10482), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14162 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12341), .B1(
        n10436), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14163 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12343), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11087) );
  NAND2_X1 U14164 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11086) );
  NAND4_X1 U14165 ( .A1(n11089), .A2(n11088), .A3(n11087), .A4(n11086), .ZN(
        n11090) );
  INV_X1 U14166 ( .A(n12223), .ZN(n13011) );
  OAI22_X1 U14167 ( .A1(n11210), .A2(n11092), .B1(n11150), .B2(n13011), .ZN(
        n11093) );
  AOI211_X1 U14168 ( .C1(n11207), .C2(P2_EAX_REG_8__SCAN_IN), .A(n11094), .B(
        n11093), .ZN(n15981) );
  AOI22_X1 U14169 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10428), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14170 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12332), .B1(
        n12333), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11096) );
  NAND2_X1 U14171 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11095) );
  AND2_X1 U14172 ( .A1(n11096), .A2(n11095), .ZN(n11099) );
  AOI22_X1 U14173 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14174 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10482), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11097) );
  NAND4_X1 U14175 ( .A1(n11100), .A2(n11099), .A3(n11098), .A4(n11097), .ZN(
        n11106) );
  AOI22_X1 U14176 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10382), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14177 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12341), .B1(
        n10436), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11103) );
  AOI22_X1 U14178 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12343), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U14179 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11101) );
  NAND4_X1 U14180 ( .A1(n11104), .A2(n11103), .A3(n11102), .A4(n11101), .ZN(
        n11105) );
  AOI22_X1 U14181 ( .A1(n11294), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n11180), 
        .B2(n12948), .ZN(n11108) );
  AOI22_X1 U14182 ( .A1(n11207), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11076), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11107) );
  NAND2_X1 U14183 ( .A1(n11108), .A2(n11107), .ZN(n12825) );
  NAND2_X1 U14184 ( .A1(n11294), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U14185 ( .A1(n11207), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U14186 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10511), .B1(
        n10428), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14187 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12332), .B1(
        n12333), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11110) );
  NAND2_X1 U14188 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11109) );
  AND2_X1 U14189 ( .A1(n11110), .A2(n11109), .ZN(n11113) );
  AOI22_X1 U14190 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14191 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11111) );
  NAND4_X1 U14192 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(
        n11120) );
  AOI22_X1 U14193 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14194 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10436), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14195 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11116) );
  NAND2_X1 U14196 ( .A1(n12341), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11115) );
  NAND4_X1 U14197 ( .A1(n11118), .A2(n11117), .A3(n11116), .A4(n11115), .ZN(
        n11119) );
  NAND2_X1 U14198 ( .A1(n11180), .A2(n12951), .ZN(n11121) );
  AOI22_X1 U14199 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14200 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11125) );
  NAND2_X1 U14201 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11124) );
  AND2_X1 U14202 ( .A1(n11125), .A2(n11124), .ZN(n11128) );
  AOI22_X1 U14203 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11127) );
  AOI22_X1 U14204 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11126) );
  NAND4_X1 U14205 ( .A1(n11129), .A2(n11128), .A3(n11127), .A4(n11126), .ZN(
        n11135) );
  AOI22_X1 U14206 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U14207 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U14208 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11131) );
  NAND2_X1 U14209 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11130) );
  NAND4_X1 U14210 ( .A1(n11133), .A2(n11132), .A3(n11131), .A4(n11130), .ZN(
        n11134) );
  AOI22_X1 U14211 ( .A1(n11294), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11180), 
        .B2(n13065), .ZN(n11137) );
  AOI22_X1 U14212 ( .A1(n11207), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14213 ( .A1(n11137), .A2(n11136), .ZN(n15284) );
  NOR2_X1 U14214 ( .A1(n11185), .A2(n15972), .ZN(n11153) );
  AOI22_X1 U14215 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14216 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U14217 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11138) );
  AND2_X1 U14218 ( .A1(n11139), .A2(n11138), .ZN(n11142) );
  AOI22_X1 U14219 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10382), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U14220 ( .A1(n10431), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11140) );
  NAND4_X1 U14221 ( .A1(n11143), .A2(n11142), .A3(n11141), .A4(n11140), .ZN(
        n11149) );
  AOI22_X1 U14222 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14223 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11146) );
  AOI22_X1 U14224 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U14225 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11144) );
  NAND4_X1 U14226 ( .A1(n11147), .A2(n11146), .A3(n11145), .A4(n11144), .ZN(
        n11148) );
  INV_X1 U14227 ( .A(n12226), .ZN(n13143) );
  OAI22_X1 U14228 ( .A1(n11210), .A2(n11151), .B1(n11150), .B2(n13143), .ZN(
        n11152) );
  AOI211_X1 U14229 ( .C1(n11207), .C2(P2_EAX_REG_12__SCAN_IN), .A(n11153), .B(
        n11152), .ZN(n13150) );
  AOI22_X1 U14230 ( .A1(n11294), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11207), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14231 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11159) );
  AOI22_X1 U14232 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11155) );
  NAND2_X1 U14233 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11154) );
  AND2_X1 U14234 ( .A1(n11155), .A2(n11154), .ZN(n11158) );
  AOI22_X1 U14235 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U14236 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11156) );
  NAND4_X1 U14237 ( .A1(n11159), .A2(n11158), .A3(n11157), .A4(n11156), .ZN(
        n11165) );
  AOI22_X1 U14238 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14239 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14240 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14241 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11160) );
  NAND4_X1 U14242 ( .A1(n11163), .A2(n11162), .A3(n11161), .A4(n11160), .ZN(
        n11164) );
  AOI22_X1 U14243 ( .A1(n11180), .A2(n13377), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11076), .ZN(n11166) );
  NAND2_X1 U14244 ( .A1(n11167), .A2(n11166), .ZN(n13179) );
  AOI22_X1 U14245 ( .A1(n11294), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11076), .ZN(n11182) );
  AOI22_X1 U14246 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11173) );
  AOI22_X1 U14247 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11169) );
  NAND2_X1 U14248 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11168) );
  AND2_X1 U14249 ( .A1(n11169), .A2(n11168), .ZN(n11172) );
  AOI22_X1 U14250 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14251 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11170) );
  NAND4_X1 U14252 ( .A1(n11173), .A2(n11172), .A3(n11171), .A4(n11170), .ZN(
        n11179) );
  AOI22_X1 U14253 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14254 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14255 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11175) );
  NAND2_X1 U14256 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11174) );
  NAND4_X1 U14257 ( .A1(n11177), .A2(n11176), .A3(n11175), .A4(n11174), .ZN(
        n11178) );
  AOI22_X1 U14258 ( .A1(n11180), .A2(n13565), .B1(n11207), .B2(
        P2_EAX_REG_15__SCAN_IN), .ZN(n11181) );
  NAND2_X1 U14259 ( .A1(n11182), .A2(n11181), .ZN(n13438) );
  NAND2_X1 U14260 ( .A1(n11294), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U14261 ( .A1(n11207), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11183) );
  INV_X1 U14262 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13608) );
  OAI222_X1 U14263 ( .A1(n11210), .A2(n19656), .B1(n11186), .B2(n13608), .C1(
        n15009), .C2(n11185), .ZN(n13606) );
  NAND2_X1 U14264 ( .A1(n11294), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14265 ( .A1(n11207), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11187) );
  AND2_X1 U14266 ( .A1(n11188), .A2(n11187), .ZN(n13680) );
  OR2_X2 U14267 ( .A1(n13681), .A2(n13680), .ZN(n14855) );
  NAND2_X1 U14268 ( .A1(n11294), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14269 ( .A1(n11207), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14270 ( .A1(n11207), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11191) );
  OAI21_X1 U14271 ( .B1(n19661), .B2(n11210), .A(n11191), .ZN(n15173) );
  AOI22_X1 U14272 ( .A1(n11207), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11192) );
  OAI21_X1 U14273 ( .B1(n20723), .B2(n11210), .A(n11192), .ZN(n12565) );
  NAND2_X1 U14274 ( .A1(n11294), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14275 ( .A1(n11207), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U14276 ( .A1(n11294), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14277 ( .A1(n11207), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11195) );
  AND2_X1 U14278 ( .A1(n11196), .A2(n11195), .ZN(n12574) );
  OR2_X2 U14279 ( .A1(n9645), .A2(n12574), .ZN(n14831) );
  NAND2_X1 U14280 ( .A1(n11294), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14281 ( .A1(n11207), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11197) );
  NOR2_X2 U14282 ( .A1(n14831), .A2(n14832), .ZN(n14830) );
  AOI22_X1 U14283 ( .A1(n11207), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11199) );
  OAI21_X1 U14284 ( .B1(n11210), .B2(n19669), .A(n11199), .ZN(n14823) );
  NAND2_X1 U14285 ( .A1(n14830), .A2(n14823), .ZN(n14825) );
  NAND2_X1 U14286 ( .A1(n11294), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14287 ( .A1(n11207), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11200) );
  NAND2_X1 U14288 ( .A1(n11294), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14289 ( .A1(n11207), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14290 ( .A1(n11207), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11205) );
  NAND2_X1 U14291 ( .A1(n11294), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11204) );
  NAND2_X1 U14292 ( .A1(n11205), .A2(n11204), .ZN(n14794) );
  AOI22_X1 U14293 ( .A1(n11207), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11206) );
  OAI21_X1 U14294 ( .B1(n11210), .B2(n20752), .A(n11206), .ZN(n14785) );
  AOI22_X1 U14295 ( .A1(n11207), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11076), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11208) );
  OAI21_X1 U14296 ( .B1(n11210), .B2(n11209), .A(n11208), .ZN(n11212) );
  OAI21_X1 U14297 ( .B1(n11211), .B2(n11212), .A(n9640), .ZN(n11275) );
  INV_X1 U14298 ( .A(n11213), .ZN(n11214) );
  NAND2_X1 U14299 ( .A1(n11214), .A2(n13248), .ZN(n13199) );
  NAND2_X1 U14300 ( .A1(n13233), .A2(n19006), .ZN(n11216) );
  AND2_X1 U14301 ( .A1(n13199), .A2(n11216), .ZN(n11217) );
  INV_X1 U14302 ( .A(n11223), .ZN(n15809) );
  AND2_X1 U14304 ( .A1(n9641), .A2(n14890), .ZN(n11224) );
  NOR2_X1 U14305 ( .A1(n10923), .A2(n11224), .ZN(n15819) );
  NAND2_X1 U14306 ( .A1(n9694), .A2(n14900), .ZN(n11225) );
  AND2_X1 U14307 ( .A1(n9641), .A2(n11225), .ZN(n15831) );
  OR2_X1 U14308 ( .A1(n11228), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11227) );
  AND2_X1 U14309 ( .A1(n11227), .A2(n9694), .ZN(n15842) );
  INV_X1 U14310 ( .A(n11228), .ZN(n11231) );
  NAND2_X1 U14311 ( .A1(n11234), .A2(n11229), .ZN(n11230) );
  NAND2_X1 U14312 ( .A1(n11231), .A2(n11230), .ZN(n14919) );
  INV_X1 U14313 ( .A(n14919), .ZN(n15851) );
  INV_X1 U14314 ( .A(n11234), .ZN(n11235) );
  AOI21_X1 U14315 ( .B1(n14928), .B2(n11233), .A(n11235), .ZN(n14926) );
  INV_X1 U14316 ( .A(n11236), .ZN(n11237) );
  OAI21_X1 U14317 ( .B1(n11237), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n11233), .ZN(n14943) );
  INV_X1 U14318 ( .A(n14943), .ZN(n15573) );
  OAI21_X1 U14319 ( .B1(n11238), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n11236), .ZN(n11239) );
  INV_X1 U14320 ( .A(n11239), .ZN(n14970) );
  INV_X1 U14321 ( .A(n11240), .ZN(n11243) );
  INV_X1 U14322 ( .A(n11238), .ZN(n11241) );
  OAI21_X1 U14323 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11243), .A(
        n11241), .ZN(n14986) );
  INV_X1 U14324 ( .A(n14986), .ZN(n18624) );
  INV_X1 U14325 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11244) );
  INV_X1 U14326 ( .A(n11242), .ZN(n11247) );
  AOI21_X1 U14327 ( .B1(n11244), .B2(n11247), .A(n11243), .ZN(n18632) );
  NAND2_X1 U14328 ( .A1(n10596), .A2(n11245), .ZN(n11246) );
  NAND2_X1 U14329 ( .A1(n11247), .A2(n11246), .ZN(n15007) );
  INV_X1 U14330 ( .A(n15007), .ZN(n18642) );
  INV_X1 U14331 ( .A(n11248), .ZN(n11250) );
  AOI21_X1 U14332 ( .B1(n15031), .B2(n11250), .A(n11249), .ZN(n18664) );
  AND2_X1 U14333 ( .A1(n11251), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11267) );
  OAI21_X1 U14334 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11267), .A(
        n11252), .ZN(n18688) );
  INV_X1 U14335 ( .A(n18688), .ZN(n11269) );
  INV_X1 U14336 ( .A(n11251), .ZN(n11268) );
  OAI21_X1 U14337 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11253), .A(
        n11268), .ZN(n18710) );
  INV_X1 U14338 ( .A(n18710), .ZN(n11266) );
  OAI21_X1 U14339 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11254), .A(
        n11255), .ZN(n15921) );
  INV_X1 U14340 ( .A(n15921), .ZN(n18734) );
  INV_X1 U14341 ( .A(n11257), .ZN(n11258) );
  AOI21_X1 U14342 ( .B1(n18756), .B2(n11256), .A(n11258), .ZN(n18753) );
  AOI21_X1 U14343 ( .B1(n15954), .B2(n11259), .A(n11260), .ZN(n18782) );
  NOR2_X1 U14344 ( .A1(n13547), .A2(n11261), .ZN(n11264) );
  AOI21_X1 U14345 ( .B1(n13547), .B2(n11261), .A(n11264), .ZN(n18814) );
  AOI21_X1 U14346 ( .B1(n12684), .B2(n11262), .A(n11263), .ZN(n13522) );
  AOI22_X1 U14347 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18596), .ZN(n18837) );
  AOI22_X1 U14348 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n12684), .B2(n18596), .ZN(
        n12545) );
  NAND2_X1 U14349 ( .A1(n18837), .A2(n12545), .ZN(n13520) );
  NOR2_X1 U14350 ( .A1(n13522), .A2(n13520), .ZN(n13571) );
  OAI21_X1 U14351 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11263), .A(
        n11261), .ZN(n13572) );
  NAND2_X1 U14352 ( .A1(n13571), .A2(n13572), .ZN(n18810) );
  NOR2_X1 U14353 ( .A1(n18814), .A2(n18810), .ZN(n18792) );
  OAI21_X1 U14354 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11264), .A(
        n11259), .ZN(n18794) );
  NAND2_X1 U14355 ( .A1(n18792), .A2(n18794), .ZN(n18780) );
  NOR2_X1 U14356 ( .A1(n18782), .A2(n18780), .ZN(n18763) );
  OAI21_X1 U14357 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11260), .A(
        n11256), .ZN(n18766) );
  NAND2_X1 U14358 ( .A1(n18763), .A2(n18766), .ZN(n18751) );
  NOR2_X1 U14359 ( .A1(n18753), .A2(n18751), .ZN(n18743) );
  AOI21_X1 U14360 ( .B1(n18741), .B2(n11257), .A(n11254), .ZN(n15923) );
  INV_X1 U14361 ( .A(n15923), .ZN(n18744) );
  NAND2_X1 U14362 ( .A1(n18743), .A2(n18744), .ZN(n18732) );
  NOR2_X1 U14363 ( .A1(n18734), .A2(n18732), .ZN(n18719) );
  AOI21_X1 U14364 ( .B1(n15914), .B2(n11255), .A(n11253), .ZN(n18720) );
  INV_X1 U14365 ( .A(n18720), .ZN(n11265) );
  NAND2_X1 U14366 ( .A1(n18719), .A2(n11265), .ZN(n18708) );
  NOR2_X1 U14367 ( .A1(n11266), .A2(n18708), .ZN(n18699) );
  INV_X1 U14368 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18697) );
  AOI21_X1 U14369 ( .B1(n18697), .B2(n11268), .A(n11267), .ZN(n15903) );
  INV_X1 U14370 ( .A(n15903), .ZN(n18701) );
  NAND2_X1 U14371 ( .A1(n18699), .A2(n18701), .ZN(n18686) );
  NOR2_X1 U14372 ( .A1(n11269), .A2(n18686), .ZN(n18675) );
  AOI21_X1 U14373 ( .B1(n11252), .B2(n18685), .A(n11248), .ZN(n15044) );
  INV_X1 U14374 ( .A(n15044), .ZN(n18678) );
  NAND2_X1 U14375 ( .A1(n18675), .A2(n18678), .ZN(n18662) );
  NOR2_X1 U14376 ( .A1(n18664), .A2(n18662), .ZN(n18651) );
  OAI21_X1 U14377 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n11249), .A(
        n11245), .ZN(n18661) );
  NOR2_X1 U14378 ( .A1(n14970), .A2(n12561), .ZN(n12560) );
  NOR2_X1 U14379 ( .A1(n18764), .A2(n12560), .ZN(n15572) );
  NOR2_X1 U14380 ( .A1(n15573), .A2(n15572), .ZN(n15571) );
  NOR2_X1 U14381 ( .A1(n18764), .A2(n15850), .ZN(n15843) );
  NOR2_X1 U14382 ( .A1(n15842), .A2(n15843), .ZN(n15841) );
  NOR2_X1 U14383 ( .A1(n18676), .A2(n15841), .ZN(n15830) );
  NOR2_X1 U14384 ( .A1(n15831), .A2(n15830), .ZN(n15829) );
  INV_X1 U14385 ( .A(n10922), .ZN(n11272) );
  INV_X1 U14386 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11271) );
  AOI21_X1 U14387 ( .B1(n11272), .B2(n11271), .A(n11270), .ZN(n15794) );
  XNOR2_X1 U14388 ( .A(n11270), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15788) );
  XNOR2_X1 U14389 ( .A(n11273), .B(n15788), .ZN(n11274) );
  NOR4_X1 U14390 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n10711), .ZN(n11284) );
  NAND2_X1 U14391 ( .A1(n11274), .A2(n18819), .ZN(n11293) );
  NAND2_X1 U14392 ( .A1(n11282), .A2(n12613), .ZN(n12550) );
  NOR2_X1 U14393 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12603), .ZN(n11276) );
  INV_X1 U14394 ( .A(n19617), .ZN(n19633) );
  NOR2_X1 U14395 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19633), .ZN(n11277) );
  INV_X1 U14396 ( .A(n11276), .ZN(n13271) );
  AND2_X1 U14397 ( .A1(n18958), .A2(n13271), .ZN(n15785) );
  INV_X1 U14398 ( .A(n11277), .ZN(n11280) );
  INV_X1 U14399 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15861) );
  NAND2_X1 U14400 ( .A1(n11280), .A2(n15861), .ZN(n11278) );
  NOR2_X1 U14401 ( .A1(n12580), .A2(n11278), .ZN(n11279) );
  OR2_X2 U14402 ( .A1(n15785), .A2(n11279), .ZN(n18803) );
  AND2_X1 U14403 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n11280), .ZN(n11281) );
  NAND2_X1 U14404 ( .A1(n13233), .A2(n11282), .ZN(n12585) );
  NAND2_X1 U14405 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13409), .ZN(n13494) );
  NOR2_X1 U14406 ( .A1(n11283), .A2(n13494), .ZN(n16001) );
  NAND2_X1 U14407 ( .A1(n18970), .A2(n18811), .ZN(n11285) );
  AOI22_X1 U14408 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18802), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18807), .ZN(n11286) );
  OAI21_X1 U14409 ( .B1(n11287), .B2(n18822), .A(n11286), .ZN(n11288) );
  AOI21_X1 U14410 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n18803), .A(n11288), .ZN(
        n11289) );
  NAND2_X1 U14411 ( .A1(n11293), .A2(n11292), .ZN(P2_U2825) );
  AOI222_X1 U14412 ( .A1(n11294), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11207), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11076), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11295) );
  XNOR2_X2 U14413 ( .A(n9640), .B(n11295), .ZN(n15786) );
  NAND3_X1 U14414 ( .A1(n11296), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15267), .ZN(n11301) );
  INV_X1 U14415 ( .A(n11297), .ZN(n11300) );
  INV_X2 U14416 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11305) );
  AND2_X2 U14417 ( .A1(n11305), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11307) );
  AND2_X2 U14418 ( .A1(n11307), .A2(n11314), .ZN(n11332) );
  NOR2_X4 U14419 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13116) );
  AND2_X2 U14420 ( .A1(n11314), .A2(n13116), .ZN(n11462) );
  AOI22_X1 U14421 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11311) );
  NOR2_X2 U14422 ( .A1(n11306), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11313) );
  AOI22_X1 U14423 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11563), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11310) );
  NOR2_X4 U14424 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11316) );
  AND2_X2 U14425 ( .A1(n11316), .A2(n13115), .ZN(n11483) );
  AOI22_X1 U14426 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14427 ( .A1(n11342), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11308) );
  INV_X1 U14428 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11312) );
  AND2_X2 U14429 ( .A1(n11312), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11315) );
  AOI22_X1 U14430 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11468), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11320) );
  AND2_X2 U14431 ( .A1(n11314), .A2(n13115), .ZN(n12046) );
  AOI22_X1 U14432 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14433 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11318) );
  AND2_X2 U14434 ( .A1(n13116), .A2(n11316), .ZN(n11470) );
  AOI22_X1 U14435 ( .A1(n11377), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11317) );
  NAND2_X2 U14436 ( .A1(n11321), .A2(n9646), .ZN(n11437) );
  AOI22_X1 U14437 ( .A1(n11468), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14438 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11377), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14439 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14440 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11322) );
  NAND4_X1 U14441 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11331) );
  AOI22_X1 U14442 ( .A1(n11342), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11563), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14443 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11351), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14444 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14445 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11470), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11326) );
  NAND4_X1 U14446 ( .A1(n11329), .A2(n11328), .A3(n11327), .A4(n11326), .ZN(
        n11330) );
  AOI22_X1 U14447 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11342), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14448 ( .A1(n11468), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12046), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14449 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14450 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14451 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11563), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14452 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11377), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14453 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14454 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14455 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14456 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11563), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14457 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14458 ( .A1(n11342), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14459 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11468), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14460 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14461 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14462 ( .A1(n11377), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14463 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11468), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14464 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11351), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14465 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14466 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11352) );
  NAND4_X1 U14467 ( .A1(n11355), .A2(n11354), .A3(n11353), .A4(n11352), .ZN(
        n11361) );
  AOI22_X1 U14468 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14469 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11563), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14470 ( .A1(n11342), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14471 ( .A1(n11377), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11356) );
  NAND4_X1 U14472 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11360) );
  AOI22_X1 U14473 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11468), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14474 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11362) );
  NAND2_X1 U14475 ( .A1(n11363), .A2(n11362), .ZN(n11367) );
  AOI22_X1 U14476 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14477 ( .A1(n11377), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11364) );
  NAND2_X1 U14478 ( .A1(n11365), .A2(n11364), .ZN(n11366) );
  AOI22_X1 U14479 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14480 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11563), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14481 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11369) );
  AOI22_X1 U14482 ( .A1(n11342), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11368) );
  NAND2_X1 U14483 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11376) );
  NAND2_X1 U14484 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11375) );
  NAND2_X1 U14485 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11374) );
  NAND2_X1 U14486 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11373) );
  NAND2_X1 U14487 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11381) );
  NAND2_X1 U14488 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11380) );
  NAND2_X1 U14489 ( .A1(n11377), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11379) );
  NAND2_X1 U14490 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11378) );
  NAND2_X1 U14491 ( .A1(n11468), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11385) );
  NAND2_X1 U14492 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U14493 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11383) );
  NAND2_X1 U14494 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11382) );
  NAND2_X1 U14495 ( .A1(n11563), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11389) );
  NAND2_X1 U14496 ( .A1(n11342), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U14497 ( .A1(n11986), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11387) );
  NAND2_X1 U14498 ( .A1(n11483), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11386) );
  INV_X1 U14499 ( .A(n12156), .ZN(n11415) );
  NAND2_X1 U14500 ( .A1(n12072), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11397) );
  NAND2_X1 U14501 ( .A1(n11468), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11396) );
  NAND2_X1 U14502 ( .A1(n11377), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11395) );
  NAND2_X1 U14503 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11394) );
  NAND2_X1 U14504 ( .A1(n11342), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11401) );
  NAND2_X1 U14505 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11400) );
  NAND2_X1 U14506 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11399) );
  NAND2_X1 U14507 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11398) );
  NAND2_X1 U14508 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11406) );
  NAND2_X1 U14509 ( .A1(n11563), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11405) );
  NAND2_X1 U14510 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11404) );
  NAND2_X1 U14511 ( .A1(n11402), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11403) );
  NAND2_X1 U14512 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11410) );
  NAND2_X1 U14513 ( .A1(n11498), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11409) );
  NAND2_X1 U14514 ( .A1(n11483), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11408) );
  NAND2_X1 U14515 ( .A1(n11986), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11407) );
  NAND4_X2 U14516 ( .A1(n11414), .A2(n11413), .A3(n11412), .A4(n11411), .ZN(
        n11424) );
  NAND2_X1 U14517 ( .A1(n11415), .A2(n11424), .ZN(n11423) );
  INV_X1 U14518 ( .A(n11417), .ZN(n11416) );
  NAND2_X1 U14519 ( .A1(n11421), .A2(n11630), .ZN(n11436) );
  INV_X1 U14520 ( .A(n11436), .ZN(n11441) );
  NAND2_X1 U14521 ( .A1(n11416), .A2(n11441), .ZN(n11818) );
  NAND2_X1 U14522 ( .A1(n11818), .A2(n19954), .ZN(n11420) );
  INV_X2 U14523 ( .A(n11630), .ZN(n19968) );
  NAND3_X1 U14524 ( .A1(n9937), .A2(n11421), .A3(n19968), .ZN(n11419) );
  NAND2_X1 U14525 ( .A1(n11426), .A2(n11417), .ZN(n11418) );
  NOR2_X1 U14526 ( .A1(n11432), .A2(n19932), .ZN(n11422) );
  NAND2_X1 U14527 ( .A1(n11423), .A2(n12766), .ZN(n12898) );
  XNOR2_X1 U14528 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12696) );
  NOR2_X1 U14529 ( .A1(n19932), .A2(n11424), .ZN(n11425) );
  NAND3_X1 U14530 ( .A1(n11425), .A2(n12116), .A3(n13124), .ZN(n12786) );
  NOR2_X1 U14531 ( .A1(n12898), .A2(n11429), .ZN(n11515) );
  NAND2_X1 U14532 ( .A1(n11432), .A2(n19949), .ZN(n11430) );
  AND2_X2 U14533 ( .A1(n11431), .A2(n11430), .ZN(n12785) );
  INV_X1 U14534 ( .A(n13124), .ZN(n12778) );
  NAND2_X1 U14535 ( .A1(n12785), .A2(n12778), .ZN(n11444) );
  INV_X1 U14536 ( .A(n11432), .ZN(n12111) );
  AND2_X1 U14537 ( .A1(n19949), .A2(n19932), .ZN(n11433) );
  AOI21_X2 U14538 ( .B1(n12111), .B2(n12643), .A(n11433), .ZN(n11458) );
  NAND2_X1 U14539 ( .A1(n11434), .A2(n19932), .ZN(n13342) );
  NAND2_X2 U14540 ( .A1(n13342), .A2(n11448), .ZN(n13081) );
  INV_X1 U14541 ( .A(n12881), .ZN(n12159) );
  NAND2_X1 U14542 ( .A1(n13081), .A2(n12159), .ZN(n11435) );
  AND2_X2 U14543 ( .A1(n11458), .A2(n11435), .ZN(n12905) );
  OR2_X1 U14544 ( .A1(n13073), .A2(n11437), .ZN(n11440) );
  NAND2_X1 U14545 ( .A1(n12116), .A2(n19968), .ZN(n11439) );
  AND2_X1 U14546 ( .A1(n11439), .A2(n11438), .ZN(n11455) );
  NAND2_X1 U14547 ( .A1(n11441), .A2(n12756), .ZN(n11442) );
  NAND2_X1 U14548 ( .A1(n11442), .A2(n11437), .ZN(n11451) );
  NAND2_X1 U14549 ( .A1(n13280), .A2(n13289), .ZN(n13293) );
  NAND4_X1 U14550 ( .A1(n12905), .A2(n12779), .A3(n11451), .A4(n13293), .ZN(
        n11443) );
  AOI21_X1 U14551 ( .B1(n11444), .B2(n13280), .A(n11443), .ZN(n11445) );
  INV_X1 U14552 ( .A(n15611), .ZN(n11559) );
  NAND2_X1 U14553 ( .A1(n15606), .A2(n20357), .ZN(n20611) );
  MUX2_X1 U14554 ( .A(n11559), .B(n11560), .S(n20397), .Z(n11446) );
  INV_X1 U14555 ( .A(n12785), .ZN(n11453) );
  NAND2_X1 U14556 ( .A1(n13073), .A2(n19954), .ZN(n11449) );
  NAND2_X1 U14557 ( .A1(n11449), .A2(n13977), .ZN(n11450) );
  NAND2_X1 U14558 ( .A1(n11451), .A2(n11450), .ZN(n11452) );
  MUX2_X1 U14559 ( .A(n11453), .B(n11452), .S(n13309), .Z(n11454) );
  INV_X1 U14560 ( .A(n11454), .ZN(n11460) );
  AND2_X1 U14561 ( .A1(n20357), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13284) );
  AND2_X1 U14562 ( .A1(n13293), .A2(n13284), .ZN(n11457) );
  OR2_X1 U14563 ( .A1(n12778), .A2(n19968), .ZN(n12903) );
  INV_X1 U14564 ( .A(n11455), .ZN(n11456) );
  NAND2_X1 U14565 ( .A1(n11456), .A2(n19932), .ZN(n12758) );
  INV_X1 U14566 ( .A(n11462), .ZN(n11579) );
  AOI22_X1 U14567 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11467) );
  AOI22_X1 U14568 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11466) );
  INV_X1 U14569 ( .A(n11498), .ZN(n11477) );
  AOI22_X1 U14570 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12080), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14571 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11464) );
  NAND4_X1 U14572 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(
        n11476) );
  AOI22_X1 U14573 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12082), .B1(
        n12051), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14574 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11968), .B1(
        n12046), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14576 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n11469), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14577 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11916), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11471) );
  NAND4_X1 U14578 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n11475) );
  NAND2_X1 U14579 ( .A1(n12901), .A2(n11681), .ZN(n11491) );
  AOI22_X1 U14580 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14581 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14582 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14583 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14584 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11490) );
  AOI22_X1 U14585 ( .A1(n11463), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11469), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14586 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12046), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11487) );
  INV_X1 U14587 ( .A(n11483), .ZN(n11539) );
  AOI22_X1 U14588 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14589 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11485) );
  NAND4_X1 U14590 ( .A1(n11488), .A2(n11487), .A3(n11486), .A4(n11485), .ZN(
        n11489) );
  MUX2_X1 U14591 ( .A(n13656), .B(n11491), .S(n13048), .Z(n11492) );
  INV_X1 U14592 ( .A(n11492), .ZN(n11493) );
  INV_X1 U14593 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11495) );
  AOI21_X1 U14594 ( .B1(n13280), .B2(n13048), .A(n15614), .ZN(n11494) );
  OAI211_X1 U14595 ( .C1(n12757), .C2(n11495), .A(n11494), .B(n13656), .ZN(
        n11629) );
  NAND2_X1 U14596 ( .A1(n12901), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11550) );
  INV_X1 U14597 ( .A(n11550), .ZN(n11520) );
  NAND2_X1 U14598 ( .A1(n13280), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11551) );
  INV_X1 U14599 ( .A(n11551), .ZN(n11509) );
  AOI22_X1 U14600 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14601 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14602 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14603 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11499) );
  NAND4_X1 U14604 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11508) );
  AOI22_X1 U14605 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14606 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14607 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14608 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11503) );
  NAND4_X1 U14609 ( .A1(n11506), .A2(n11505), .A3(n11504), .A4(n11503), .ZN(
        n11507) );
  AOI22_X1 U14610 ( .A1(n11520), .A2(n11681), .B1(n11509), .B2(n13049), .ZN(
        n11511) );
  NAND2_X1 U14611 ( .A1(n12138), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11510) );
  INV_X1 U14612 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11512) );
  NAND2_X1 U14613 ( .A1(n20467), .A2(n20397), .ZN(n20351) );
  NAND2_X1 U14614 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20317) );
  NAND2_X1 U14615 ( .A1(n20351), .A2(n20317), .ZN(n20275) );
  OR2_X1 U14616 ( .A1(n15611), .A2(n20467), .ZN(n11528) );
  OAI21_X1 U14617 ( .B1(n12938), .B2(n20275), .A(n11528), .ZN(n11513) );
  INV_X1 U14618 ( .A(n11513), .ZN(n11514) );
  INV_X1 U14619 ( .A(n11515), .ZN(n11516) );
  OR2_X2 U14620 ( .A1(n20050), .A2(n11519), .ZN(n20399) );
  NAND2_X1 U14621 ( .A1(n11520), .A2(n13049), .ZN(n11521) );
  OAI21_X2 U14622 ( .B1(n13879), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11521), 
        .ZN(n11522) );
  NAND2_X1 U14623 ( .A1(n11621), .A2(n12880), .ZN(n11527) );
  INV_X1 U14624 ( .A(n11523), .ZN(n11524) );
  INV_X1 U14625 ( .A(n11614), .ZN(n11556) );
  INV_X1 U14626 ( .A(n11528), .ZN(n11531) );
  INV_X1 U14627 ( .A(n11529), .ZN(n11530) );
  OAI21_X1 U14628 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11531), .A(
        n11530), .ZN(n11532) );
  NAND2_X1 U14629 ( .A1(n11533), .A2(n11532), .ZN(n11538) );
  XNOR2_X1 U14630 ( .A(n20317), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19940) );
  NAND2_X1 U14631 ( .A1(n11560), .A2(n19940), .ZN(n11535) );
  AOI22_X1 U14632 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14633 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14634 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14635 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11540) );
  NAND4_X1 U14636 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11549) );
  AOI22_X1 U14637 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14638 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14639 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14640 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U14641 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  INV_X1 U14642 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11552) );
  OAI22_X1 U14643 ( .A1(n12145), .A2(n11552), .B1(n11551), .B2(n13051), .ZN(
        n11553) );
  INV_X1 U14644 ( .A(n11553), .ZN(n11554) );
  OAI21_X1 U14645 ( .B1(n20317), .B2(n20220), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11558) );
  INV_X1 U14646 ( .A(n20317), .ZN(n20465) );
  NAND2_X1 U14647 ( .A1(n20276), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20150) );
  INV_X1 U14648 ( .A(n20150), .ZN(n11557) );
  NAND2_X1 U14649 ( .A1(n20465), .A2(n11557), .ZN(n20206) );
  NAND2_X1 U14650 ( .A1(n11558), .A2(n20206), .ZN(n20222) );
  AOI22_X1 U14651 ( .A1(n11560), .A2(n20222), .B1(n11559), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11561) );
  INV_X1 U14652 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14653 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11568) );
  INV_X1 U14654 ( .A(n11563), .ZN(n11564) );
  INV_X2 U14655 ( .A(n11564), .ZN(n12074) );
  AOI22_X1 U14656 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14657 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14658 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11565) );
  NAND4_X1 U14659 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n11574) );
  AOI22_X1 U14660 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14661 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14662 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14663 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11569) );
  NAND4_X1 U14664 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(
        n11573) );
  INV_X1 U14665 ( .A(n13089), .ZN(n11575) );
  OAI22_X1 U14666 ( .A1(n11576), .A2(n12145), .B1(n12118), .B2(n11575), .ZN(
        n11577) );
  INV_X1 U14667 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14668 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14669 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11582) );
  INV_X2 U14670 ( .A(n11477), .ZN(n12080) );
  AOI22_X1 U14671 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14672 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11580) );
  NAND4_X1 U14673 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11590) );
  AOI22_X1 U14674 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14675 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14676 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14677 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U14678 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11589) );
  OR2_X1 U14679 ( .A1(n12118), .A2(n13323), .ZN(n11591) );
  OAI21_X1 U14680 ( .B1(n12145), .B2(n11592), .A(n11591), .ZN(n11645) );
  INV_X1 U14681 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14682 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14683 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14684 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14685 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11593) );
  NAND4_X1 U14686 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n11602) );
  AOI22_X1 U14687 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14688 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14689 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14690 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11597) );
  NAND4_X1 U14691 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n11601) );
  OR2_X1 U14692 ( .A1(n12118), .A2(n13327), .ZN(n11603) );
  OAI21_X1 U14693 ( .B1(n12145), .B2(n11604), .A(n11603), .ZN(n11606) );
  INV_X1 U14694 ( .A(n11606), .ZN(n11605) );
  NAND2_X1 U14695 ( .A1(n11607), .A2(n11605), .ZN(n11608) );
  INV_X2 U14696 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11609) );
  INV_X1 U14697 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11611) );
  NAND2_X1 U14698 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11615) );
  XNOR2_X1 U14699 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B(n11673), .ZN(
        n19812) );
  AOI22_X1 U14700 ( .A1(n12096), .A2(n19812), .B1(n12097), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11610) );
  OAI21_X1 U14701 ( .B1(n10121), .B2(n11611), .A(n11610), .ZN(n11612) );
  XNOR2_X1 U14702 ( .A(n11614), .B(n11613), .ZN(n13047) );
  NAND2_X1 U14703 ( .A1(n13047), .A2(n11800), .ZN(n11620) );
  NAND2_X1 U14704 ( .A1(n11427), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11641) );
  NAND2_X1 U14705 ( .A1(n12098), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11617) );
  OAI21_X1 U14706 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n11615), .ZN(n13354) );
  OAI21_X1 U14707 ( .B1(n13354), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n11609), 
        .ZN(n11616) );
  OAI211_X1 U14708 ( .C1(n11641), .C2(n13112), .A(n11617), .B(n11616), .ZN(
        n11618) );
  INV_X1 U14709 ( .A(n11618), .ZN(n11619) );
  NAND2_X1 U14710 ( .A1(n12097), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13075) );
  NAND2_X1 U14711 ( .A1(n13138), .A2(n11800), .ZN(n11626) );
  INV_X2 U14712 ( .A(n10121), .ZN(n12098) );
  AOI22_X1 U14713 ( .A1(n12098), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11609), .ZN(n11624) );
  INV_X1 U14714 ( .A(n11641), .ZN(n11647) );
  NAND2_X1 U14715 ( .A1(n11647), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11623) );
  AND2_X1 U14716 ( .A1(n11624), .A2(n11623), .ZN(n11625) );
  NAND2_X1 U14717 ( .A1(n11626), .A2(n11625), .ZN(n12831) );
  AOI21_X1 U14718 ( .B1(n20009), .B2(n11630), .A(n11609), .ZN(n12933) );
  NAND2_X1 U14719 ( .A1(n11609), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11633) );
  NAND2_X1 U14720 ( .A1(n12098), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11632) );
  OAI211_X1 U14721 ( .C1(n11641), .C2(n12794), .A(n11633), .B(n11632), .ZN(
        n11634) );
  AOI21_X1 U14722 ( .B1(n11631), .B2(n11800), .A(n11634), .ZN(n12932) );
  MUX2_X1 U14723 ( .A(n12933), .B(n12096), .S(n12932), .Z(n12830) );
  NAND2_X1 U14724 ( .A1(n12831), .A2(n12830), .ZN(n12864) );
  NAND2_X1 U14725 ( .A1(n12862), .A2(n13075), .ZN(n11644) );
  INV_X1 U14726 ( .A(n11800), .ZN(n11762) );
  OAI21_X1 U14727 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11638), .A(
        n11649), .ZN(n13370) );
  AOI22_X1 U14728 ( .A1(n12096), .A2(n13370), .B1(n12097), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11640) );
  NAND2_X1 U14729 ( .A1(n12098), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11639) );
  OAI211_X1 U14730 ( .C1(n11641), .C2(n11305), .A(n11640), .B(n11639), .ZN(
        n11642) );
  INV_X1 U14731 ( .A(n11642), .ZN(n11643) );
  OAI21_X1 U14732 ( .B1(n13137), .B2(n11762), .A(n11643), .ZN(n13077) );
  NAND2_X1 U14733 ( .A1(n11644), .A2(n13077), .ZN(n13078) );
  XNOR2_X1 U14734 ( .A(n11646), .B(n11645), .ZN(n13158) );
  NAND2_X1 U14735 ( .A1(n11647), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11651) );
  AOI21_X1 U14736 ( .B1(n13433), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11648) );
  AOI21_X1 U14737 ( .B1(n12098), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11648), .ZN(
        n11650) );
  AOI21_X1 U14738 ( .B1(n13433), .B2(n11649), .A(n11673), .ZN(n19823) );
  AOI22_X1 U14739 ( .A1(n11651), .A2(n11650), .B1(n12096), .B2(n19823), .ZN(
        n11652) );
  AOI21_X1 U14740 ( .B1(n13158), .B2(n11800), .A(n11652), .ZN(n13193) );
  INV_X1 U14741 ( .A(n11671), .ZN(n11669) );
  INV_X1 U14742 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14743 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14744 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14745 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14746 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11655) );
  NAND4_X1 U14747 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(
        n11664) );
  AOI22_X1 U14748 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14749 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14750 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14751 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11659) );
  NAND4_X1 U14752 ( .A1(n11662), .A2(n11661), .A3(n11660), .A4(n11659), .ZN(
        n11663) );
  INV_X1 U14753 ( .A(n13648), .ZN(n11665) );
  OR2_X1 U14754 ( .A1(n12118), .A2(n11665), .ZN(n11666) );
  OAI21_X1 U14755 ( .B1(n12145), .B2(n11667), .A(n11666), .ZN(n11668) );
  INV_X1 U14756 ( .A(n11668), .ZN(n11670) );
  NAND2_X1 U14757 ( .A1(n11671), .A2(n11670), .ZN(n11672) );
  INV_X1 U14758 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11679) );
  INV_X1 U14759 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11676) );
  INV_X1 U14760 ( .A(n11674), .ZN(n11675) );
  NAND2_X1 U14761 ( .A1(n11676), .A2(n11675), .ZN(n11677) );
  NAND2_X1 U14762 ( .A1(n11684), .A2(n11677), .ZN(n19800) );
  INV_X2 U14763 ( .A(n12065), .ZN(n12096) );
  AOI22_X1 U14764 ( .A1(n19800), .A2(n12096), .B1(n12097), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11678) );
  OAI21_X1 U14765 ( .B1(n10121), .B2(n11679), .A(n11678), .ZN(n11680) );
  NOR2_X2 U14766 ( .A1(n13359), .A2(n13386), .ZN(n13387) );
  INV_X1 U14767 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11682) );
  OAI22_X1 U14768 ( .A1(n11682), .A2(n12145), .B1(n12118), .B2(n11681), .ZN(
        n11683) );
  NAND2_X1 U14769 ( .A1(n13646), .A2(n11800), .ZN(n11689) );
  AND2_X1 U14770 ( .A1(n11684), .A2(n19781), .ZN(n11685) );
  OR2_X1 U14771 ( .A1(n11685), .A2(n11714), .ZN(n19787) );
  NAND2_X1 U14772 ( .A1(n19787), .A2(n12096), .ZN(n11686) );
  OAI21_X1 U14773 ( .B1(n19781), .B2(n11804), .A(n11686), .ZN(n11687) );
  AOI21_X1 U14774 ( .B1(n12098), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11687), .ZN(
        n11688) );
  NAND2_X1 U14775 ( .A1(n11689), .A2(n11688), .ZN(n13472) );
  AOI22_X1 U14776 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14777 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14778 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14779 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11690) );
  NAND4_X1 U14780 ( .A1(n11693), .A2(n11692), .A3(n11691), .A4(n11690), .ZN(
        n11699) );
  AOI22_X1 U14781 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14782 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14783 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14784 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11694) );
  NAND4_X1 U14785 ( .A1(n11697), .A2(n11696), .A3(n11695), .A4(n11694), .ZN(
        n11698) );
  NOR2_X1 U14786 ( .A1(n11699), .A2(n11698), .ZN(n11703) );
  XOR2_X1 U14787 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11714), .Z(n13673) );
  INV_X1 U14788 ( .A(n13673), .ZN(n11700) );
  AOI22_X1 U14789 ( .A1(n12097), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12096), .B2(n11700), .ZN(n11702) );
  NAND2_X1 U14790 ( .A1(n12098), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11701) );
  OAI211_X1 U14791 ( .C1(n11762), .C2(n11703), .A(n11702), .B(n11701), .ZN(
        n13473) );
  INV_X1 U14792 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U14793 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14794 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14795 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14796 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11704) );
  NAND4_X1 U14797 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n11713) );
  AOI22_X1 U14798 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14799 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11469), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14800 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14801 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11708) );
  NAND4_X1 U14802 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11712) );
  OAI21_X1 U14803 ( .B1(n11713), .B2(n11712), .A(n11800), .ZN(n11717) );
  INV_X1 U14804 ( .A(n11718), .ZN(n11715) );
  XNOR2_X1 U14805 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11715), .ZN(
        n19770) );
  AOI22_X1 U14806 ( .A1(n12096), .A2(n19770), .B1(n12097), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11716) );
  OAI211_X1 U14807 ( .C1(n10121), .C2(n13600), .A(n11717), .B(n11716), .ZN(
        n13555) );
  XOR2_X1 U14808 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n11732), .Z(
        n15680) );
  AOI22_X1 U14809 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11469), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14810 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14811 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14812 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11719) );
  NAND4_X1 U14813 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11728) );
  AOI22_X1 U14814 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14815 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14816 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14817 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11723) );
  NAND4_X1 U14818 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11727) );
  OR2_X1 U14819 ( .A1(n11728), .A2(n11727), .ZN(n11729) );
  AOI22_X1 U14820 ( .A1(n11800), .A2(n11729), .B1(n12097), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11731) );
  NAND2_X1 U14821 ( .A1(n12098), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11730) );
  XNOR2_X1 U14822 ( .A(n11758), .B(n11757), .ZN(n14496) );
  INV_X1 U14823 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19864) );
  OAI22_X1 U14824 ( .A1(n10121), .A2(n19864), .B1(n11804), .B2(n11757), .ZN(
        n11733) );
  AOI21_X1 U14825 ( .B1(n14496), .B2(n12096), .A(n11733), .ZN(n11746) );
  AOI22_X1 U14826 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14827 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14828 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14829 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14830 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11743) );
  AOI22_X1 U14831 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14832 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14833 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14834 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11738) );
  NAND4_X1 U14835 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11742) );
  OR2_X1 U14836 ( .A1(n11743), .A2(n11742), .ZN(n11744) );
  NAND2_X1 U14837 ( .A1(n11800), .A2(n11744), .ZN(n13718) );
  AOI22_X1 U14838 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14839 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14840 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U14841 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11747) );
  NAND4_X1 U14842 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11756) );
  AOI22_X1 U14843 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U14844 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14845 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14846 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11751) );
  NAND4_X1 U14847 ( .A1(n11754), .A2(n11753), .A3(n11752), .A4(n11751), .ZN(
        n11755) );
  NOR2_X1 U14848 ( .A1(n11756), .A2(n11755), .ZN(n11761) );
  XNOR2_X1 U14849 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11776), .ZN(
        n15663) );
  AOI22_X1 U14850 ( .A1(n12096), .A2(n15663), .B1(n12097), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11760) );
  NAND2_X1 U14851 ( .A1(n12098), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11759) );
  OAI211_X1 U14852 ( .C1(n11762), .C2(n11761), .A(n11760), .B(n11759), .ZN(
        n13735) );
  INV_X1 U14853 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14854 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14855 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14856 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U14857 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11764) );
  NAND4_X1 U14858 ( .A1(n11767), .A2(n11766), .A3(n11765), .A4(n11764), .ZN(
        n11773) );
  AOI22_X1 U14859 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14860 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14861 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14862 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11768) );
  NAND4_X1 U14863 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n11772) );
  OAI21_X1 U14864 ( .B1(n11773), .B2(n11772), .A(n11800), .ZN(n11774) );
  OAI21_X1 U14865 ( .B1(n11804), .B2(n11775), .A(n11774), .ZN(n11778) );
  XNOR2_X1 U14866 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11779), .ZN(
        n15657) );
  NOR2_X1 U14867 ( .A1(n15657), .A2(n12065), .ZN(n11777) );
  AOI211_X1 U14868 ( .C1(n12098), .C2(P1_EAX_REG_13__SCAN_IN), .A(n11778), .B(
        n11777), .ZN(n14199) );
  INV_X1 U14869 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14164) );
  XNOR2_X1 U14870 ( .A(n11805), .B(n14164), .ZN(n14162) );
  AOI22_X1 U14871 ( .A1(n12098), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n12097), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14872 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14873 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14874 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14875 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11780) );
  NAND4_X1 U14876 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11789) );
  AOI22_X1 U14877 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14878 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14879 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14880 ( .A1(n11484), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U14881 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11788) );
  OAI21_X1 U14882 ( .B1(n11789), .B2(n11788), .A(n11800), .ZN(n11790) );
  OAI211_X1 U14883 ( .C1(n14162), .C2(n12065), .A(n11791), .B(n11790), .ZN(
        n14159) );
  AOI22_X1 U14884 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U14885 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9597), .B1(
        n11469), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14886 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12079), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14887 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12082), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11792) );
  NAND4_X1 U14888 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11802) );
  AOI22_X1 U14889 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12051), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14890 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14891 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14892 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U14893 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11801) );
  OAI21_X1 U14894 ( .B1(n11802), .B2(n11801), .A(n11800), .ZN(n11803) );
  OAI21_X1 U14895 ( .B1(n11804), .B2(n15643), .A(n11803), .ZN(n11807) );
  XNOR2_X1 U14896 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11808), .ZN(
        n15640) );
  NOR2_X1 U14897 ( .A1(n15640), .A2(n12065), .ZN(n11806) );
  AOI211_X1 U14898 ( .C1(n12098), .C2(P1_EAX_REG_15__SCAN_IN), .A(n11807), .B(
        n11806), .ZN(n14190) );
  INV_X1 U14899 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14442) );
  XNOR2_X1 U14900 ( .A(n11838), .B(n14442), .ZN(n14451) );
  AOI21_X1 U14901 ( .B1(n14442), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11809) );
  AOI21_X1 U14902 ( .B1(n12098), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11809), .ZN(
        n11822) );
  AOI22_X1 U14903 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14904 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14905 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U14906 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11810) );
  NAND4_X1 U14907 ( .A1(n11813), .A2(n11812), .A3(n11811), .A4(n11810), .ZN(
        n11820) );
  AOI22_X1 U14908 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U14909 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11816) );
  INV_X1 U14910 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20766) );
  AOI22_X1 U14911 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14912 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11814) );
  NAND4_X1 U14913 ( .A1(n11817), .A2(n11816), .A3(n11815), .A4(n11814), .ZN(
        n11819) );
  OAI21_X1 U14914 ( .B1(n11820), .B2(n11819), .A(n12092), .ZN(n11821) );
  AOI22_X1 U14915 ( .A1(n14451), .A2(n12096), .B1(n11822), .B2(n11821), .ZN(
        n14146) );
  NAND2_X1 U14916 ( .A1(n11838), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11823) );
  XNOR2_X1 U14917 ( .A(n11823), .B(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14436) );
  AOI22_X1 U14918 ( .A1(n12098), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12097), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14919 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14920 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14921 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14922 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11824) );
  NAND4_X1 U14923 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11833) );
  AOI22_X1 U14924 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14925 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14926 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14927 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11828) );
  NAND4_X1 U14928 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(
        n11832) );
  OAI21_X1 U14929 ( .B1(n11833), .B2(n11832), .A(n12092), .ZN(n11834) );
  OAI211_X1 U14930 ( .C1(n14436), .C2(n12065), .A(n11835), .B(n11834), .ZN(
        n11836) );
  INV_X1 U14931 ( .A(n11836), .ZN(n14135) );
  AOI21_X1 U14932 ( .B1(n20756), .B2(n11839), .A(n11853), .ZN(n14426) );
  AOI21_X1 U14933 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20756), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11840) );
  AOI21_X1 U14934 ( .B1(n12098), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11840), .ZN(
        n11852) );
  AOI22_X1 U14935 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14936 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14937 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14938 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11841) );
  NAND4_X1 U14939 ( .A1(n11844), .A2(n11843), .A3(n11842), .A4(n11841), .ZN(
        n11850) );
  AOI22_X1 U14940 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12080), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14941 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14942 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14943 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11845) );
  NAND4_X1 U14944 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11849) );
  OAI21_X1 U14945 ( .B1(n11850), .B2(n11849), .A(n12092), .ZN(n11851) );
  AOI22_X1 U14946 ( .A1(n14426), .A2(n12096), .B1(n11852), .B2(n11851), .ZN(
        n14124) );
  INV_X1 U14947 ( .A(n11853), .ZN(n11854) );
  INV_X1 U14948 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U14949 ( .A1(n11854), .A2(n14114), .ZN(n11855) );
  NAND2_X1 U14950 ( .A1(n11883), .A2(n11855), .ZN(n14416) );
  INV_X1 U14951 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14248) );
  AOI22_X1 U14952 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14953 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11469), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14954 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14955 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11856) );
  NAND4_X1 U14956 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(
        n11865) );
  AOI22_X1 U14957 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14958 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14959 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14960 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11860) );
  NAND4_X1 U14961 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11864) );
  OAI21_X1 U14962 ( .B1(n11865), .B2(n11864), .A(n12092), .ZN(n11867) );
  OAI21_X1 U14963 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20429), .A(
        n11609), .ZN(n11866) );
  OAI211_X1 U14964 ( .C1(n10121), .C2(n14248), .A(n11867), .B(n11866), .ZN(
        n11868) );
  OAI21_X1 U14965 ( .B1(n14416), .B2(n12065), .A(n11868), .ZN(n14108) );
  XNOR2_X1 U14966 ( .A(n11883), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14402) );
  INV_X1 U14967 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11882) );
  AOI21_X1 U14968 ( .B1(n11882), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11869) );
  AOI21_X1 U14969 ( .B1(n12098), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11869), .ZN(
        n11881) );
  AOI22_X1 U14970 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14971 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14972 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14973 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11870) );
  NAND4_X1 U14974 ( .A1(n11873), .A2(n11872), .A3(n11871), .A4(n11870), .ZN(
        n11879) );
  AOI22_X1 U14975 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14976 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11968), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14977 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14978 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11874) );
  NAND4_X1 U14979 ( .A1(n11877), .A2(n11876), .A3(n11875), .A4(n11874), .ZN(
        n11878) );
  OAI21_X1 U14980 ( .B1(n11879), .B2(n11878), .A(n12092), .ZN(n11880) );
  AOI22_X1 U14981 ( .A1(n14402), .A2(n12096), .B1(n11881), .B2(n11880), .ZN(
        n14098) );
  NAND2_X1 U14982 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  NAND2_X1 U14983 ( .A1(n11914), .A2(n11886), .ZN(n14395) );
  INV_X1 U14984 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U14985 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14986 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14987 ( .A1(n11985), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U14988 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11887) );
  NAND4_X1 U14989 ( .A1(n11890), .A2(n11889), .A3(n11888), .A4(n11887), .ZN(
        n11896) );
  AOI22_X1 U14990 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14991 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11584), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14992 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U14993 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11891) );
  NAND4_X1 U14994 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n11895) );
  OAI21_X1 U14995 ( .B1(n11896), .B2(n11895), .A(n12092), .ZN(n11898) );
  AOI21_X1 U14996 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11609), .A(
        n12096), .ZN(n11897) );
  OAI211_X1 U14997 ( .C1(n10121), .C2(n14239), .A(n11898), .B(n11897), .ZN(
        n11899) );
  OAI21_X1 U14998 ( .B1(n14395), .B2(n12065), .A(n11899), .ZN(n14085) );
  XNOR2_X1 U14999 ( .A(n11914), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14384) );
  NOR2_X1 U15000 ( .A1(n14386), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11900) );
  AOI211_X1 U15001 ( .C1(n12098), .C2(P1_EAX_REG_22__SCAN_IN), .A(n12096), .B(
        n11900), .ZN(n11913) );
  AOI22_X1 U15002 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15003 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U15004 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U15005 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11902) );
  NAND4_X1 U15006 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n11911) );
  AOI22_X1 U15007 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U15008 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11469), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U15009 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U15010 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11906) );
  NAND4_X1 U15011 ( .A1(n11909), .A2(n11908), .A3(n11907), .A4(n11906), .ZN(
        n11910) );
  OAI21_X1 U15012 ( .B1(n11911), .B2(n11910), .A(n12092), .ZN(n11912) );
  AOI22_X1 U15013 ( .A1(n14384), .A2(n12096), .B1(n11913), .B2(n11912), .ZN(
        n14073) );
  OAI21_X1 U15014 ( .B1(n11915), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n11958), .ZN(n14377) );
  INV_X1 U15015 ( .A(n12092), .ZN(n12062) );
  AOI22_X1 U15016 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U15017 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12082), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15018 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12051), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15019 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11917) );
  NAND4_X1 U15020 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n11927) );
  AOI22_X1 U15021 ( .A1(n11921), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15022 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15023 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U15024 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11922) );
  NAND4_X1 U15025 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11926) );
  NOR2_X1 U15026 ( .A1(n11927), .A2(n11926), .ZN(n11954) );
  AOI22_X1 U15027 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U15028 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11469), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15029 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15030 ( .A1(n11478), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11928) );
  NAND4_X1 U15031 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11937) );
  AOI22_X1 U15032 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U15033 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15034 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15035 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11932) );
  NAND4_X1 U15036 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11936) );
  NOR2_X1 U15037 ( .A1(n11937), .A2(n11936), .ZN(n11953) );
  XNOR2_X1 U15038 ( .A(n11954), .B(n11953), .ZN(n11940) );
  OAI21_X1 U15039 ( .B1(n20429), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n11609), .ZN(n11939) );
  NAND2_X1 U15040 ( .A1(n12098), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n11938) );
  OAI211_X1 U15041 ( .C1(n12062), .C2(n11940), .A(n11939), .B(n11938), .ZN(
        n11941) );
  OAI21_X1 U15042 ( .B1(n14377), .B2(n12065), .A(n11941), .ZN(n14062) );
  XNOR2_X1 U15043 ( .A(n11958), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14368) );
  INV_X1 U15044 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14053) );
  NOR2_X1 U15045 ( .A1(n14053), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11942) );
  AOI211_X1 U15046 ( .C1(n12098), .C2(P1_EAX_REG_24__SCAN_IN), .A(n12096), .B(
        n11942), .ZN(n11957) );
  AOI22_X1 U15047 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11478), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U15048 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15049 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11944) );
  INV_X1 U15050 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n20790) );
  AOI22_X1 U15051 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11943) );
  NAND4_X1 U15052 ( .A1(n11946), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11952) );
  AOI22_X1 U15053 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15054 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15055 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15056 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U15057 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11951) );
  NOR2_X1 U15058 ( .A1(n11954), .A2(n11953), .ZN(n11976) );
  XOR2_X1 U15059 ( .A(n11975), .B(n11976), .Z(n11955) );
  NAND2_X1 U15060 ( .A1(n11955), .A2(n12092), .ZN(n11956) );
  AOI22_X1 U15061 ( .A1(n14368), .A2(n12096), .B1(n11957), .B2(n11956), .ZN(
        n14051) );
  INV_X1 U15062 ( .A(n11958), .ZN(n11959) );
  INV_X1 U15063 ( .A(n11960), .ZN(n11962) );
  INV_X1 U15064 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11961) );
  NAND2_X1 U15065 ( .A1(n11962), .A2(n11961), .ZN(n11963) );
  NAND2_X1 U15066 ( .A1(n12002), .A2(n11963), .ZN(n14360) );
  AOI22_X1 U15067 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15068 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12079), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15069 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15070 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11964) );
  NAND4_X1 U15071 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11974) );
  AOI22_X1 U15072 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9597), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15073 ( .A1(n11968), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15074 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U15075 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11402), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11969) );
  NAND4_X1 U15076 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11973) );
  NOR2_X1 U15077 ( .A1(n11974), .A2(n11973), .ZN(n11996) );
  NAND2_X1 U15078 ( .A1(n11976), .A2(n11975), .ZN(n11995) );
  XNOR2_X1 U15079 ( .A(n11996), .B(n11995), .ZN(n11979) );
  OAI21_X1 U15080 ( .B1(n20429), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n11609), .ZN(n11978) );
  NAND2_X1 U15081 ( .A1(n12098), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n11977) );
  OAI211_X1 U15082 ( .C1(n11979), .C2(n12062), .A(n11978), .B(n11977), .ZN(
        n11980) );
  OAI21_X1 U15083 ( .B1(n14360), .B2(n12065), .A(n11980), .ZN(n14039) );
  XNOR2_X1 U15084 ( .A(n12002), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14347) );
  INV_X1 U15085 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11981) );
  NOR2_X1 U15086 ( .A1(n11579), .A2(n11981), .ZN(n11984) );
  INV_X1 U15087 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11982) );
  OAI22_X1 U15088 ( .A1(n11477), .A2(n11982), .B1(n11539), .B2(n11576), .ZN(
        n11983) );
  AOI211_X1 U15089 ( .C1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .C2(n11985), .A(
        n11984), .B(n11983), .ZN(n11994) );
  AOI22_X1 U15090 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11986), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15091 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15092 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15093 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15094 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15095 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11987) );
  AND4_X1 U15096 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11991) );
  NAND4_X1 U15097 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n12018) );
  NOR2_X1 U15098 ( .A1(n11996), .A2(n11995), .ZN(n12019) );
  XOR2_X1 U15099 ( .A(n12018), .B(n12019), .Z(n12000) );
  INV_X1 U15100 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n11998) );
  NOR2_X1 U15101 ( .A1(n20429), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11997) );
  OAI22_X1 U15102 ( .A1(n10121), .A2(n11998), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11997), .ZN(n11999) );
  AOI21_X1 U15103 ( .B1(n12000), .B2(n12092), .A(n11999), .ZN(n12001) );
  AOI21_X1 U15104 ( .B1(n14347), .B2(n12096), .A(n12001), .ZN(n14028) );
  INV_X1 U15105 ( .A(n12002), .ZN(n12003) );
  INV_X1 U15106 ( .A(n12004), .ZN(n12006) );
  INV_X1 U15107 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12005) );
  NAND2_X1 U15108 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  NAND2_X1 U15109 ( .A1(n12040), .A2(n12007), .ZN(n14339) );
  AOI22_X1 U15110 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15111 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15112 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U15113 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12008) );
  NAND4_X1 U15114 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n12017) );
  AOI22_X1 U15115 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15116 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12046), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15117 ( .A1(n11462), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11484), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15118 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U15119 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12016) );
  NOR2_X1 U15120 ( .A1(n12017), .A2(n12016), .ZN(n12036) );
  NAND2_X1 U15121 ( .A1(n12019), .A2(n12018), .ZN(n12035) );
  XNOR2_X1 U15122 ( .A(n12036), .B(n12035), .ZN(n12022) );
  AOI21_X1 U15123 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n11609), .A(
        n12096), .ZN(n12021) );
  NAND2_X1 U15124 ( .A1(n12098), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12020) );
  OAI211_X1 U15125 ( .C1(n12022), .C2(n12062), .A(n12021), .B(n12020), .ZN(
        n12023) );
  OAI21_X1 U15126 ( .B1(n14339), .B2(n12065), .A(n12023), .ZN(n14014) );
  XNOR2_X1 U15127 ( .A(n12040), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14328) );
  INV_X1 U15128 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14330) );
  NOR2_X1 U15129 ( .A1(n14330), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12024) );
  AOI211_X1 U15130 ( .C1(n12098), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12096), .B(
        n12024), .ZN(n12039) );
  AOI22_X1 U15131 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15132 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15133 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15134 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12025) );
  NAND4_X1 U15135 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12034) );
  AOI22_X1 U15136 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12082), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15137 ( .A1(n12079), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15138 ( .A1(n11469), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15139 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12029) );
  NAND4_X1 U15140 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12033) );
  OR2_X1 U15141 ( .A1(n12034), .A2(n12033), .ZN(n12058) );
  NOR2_X1 U15142 ( .A1(n12036), .A2(n12035), .ZN(n12059) );
  XOR2_X1 U15143 ( .A(n12058), .B(n12059), .Z(n12037) );
  NAND2_X1 U15144 ( .A1(n12037), .A2(n12092), .ZN(n12038) );
  INV_X1 U15145 ( .A(n12040), .ZN(n12041) );
  INV_X1 U15146 ( .A(n12042), .ZN(n12044) );
  INV_X1 U15147 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12043) );
  NAND2_X1 U15148 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  NAND2_X1 U15149 ( .A1(n13282), .A2(n12045), .ZN(n14320) );
  AOI22_X1 U15150 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12074), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15151 ( .A1(n12046), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15152 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15153 ( .A1(n12082), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15154 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12057) );
  AOI22_X1 U15155 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15156 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15157 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15158 ( .A1(n11584), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12052) );
  NAND4_X1 U15159 ( .A1(n12055), .A2(n12054), .A3(n12053), .A4(n12052), .ZN(
        n12056) );
  NOR2_X1 U15160 ( .A1(n12057), .A2(n12056), .ZN(n12068) );
  NAND2_X1 U15161 ( .A1(n12059), .A2(n12058), .ZN(n12067) );
  XNOR2_X1 U15162 ( .A(n12068), .B(n12067), .ZN(n12063) );
  AOI21_X1 U15163 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n11609), .A(
        n12096), .ZN(n12061) );
  NAND2_X1 U15164 ( .A1(n12098), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12060) );
  OAI211_X1 U15165 ( .C1(n12063), .C2(n12062), .A(n12061), .B(n12060), .ZN(
        n12064) );
  OAI21_X1 U15166 ( .B1(n14320), .B2(n12065), .A(n12064), .ZN(n13990) );
  XNOR2_X1 U15167 ( .A(n13282), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13980) );
  INV_X1 U15168 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13281) );
  NOR2_X1 U15169 ( .A1(n13281), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12066) );
  AOI211_X1 U15170 ( .C1(n12098), .C2(P1_EAX_REG_30__SCAN_IN), .A(n12066), .B(
        n12096), .ZN(n12095) );
  NOR2_X1 U15171 ( .A1(n12068), .A2(n12067), .ZN(n12091) );
  AOI22_X1 U15172 ( .A1(n12069), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11462), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15173 ( .A1(n12071), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12070), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15174 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12072), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15175 ( .A1(n12074), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12073), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12075) );
  NAND4_X1 U15176 ( .A1(n12078), .A2(n12077), .A3(n12076), .A4(n12075), .ZN(
        n12089) );
  AOI22_X1 U15177 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12079), .B1(
        n11469), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15178 ( .A1(n12080), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11483), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15179 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n12082), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15180 ( .A1(n9597), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12083), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12084) );
  NAND4_X1 U15181 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(
        n12088) );
  NOR2_X1 U15182 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  XNOR2_X1 U15183 ( .A(n12091), .B(n12090), .ZN(n12093) );
  NAND2_X1 U15184 ( .A1(n12093), .A2(n12092), .ZN(n12094) );
  AOI22_X1 U15185 ( .A1(n12098), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12097), .ZN(n12099) );
  INV_X1 U15186 ( .A(n12099), .ZN(n12100) );
  NAND2_X1 U15187 ( .A1(n20467), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12102) );
  NAND2_X1 U15188 ( .A1(n11512), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12101) );
  NAND2_X1 U15189 ( .A1(n12102), .A2(n12101), .ZN(n12119) );
  NAND2_X1 U15190 ( .A1(n12789), .A2(n20397), .ZN(n12120) );
  NAND2_X1 U15191 ( .A1(n12121), .A2(n12102), .ZN(n12108) );
  NAND2_X1 U15192 ( .A1(n13112), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12103) );
  NAND2_X1 U15193 ( .A1(n12108), .A2(n12107), .ZN(n12106) );
  NAND2_X1 U15194 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12147), .ZN(
        n12105) );
  INV_X1 U15195 ( .A(n12118), .ZN(n12148) );
  OAI21_X1 U15196 ( .B1(n12108), .B2(n12107), .A(n12106), .ZN(n12163) );
  INV_X1 U15197 ( .A(n12163), .ZN(n12109) );
  NAND2_X1 U15198 ( .A1(n12148), .A2(n12109), .ZN(n12136) );
  NAND2_X1 U15199 ( .A1(n12979), .A2(n11421), .ZN(n12126) );
  INV_X1 U15200 ( .A(n12126), .ZN(n12110) );
  OAI21_X1 U15201 ( .B1(n12789), .B2(n20397), .A(n12120), .ZN(n12113) );
  NOR2_X1 U15202 ( .A1(n12118), .A2(n12113), .ZN(n12115) );
  NAND2_X1 U15203 ( .A1(n19932), .A2(n12111), .ZN(n12112) );
  NAND2_X1 U15204 ( .A1(n10116), .A2(n12112), .ZN(n12114) );
  OAI22_X1 U15205 ( .A1(n12150), .A2(n12115), .B1(n12114), .B2(n12113), .ZN(
        n12131) );
  NAND2_X1 U15206 ( .A1(n12116), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12117) );
  NAND2_X1 U15207 ( .A1(n12118), .A2(n12117), .ZN(n12127) );
  INV_X1 U15208 ( .A(n12119), .ZN(n12123) );
  INV_X1 U15209 ( .A(n12120), .ZN(n12122) );
  OAI21_X1 U15210 ( .B1(n12123), .B2(n12122), .A(n12121), .ZN(n12161) );
  NAND2_X1 U15211 ( .A1(n12140), .A2(n12161), .ZN(n12124) );
  INV_X1 U15212 ( .A(n12124), .ZN(n12130) );
  INV_X1 U15213 ( .A(n12131), .ZN(n12125) );
  NOR2_X1 U15214 ( .A1(n12125), .A2(n12124), .ZN(n12129) );
  AOI22_X1 U15215 ( .A1(n12138), .A2(n12161), .B1(n12127), .B2(n12126), .ZN(
        n12128) );
  OAI222_X1 U15216 ( .A1(n12136), .A2(n10116), .B1(n12131), .B2(n12130), .C1(
        n12129), .C2(n12128), .ZN(n12143) );
  AOI21_X1 U15217 ( .B1(n12134), .B2(n12133), .A(n12132), .ZN(n12135) );
  INV_X1 U15218 ( .A(n12135), .ZN(n12162) );
  AOI21_X1 U15219 ( .B1(n10116), .B2(n12136), .A(n12162), .ZN(n12137) );
  AOI21_X1 U15220 ( .B1(n12138), .B2(n12163), .A(n12137), .ZN(n12139) );
  INV_X1 U15221 ( .A(n12139), .ZN(n12142) );
  INV_X1 U15222 ( .A(n12140), .ZN(n12141) );
  AOI222_X1 U15223 ( .A1(n12143), .A2(n12142), .B1(n12164), .B2(n12141), .C1(
        n12162), .C2(n12150), .ZN(n12144) );
  AOI21_X1 U15224 ( .B1(n12164), .B2(n12145), .A(n12144), .ZN(n12146) );
  AOI222_X1 U15225 ( .A1(n12147), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n12147), .B2(n12771), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n12771), .ZN(n12165) );
  NAND2_X1 U15226 ( .A1(n12165), .A2(n12148), .ZN(n12149) );
  NAND2_X1 U15227 ( .A1(n12153), .A2(n12149), .ZN(n12152) );
  INV_X1 U15228 ( .A(n12150), .ZN(n12151) );
  NAND2_X1 U15229 ( .A1(n12152), .A2(n12151), .ZN(n12155) );
  NAND2_X1 U15230 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20623) );
  AND2_X1 U15231 ( .A1(n11424), .A2(n20623), .ZN(n12158) );
  INV_X1 U15232 ( .A(n12936), .ZN(n12699) );
  NOR2_X1 U15233 ( .A1(n12159), .A2(n13309), .ZN(n12160) );
  NAND2_X1 U15234 ( .A1(n14710), .A2(n12160), .ZN(n12754) );
  NOR4_X1 U15235 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .ZN(
        n12166) );
  NOR2_X1 U15236 ( .A1(n12166), .A2(n12165), .ZN(n12887) );
  NOR2_X1 U15237 ( .A1(n11424), .A2(n20631), .ZN(n12167) );
  NAND2_X1 U15238 ( .A1(n19739), .A2(n12167), .ZN(n12762) );
  NAND4_X1 U15239 ( .A1(n13124), .A2(n12168), .A3(n14209), .A4(n19968), .ZN(
        n12826) );
  OR2_X1 U15240 ( .A1(n12826), .A2(n13309), .ZN(n12169) );
  OAI211_X1 U15241 ( .C1(n12699), .C2(n12754), .A(n12762), .B(n12169), .ZN(
        n12170) );
  NAND2_X1 U15242 ( .A1(n12170), .A2(n12937), .ZN(n12171) );
  AND2_X1 U15243 ( .A1(n14270), .A2(n14209), .ZN(n12173) );
  NAND2_X1 U15244 ( .A1(n13885), .A2(n12173), .ZN(n12190) );
  NOR4_X1 U15245 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12177) );
  NOR4_X1 U15246 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12176) );
  NOR4_X1 U15247 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12175) );
  NOR4_X1 U15248 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12174) );
  AND4_X1 U15249 ( .A1(n12177), .A2(n12176), .A3(n12175), .A4(n12174), .ZN(
        n12182) );
  NOR4_X1 U15250 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12180) );
  NOR4_X1 U15251 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12179) );
  NOR4_X1 U15252 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12178) );
  INV_X1 U15253 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20546) );
  AND4_X1 U15254 ( .A1(n12180), .A2(n12179), .A3(n12178), .A4(n20546), .ZN(
        n12181) );
  NAND2_X1 U15255 ( .A1(n12182), .A2(n12181), .ZN(n12183) );
  INV_X1 U15256 ( .A(n19925), .ZN(n19923) );
  NOR2_X1 U15257 ( .A1(n11426), .A2(n19923), .ZN(n12184) );
  INV_X1 U15258 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16086) );
  NOR2_X1 U15259 ( .A1(n14263), .A2(n16086), .ZN(n12188) );
  NOR3_X1 U15260 ( .A1(n14275), .A2(n19925), .A3(n11426), .ZN(n12185) );
  AOI22_X1 U15261 ( .A1(n14268), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14275), .ZN(n12186) );
  INV_X1 U15262 ( .A(n12186), .ZN(n12187) );
  NOR2_X1 U15263 ( .A1(n12188), .A2(n12187), .ZN(n12189) );
  NAND2_X1 U15264 ( .A1(n12190), .A2(n12189), .ZN(P1_U2873) );
  NAND2_X1 U15265 ( .A1(n19033), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12191) );
  NAND2_X1 U15266 ( .A1(n19368), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18996) );
  NAND2_X1 U15267 ( .A1(n18996), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12192) );
  NAND2_X1 U15268 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n13264), .ZN(
        n19170) );
  NAND2_X1 U15269 ( .A1(n19368), .A2(n19212), .ZN(n19281) );
  NAND2_X1 U15270 ( .A1(n12192), .A2(n19281), .ZN(n12193) );
  AND2_X1 U15271 ( .A1(n12193), .A2(n19688), .ZN(n19412) );
  AOI21_X1 U15272 ( .B1(n12215), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19412), .ZN(n12194) );
  INV_X1 U15273 ( .A(n12209), .ZN(n12200) );
  INV_X1 U15274 ( .A(n19368), .ZN(n12212) );
  NAND2_X1 U15275 ( .A1(n10562), .A2(n19720), .ZN(n19278) );
  AND2_X1 U15276 ( .A1(n19213), .A2(n19688), .ZN(n19208) );
  AOI21_X1 U15277 ( .B1(n12215), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19208), .ZN(n12198) );
  AOI22_X1 U15278 ( .A1(n12215), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19688), .B2(n19720), .ZN(n12201) );
  INV_X1 U15279 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12203) );
  XNOR2_X1 U15280 ( .A(n12204), .B(n12205), .ZN(n12546) );
  NAND2_X1 U15281 ( .A1(n12547), .A2(n12546), .ZN(n12548) );
  INV_X1 U15282 ( .A(n12205), .ZN(n12206) );
  OR2_X1 U15283 ( .A1(n12204), .A2(n12206), .ZN(n12207) );
  INV_X1 U15284 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12208) );
  NAND2_X1 U15285 ( .A1(n12210), .A2(n12200), .ZN(n12217) );
  INV_X1 U15286 ( .A(n19688), .ZN(n19692) );
  NAND2_X1 U15287 ( .A1(n12212), .A2(n12211), .ZN(n12213) );
  NAND2_X1 U15288 ( .A1(n18996), .A2(n12213), .ZN(n19138) );
  NOR2_X1 U15289 ( .A1(n19692), .A2(n19138), .ZN(n12214) );
  AOI21_X1 U15290 ( .B1(n12215), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12214), .ZN(n12216) );
  NAND2_X1 U15291 ( .A1(n12725), .A2(n12723), .ZN(n12218) );
  INV_X1 U15292 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12220) );
  AND4_X1 U15293 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__6__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U15294 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  NOR2_X1 U15295 ( .A1(n12413), .A2(n12224), .ZN(n12225) );
  AND2_X1 U15296 ( .A1(n13377), .A2(n13376), .ZN(n12227) );
  AOI22_X1 U15297 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n10428), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15298 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12332), .B1(
        n12333), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U15299 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12229) );
  AND2_X1 U15300 ( .A1(n12230), .A2(n12229), .ZN(n12233) );
  AOI22_X1 U15301 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15302 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10482), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12231) );
  NAND4_X1 U15303 ( .A1(n12234), .A2(n12233), .A3(n12232), .A4(n12231), .ZN(
        n12240) );
  AOI22_X1 U15304 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n10382), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15305 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10436), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15306 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12343), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12236) );
  NAND2_X1 U15307 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12235) );
  NAND4_X1 U15308 ( .A1(n12238), .A2(n12237), .A3(n12236), .A4(n12235), .ZN(
        n12239) );
  AOI22_X1 U15309 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10388), .B1(
        n10428), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15310 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12332), .B1(
        n12333), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12242) );
  NAND2_X1 U15311 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12241) );
  AND2_X1 U15312 ( .A1(n12242), .A2(n12241), .ZN(n12245) );
  AOI22_X1 U15313 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15314 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10482), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12243) );
  NAND4_X1 U15315 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(
        n12252) );
  AOI22_X1 U15316 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10382), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15317 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10436), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15318 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12342), .B1(
        n12343), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12248) );
  NAND2_X1 U15319 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12247) );
  NAND4_X1 U15320 ( .A1(n12250), .A2(n12249), .A3(n12248), .A4(n12247), .ZN(
        n12251) );
  NOR2_X1 U15321 ( .A1(n12252), .A2(n12251), .ZN(n13604) );
  INV_X1 U15322 ( .A(n13604), .ZN(n12253) );
  AOI22_X1 U15323 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10388), .B1(
        n10428), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15324 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12333), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12255) );
  NAND2_X1 U15325 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12254) );
  AND2_X1 U15326 ( .A1(n12255), .A2(n12254), .ZN(n12258) );
  AOI22_X1 U15327 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15328 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10431), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12256) );
  NAND4_X1 U15329 ( .A1(n12259), .A2(n12258), .A3(n12257), .A4(n12256), .ZN(
        n12265) );
  AOI22_X1 U15330 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15331 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15332 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12343), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12261) );
  NAND2_X1 U15333 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12260) );
  NAND4_X1 U15334 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12264) );
  NOR2_X1 U15335 ( .A1(n12265), .A2(n12264), .ZN(n13688) );
  AOI22_X1 U15336 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15337 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12267) );
  NAND2_X1 U15338 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12266) );
  AND2_X1 U15339 ( .A1(n12267), .A2(n12266), .ZN(n12270) );
  AOI22_X1 U15340 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15341 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12268) );
  NAND4_X1 U15342 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12277) );
  AOI22_X1 U15343 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15344 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15345 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12273) );
  NAND2_X1 U15346 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12272) );
  NAND4_X1 U15347 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        n12276) );
  OR2_X1 U15348 ( .A1(n12277), .A2(n12276), .ZN(n14779) );
  AOI22_X1 U15349 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15350 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12279) );
  NAND2_X1 U15351 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12278) );
  AND2_X1 U15352 ( .A1(n12279), .A2(n12278), .ZN(n12282) );
  AOI22_X1 U15353 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15354 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12280) );
  NAND4_X1 U15355 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12289) );
  AOI22_X1 U15356 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15357 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15358 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U15359 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12284) );
  NAND4_X1 U15360 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12288) );
  AOI22_X1 U15361 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15362 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12291) );
  NAND2_X1 U15363 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12290) );
  AND2_X1 U15364 ( .A1(n12291), .A2(n12290), .ZN(n12294) );
  AOI22_X1 U15365 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15366 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12292) );
  NAND4_X1 U15367 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n12301) );
  AOI22_X1 U15368 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15369 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15370 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12297) );
  NAND2_X1 U15371 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12296) );
  NAND4_X1 U15372 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12300) );
  NOR2_X1 U15373 ( .A1(n12301), .A2(n12300), .ZN(n14773) );
  INV_X1 U15374 ( .A(n14773), .ZN(n12302) );
  AOI22_X1 U15375 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15376 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12304) );
  NAND2_X1 U15377 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12303) );
  AND2_X1 U15378 ( .A1(n12304), .A2(n12303), .ZN(n12307) );
  AOI22_X1 U15379 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15380 ( .A1(n10482), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12305) );
  NAND4_X1 U15381 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(
        n12314) );
  AOI22_X1 U15382 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12340), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15383 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15384 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12310) );
  NAND2_X1 U15385 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12309) );
  NAND4_X1 U15386 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(
        n12313) );
  NOR2_X1 U15387 ( .A1(n12314), .A2(n12313), .ZN(n15866) );
  AOI22_X1 U15388 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12486), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12322) );
  AND2_X1 U15389 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12316) );
  OR2_X1 U15390 ( .A1(n12316), .A2(n12315), .ZN(n12491) );
  INV_X1 U15391 ( .A(n12491), .ZN(n12456) );
  NAND2_X1 U15392 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12318) );
  NAND2_X1 U15393 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12317) );
  AND3_X1 U15394 ( .A1(n12456), .A2(n12318), .A3(n12317), .ZN(n12321) );
  AOI22_X1 U15395 ( .A1(n12483), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15396 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12319) );
  NAND4_X1 U15397 ( .A1(n12322), .A2(n12321), .A3(n12320), .A4(n12319), .ZN(
        n12330) );
  AOI22_X1 U15398 ( .A1(n12483), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12486), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15399 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10208), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15400 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U15401 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12324) );
  NAND2_X1 U15402 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12323) );
  AND3_X1 U15403 ( .A1(n12324), .A2(n12491), .A3(n12323), .ZN(n12325) );
  NAND4_X1 U15404 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12329) );
  NAND2_X1 U15405 ( .A1(n19006), .A2(n12371), .ZN(n12350) );
  AOI22_X1 U15406 ( .A1(n12331), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15407 ( .A1(n12333), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12332), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12335) );
  NAND2_X1 U15408 ( .A1(n10428), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12334) );
  AND2_X1 U15409 ( .A1(n12335), .A2(n12334), .ZN(n12338) );
  AOI22_X1 U15410 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10431), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U15411 ( .A1(n10382), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13224), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12336) );
  NAND4_X1 U15412 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12349) );
  AOI22_X1 U15413 ( .A1(n12340), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15414 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12341), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15415 ( .A1(n12343), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12342), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12345) );
  NAND2_X1 U15416 ( .A1(n10436), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12344) );
  NAND4_X1 U15417 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12348) );
  XNOR2_X1 U15418 ( .A(n12350), .B(n12368), .ZN(n12374) );
  NAND2_X1 U15419 ( .A1(n9600), .A2(n12371), .ZN(n14843) );
  AOI22_X1 U15420 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12483), .B1(
        n9602), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15421 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10208), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15422 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12479), .B1(
        n12461), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12357) );
  NAND2_X1 U15423 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12355) );
  NAND2_X1 U15424 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12354) );
  AND3_X1 U15425 ( .A1(n12355), .A2(n12491), .A3(n12354), .ZN(n12356) );
  NAND4_X1 U15426 ( .A1(n12359), .A2(n12358), .A3(n12357), .A4(n12356), .ZN(
        n12367) );
  AOI22_X1 U15427 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12365) );
  NAND2_X1 U15428 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12361) );
  NAND2_X1 U15429 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12360) );
  AND3_X1 U15430 ( .A1(n12456), .A2(n12361), .A3(n12360), .ZN(n12364) );
  AOI22_X1 U15431 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10208), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15432 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12362) );
  NAND4_X1 U15433 ( .A1(n12365), .A2(n12364), .A3(n12363), .A4(n12362), .ZN(
        n12366) );
  NAND2_X1 U15434 ( .A1(n12367), .A2(n12366), .ZN(n12375) );
  NAND2_X1 U15435 ( .A1(n12368), .A2(n12371), .ZN(n12376) );
  XOR2_X1 U15436 ( .A(n12375), .B(n12376), .Z(n12369) );
  NAND2_X1 U15437 ( .A1(n12369), .A2(n12854), .ZN(n14764) );
  INV_X1 U15438 ( .A(n12375), .ZN(n12370) );
  NAND2_X1 U15439 ( .A1(n9600), .A2(n12370), .ZN(n14767) );
  INV_X1 U15440 ( .A(n12371), .ZN(n12372) );
  NOR2_X1 U15441 ( .A1(n14767), .A2(n12372), .ZN(n12373) );
  NOR2_X1 U15442 ( .A1(n12376), .A2(n12375), .ZN(n12391) );
  AOI22_X1 U15443 ( .A1(n12483), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12486), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12382) );
  NAND2_X1 U15444 ( .A1(n12489), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12378) );
  NAND2_X1 U15445 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12377) );
  AND3_X1 U15446 ( .A1(n12456), .A2(n12378), .A3(n12377), .ZN(n12381) );
  AOI22_X1 U15447 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10208), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15448 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12379) );
  NAND4_X1 U15449 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12390) );
  INV_X1 U15450 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20737) );
  AOI22_X1 U15451 ( .A1(n12483), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12486), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12388) );
  INV_X1 U15452 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n19058) );
  AOI22_X1 U15453 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15454 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12386) );
  NAND2_X1 U15455 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12384) );
  NAND2_X1 U15456 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12383) );
  AND3_X1 U15457 ( .A1(n12384), .A2(n12383), .A3(n12491), .ZN(n12385) );
  NAND4_X1 U15458 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n12385), .ZN(
        n12389) );
  AND2_X1 U15459 ( .A1(n12390), .A2(n12389), .ZN(n12392) );
  NAND2_X1 U15460 ( .A1(n12391), .A2(n12392), .ZN(n12414) );
  OAI211_X1 U15461 ( .C1(n12391), .C2(n12392), .A(n12854), .B(n12414), .ZN(
        n12395) );
  INV_X1 U15462 ( .A(n12392), .ZN(n12393) );
  NOR2_X1 U15463 ( .A1(n19006), .A2(n12393), .ZN(n14755) );
  INV_X1 U15464 ( .A(n12394), .ZN(n12397) );
  AOI22_X1 U15465 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15466 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10344), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15467 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U15468 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12400) );
  NAND2_X1 U15469 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12399) );
  AND3_X1 U15470 ( .A1(n12400), .A2(n12491), .A3(n12399), .ZN(n12401) );
  NAND4_X1 U15471 ( .A1(n12404), .A2(n12403), .A3(n12402), .A4(n12401), .ZN(
        n12412) );
  AOI22_X1 U15472 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12410) );
  NAND2_X1 U15473 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12406) );
  NAND2_X1 U15474 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12405) );
  AND3_X1 U15475 ( .A1(n12456), .A2(n12406), .A3(n12405), .ZN(n12409) );
  AOI22_X1 U15476 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10208), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15477 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12407) );
  NAND4_X1 U15478 ( .A1(n12410), .A2(n12409), .A3(n12408), .A4(n12407), .ZN(
        n12411) );
  NAND2_X1 U15479 ( .A1(n12412), .A2(n12411), .ZN(n12416) );
  AOI21_X1 U15480 ( .B1(n12414), .B2(n12416), .A(n12413), .ZN(n12415) );
  OR2_X1 U15481 ( .A1(n12414), .A2(n12416), .ZN(n12435) );
  INV_X1 U15482 ( .A(n12416), .ZN(n12417) );
  NAND2_X1 U15483 ( .A1(n9600), .A2(n12417), .ZN(n14750) );
  AOI22_X1 U15484 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15485 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10344), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15486 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12424) );
  NAND2_X1 U15487 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12422) );
  NAND2_X1 U15488 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12421) );
  AND3_X1 U15489 ( .A1(n12422), .A2(n12491), .A3(n12421), .ZN(n12423) );
  NAND4_X1 U15490 ( .A1(n12426), .A2(n12425), .A3(n12424), .A4(n12423), .ZN(
        n12434) );
  AOI22_X1 U15491 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12432) );
  NAND2_X1 U15492 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12428) );
  NAND2_X1 U15493 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12427) );
  AND3_X1 U15494 ( .A1(n12456), .A2(n12428), .A3(n12427), .ZN(n12431) );
  AOI22_X1 U15495 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U15496 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12429) );
  NAND4_X1 U15497 ( .A1(n12432), .A2(n12431), .A3(n12430), .A4(n12429), .ZN(
        n12433) );
  NAND2_X1 U15498 ( .A1(n12434), .A2(n12433), .ZN(n12439) );
  INV_X1 U15499 ( .A(n12439), .ZN(n12437) );
  INV_X1 U15500 ( .A(n12435), .ZN(n12436) );
  OR2_X1 U15501 ( .A1(n12435), .A2(n12439), .ZN(n12470) );
  OAI211_X1 U15502 ( .C1(n12437), .C2(n12436), .A(n12854), .B(n12470), .ZN(
        n12438) );
  NOR2_X1 U15503 ( .A1(n19006), .A2(n12439), .ZN(n14741) );
  NAND2_X1 U15504 ( .A1(n14742), .A2(n14741), .ZN(n14740) );
  AOI22_X1 U15505 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15506 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15507 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12443) );
  NAND2_X1 U15508 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12441) );
  NAND2_X1 U15509 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12440) );
  AND3_X1 U15510 ( .A1(n12441), .A2(n12491), .A3(n12440), .ZN(n12442) );
  NAND4_X1 U15511 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n12453) );
  AOI22_X1 U15512 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12451) );
  NAND2_X1 U15513 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12447) );
  NAND2_X1 U15514 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12446) );
  AND3_X1 U15515 ( .A1(n12456), .A2(n12447), .A3(n12446), .ZN(n12450) );
  AOI22_X1 U15516 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10344), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15517 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12448) );
  NAND4_X1 U15518 ( .A1(n12451), .A2(n12450), .A3(n12449), .A4(n12448), .ZN(
        n12452) );
  NAND2_X1 U15519 ( .A1(n12453), .A2(n12452), .ZN(n12471) );
  AOI22_X1 U15520 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12460) );
  NAND2_X1 U15521 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12455) );
  NAND2_X1 U15522 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12454) );
  AND3_X1 U15523 ( .A1(n12456), .A2(n12455), .A3(n12454), .ZN(n12459) );
  AOI22_X1 U15524 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15525 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U15526 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12469) );
  AOI22_X1 U15527 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U15528 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12466) );
  AOI22_X1 U15529 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12465) );
  NAND2_X1 U15530 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12463) );
  NAND2_X1 U15531 ( .A1(n12485), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12462) );
  AND3_X1 U15532 ( .A1(n12463), .A2(n12491), .A3(n12462), .ZN(n12464) );
  NAND4_X1 U15533 ( .A1(n12467), .A2(n12466), .A3(n12465), .A4(n12464), .ZN(
        n12468) );
  NAND2_X1 U15534 ( .A1(n12469), .A2(n12468), .ZN(n12474) );
  INV_X1 U15535 ( .A(n12470), .ZN(n14735) );
  INV_X1 U15536 ( .A(n12471), .ZN(n14736) );
  AND2_X1 U15537 ( .A1(n19006), .A2(n14736), .ZN(n12472) );
  NAND2_X1 U15538 ( .A1(n14735), .A2(n12472), .ZN(n12473) );
  NOR2_X1 U15539 ( .A1(n12473), .A2(n12474), .ZN(n12475) );
  AOI21_X1 U15540 ( .B1(n12474), .B2(n12473), .A(n12475), .ZN(n14729) );
  INV_X1 U15541 ( .A(n12475), .ZN(n12476) );
  AOI22_X1 U15542 ( .A1(n9602), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12486), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15543 ( .A1(n12483), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12490), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12477) );
  NAND2_X1 U15544 ( .A1(n12478), .A2(n12477), .ZN(n12498) );
  INV_X1 U15545 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12482) );
  AOI21_X1 U15546 ( .B1(n12485), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n12491), .ZN(n12481) );
  AOI22_X1 U15547 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12479), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12480) );
  OAI211_X1 U15548 ( .C1(n10336), .C2(n12482), .A(n12481), .B(n12480), .ZN(
        n12497) );
  AOI22_X1 U15549 ( .A1(n12484), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12483), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15550 ( .A1(n12486), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12485), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12487) );
  NAND2_X1 U15551 ( .A1(n12488), .A2(n12487), .ZN(n12496) );
  AOI22_X1 U15552 ( .A1(n12461), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12489), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12494) );
  NAND2_X1 U15553 ( .A1(n12490), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12493) );
  NAND2_X1 U15554 ( .A1(n10335), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12492) );
  NAND4_X1 U15555 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12495) );
  OAI22_X1 U15556 ( .A1(n12498), .A2(n12497), .B1(n12496), .B2(n12495), .ZN(
        n12499) );
  INV_X1 U15557 ( .A(n13236), .ZN(n12500) );
  NAND2_X1 U15558 ( .A1(n12500), .A2(n13237), .ZN(n12503) );
  NAND2_X1 U15559 ( .A1(n12501), .A2(n19617), .ZN(n12582) );
  OR2_X1 U15560 ( .A1(n12585), .A2(n12582), .ZN(n12502) );
  INV_X1 U15561 ( .A(n12504), .ZN(n12505) );
  NAND2_X1 U15562 ( .A1(n12505), .A2(n10118), .ZN(n12506) );
  NAND2_X1 U15563 ( .A1(n12535), .A2(n18884), .ZN(n12531) );
  OR2_X1 U15564 ( .A1(n18881), .A2(n12508), .ZN(n12731) );
  NOR2_X1 U15565 ( .A1(n12731), .A2(n12509), .ZN(n12520) );
  NOR4_X1 U15566 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12513) );
  NOR4_X1 U15567 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12512) );
  NOR4_X1 U15568 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12511) );
  NOR4_X1 U15569 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12510) );
  NAND4_X1 U15570 ( .A1(n12513), .A2(n12512), .A3(n12511), .A4(n12510), .ZN(
        n12518) );
  NOR4_X1 U15571 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12516) );
  NOR4_X1 U15572 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12515) );
  NOR4_X1 U15573 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n12514) );
  NAND4_X1 U15574 ( .A1(n12516), .A2(n12515), .A3(n12514), .A4(n19643), .ZN(
        n12517) );
  INV_X1 U15575 ( .A(n18858), .ZN(n14835) );
  INV_X1 U15576 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U15577 ( .A1(n12521), .A2(n19044), .ZN(n12522) );
  OR2_X1 U15578 ( .A1(n18881), .A2(n12522), .ZN(n14859) );
  NAND2_X1 U15579 ( .A1(n14847), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12525) );
  INV_X1 U15580 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12523) );
  OR2_X1 U15581 ( .A1(n14847), .A2(n12523), .ZN(n12524) );
  NAND2_X1 U15582 ( .A1(n12525), .A2(n12524), .ZN(n18954) );
  AOI22_X1 U15583 ( .A1(n18857), .A2(n18954), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n18881), .ZN(n12526) );
  OAI21_X1 U15584 ( .B1(n14835), .B2(n12527), .A(n12526), .ZN(n12528) );
  AOI21_X1 U15585 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n18859), .A(n12528), .ZN(
        n12529) );
  NAND2_X1 U15586 ( .A1(n12531), .A2(n10123), .ZN(P2_U2889) );
  INV_X1 U15587 ( .A(n13237), .ZN(n12532) );
  INV_X1 U15588 ( .A(n13199), .ZN(n13231) );
  NAND2_X1 U15589 ( .A1(n12532), .A2(n13231), .ZN(n12606) );
  INV_X1 U15590 ( .A(n12533), .ZN(n13201) );
  NAND2_X1 U15591 ( .A1(n12606), .A2(n13201), .ZN(n12534) );
  NAND2_X1 U15592 ( .A1(n18843), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12536) );
  NAND2_X1 U15593 ( .A1(n12539), .A2(n12538), .ZN(P2_U2857) );
  NOR2_X1 U15594 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .ZN(n12541) );
  NOR4_X1 U15595 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_BE_N_REG_3__SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12540) );
  NAND4_X1 U15596 ( .A1(n12541), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n12540), .ZN(n12544) );
  INV_X1 U15597 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20622) );
  NOR3_X1 U15598 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20622), .ZN(n12543) );
  NOR4_X1 U15599 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12542) );
  NAND4_X1 U15600 ( .A1(n19925), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12543), .A4(
        n12542), .ZN(U214) );
  NAND2_X1 U15601 ( .A1(n16085), .A2(U214), .ZN(U212) );
  NAND2_X1 U15602 ( .A1(n18819), .A2(n18676), .ZN(n18660) );
  OAI211_X1 U15603 ( .C1(n18837), .C2(n12545), .A(n9969), .B(n13520), .ZN(
        n15339) );
  OAI22_X1 U15604 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18660), .B1(
        n15339), .B2(n18811), .ZN(n12559) );
  OR2_X1 U15605 ( .A1(n12614), .A2(n12550), .ZN(n13583) );
  NOR2_X1 U15606 ( .A1(n18992), .A2(n13583), .ZN(n12558) );
  INV_X1 U15607 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19640) );
  OAI22_X1 U15608 ( .A1(n12684), .A2(n18833), .B1(n19640), .B2(n18825), .ZN(
        n12557) );
  INV_X1 U15609 ( .A(n12679), .ZN(n12551) );
  AOI22_X1 U15610 ( .A1(n18803), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n18775), .B2(
        n12551), .ZN(n12555) );
  XNOR2_X1 U15611 ( .A(n12553), .B(n12552), .ZN(n19711) );
  NAND2_X1 U15612 ( .A1(n19711), .A2(n18759), .ZN(n12554) );
  OAI211_X1 U15613 ( .C1(n9592), .C2(n18796), .A(n12555), .B(n12554), .ZN(
        n12556) );
  AOI211_X1 U15614 ( .C1(n14970), .C2(n12561), .A(n12560), .B(n18811), .ZN(
        n12569) );
  INV_X1 U15615 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14968) );
  OAI22_X1 U15616 ( .A1(n14968), .A2(n18833), .B1(n20723), .B2(n18825), .ZN(
        n12568) );
  INV_X1 U15617 ( .A(n18803), .ZN(n18828) );
  OAI22_X1 U15618 ( .A1(n18828), .A2(n10803), .B1(n12562), .B2(n18822), .ZN(
        n12567) );
  INV_X1 U15619 ( .A(n14983), .ZN(n12564) );
  OAI21_X1 U15620 ( .B1(n12564), .B2(n10050), .A(n14939), .ZN(n15161) );
  OAI21_X1 U15621 ( .B1(n15176), .B2(n12565), .A(n9675), .ZN(n15168) );
  OAI22_X1 U15622 ( .A1(n15161), .A2(n18796), .B1(n15168), .B2(n18823), .ZN(
        n12566) );
  OR4_X1 U15623 ( .A1(n12569), .A2(n12568), .A3(n12567), .A4(n12566), .ZN(
        P2_U2834) );
  AOI211_X1 U15624 ( .C1(n14926), .C2(n12571), .A(n18811), .B(n12570), .ZN(
        n12579) );
  OAI22_X1 U15625 ( .A1(n14928), .A2(n18833), .B1(n19665), .B2(n18825), .ZN(
        n12578) );
  OAI22_X1 U15626 ( .A1(n18828), .A2(n10860), .B1(n12572), .B2(n18822), .ZN(
        n12577) );
  AOI21_X1 U15627 ( .B1(n12573), .B2(n14941), .A(n14769), .ZN(n14930) );
  INV_X1 U15628 ( .A(n14930), .ZN(n15865) );
  INV_X1 U15629 ( .A(n9645), .ZN(n15146) );
  INV_X1 U15630 ( .A(n12574), .ZN(n12575) );
  OAI21_X1 U15631 ( .B1(n15146), .B2(n12575), .A(n14831), .ZN(n15140) );
  OAI22_X1 U15632 ( .A1(n15865), .A2(n18796), .B1(n15140), .B2(n18823), .ZN(
        n12576) );
  OR4_X1 U15633 ( .A1(n12579), .A2(n12578), .A3(n12577), .A4(n12576), .ZN(
        P2_U2832) );
  INV_X1 U15634 ( .A(n13583), .ZN(n18834) );
  INV_X1 U15635 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19737) );
  OAI211_X1 U15636 ( .C1(n18834), .C2(n19737), .A(n18595), .B(n12580), .ZN(
        P2_U2814) );
  NOR2_X1 U15637 ( .A1(n18598), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12581)
         );
  AOI22_X1 U15638 ( .A1(n12581), .A2(n18595), .B1(n12591), .B2(n18598), .ZN(
        P2_U3612) );
  INV_X1 U15639 ( .A(n12582), .ZN(n12583) );
  NOR3_X1 U15640 ( .A1(n12585), .A2(n12584), .A3(n12583), .ZN(n13242) );
  NOR2_X1 U15641 ( .A1(n13242), .A2(n16003), .ZN(n19723) );
  OAI21_X1 U15642 ( .B1(n12611), .B2(n19723), .A(n12586), .ZN(P2_U2819) );
  NOR2_X1 U15643 ( .A1(n12587), .A2(n13409), .ZN(n13274) );
  OAI22_X1 U15644 ( .A1(n19633), .A2(n18909), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n13274), .ZN(n12588) );
  NOR2_X1 U15645 ( .A1(n18598), .A2(n12588), .ZN(n12594) );
  INV_X1 U15646 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19629) );
  AOI21_X1 U15647 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19617), .A(n15994), 
        .ZN(n12589) );
  NOR2_X1 U15648 ( .A1(n12594), .A2(n12589), .ZN(n12593) );
  OAI21_X1 U15649 ( .B1(n13457), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19623), 
        .ZN(n12590) );
  NAND3_X1 U15650 ( .A1(n12591), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12590), 
        .ZN(n12592) );
  AOI22_X1 U15651 ( .A1(n12594), .A2(n19629), .B1(n12593), .B2(n12592), .ZN(
        P2_U3610) );
  INV_X1 U15652 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n12597) );
  INV_X1 U15653 ( .A(n18954), .ZN(n12596) );
  INV_X1 U15654 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12625) );
  OAI222_X1 U15655 ( .A1(n12597), .A2(n12650), .B1(n18961), .B2(n12596), .C1(
        n12666), .C2(n12625), .ZN(P2_U2966) );
  OR2_X1 U15656 ( .A1(n12614), .A2(n16003), .ZN(n12598) );
  OAI21_X1 U15657 ( .B1(n12599), .B2(n12598), .A(n12666), .ZN(n12600) );
  NAND2_X1 U15658 ( .A1(n18894), .A2(n12601), .ZN(n12639) );
  INV_X1 U15659 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14839) );
  INV_X1 U15660 ( .A(n18909), .ZN(n18924) );
  INV_X1 U15661 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16154) );
  INV_X1 U15662 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n20656) );
  OAI222_X1 U15663 ( .A1(n12639), .A2(n14839), .B1(n18911), .B2(n16154), .C1(
        n20656), .C2(n18909), .ZN(P2_U2928) );
  INV_X1 U15664 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n20726) );
  INV_X1 U15665 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n12602) );
  OAI222_X1 U15666 ( .A1(n12639), .A2(n13608), .B1(n18911), .B2(n20726), .C1(
        n12602), .C2(n18909), .ZN(P2_U2934) );
  NOR2_X1 U15667 ( .A1(n12614), .A2(n12603), .ZN(n12604) );
  NAND2_X1 U15668 ( .A1(n12605), .A2(n12604), .ZN(n12609) );
  NAND4_X1 U15669 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n13229) );
  NOR2_X1 U15670 ( .A1(n18596), .A2(n12610), .ZN(n15632) );
  INV_X1 U15671 ( .A(n15632), .ZN(n15993) );
  OAI22_X1 U15672 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19544), .B1(n12611), 
        .B2(n15993), .ZN(n12612) );
  AOI21_X1 U15673 ( .B1(n13229), .B2(n12613), .A(n12612), .ZN(n15356) );
  INV_X1 U15674 ( .A(n15356), .ZN(n12616) );
  NOR2_X1 U15675 ( .A1(n12614), .A2(n19006), .ZN(n13241) );
  NAND4_X1 U15676 ( .A1(n12616), .A2(n13241), .A3(n13240), .A4(n15342), .ZN(
        n12615) );
  OAI21_X1 U15677 ( .B1(n12220), .B2(n12616), .A(n12615), .ZN(P2_U3595) );
  INV_X1 U15678 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20636) );
  INV_X1 U15679 ( .A(n12976), .ZN(n19740) );
  AND2_X1 U15680 ( .A1(n20398), .A2(n15606), .ZN(n12644) );
  INV_X1 U15681 ( .A(n12644), .ZN(n12617) );
  OAI211_X1 U15682 ( .C1(n12642), .C2(n20636), .A(n19740), .B(n12617), .ZN(
        P1_U2801) );
  INV_X1 U15683 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15684 ( .A1(n18924), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12618) );
  OAI21_X1 U15685 ( .B1(n12660), .B2(n12639), .A(n12618), .ZN(P2_U2925) );
  INV_X1 U15686 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15687 ( .A1(n12636), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12619) );
  OAI21_X1 U15688 ( .B1(n12663), .B2(n12639), .A(n12619), .ZN(P2_U2924) );
  INV_X1 U15689 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15690 ( .A1(n12636), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12620) );
  OAI21_X1 U15691 ( .B1(n12621), .B2(n12639), .A(n12620), .ZN(P2_U2923) );
  INV_X1 U15692 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15693 ( .A1(n12636), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12622) );
  OAI21_X1 U15694 ( .B1(n12623), .B2(n12639), .A(n12622), .ZN(P2_U2922) );
  AOI22_X1 U15695 ( .A1(n18924), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12624) );
  OAI21_X1 U15696 ( .B1(n12625), .B2(n12639), .A(n12624), .ZN(P2_U2921) );
  INV_X1 U15697 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U15698 ( .A1(n12636), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12626) );
  OAI21_X1 U15699 ( .B1(n12627), .B2(n12639), .A(n12626), .ZN(P2_U2931) );
  INV_X1 U15700 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15701 ( .A1(n12636), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12628) );
  OAI21_X1 U15702 ( .B1(n12629), .B2(n12639), .A(n12628), .ZN(P2_U2930) );
  INV_X1 U15703 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15704 ( .A1(n12636), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12630) );
  OAI21_X1 U15705 ( .B1(n12631), .B2(n12639), .A(n12630), .ZN(P2_U2929) );
  INV_X1 U15706 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12657) );
  AOI22_X1 U15707 ( .A1(n12636), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12632) );
  OAI21_X1 U15708 ( .B1(n12657), .B2(n12639), .A(n12632), .ZN(P2_U2927) );
  INV_X1 U15709 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15710 ( .A1(n12636), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12633) );
  OAI21_X1 U15711 ( .B1(n12634), .B2(n12639), .A(n12633), .ZN(P2_U2935) );
  INV_X1 U15712 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13683) );
  AOI22_X1 U15713 ( .A1(n12636), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12635) );
  OAI21_X1 U15714 ( .B1(n13683), .B2(n12639), .A(n12635), .ZN(P2_U2933) );
  INV_X1 U15715 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14857) );
  AOI22_X1 U15716 ( .A1(n12636), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12637) );
  OAI21_X1 U15717 ( .B1(n14857), .B2(n12639), .A(n12637), .ZN(P2_U2932) );
  INV_X1 U15718 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U15719 ( .A1(n18924), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12638) );
  OAI21_X1 U15720 ( .B1(n12640), .B2(n12639), .A(n12638), .ZN(P2_U2926) );
  MUX2_X1 U15721 ( .A(n10726), .B(n9592), .S(n18851), .Z(n12641) );
  OAI21_X1 U15722 ( .B1(n18992), .B2(n18844), .A(n12641), .ZN(P2_U2886) );
  CLKBUF_X3 U15723 ( .A(n12643), .Z(n13951) );
  NOR2_X1 U15724 ( .A1(n11425), .A2(n13951), .ZN(n12646) );
  OAI21_X1 U15725 ( .B1(n12644), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20628), 
        .ZN(n12645) );
  OAI21_X1 U15726 ( .B1(n20628), .B2(n12646), .A(n12645), .ZN(P1_U3487) );
  INV_X1 U15727 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18901) );
  NAND2_X1 U15728 ( .A1(n18959), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12649) );
  INV_X1 U15729 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16113) );
  OR2_X1 U15730 ( .A1(n14847), .A2(n16113), .ZN(n12648) );
  NAND2_X1 U15731 ( .A1(n14847), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U15732 ( .A1(n12648), .A2(n12647), .ZN(n18871) );
  NAND2_X1 U15733 ( .A1(n18955), .A2(n18871), .ZN(n12661) );
  OAI211_X1 U15734 ( .C1(n18901), .C2(n12666), .A(n12649), .B(n12661), .ZN(
        P2_U2978) );
  INV_X1 U15735 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n18903) );
  INV_X2 U15736 ( .A(n12650), .ZN(n18959) );
  NAND2_X1 U15737 ( .A1(n18959), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12653) );
  INV_X1 U15738 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20765) );
  OR2_X1 U15739 ( .A1(n14847), .A2(n20765), .ZN(n12652) );
  NAND2_X1 U15740 ( .A1(n14847), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12651) );
  NAND2_X1 U15741 ( .A1(n12652), .A2(n12651), .ZN(n18874) );
  NAND2_X1 U15742 ( .A1(n18955), .A2(n18874), .ZN(n12658) );
  OAI211_X1 U15743 ( .C1(n18903), .C2(n12666), .A(n12653), .B(n12658), .ZN(
        P2_U2977) );
  NAND2_X1 U15744 ( .A1(n18959), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12656) );
  INV_X1 U15745 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16117) );
  OR2_X1 U15746 ( .A1(n14847), .A2(n16117), .ZN(n12655) );
  NAND2_X1 U15747 ( .A1(n14847), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U15748 ( .A1(n12655), .A2(n12654), .ZN(n18878) );
  NAND2_X1 U15749 ( .A1(n18955), .A2(n18878), .ZN(n12664) );
  OAI211_X1 U15750 ( .C1(n12657), .C2(n12666), .A(n12656), .B(n12664), .ZN(
        P2_U2960) );
  NAND2_X1 U15751 ( .A1(n18959), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12659) );
  OAI211_X1 U15752 ( .C1(n12660), .C2(n12666), .A(n12659), .B(n12658), .ZN(
        P2_U2962) );
  NAND2_X1 U15753 ( .A1(n18959), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12662) );
  OAI211_X1 U15754 ( .C1(n12666), .C2(n12663), .A(n12662), .B(n12661), .ZN(
        P2_U2963) );
  INV_X1 U15755 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n18907) );
  NAND2_X1 U15756 ( .A1(n18959), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12665) );
  OAI211_X1 U15757 ( .C1(n18907), .C2(n12666), .A(n12665), .B(n12664), .ZN(
        P2_U2975) );
  OAI21_X1 U15758 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n12668), .A(
        n12667), .ZN(n12716) );
  INV_X1 U15759 ( .A(n12716), .ZN(n12671) );
  INV_X1 U15760 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18826) );
  NOR2_X1 U15761 ( .A1(n18970), .A2(n18826), .ZN(n12719) );
  OR2_X1 U15762 ( .A1(n18820), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12669) );
  NAND2_X1 U15763 ( .A1(n12678), .A2(n12669), .ZN(n12717) );
  NOR2_X1 U15764 ( .A1(n15946), .A2(n12717), .ZN(n12670) );
  AOI211_X1 U15765 ( .C1(n12671), .C2(n15939), .A(n12719), .B(n12670), .ZN(
        n12674) );
  OAI21_X1 U15766 ( .B1(n15915), .B2(n12672), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12673) );
  OAI211_X1 U15767 ( .C1(n15063), .C2(n12202), .A(n12674), .B(n12673), .ZN(
        P2_U3014) );
  AOI21_X1 U15768 ( .B1(n15340), .B2(n12676), .A(n12675), .ZN(n12746) );
  INV_X1 U15769 ( .A(n12746), .ZN(n12682) );
  OAI21_X1 U15770 ( .B1(n12679), .B2(n12678), .A(n12677), .ZN(n12680) );
  XNOR2_X1 U15771 ( .A(n12680), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12740) );
  AOI22_X1 U15772 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n15915), .B1(
        n10903), .B2(n12740), .ZN(n12681) );
  OR2_X1 U15773 ( .A1(n15891), .A2(n19640), .ZN(n12738) );
  OAI211_X1 U15774 ( .C1(n15947), .C2(n12682), .A(n12681), .B(n12738), .ZN(
        n12683) );
  AOI21_X1 U15775 ( .B1(n15944), .B2(n12684), .A(n12683), .ZN(n12685) );
  OAI21_X1 U15776 ( .B1(n9592), .B2(n15063), .A(n12685), .ZN(P2_U3013) );
  NAND2_X1 U15777 ( .A1(n12687), .A2(n12686), .ZN(n18974) );
  AND3_X1 U15778 ( .A1(n10903), .A2(n18975), .A3(n18974), .ZN(n12694) );
  INV_X1 U15779 ( .A(n13522), .ZN(n12692) );
  AOI21_X1 U15780 ( .B1(n12690), .B2(n12689), .A(n12688), .ZN(n18976) );
  AOI22_X1 U15781 ( .A1(n15939), .A2(n18976), .B1(P2_REIP_REG_2__SCAN_IN), 
        .B2(n18791), .ZN(n12691) );
  OAI21_X1 U15782 ( .B1(n15922), .B2(n12692), .A(n12691), .ZN(n12693) );
  AOI211_X1 U15783 ( .C1(n15915), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n12694), .B(n12693), .ZN(n12695) );
  OAI21_X1 U15784 ( .B1(n12729), .B2(n15063), .A(n12695), .ZN(P2_U3012) );
  INV_X1 U15785 ( .A(n12696), .ZN(n12698) );
  INV_X1 U15786 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12697) );
  NAND2_X1 U15787 ( .A1(n12698), .A2(n12697), .ZN(n15627) );
  NAND2_X1 U15788 ( .A1(n13945), .A2(n15627), .ZN(n12753) );
  NOR2_X1 U15789 ( .A1(n12753), .A2(n11425), .ZN(n20625) );
  NAND2_X1 U15790 ( .A1(n12699), .A2(n13309), .ZN(n12701) );
  NAND2_X1 U15791 ( .A1(n19742), .A2(n12156), .ZN(n12700) );
  OAI211_X1 U15792 ( .C1(n20631), .C2(n20625), .A(n12701), .B(n12700), .ZN(
        n15593) );
  AND2_X1 U15793 ( .A1(n15593), .A2(n12937), .ZN(n19750) );
  INV_X1 U15794 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15594) );
  NAND2_X1 U15795 ( .A1(n14710), .A2(n12881), .ZN(n12704) );
  INV_X1 U15796 ( .A(n12904), .ZN(n12702) );
  NAND2_X1 U15797 ( .A1(n12704), .A2(n12702), .ZN(n12703) );
  NAND2_X1 U15798 ( .A1(n12703), .A2(n12779), .ZN(n12761) );
  NOR2_X1 U15799 ( .A1(n12761), .A2(n11432), .ZN(n12935) );
  INV_X1 U15800 ( .A(n12754), .ZN(n13104) );
  NOR2_X1 U15801 ( .A1(n12935), .A2(n13104), .ZN(n12900) );
  NOR2_X1 U15802 ( .A1(n12704), .A2(n13945), .ZN(n13105) );
  NAND2_X1 U15803 ( .A1(n12936), .A2(n13105), .ZN(n12705) );
  OAI21_X1 U15804 ( .B1(n12936), .B2(n12900), .A(n12705), .ZN(n12707) );
  INV_X1 U15805 ( .A(n12752), .ZN(n12760) );
  OAI22_X1 U15806 ( .A1(n12936), .A2(n12156), .B1(n12887), .B2(n12760), .ZN(
        n12706) );
  OR2_X1 U15807 ( .A1(n12707), .A2(n12706), .ZN(n15595) );
  NAND2_X1 U15808 ( .A1(n19750), .A2(n15595), .ZN(n12708) );
  OAI21_X1 U15809 ( .B1(n19750), .B2(n15594), .A(n12708), .ZN(P1_U3484) );
  AOI21_X1 U15810 ( .B1(n19006), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12709) );
  AND2_X1 U15811 ( .A1(n12710), .A2(n12709), .ZN(n12711) );
  MUX2_X1 U15812 ( .A(n12202), .B(n18827), .S(n18843), .Z(n12712) );
  OAI21_X1 U15813 ( .B1(n19715), .B2(n18844), .A(n12712), .ZN(P2_U2887) );
  INV_X1 U15814 ( .A(n15203), .ZN(n15221) );
  INV_X1 U15815 ( .A(n12713), .ZN(n12715) );
  XNOR2_X1 U15816 ( .A(n12715), .B(n12714), .ZN(n12772) );
  INV_X1 U15817 ( .A(n12772), .ZN(n18824) );
  OAI22_X1 U15818 ( .A1(n15978), .A2(n12716), .B1(n18986), .B2(n18824), .ZN(
        n12721) );
  NOR2_X1 U15819 ( .A1(n15330), .A2(n12202), .ZN(n12720) );
  OAI22_X1 U15820 ( .A1(n15336), .A2(n12743), .B1(n15309), .B2(n12717), .ZN(
        n12718) );
  NOR4_X1 U15821 ( .A1(n12721), .A2(n12720), .A3(n12719), .A4(n12718), .ZN(
        n12722) );
  OAI21_X1 U15822 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15221), .A(
        n12722), .ZN(P2_U3046) );
  INV_X1 U15823 ( .A(n12723), .ZN(n12724) );
  XNOR2_X1 U15824 ( .A(n12725), .B(n12724), .ZN(n12727) );
  MUX2_X1 U15825 ( .A(n12729), .B(n12728), .S(n18843), .Z(n12730) );
  OAI21_X1 U15826 ( .B1(n19139), .B2(n18844), .A(n12730), .ZN(P2_U2885) );
  INV_X1 U15827 ( .A(n12731), .ZN(n12732) );
  OAI22_X1 U15828 ( .A1(n14847), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14848), .ZN(n19034) );
  XNOR2_X1 U15829 ( .A(n12734), .B(n12733), .ZN(n18787) );
  INV_X1 U15830 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18913) );
  OAI222_X1 U15831 ( .A1(n13439), .A2(n19034), .B1(n18787), .B2(n18890), .C1(
        n18913), .C2(n14858), .ZN(P2_U2913) );
  AOI21_X1 U15832 ( .B1(n19715), .B2(n18884), .A(n18852), .ZN(n12737) );
  INV_X1 U15833 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16132) );
  INV_X1 U15834 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n17913) );
  AOI22_X1 U15835 ( .A1(n14848), .A2(n16132), .B1(n17913), .B2(n14847), .ZN(
        n18856) );
  AOI22_X1 U15836 ( .A1(n18883), .A2(n18856), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n18881), .ZN(n12736) );
  NAND3_X1 U15837 ( .A1(n19276), .A2(n18884), .A3(n18824), .ZN(n12735) );
  OAI211_X1 U15838 ( .C1(n12737), .C2(n18824), .A(n12736), .B(n12735), .ZN(
        P2_U2919) );
  INV_X1 U15839 ( .A(n19711), .ZN(n12739) );
  OAI21_X1 U15840 ( .B1(n18986), .B2(n12739), .A(n12738), .ZN(n12745) );
  OAI211_X1 U15841 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15203), .B(n18965), .ZN(n12742) );
  NAND2_X1 U15842 ( .A1(n11303), .A2(n12740), .ZN(n12741) );
  OAI211_X1 U15843 ( .C1(n12743), .C2(n15340), .A(n12742), .B(n12741), .ZN(
        n12744) );
  AOI211_X1 U15844 ( .C1(n18977), .C2(n12746), .A(n12745), .B(n12744), .ZN(
        n12747) );
  OAI21_X1 U15845 ( .B1(n9592), .B2(n15330), .A(n12747), .ZN(P2_U3045) );
  AOI22_X1 U15846 ( .A1(n14848), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14847), .ZN(n19047) );
  OR2_X1 U15847 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  NAND2_X1 U15848 ( .A1(n12750), .A2(n15980), .ZN(n18770) );
  INV_X1 U15849 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18910) );
  OAI222_X1 U15850 ( .A1(n13439), .A2(n19047), .B1(n18770), .B2(n18890), .C1(
        n18910), .C2(n14858), .ZN(P2_U2912) );
  NAND2_X1 U15851 ( .A1(n14710), .A2(n11424), .ZN(n12751) );
  NAND2_X1 U15852 ( .A1(n12891), .A2(n12904), .ZN(n12828) );
  OAI211_X1 U15853 ( .C1(n14712), .C2(n9939), .A(n12753), .B(n20623), .ZN(
        n12755) );
  NAND2_X1 U15854 ( .A1(n12755), .A2(n12754), .ZN(n12764) );
  INV_X1 U15855 ( .A(n12756), .ZN(n13661) );
  NAND2_X1 U15856 ( .A1(n12758), .A2(n12757), .ZN(n12759) );
  MUX2_X1 U15857 ( .A(n13661), .B(n12759), .S(n13073), .Z(n12782) );
  OAI21_X1 U15858 ( .B1(n12761), .B2(n12782), .A(n12760), .ZN(n12888) );
  OAI211_X1 U15859 ( .C1(n13293), .C2(n19949), .A(n12762), .B(n12888), .ZN(
        n12763) );
  AOI21_X1 U15860 ( .B1(n12936), .B2(n12764), .A(n12763), .ZN(n12765) );
  NAND2_X1 U15861 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15781), .ZN(n15782) );
  INV_X1 U15862 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19749) );
  OAI22_X1 U15863 ( .A1(n15585), .A2(n19741), .B1(n15782), .B2(n19749), .ZN(
        n12769) );
  NOR2_X1 U15864 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20357), .ZN(n19931) );
  INV_X1 U15865 ( .A(n20613), .ZN(n12793) );
  INV_X1 U15866 ( .A(n20611), .ZN(n14722) );
  INV_X1 U15867 ( .A(n12766), .ZN(n13130) );
  INV_X1 U15868 ( .A(n20087), .ZN(n20355) );
  OR2_X1 U15869 ( .A1(n12767), .A2(n20355), .ZN(n12768) );
  XNOR2_X1 U15870 ( .A(n12768), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19815) );
  NAND4_X1 U15871 ( .A1(n12769), .A2(n14722), .A3(n13130), .A4(n19815), .ZN(
        n12770) );
  OAI21_X1 U15872 ( .B1(n12793), .B2(n12771), .A(n12770), .ZN(P1_U3468) );
  AOI22_X1 U15873 ( .A1(n14848), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14847), .ZN(n19007) );
  NOR2_X1 U15874 ( .A1(n19709), .A2(n19711), .ZN(n12923) );
  AOI21_X1 U15875 ( .B1(n19711), .B2(n19709), .A(n12923), .ZN(n12774) );
  NAND2_X1 U15876 ( .A1(n19276), .A2(n12772), .ZN(n12773) );
  NAND2_X1 U15877 ( .A1(n12774), .A2(n12773), .ZN(n12925) );
  OAI21_X1 U15878 ( .B1(n12774), .B2(n12773), .A(n12925), .ZN(n12775) );
  NAND2_X1 U15879 ( .A1(n12775), .A2(n18884), .ZN(n12777) );
  AOI22_X1 U15880 ( .A1(n18852), .A2(n19711), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n18881), .ZN(n12776) );
  OAI211_X1 U15881 ( .C1(n19007), .C2(n13439), .A(n12777), .B(n12776), .ZN(
        P2_U2918) );
  INV_X1 U15882 ( .A(n11631), .ZN(n13463) );
  NAND2_X1 U15883 ( .A1(n12779), .A2(n12778), .ZN(n12781) );
  INV_X1 U15884 ( .A(n13293), .ZN(n12780) );
  AOI22_X1 U15885 ( .A1(n12781), .A2(n13289), .B1(n12780), .B2(n11432), .ZN(
        n12784) );
  INV_X1 U15886 ( .A(n12782), .ZN(n12783) );
  OAI211_X1 U15887 ( .C1(n12785), .C2(n13309), .A(n12784), .B(n12783), .ZN(
        n12907) );
  NAND4_X1 U15888 ( .A1(n12766), .A2(n12905), .A3(n12892), .A4(n12786), .ZN(
        n12787) );
  NOR2_X1 U15889 ( .A1(n12907), .A2(n12787), .ZN(n14709) );
  OAI22_X1 U15890 ( .A1(n13463), .A2(n14709), .B1(n12789), .B2(n11818), .ZN(
        n15581) );
  INV_X1 U15891 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14715) );
  AOI22_X1 U15892 ( .A1(n15581), .A2(n14722), .B1(P1_STATE2_REG_1__SCAN_IN), 
        .B2(n14715), .ZN(n12788) );
  OAI21_X1 U15893 ( .B1(n20609), .B2(n12789), .A(n12788), .ZN(n12791) );
  INV_X1 U15894 ( .A(n14712), .ZN(n12790) );
  NOR2_X1 U15895 ( .A1(n12790), .A2(n12794), .ZN(n15580) );
  AOI22_X1 U15896 ( .A1(n12793), .A2(n12791), .B1(n14722), .B2(n15580), .ZN(
        n12792) );
  OAI21_X1 U15897 ( .B1(n12794), .B2(n12793), .A(n12792), .ZN(P1_U3474) );
  NAND2_X1 U15898 ( .A1(n12976), .A2(n12979), .ZN(n12796) );
  NAND3_X1 U15899 ( .A1(n12936), .A2(n12937), .A3(n14712), .ZN(n12795) );
  NAND2_X1 U15900 ( .A1(n12796), .A2(n12795), .ZN(n12797) );
  INV_X1 U15901 ( .A(n15627), .ZN(n15603) );
  NAND2_X1 U15902 ( .A1(n15614), .A2(n15781), .ZN(n20630) );
  INV_X2 U15903 ( .A(n20630), .ZN(n19883) );
  NOR2_X4 U15904 ( .A1(n19860), .A2(n19883), .ZN(n19882) );
  AOI22_X1 U15905 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12798) );
  OAI21_X1 U15906 ( .B1(n14239), .B2(n19851), .A(n12798), .ZN(P1_U2915) );
  AOI22_X1 U15907 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12799) );
  OAI21_X1 U15908 ( .B1(n14248), .B2(n19851), .A(n12799), .ZN(P1_U2917) );
  INV_X1 U15909 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U15910 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12800) );
  OAI21_X1 U15911 ( .B1(n12801), .B2(n19851), .A(n12800), .ZN(P1_U2918) );
  INV_X1 U15912 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U15913 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12802) );
  OAI21_X1 U15914 ( .B1(n12803), .B2(n19851), .A(n12802), .ZN(P1_U2906) );
  INV_X1 U15915 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n20747) );
  AOI22_X1 U15916 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12804) );
  OAI21_X1 U15917 ( .B1(n20747), .B2(n19851), .A(n12804), .ZN(P1_U2907) );
  INV_X1 U15918 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14230) );
  AOI22_X1 U15919 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12805) );
  OAI21_X1 U15920 ( .B1(n14230), .B2(n19851), .A(n12805), .ZN(P1_U2913) );
  INV_X1 U15921 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U15922 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12806) );
  OAI21_X1 U15923 ( .B1(n12807), .B2(n19851), .A(n12806), .ZN(P1_U2914) );
  INV_X1 U15924 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U15925 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12808) );
  OAI21_X1 U15926 ( .B1(n12809), .B2(n19851), .A(n12808), .ZN(P1_U2908) );
  INV_X1 U15927 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U15928 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12810) );
  OAI21_X1 U15929 ( .B1(n12811), .B2(n19851), .A(n12810), .ZN(P1_U2909) );
  INV_X1 U15930 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U15931 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12812) );
  OAI21_X1 U15932 ( .B1(n12813), .B2(n19851), .A(n12812), .ZN(P1_U2919) );
  INV_X1 U15933 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U15934 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12814) );
  OAI21_X1 U15935 ( .B1(n12815), .B2(n19851), .A(n12814), .ZN(P1_U2911) );
  INV_X1 U15936 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12817) );
  AOI22_X1 U15937 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12816) );
  OAI21_X1 U15938 ( .B1(n12817), .B2(n19851), .A(n12816), .ZN(P1_U2912) );
  INV_X1 U15939 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U15940 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12818) );
  OAI21_X1 U15941 ( .B1(n12819), .B2(n19851), .A(n12818), .ZN(P1_U2920) );
  INV_X1 U15942 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U15943 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12820) );
  OAI21_X1 U15944 ( .B1(n12821), .B2(n19851), .A(n12820), .ZN(P1_U2916) );
  INV_X1 U15945 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12822) );
  OR2_X1 U15946 ( .A1(n14847), .A2(n12822), .ZN(n12824) );
  NAND2_X1 U15947 ( .A1(n14847), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12823) );
  AND2_X1 U15948 ( .A1(n12824), .A2(n12823), .ZN(n18949) );
  OAI21_X1 U15949 ( .B1(n15979), .B2(n12825), .A(n15304), .ZN(n18750) );
  INV_X1 U15950 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18905) );
  OAI222_X1 U15951 ( .A1(n13439), .A2(n18949), .B1(n18750), .B2(n18890), .C1(
        n18905), .C2(n14858), .ZN(P2_U2910) );
  NAND2_X1 U15952 ( .A1(n12828), .A2(n12827), .ZN(n12829) );
  OR2_X1 U15953 ( .A1(n12831), .A2(n12830), .ZN(n12832) );
  AND2_X1 U15954 ( .A1(n12864), .A2(n12832), .ZN(n19841) );
  INV_X1 U15955 ( .A(n19841), .ZN(n13413) );
  AND2_X2 U15956 ( .A1(n13951), .A2(n13949), .ZN(n13943) );
  INV_X1 U15957 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12834) );
  NAND2_X1 U15958 ( .A1(n13943), .A2(n12834), .ZN(n12838) );
  INV_X1 U15959 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12833) );
  NAND2_X1 U15960 ( .A1(n13938), .A2(n12833), .ZN(n12836) );
  NAND2_X1 U15961 ( .A1(n13949), .A2(n12834), .ZN(n12835) );
  NAND3_X1 U15962 ( .A1(n12836), .A2(n13977), .A3(n12835), .ZN(n12837) );
  NAND2_X1 U15963 ( .A1(n13938), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12839) );
  OAI21_X1 U15964 ( .B1(n13951), .B2(P1_EBX_REG_0__SCAN_IN), .A(n12839), .ZN(
        n13100) );
  XNOR2_X1 U15965 ( .A(n12866), .B(n13100), .ZN(n19831) );
  OR2_X1 U15966 ( .A1(n19831), .A2(n13949), .ZN(n12840) );
  NAND2_X1 U15967 ( .A1(n19831), .A2(n13949), .ZN(n12867) );
  AND2_X1 U15968 ( .A1(n12840), .A2(n12867), .ZN(n12913) );
  INV_X1 U15969 ( .A(n12913), .ZN(n12841) );
  AOI22_X1 U15970 ( .A1(n19845), .A2(n12841), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14197), .ZN(n12842) );
  OAI21_X1 U15971 ( .B1(n14196), .B2(n13413), .A(n12842), .ZN(P1_U2871) );
  NOR2_X1 U15972 ( .A1(n12845), .A2(n18843), .ZN(n12846) );
  AOI21_X1 U15973 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n18843), .A(n12846), .ZN(
        n12847) );
  OAI21_X1 U15974 ( .B1(n19277), .B2(n18844), .A(n12847), .ZN(P2_U2884) );
  XOR2_X1 U15975 ( .A(n12848), .B(n12948), .Z(n12853) );
  OR2_X1 U15976 ( .A1(n13009), .A2(n12849), .ZN(n12850) );
  AND2_X1 U15977 ( .A1(n12850), .A2(n12953), .ZN(n18747) );
  NOR2_X1 U15978 ( .A1(n18851), .A2(n9834), .ZN(n12851) );
  AOI21_X1 U15979 ( .B1(n18747), .B2(n18851), .A(n12851), .ZN(n12852) );
  OAI21_X1 U15980 ( .B1(n12853), .B2(n18844), .A(n12852), .ZN(P2_U2878) );
  AND2_X1 U15981 ( .A1(n12854), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13419) );
  NAND2_X1 U15982 ( .A1(n12855), .A2(n13419), .ZN(n13422) );
  XOR2_X1 U15983 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13422), .Z(n12861)
         );
  OAI21_X1 U15984 ( .B1(n12856), .B2(n12858), .A(n12857), .ZN(n18795) );
  NOR2_X1 U15985 ( .A1(n18795), .A2(n18843), .ZN(n12859) );
  AOI21_X1 U15986 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n18843), .A(n12859), .ZN(
        n12860) );
  OAI21_X1 U15987 ( .B1(n12861), .B2(n18844), .A(n12860), .ZN(P2_U2882) );
  NAND2_X1 U15988 ( .A1(n12863), .A2(n12864), .ZN(n12865) );
  INV_X1 U15989 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12875) );
  NAND2_X1 U15990 ( .A1(n13943), .A2(n12875), .ZN(n12871) );
  INV_X1 U15991 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13046) );
  NAND2_X1 U15992 ( .A1(n13938), .A2(n13046), .ZN(n12869) );
  NAND2_X1 U15993 ( .A1(n13949), .A2(n12875), .ZN(n12868) );
  NAND3_X1 U15994 ( .A1(n12869), .A2(n13977), .A3(n12868), .ZN(n12870) );
  AND2_X1 U15995 ( .A1(n12871), .A2(n12870), .ZN(n12872) );
  NAND2_X1 U15996 ( .A1(n12873), .A2(n12872), .ZN(n12874) );
  NAND2_X1 U15997 ( .A1(n13084), .A2(n12874), .ZN(n13312) );
  OAI22_X1 U15998 ( .A1(n14206), .A2(n13312), .B1(n12875), .B2(n19850), .ZN(
        n12876) );
  AOI21_X1 U15999 ( .B1(n13356), .B2(n19846), .A(n12876), .ZN(n12877) );
  INV_X1 U16000 ( .A(n12877), .ZN(P1_U2870) );
  NAND2_X1 U16001 ( .A1(n13280), .A2(n19954), .ZN(n13052) );
  OAI21_X1 U16002 ( .B1(n12756), .B2(n13048), .A(n13052), .ZN(n12878) );
  INV_X1 U16003 ( .A(n12878), .ZN(n12879) );
  NAND2_X1 U16004 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13041) );
  NAND2_X1 U16005 ( .A1(n12880), .A2(n13289), .ZN(n12885) );
  XNOR2_X1 U16006 ( .A(n13049), .B(n13048), .ZN(n12882) );
  OAI211_X1 U16007 ( .C1(n12882), .C2(n12756), .A(n12881), .B(n11421), .ZN(
        n12883) );
  INV_X1 U16008 ( .A(n12883), .ZN(n12884) );
  XNOR2_X1 U16009 ( .A(n13041), .B(n13042), .ZN(n13040) );
  XNOR2_X1 U16010 ( .A(n13040), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13418) );
  NAND2_X1 U16011 ( .A1(n11424), .A2(n15627), .ZN(n12886) );
  NAND4_X1 U16012 ( .A1(n12887), .A2(n19949), .A3(n20623), .A4(n12886), .ZN(
        n12889) );
  NAND2_X1 U16013 ( .A1(n12889), .A2(n12888), .ZN(n12890) );
  OAI21_X1 U16014 ( .B1(n12891), .B2(n12890), .A(n12937), .ZN(n12897) );
  OAI21_X1 U16015 ( .B1(n12892), .B2(n20631), .A(n19932), .ZN(n12893) );
  OAI21_X1 U16016 ( .B1(n15603), .B2(n12756), .A(n12893), .ZN(n12894) );
  NAND2_X1 U16017 ( .A1(n12894), .A2(n11426), .ZN(n12895) );
  NAND4_X1 U16018 ( .A1(n12936), .A2(n9937), .A3(n12937), .A4(n12895), .ZN(
        n12896) );
  INV_X1 U16019 ( .A(n12898), .ZN(n12899) );
  OAI211_X1 U16020 ( .C1(n12901), .C2(n12911), .A(n12900), .B(n12899), .ZN(
        n12902) );
  OAI21_X1 U16021 ( .B1(n12905), .B2(n12904), .A(n12903), .ZN(n12906) );
  OR2_X1 U16022 ( .A1(n12907), .A2(n12906), .ZN(n12908) );
  NAND2_X1 U16023 ( .A1(n12915), .A2(n12908), .ZN(n19914) );
  OR2_X1 U16024 ( .A1(n19914), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12910) );
  OR2_X1 U16025 ( .A1(n12915), .A2(n19819), .ZN(n12909) );
  OAI21_X1 U16026 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19915), .A(
        n14520), .ZN(n19917) );
  OR2_X1 U16027 ( .A1(n12156), .A2(n13289), .ZN(n15605) );
  OAI21_X1 U16028 ( .B1(n12911), .B2(n11437), .A(n15605), .ZN(n12912) );
  INV_X2 U16029 ( .A(n19819), .ZN(n19921) );
  INV_X1 U16030 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20547) );
  OAI22_X1 U16031 ( .A1(n12913), .A2(n15775), .B1(n19921), .B2(n20547), .ZN(
        n12914) );
  AOI21_X1 U16032 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n19917), .A(
        n12914), .ZN(n12918) );
  NAND2_X1 U16033 ( .A1(n12915), .A2(n14712), .ZN(n14679) );
  INV_X1 U16034 ( .A(n14660), .ZN(n14536) );
  INV_X1 U16035 ( .A(n13061), .ZN(n12916) );
  NAND3_X1 U16036 ( .A1(n14536), .A2(n12833), .A3(n12916), .ZN(n12917) );
  OAI211_X1 U16037 ( .C1(n13418), .C2(n14704), .A(n12918), .B(n12917), .ZN(
        P1_U3030) );
  NAND2_X1 U16038 ( .A1(n12920), .A2(n12919), .ZN(n12922) );
  AND2_X1 U16039 ( .A1(n12922), .A2(n10062), .ZN(n18987) );
  INV_X1 U16040 ( .A(n19139), .ZN(n19701) );
  INV_X1 U16041 ( .A(n18987), .ZN(n19699) );
  NOR2_X1 U16042 ( .A1(n19701), .A2(n19699), .ZN(n13182) );
  AOI21_X1 U16043 ( .B1(n19701), .B2(n19699), .A(n13182), .ZN(n12927) );
  INV_X1 U16044 ( .A(n12923), .ZN(n12924) );
  NAND2_X1 U16045 ( .A1(n12925), .A2(n12924), .ZN(n12926) );
  NAND2_X1 U16046 ( .A1(n12927), .A2(n12926), .ZN(n13184) );
  OAI21_X1 U16047 ( .B1(n12927), .B2(n12926), .A(n13184), .ZN(n12928) );
  NAND2_X1 U16048 ( .A1(n12928), .A2(n18884), .ZN(n12931) );
  AOI22_X1 U16049 ( .A1(n14848), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14847), .ZN(n19011) );
  INV_X1 U16050 ( .A(n19011), .ZN(n12929) );
  AOI22_X1 U16051 ( .A1(n18883), .A2(n12929), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n18881), .ZN(n12930) );
  OAI211_X1 U16052 ( .C1(n18987), .C2(n18862), .A(n12931), .B(n12930), .ZN(
        P2_U2917) );
  XNOR2_X1 U16053 ( .A(n12933), .B(n12932), .ZN(n13470) );
  INV_X1 U16054 ( .A(n13470), .ZN(n13101) );
  NAND3_X1 U16055 ( .A1(n15614), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15776) );
  INV_X1 U16056 ( .A(n15776), .ZN(n12934) );
  INV_X1 U16057 ( .A(n20398), .ZN(n20469) );
  AND2_X1 U16058 ( .A1(n12938), .A2(n20469), .ZN(n20629) );
  INV_X1 U16059 ( .A(n20629), .ZN(n12939) );
  NAND2_X1 U16060 ( .A1(n12939), .A2(n15614), .ZN(n12940) );
  NAND2_X1 U16061 ( .A1(n15614), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12942) );
  NAND2_X1 U16062 ( .A1(n20429), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12941) );
  AND2_X1 U16063 ( .A1(n12942), .A2(n12941), .ZN(n13351) );
  NAND2_X1 U16064 ( .A1(n14459), .A2(n13351), .ZN(n12946) );
  OAI21_X1 U16065 ( .B1(n12943), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13041), .ZN(n19908) );
  INV_X1 U16066 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n12944) );
  OAI22_X1 U16067 ( .A1(n19748), .A2(n19908), .B1(n19921), .B2(n12944), .ZN(
        n12945) );
  AOI21_X1 U16068 ( .B1(n12946), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n12945), .ZN(n12947) );
  OAI21_X1 U16069 ( .B1(n13101), .B2(n19924), .A(n12947), .ZN(P1_U2999) );
  INV_X1 U16070 ( .A(n12948), .ZN(n12949) );
  NOR2_X1 U16071 ( .A1(n12848), .A2(n12949), .ZN(n12952) );
  OAI211_X1 U16072 ( .C1(n12952), .C2(n12951), .A(n18848), .B(n12950), .ZN(
        n12958) );
  NAND2_X1 U16073 ( .A1(n12954), .A2(n12953), .ZN(n12956) );
  INV_X1 U16074 ( .A(n13066), .ZN(n12955) );
  AND2_X1 U16075 ( .A1(n12956), .A2(n12955), .ZN(n18736) );
  NAND2_X1 U16076 ( .A1(n18736), .A2(n18851), .ZN(n12957) );
  OAI211_X1 U16077 ( .C1(n18851), .C2(n12959), .A(n12958), .B(n12957), .ZN(
        P2_U2877) );
  INV_X1 U16078 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12960) );
  NOR3_X1 U16079 ( .A1(n13422), .A2(n12967), .A3(n12960), .ZN(n12968) );
  XNOR2_X1 U16080 ( .A(n12968), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12966) );
  NAND2_X1 U16081 ( .A1(n12961), .A2(n12962), .ZN(n12963) );
  NAND2_X1 U16082 ( .A1(n13008), .A2(n12963), .ZN(n18769) );
  INV_X1 U16083 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12964) );
  MUX2_X1 U16084 ( .A(n18769), .B(n12964), .S(n18843), .Z(n12965) );
  OAI21_X1 U16085 ( .B1(n12966), .B2(n18844), .A(n12965), .ZN(P2_U2880) );
  NOR2_X1 U16086 ( .A1(n13422), .A2(n12967), .ZN(n12969) );
  INV_X1 U16087 ( .A(n12968), .ZN(n13013) );
  OAI211_X1 U16088 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n12969), .A(
        n13013), .B(n18848), .ZN(n12973) );
  NAND2_X1 U16089 ( .A1(n12857), .A2(n12970), .ZN(n12971) );
  AND2_X1 U16090 ( .A1(n12961), .A2(n12971), .ZN(n18783) );
  NAND2_X1 U16091 ( .A1(n18783), .A2(n18851), .ZN(n12972) );
  OAI211_X1 U16092 ( .C1(n18851), .C2(n12974), .A(n12973), .B(n12972), .ZN(
        P2_U2881) );
  NAND2_X1 U16093 ( .A1(n12756), .A2(n20631), .ZN(n12975) );
  NOR2_X2 U16094 ( .A1(n19904), .A2(n12979), .ZN(n19892) );
  INV_X1 U16095 ( .A(DATAI_4_), .ZN(n12978) );
  NAND2_X1 U16096 ( .A1(n19925), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U16097 ( .B1(n19925), .B2(n12978), .A(n12977), .ZN(n14245) );
  NAND2_X1 U16098 ( .A1(n19892), .A2(n14245), .ZN(n13021) );
  AND2_X2 U16099 ( .A1(n13006), .A2(n12979), .ZN(n19905) );
  AOI22_X1 U16100 ( .A1(n19905), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U16101 ( .A1(n13021), .A2(n12980), .ZN(P1_U2941) );
  MUX2_X1 U16102 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n19925), .Z(
        n14217) );
  NAND2_X1 U16103 ( .A1(n19892), .A2(n14217), .ZN(n13037) );
  AOI22_X1 U16104 ( .A1(n19905), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n12981) );
  NAND2_X1 U16105 ( .A1(n13037), .A2(n12981), .ZN(P1_U2963) );
  INV_X1 U16106 ( .A(DATAI_1_), .ZN(n12983) );
  NAND2_X1 U16107 ( .A1(n19925), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12982) );
  OAI21_X1 U16108 ( .B1(n19925), .B2(n12983), .A(n12982), .ZN(n14258) );
  NAND2_X1 U16109 ( .A1(n19892), .A2(n14258), .ZN(n13039) );
  AOI22_X1 U16110 ( .A1(n19905), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n12984) );
  NAND2_X1 U16111 ( .A1(n13039), .A2(n12984), .ZN(P1_U2938) );
  NAND2_X1 U16112 ( .A1(n19923), .A2(DATAI_2_), .ZN(n12986) );
  NAND2_X1 U16113 ( .A1(n19925), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12985) );
  AND2_X1 U16114 ( .A1(n12986), .A2(n12985), .ZN(n19951) );
  INV_X1 U16115 ( .A(n19951), .ZN(n14254) );
  NAND2_X1 U16116 ( .A1(n19892), .A2(n14254), .ZN(n13035) );
  AOI22_X1 U16117 ( .A1(n19905), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n12987) );
  NAND2_X1 U16118 ( .A1(n13035), .A2(n12987), .ZN(P1_U2939) );
  INV_X1 U16119 ( .A(DATAI_5_), .ZN(n12989) );
  NAND2_X1 U16120 ( .A1(n19925), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12988) );
  OAI21_X1 U16121 ( .B1(n19925), .B2(n12989), .A(n12988), .ZN(n14241) );
  NAND2_X1 U16122 ( .A1(n19892), .A2(n14241), .ZN(n13019) );
  AOI22_X1 U16123 ( .A1(n19905), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n12990) );
  NAND2_X1 U16124 ( .A1(n13019), .A2(n12990), .ZN(P1_U2942) );
  INV_X1 U16125 ( .A(DATAI_6_), .ZN(n12992) );
  NAND2_X1 U16126 ( .A1(n19925), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12991) );
  OAI21_X1 U16127 ( .B1(n19925), .B2(n12992), .A(n12991), .ZN(n14236) );
  NAND2_X1 U16128 ( .A1(n19892), .A2(n14236), .ZN(n13031) );
  AOI22_X1 U16129 ( .A1(n19905), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n12993) );
  NAND2_X1 U16130 ( .A1(n13031), .A2(n12993), .ZN(P1_U2943) );
  NAND2_X1 U16131 ( .A1(n19923), .A2(DATAI_0_), .ZN(n12995) );
  NAND2_X1 U16132 ( .A1(n19925), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12994) );
  AND2_X1 U16133 ( .A1(n12995), .A2(n12994), .ZN(n19938) );
  INV_X1 U16134 ( .A(n19938), .ZN(n12996) );
  NAND2_X1 U16135 ( .A1(n19892), .A2(n12996), .ZN(n13033) );
  AOI22_X1 U16136 ( .A1(n19905), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n12997) );
  NAND2_X1 U16137 ( .A1(n13033), .A2(n12997), .ZN(P1_U2937) );
  INV_X1 U16138 ( .A(DATAI_3_), .ZN(n12999) );
  NAND2_X1 U16139 ( .A1(n19925), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12998) );
  OAI21_X1 U16140 ( .B1(n19925), .B2(n12999), .A(n12998), .ZN(n14250) );
  NAND2_X1 U16141 ( .A1(n19892), .A2(n14250), .ZN(n13027) );
  AOI22_X1 U16142 ( .A1(n19905), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U16143 ( .A1(n13027), .A2(n13000), .ZN(P1_U2940) );
  INV_X1 U16144 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19854) );
  INV_X1 U16145 ( .A(n19892), .ZN(n13003) );
  INV_X1 U16146 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13001) );
  NOR2_X1 U16147 ( .A1(n19923), .A2(n13001), .ZN(n13002) );
  AOI21_X1 U16148 ( .B1(DATAI_15_), .B2(n19923), .A(n13002), .ZN(n14271) );
  INV_X1 U16149 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19855) );
  OAI222_X1 U16150 ( .A1(n13017), .A2(n19854), .B1(n13003), .B2(n14271), .C1(
        n13006), .C2(n19855), .ZN(P1_U2967) );
  MUX2_X1 U16151 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n19925), .Z(
        n14276) );
  NAND2_X1 U16152 ( .A1(n19892), .A2(n14276), .ZN(n19902) );
  NAND2_X1 U16153 ( .A1(n19904), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13004) );
  OAI211_X1 U16154 ( .C1(n20747), .C2(n13017), .A(n19902), .B(n13004), .ZN(
        P1_U2950) );
  INV_X1 U16155 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n20677) );
  MUX2_X1 U16156 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n19925), .Z(
        n14221) );
  NAND2_X1 U16157 ( .A1(n19892), .A2(n14221), .ZN(n19898) );
  NAND2_X1 U16158 ( .A1(n19905), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13005) );
  OAI211_X1 U16159 ( .C1(n13006), .C2(n20677), .A(n19898), .B(n13005), .ZN(
        P1_U2947) );
  AND2_X1 U16160 ( .A1(n13008), .A2(n13007), .ZN(n13010) );
  OR2_X1 U16161 ( .A1(n13010), .A2(n13009), .ZN(n15929) );
  INV_X1 U16162 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13012) );
  OAI21_X1 U16163 ( .B1(n13013), .B2(n13012), .A(n13011), .ZN(n13014) );
  NAND3_X1 U16164 ( .A1(n13014), .A2(n18848), .A3(n12848), .ZN(n13016) );
  NAND2_X1 U16165 ( .A1(n18843), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13015) );
  OAI211_X1 U16166 ( .C1(n15929), .C2(n18843), .A(n13016), .B(n13015), .ZN(
        P2_U2879) );
  AOI22_X1 U16167 ( .A1(n19905), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13018) );
  NAND2_X1 U16168 ( .A1(n13019), .A2(n13018), .ZN(P1_U2957) );
  AOI22_X1 U16169 ( .A1(n19905), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13020) );
  NAND2_X1 U16170 ( .A1(n13021), .A2(n13020), .ZN(P1_U2956) );
  MUX2_X1 U16171 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n19925), .Z(
        n14224) );
  NAND2_X1 U16172 ( .A1(n19892), .A2(n14224), .ZN(n19896) );
  AOI22_X1 U16173 ( .A1(n19905), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U16174 ( .A1(n19896), .A2(n13022), .ZN(P1_U2946) );
  INV_X1 U16175 ( .A(DATAI_7_), .ZN(n13024) );
  NAND2_X1 U16176 ( .A1(n19925), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13023) );
  OAI21_X1 U16177 ( .B1(n19925), .B2(n13024), .A(n13023), .ZN(n19977) );
  NAND2_X1 U16178 ( .A1(n19892), .A2(n19977), .ZN(n13029) );
  AOI22_X1 U16179 ( .A1(n19905), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13025) );
  NAND2_X1 U16180 ( .A1(n13029), .A2(n13025), .ZN(P1_U2959) );
  AOI22_X1 U16181 ( .A1(n19905), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13026) );
  NAND2_X1 U16182 ( .A1(n13027), .A2(n13026), .ZN(P1_U2955) );
  AOI22_X1 U16183 ( .A1(n19905), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13028) );
  NAND2_X1 U16184 ( .A1(n13029), .A2(n13028), .ZN(P1_U2944) );
  AOI22_X1 U16185 ( .A1(n19905), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U16186 ( .A1(n13031), .A2(n13030), .ZN(P1_U2958) );
  AOI22_X1 U16187 ( .A1(n19905), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13032) );
  NAND2_X1 U16188 ( .A1(n13033), .A2(n13032), .ZN(P1_U2952) );
  AOI22_X1 U16189 ( .A1(n19905), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13034) );
  NAND2_X1 U16190 ( .A1(n13035), .A2(n13034), .ZN(P1_U2954) );
  AOI22_X1 U16191 ( .A1(n19905), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13036) );
  NAND2_X1 U16192 ( .A1(n13037), .A2(n13036), .ZN(P1_U2948) );
  AOI22_X1 U16193 ( .A1(n19905), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U16194 ( .A1(n13039), .A2(n13038), .ZN(P1_U2953) );
  NAND2_X1 U16195 ( .A1(n13040), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13045) );
  INV_X1 U16196 ( .A(n13041), .ZN(n13043) );
  NAND2_X1 U16197 ( .A1(n13043), .A2(n13042), .ZN(n13044) );
  INV_X1 U16198 ( .A(n13655), .ZN(n13645) );
  NAND2_X1 U16199 ( .A1(n13049), .A2(n13048), .ZN(n13050) );
  NAND2_X1 U16200 ( .A1(n13050), .A2(n13051), .ZN(n13088) );
  OAI21_X1 U16201 ( .B1(n13051), .B2(n13050), .A(n13088), .ZN(n13054) );
  INV_X1 U16202 ( .A(n13052), .ZN(n13053) );
  AOI21_X1 U16203 ( .B1(n13054), .B2(n13661), .A(n13053), .ZN(n13055) );
  NAND2_X1 U16204 ( .A1(n13056), .A2(n13055), .ZN(n13091) );
  XNOR2_X1 U16205 ( .A(n13092), .B(n13091), .ZN(n13358) );
  INV_X1 U16206 ( .A(n15740), .ZN(n14658) );
  NAND2_X1 U16207 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14505) );
  AOI21_X1 U16208 ( .B1(n14658), .B2(n14505), .A(n15735), .ZN(n14699) );
  INV_X1 U16209 ( .A(n14699), .ZN(n13060) );
  INV_X1 U16210 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20548) );
  NOR2_X1 U16211 ( .A1(n19921), .A2(n20548), .ZN(n13352) );
  NOR2_X1 U16212 ( .A1(n14715), .A2(n12833), .ZN(n13057) );
  OAI21_X1 U16213 ( .B1(n14715), .B2(n12833), .A(n13046), .ZN(n13336) );
  INV_X1 U16214 ( .A(n13336), .ZN(n13095) );
  AOI21_X1 U16215 ( .B1(n13057), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13095), .ZN(n13058) );
  OAI22_X1 U16216 ( .A1(n13058), .A2(n19915), .B1(n15775), .B2(n13312), .ZN(
        n13059) );
  AOI211_X1 U16217 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13060), .A(
        n13352), .B(n13059), .ZN(n13064) );
  INV_X1 U16218 ( .A(n15730), .ZN(n13062) );
  NAND3_X1 U16219 ( .A1(n13062), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13046), .ZN(n13063) );
  OAI211_X1 U16220 ( .C1(n13358), .C2(n14704), .A(n13064), .B(n13063), .ZN(
        P1_U3029) );
  INV_X1 U16221 ( .A(n13065), .ZN(n13144) );
  XNOR2_X1 U16222 ( .A(n12950), .B(n13144), .ZN(n13072) );
  OR2_X1 U16223 ( .A1(n13067), .A2(n13066), .ZN(n13069) );
  NAND2_X1 U16224 ( .A1(n13069), .A2(n13068), .ZN(n18724) );
  MUX2_X1 U16225 ( .A(n18724), .B(n13070), .S(n18843), .Z(n13071) );
  OAI21_X1 U16226 ( .B1(n13072), .B2(n18844), .A(n13071), .ZN(P2_U2876) );
  NAND2_X1 U16227 ( .A1(n13073), .A2(n9938), .ZN(n13074) );
  INV_X1 U16228 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19886) );
  OAI222_X1 U16229 ( .A1(n14279), .A2(n13101), .B1(n14272), .B2(n19938), .C1(
        n14270), .C2(n19886), .ZN(P1_U2904) );
  INV_X1 U16230 ( .A(n13075), .ZN(n13076) );
  NOR2_X1 U16231 ( .A1(n13077), .A2(n13076), .ZN(n13079) );
  AOI21_X1 U16232 ( .B1(n13079), .B2(n12862), .A(n9794), .ZN(n13372) );
  INV_X1 U16233 ( .A(n13372), .ZN(n13087) );
  INV_X1 U16234 ( .A(n14250), .ZN(n19956) );
  INV_X1 U16235 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19877) );
  OAI222_X1 U16236 ( .A1(n13087), .A2(n14279), .B1(n14272), .B2(n19956), .C1(
        n14270), .C2(n19877), .ZN(P1_U2901) );
  INV_X1 U16237 ( .A(n13356), .ZN(n13080) );
  INV_X1 U16238 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19879) );
  OAI222_X1 U16239 ( .A1(n13080), .A2(n14279), .B1(n14272), .B2(n19951), .C1(
        n14270), .C2(n19879), .ZN(P1_U2902) );
  INV_X1 U16240 ( .A(n14258), .ZN(n19946) );
  INV_X1 U16241 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19881) );
  OAI222_X1 U16242 ( .A1(n13413), .A2(n14279), .B1(n14272), .B2(n19946), .C1(
        n14270), .C2(n19881), .ZN(P1_U2903) );
  INV_X1 U16243 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13086) );
  MUX2_X1 U16244 ( .A(n13927), .B(n13977), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13082) );
  OAI21_X1 U16245 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13081), .A(
        n13082), .ZN(n13083) );
  AND2_X1 U16246 ( .A1(n13084), .A2(n13083), .ZN(n13085) );
  NOR2_X1 U16247 ( .A1(n13169), .A2(n13085), .ZN(n13096) );
  INV_X1 U16248 ( .A(n13096), .ZN(n13295) );
  OAI222_X1 U16249 ( .A1(n13087), .A2(n14208), .B1(n13086), .B2(n19850), .C1(
        n13295), .C2(n14206), .ZN(P1_U2869) );
  NAND2_X1 U16250 ( .A1(n13088), .A2(n13089), .ZN(n13324) );
  OAI211_X1 U16251 ( .C1(n13089), .C2(n13088), .A(n13324), .B(n13661), .ZN(
        n13090) );
  INV_X1 U16252 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13163) );
  XNOR2_X1 U16253 ( .A(n13156), .B(n13163), .ZN(n13155) );
  NAND2_X1 U16254 ( .A1(n13093), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13094) );
  XNOR2_X1 U16255 ( .A(n13155), .B(n13154), .ZN(n13374) );
  OAI21_X1 U16256 ( .B1(n19915), .B2(n13336), .A(n14699), .ZN(n13173) );
  OAI21_X1 U16257 ( .B1(n14505), .B2(n15730), .A(n19915), .ZN(n15722) );
  INV_X1 U16258 ( .A(n15722), .ZN(n13667) );
  NOR2_X1 U16259 ( .A1(n13095), .A2(n13667), .ZN(n13340) );
  AOI22_X1 U16260 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13173), .B1(
        n13340), .B2(n13163), .ZN(n13098) );
  INV_X1 U16261 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20550) );
  NOR2_X1 U16262 ( .A1(n19921), .A2(n20550), .ZN(n13368) );
  AOI21_X1 U16263 ( .B1(n19911), .B2(n13096), .A(n13368), .ZN(n13097) );
  OAI211_X1 U16264 ( .C1(n14704), .C2(n13374), .A(n13098), .B(n13097), .ZN(
        P1_U3028) );
  OR2_X1 U16265 ( .A1(n13081), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13099) );
  NAND2_X1 U16266 ( .A1(n13100), .A2(n13099), .ZN(n19909) );
  INV_X1 U16267 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13464) );
  OAI222_X1 U16268 ( .A1(n19909), .A2(n14206), .B1(n13464), .B2(n19850), .C1(
        n14208), .C2(n13101), .ZN(P1_U2872) );
  NOR2_X1 U16269 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n15606), .ZN(n13133) );
  OR2_X1 U16270 ( .A1(n13102), .A2(n14709), .ZN(n13111) );
  NAND2_X1 U16271 ( .A1(n13103), .A2(n13112), .ZN(n13118) );
  AND2_X1 U16272 ( .A1(n13118), .A2(n13122), .ZN(n13106) );
  NAND3_X1 U16273 ( .A1(n14709), .A2(n13124), .A3(n13106), .ZN(n13109) );
  XNOR2_X1 U16274 ( .A(n13112), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13107) );
  OR2_X1 U16275 ( .A1(n13105), .A2(n13104), .ZN(n13120) );
  INV_X1 U16276 ( .A(n13106), .ZN(n14725) );
  AOI22_X1 U16277 ( .A1(n14712), .A2(n13107), .B1(n13120), .B2(n14725), .ZN(
        n13108) );
  AND2_X1 U16278 ( .A1(n13109), .A2(n13108), .ZN(n13110) );
  NAND2_X1 U16279 ( .A1(n13111), .A2(n13110), .ZN(n14723) );
  OR2_X1 U16280 ( .A1(n15585), .A2(n14723), .ZN(n13114) );
  NAND2_X1 U16281 ( .A1(n15585), .A2(n13112), .ZN(n13113) );
  AND2_X1 U16282 ( .A1(n13114), .A2(n13113), .ZN(n15588) );
  AOI22_X1 U16283 ( .A1(n13133), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15588), .B2(n15606), .ZN(n13128) );
  INV_X1 U16284 ( .A(n20221), .ZN(n13294) );
  MUX2_X1 U16285 ( .A(n13115), .B(n11305), .S(n11512), .Z(n13117) );
  NOR2_X1 U16286 ( .A1(n13117), .A2(n13116), .ZN(n13121) );
  XNOR2_X1 U16287 ( .A(n13118), .B(n11305), .ZN(n13119) );
  AOI22_X1 U16288 ( .A1(n14712), .A2(n13121), .B1(n13120), .B2(n13119), .ZN(
        n13126) );
  NAND2_X1 U16289 ( .A1(n13122), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13123) );
  NAND2_X1 U16290 ( .A1(n11564), .A2(n13123), .ZN(n20608) );
  NAND3_X1 U16291 ( .A1(n14709), .A2(n13124), .A3(n20608), .ZN(n13125) );
  OAI211_X1 U16292 ( .C1(n13294), .C2(n14709), .A(n13126), .B(n13125), .ZN(
        n20607) );
  MUX2_X1 U16293 ( .A(n20607), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15585), .Z(n15592) );
  AOI22_X1 U16294 ( .A1(n13133), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n15606), .B2(n15592), .ZN(n13127) );
  NOR2_X1 U16295 ( .A1(n13128), .A2(n13127), .ZN(n15598) );
  INV_X1 U16296 ( .A(n11316), .ZN(n13129) );
  NAND2_X1 U16297 ( .A1(n15598), .A2(n13129), .ZN(n14705) );
  AOI21_X1 U16298 ( .B1(n13130), .B2(n19815), .A(n15585), .ZN(n13131) );
  AOI211_X1 U16299 ( .C1(n15585), .C2(n12771), .A(P1_STATE2_REG_1__SCAN_IN), 
        .B(n13131), .ZN(n13132) );
  AOI21_X1 U16300 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13133), .A(
        n13132), .ZN(n15600) );
  NAND3_X1 U16301 ( .A1(n14705), .A2(n15600), .A3(n19749), .ZN(n13136) );
  INV_X1 U16302 ( .A(n15782), .ZN(n13135) );
  NAND2_X1 U16303 ( .A1(n11609), .A2(n15606), .ZN(n20626) );
  INV_X1 U16304 ( .A(n20626), .ZN(n13134) );
  NAND2_X1 U16305 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20357), .ZN(n14706) );
  NAND2_X1 U16306 ( .A1(n13153), .A2(n14706), .ZN(n13884) );
  NAND2_X1 U16307 ( .A1(n13153), .A2(n20398), .ZN(n13880) );
  INV_X1 U16308 ( .A(n20010), .ZN(n13881) );
  NAND2_X1 U16309 ( .A1(n20426), .A2(n13881), .ZN(n20402) );
  NAND3_X1 U16310 ( .A1(n20323), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n20402), 
        .ZN(n13139) );
  NAND2_X1 U16311 ( .A1(n20010), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20322) );
  INV_X1 U16312 ( .A(n20322), .ZN(n20194) );
  AOI22_X1 U16313 ( .A1(n13139), .A2(n9817), .B1(n20194), .B2(n20199), .ZN(
        n13140) );
  OAI222_X1 U16314 ( .A1(n13153), .A2(n20276), .B1(n13884), .B2(n13294), .C1(
        n13880), .C2(n13140), .ZN(P1_U3475) );
  AOI21_X1 U16315 ( .B1(n13141), .B2(n13068), .A(n13194), .ZN(n18715) );
  INV_X1 U16316 ( .A(n18715), .ZN(n13149) );
  INV_X1 U16317 ( .A(n13142), .ZN(n13146) );
  OAI21_X1 U16318 ( .B1(n12950), .B2(n13144), .A(n13143), .ZN(n13145) );
  NAND3_X1 U16319 ( .A1(n13146), .A2(n18848), .A3(n13145), .ZN(n13148) );
  NAND2_X1 U16320 ( .A1(n18843), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13147) );
  OAI211_X1 U16321 ( .C1(n13149), .C2(n18843), .A(n13148), .B(n13147), .ZN(
        P2_U2875) );
  AOI22_X1 U16322 ( .A1(n14848), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n14847), .ZN(n18951) );
  AOI21_X1 U16323 ( .B1(n15283), .B2(n13150), .A(n13180), .ZN(n18714) );
  INV_X1 U16324 ( .A(n18714), .ZN(n13151) );
  INV_X1 U16325 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18899) );
  OAI222_X1 U16326 ( .A1(n13439), .A2(n18951), .B1(n13151), .B2(n18890), .C1(
        n18899), .C2(n14858), .ZN(P2_U2907) );
  OAI222_X1 U16327 ( .A1(n13884), .A2(n13102), .B1(n13153), .B2(n20220), .C1(
        n13880), .C2(n13152), .ZN(P1_U3476) );
  NAND2_X1 U16328 ( .A1(n13156), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13157) );
  NAND2_X1 U16329 ( .A1(n13158), .A2(n13645), .ZN(n13162) );
  XNOR2_X1 U16330 ( .A(n13324), .B(n13159), .ZN(n13160) );
  NAND2_X1 U16331 ( .A1(n13160), .A2(n13661), .ZN(n13161) );
  NAND2_X1 U16332 ( .A1(n13162), .A2(n13161), .ZN(n13334) );
  INV_X1 U16333 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13164) );
  XNOR2_X1 U16334 ( .A(n13334), .B(n13164), .ZN(n13332) );
  XNOR2_X1 U16335 ( .A(n13333), .B(n13332), .ZN(n13437) );
  NOR2_X1 U16336 ( .A1(n13164), .A2(n13163), .ZN(n13339) );
  INV_X1 U16337 ( .A(n13339), .ZN(n14504) );
  OAI211_X1 U16338 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13340), .B(n14504), .ZN(n13175) );
  INV_X1 U16339 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n13171) );
  OAI21_X1 U16340 ( .B1(n13951), .B2(n13164), .A(n13938), .ZN(n13165) );
  OAI21_X1 U16341 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n13945), .A(n13165), .ZN(
        n13167) );
  INV_X1 U16342 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13279) );
  NAND2_X1 U16343 ( .A1(n13943), .A2(n13279), .ZN(n13166) );
  NAND2_X1 U16344 ( .A1(n13167), .A2(n13166), .ZN(n13168) );
  OR2_X1 U16345 ( .A1(n13169), .A2(n13168), .ZN(n13170) );
  NAND2_X1 U16346 ( .A1(n13347), .A2(n13170), .ZN(n19820) );
  OAI22_X1 U16347 ( .A1(n19921), .A2(n13171), .B1(n15775), .B2(n19820), .ZN(
        n13172) );
  AOI21_X1 U16348 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13173), .A(
        n13172), .ZN(n13174) );
  OAI211_X1 U16349 ( .C1(n14704), .C2(n13437), .A(n13175), .B(n13174), .ZN(
        P1_U3027) );
  INV_X1 U16350 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13176) );
  OR2_X1 U16351 ( .A1(n14847), .A2(n13176), .ZN(n13178) );
  NAND2_X1 U16352 ( .A1(n14847), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13177) );
  AND2_X1 U16353 ( .A1(n13178), .A2(n13177), .ZN(n18953) );
  INV_X1 U16354 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18897) );
  OAI21_X1 U16355 ( .B1(n13180), .B2(n13179), .A(n15957), .ZN(n18702) );
  OAI222_X1 U16356 ( .A1(n13439), .A2(n18953), .B1(n14858), .B2(n18897), .C1(
        n18890), .C2(n18702), .ZN(P2_U2906) );
  XNOR2_X1 U16357 ( .A(n13181), .B(n9699), .ZN(n13580) );
  INV_X1 U16358 ( .A(n13580), .ZN(n19694) );
  INV_X1 U16359 ( .A(n13182), .ZN(n13183) );
  NAND2_X1 U16360 ( .A1(n13184), .A2(n13183), .ZN(n13186) );
  XNOR2_X1 U16361 ( .A(n19277), .B(n13580), .ZN(n13185) );
  NAND2_X1 U16362 ( .A1(n13186), .A2(n13185), .ZN(n13425) );
  OAI21_X1 U16363 ( .B1(n13186), .B2(n13185), .A(n13425), .ZN(n13187) );
  NAND2_X1 U16364 ( .A1(n13187), .A2(n18884), .ZN(n13190) );
  AOI22_X1 U16365 ( .A1(n14848), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14847), .ZN(n19017) );
  INV_X1 U16366 ( .A(n19017), .ZN(n13188) );
  AOI22_X1 U16367 ( .A1(n18883), .A2(n13188), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n18881), .ZN(n13189) );
  OAI211_X1 U16368 ( .C1(n19694), .C2(n18862), .A(n13190), .B(n13189), .ZN(
        P2_U2916) );
  INV_X1 U16369 ( .A(n13191), .ZN(n13192) );
  AOI21_X1 U16370 ( .B1(n13193), .B2(n13078), .A(n13192), .ZN(n19824) );
  INV_X1 U16371 ( .A(n19824), .ZN(n13278) );
  INV_X1 U16372 ( .A(n14245), .ZN(n19960) );
  INV_X1 U16373 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19875) );
  OAI222_X1 U16374 ( .A1(n13278), .A2(n14279), .B1(n14272), .B2(n19960), .C1(
        n14270), .C2(n19875), .ZN(P1_U2900) );
  XNOR2_X1 U16375 ( .A(n13142), .B(n13377), .ZN(n13198) );
  OR2_X1 U16376 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  NAND2_X1 U16377 ( .A1(n13380), .A2(n13196), .ZN(n18703) );
  MUX2_X1 U16378 ( .A(n18703), .B(n10792), .S(n18843), .Z(n13197) );
  OAI21_X1 U16379 ( .B1(n13198), .B2(n18844), .A(n13197), .ZN(P2_U2874) );
  INV_X1 U16380 ( .A(n13229), .ZN(n13270) );
  NAND2_X1 U16381 ( .A1(n13199), .A2(n13236), .ZN(n13212) );
  NAND2_X1 U16382 ( .A1(n13200), .A2(n15352), .ZN(n13217) );
  NAND2_X1 U16383 ( .A1(n10336), .A2(n13217), .ZN(n13203) );
  NAND2_X1 U16384 ( .A1(n13212), .A2(n13203), .ZN(n13209) );
  NAND2_X1 U16385 ( .A1(n13202), .A2(n13201), .ZN(n13215) );
  INV_X1 U16386 ( .A(n13203), .ZN(n13204) );
  NAND2_X1 U16387 ( .A1(n13215), .A2(n13204), .ZN(n13208) );
  NOR2_X1 U16388 ( .A1(n13205), .A2(n13216), .ZN(n13206) );
  NAND2_X1 U16389 ( .A1(n13256), .A2(n13206), .ZN(n13207) );
  NAND3_X1 U16390 ( .A1(n13209), .A2(n13208), .A3(n13207), .ZN(n13210) );
  AOI21_X1 U16391 ( .B1(n18983), .B2(n13252), .A(n13210), .ZN(n15348) );
  MUX2_X1 U16392 ( .A(n15352), .B(n15348), .S(n13229), .Z(n13247) );
  OAI21_X1 U16393 ( .B1(n13247), .B2(n13211), .A(n12220), .ZN(n13269) );
  INV_X1 U16394 ( .A(n13247), .ZN(n13230) );
  INV_X1 U16395 ( .A(n13252), .ZN(n13253) );
  OR2_X1 U16396 ( .A1(n12845), .A2(n13253), .ZN(n13227) );
  NAND2_X1 U16397 ( .A1(n13212), .A2(n13217), .ZN(n13214) );
  NAND2_X1 U16398 ( .A1(n13256), .A2(n13216), .ZN(n13213) );
  NAND2_X1 U16399 ( .A1(n13214), .A2(n13213), .ZN(n13223) );
  NAND2_X1 U16400 ( .A1(n13215), .A2(n10336), .ZN(n13221) );
  INV_X1 U16401 ( .A(n13216), .ZN(n13219) );
  INV_X1 U16402 ( .A(n13217), .ZN(n13218) );
  AOI21_X1 U16403 ( .B1(n13256), .B2(n13219), .A(n13218), .ZN(n13220) );
  NAND2_X1 U16404 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  MUX2_X1 U16405 ( .A(n13223), .B(n13222), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13225) );
  NOR2_X1 U16406 ( .A1(n13225), .A2(n13224), .ZN(n13226) );
  INV_X1 U16407 ( .A(n15355), .ZN(n13228) );
  NAND3_X1 U16408 ( .A1(n13230), .A2(n13229), .A3(n13228), .ZN(n13246) );
  NAND2_X1 U16409 ( .A1(n13231), .A2(n13237), .ZN(n13235) );
  NAND2_X1 U16410 ( .A1(n13233), .A2(n13232), .ZN(n13234) );
  OAI211_X1 U16411 ( .C1(n13237), .C2(n13236), .A(n13235), .B(n13234), .ZN(
        n19730) );
  INV_X1 U16412 ( .A(n19730), .ZN(n13245) );
  AOI22_X1 U16413 ( .A1(n13241), .A2(n13240), .B1(n13239), .B2(n13238), .ZN(
        n13244) );
  OAI21_X1 U16414 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n13242), .ZN(n13243) );
  NAND4_X1 U16415 ( .A1(n13246), .A2(n13245), .A3(n13244), .A4(n13243), .ZN(
        n13268) );
  NOR2_X1 U16416 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13247), .ZN(
        n13263) );
  INV_X1 U16417 ( .A(n13248), .ZN(n13250) );
  NAND2_X1 U16418 ( .A1(n13250), .A2(n13249), .ZN(n13255) );
  MUX2_X1 U16419 ( .A(n13255), .B(n13256), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13251) );
  AOI21_X1 U16420 ( .B1(n18832), .B2(n13252), .A(n13251), .ZN(n15337) );
  AOI21_X1 U16421 ( .B1(n15337), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13260) );
  OR2_X1 U16422 ( .A1(n9592), .A2(n13253), .ZN(n13258) );
  NOR2_X1 U16423 ( .A1(n10343), .A2(n10342), .ZN(n13254) );
  AOI22_X1 U16424 ( .A1(n13256), .A2(n10330), .B1(n13255), .B2(n13254), .ZN(
        n13257) );
  NAND2_X1 U16425 ( .A1(n13258), .A2(n13257), .ZN(n15343) );
  AOI21_X1 U16426 ( .B1(n15337), .B2(n19368), .A(n13270), .ZN(n13259) );
  OAI21_X1 U16427 ( .B1(n13260), .B2(n15343), .A(n13259), .ZN(n13261) );
  AOI21_X1 U16428 ( .B1(n15355), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n13261), .ZN(n13262) );
  AOI222_X1 U16429 ( .A1(n13263), .A2(n13262), .B1(n13263), .B2(n12211), .C1(
        n13262), .C2(n12211), .ZN(n13266) );
  NAND2_X1 U16430 ( .A1(n13264), .A2(n13228), .ZN(n13265) );
  AOI21_X1 U16431 ( .B1(n13266), .B2(n13265), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n13267) );
  AOI211_X1 U16432 ( .C1(n13270), .C2(n13269), .A(n13268), .B(n13267), .ZN(
        n16004) );
  AND2_X1 U16433 ( .A1(n16004), .A2(n10711), .ZN(n13275) );
  OR3_X1 U16434 ( .A1(n13272), .A2(n13271), .A3(n19006), .ZN(n13273) );
  OAI211_X1 U16435 ( .C1(n13275), .C2(n18596), .A(n13274), .B(n13273), .ZN(
        n15996) );
  INV_X1 U16436 ( .A(n15996), .ZN(n13276) );
  NOR2_X1 U16437 ( .A1(n13276), .A2(n18596), .ZN(n13277) );
  OAI21_X1 U16438 ( .B1(n13277), .B2(n19544), .A(n15993), .ZN(P2_U3593) );
  OAI222_X1 U16439 ( .A1(n19820), .A2(n14206), .B1(n13279), .B2(n19850), .C1(
        n13278), .C2(n14208), .ZN(P1_U2868) );
  AND2_X1 U16440 ( .A1(n20623), .A2(n20429), .ZN(n15602) );
  OAI21_X1 U16441 ( .B1(n13289), .B2(n15603), .A(n15602), .ZN(n13298) );
  OR2_X2 U16442 ( .A1(n13300), .A2(n13298), .ZN(n13958) );
  AND2_X1 U16444 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n15614), .ZN(n13286) );
  NOR3_X1 U16445 ( .A1(n13284), .A2(n19931), .A3(n20626), .ZN(n13285) );
  AOI21_X1 U16446 ( .B1(n12096), .B2(n13286), .A(n13285), .ZN(n13287) );
  INV_X1 U16447 ( .A(n13308), .ZN(n13288) );
  INV_X1 U16448 ( .A(n13370), .ZN(n13307) );
  INV_X1 U16449 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13303) );
  NAND2_X1 U16450 ( .A1(n13289), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13297) );
  INV_X1 U16451 ( .A(n13297), .ZN(n13291) );
  INV_X1 U16452 ( .A(n15602), .ZN(n13290) );
  NAND2_X1 U16453 ( .A1(n13291), .A2(n13290), .ZN(n13292) );
  OR2_X1 U16454 ( .A1(n20628), .A2(n13293), .ZN(n19814) );
  OAI22_X1 U16455 ( .A1(n19791), .A2(n13295), .B1(n13294), .B2(n19814), .ZN(
        n13296) );
  INV_X1 U16456 ( .A(n13296), .ZN(n13302) );
  NAND2_X1 U16457 ( .A1(n13298), .A2(n13297), .ZN(n13299) );
  NAND2_X1 U16458 ( .A1(n19834), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n13301) );
  OAI211_X1 U16459 ( .C1(n19782), .C2(n13303), .A(n13302), .B(n13301), .ZN(
        n13306) );
  NAND2_X1 U16460 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n19837), .ZN(n19802) );
  NAND2_X1 U16461 ( .A1(n19802), .A2(n19801), .ZN(n13317) );
  NOR2_X1 U16462 ( .A1(n13317), .A2(n20550), .ZN(n13305) );
  AOI211_X1 U16463 ( .C1(n19822), .C2(n13307), .A(n13306), .B(n13305), .ZN(
        n13311) );
  OAI21_X1 U16464 ( .B1(n20628), .B2(n13309), .A(n19771), .ZN(n19840) );
  NAND2_X1 U16465 ( .A1(n13372), .A2(n19840), .ZN(n13310) );
  OAI211_X1 U16466 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(n19817), .A(n13311), .B(
        n13310), .ZN(P1_U2837) );
  OAI22_X1 U16467 ( .A1(n19791), .A2(n13312), .B1(n13102), .B2(n19814), .ZN(
        n13313) );
  INV_X1 U16468 ( .A(n13313), .ZN(n13315) );
  AOI22_X1 U16469 ( .A1(n19834), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n19830), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13314) );
  OAI211_X1 U16470 ( .C1(n19843), .C2(n13354), .A(n13315), .B(n13314), .ZN(
        n13320) );
  NOR2_X1 U16471 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n13316), .ZN(n13318) );
  NOR2_X1 U16472 ( .A1(n13318), .A2(n13317), .ZN(n13319) );
  AOI211_X1 U16473 ( .C1(n13356), .C2(n19840), .A(n13320), .B(n13319), .ZN(
        n13321) );
  INV_X1 U16474 ( .A(n13321), .ZN(P1_U2838) );
  NAND2_X1 U16475 ( .A1(n13322), .A2(n13645), .ZN(n13331) );
  NOR2_X1 U16476 ( .A1(n13324), .A2(n13323), .ZN(n13326) );
  NAND2_X1 U16477 ( .A1(n13326), .A2(n13325), .ZN(n13647) );
  INV_X1 U16478 ( .A(n13326), .ZN(n13328) );
  AOI21_X1 U16479 ( .B1(n13328), .B2(n13327), .A(n12756), .ZN(n13329) );
  NAND2_X1 U16480 ( .A1(n13647), .A2(n13329), .ZN(n13330) );
  NAND2_X1 U16481 ( .A1(n13331), .A2(n13330), .ZN(n13482) );
  INV_X1 U16482 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14506) );
  XNOR2_X1 U16483 ( .A(n13482), .B(n14506), .ZN(n13480) );
  NAND2_X1 U16484 ( .A1(n13334), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13335) );
  XNOR2_X1 U16485 ( .A(n13480), .B(n13481), .ZN(n13367) );
  NAND3_X1 U16486 ( .A1(n13339), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n13336), .ZN(n15737) );
  AOI21_X1 U16487 ( .B1(n15736), .B2(n15737), .A(n15735), .ZN(n13338) );
  NAND2_X1 U16488 ( .A1(n14658), .A2(n14505), .ZN(n13337) );
  OAI211_X1 U16489 ( .C1(n15740), .C2(n13339), .A(n13338), .B(n13337), .ZN(
        n13665) );
  NOR2_X1 U16490 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14504), .ZN(
        n13666) );
  AOI22_X1 U16491 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13665), .B1(
        n13666), .B2(n13340), .ZN(n13350) );
  INV_X1 U16492 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13341) );
  NAND2_X1 U16493 ( .A1(n13937), .A2(n13341), .ZN(n13345) );
  NAND2_X1 U16494 ( .A1(n13949), .A2(n13341), .ZN(n13343) );
  OAI211_X1 U16495 ( .C1(n13951), .C2(n14506), .A(n13343), .B(n13938), .ZN(
        n13344) );
  NAND2_X1 U16496 ( .A1(n13345), .A2(n13344), .ZN(n13346) );
  NAND2_X1 U16497 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  AND2_X1 U16498 ( .A1(n13444), .A2(n13348), .ZN(n19803) );
  INV_X1 U16499 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20554) );
  NOR2_X1 U16500 ( .A1(n19921), .A2(n20554), .ZN(n13363) );
  AOI21_X1 U16501 ( .B1(n19911), .B2(n19803), .A(n13363), .ZN(n13349) );
  OAI211_X1 U16502 ( .C1(n14704), .C2(n13367), .A(n13350), .B(n13349), .ZN(
        P1_U3026) );
  INV_X1 U16503 ( .A(n19924), .ZN(n15693) );
  AOI21_X1 U16504 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13352), .ZN(n13353) );
  OAI21_X1 U16505 ( .B1(n15696), .B2(n13354), .A(n13353), .ZN(n13355) );
  AOI21_X1 U16506 ( .B1(n13356), .B2(n15693), .A(n13355), .ZN(n13357) );
  OAI21_X1 U16507 ( .B1(n19748), .B2(n13358), .A(n13357), .ZN(P1_U2997) );
  INV_X1 U16508 ( .A(n13359), .ZN(n13360) );
  AOI21_X1 U16509 ( .B1(n13361), .B2(n13191), .A(n13360), .ZN(n19809) );
  INV_X1 U16510 ( .A(n19809), .ZN(n13385) );
  AOI22_X1 U16511 ( .A1(n19845), .A2(n19803), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14197), .ZN(n13362) );
  OAI21_X1 U16512 ( .B1(n13385), .B2(n14196), .A(n13362), .ZN(P1_U2867) );
  AOI21_X1 U16513 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13363), .ZN(n13364) );
  OAI21_X1 U16514 ( .B1(n15696), .B2(n19812), .A(n13364), .ZN(n13365) );
  AOI21_X1 U16515 ( .B1(n19809), .B2(n15693), .A(n13365), .ZN(n13366) );
  OAI21_X1 U16516 ( .B1(n19748), .B2(n13367), .A(n13366), .ZN(P1_U2994) );
  AOI21_X1 U16517 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13368), .ZN(n13369) );
  OAI21_X1 U16518 ( .B1(n15696), .B2(n13370), .A(n13369), .ZN(n13371) );
  AOI21_X1 U16519 ( .B1(n13372), .B2(n15693), .A(n13371), .ZN(n13373) );
  OAI21_X1 U16520 ( .B1(n19748), .B2(n13374), .A(n13373), .ZN(P1_U2996) );
  AOI21_X1 U16521 ( .B1(n13142), .B2(n13377), .A(n13376), .ZN(n13378) );
  OR3_X1 U16522 ( .A1(n10007), .A2(n13378), .A3(n18844), .ZN(n13383) );
  NAND2_X1 U16523 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  NAND2_X1 U16524 ( .A1(n18692), .A2(n18851), .ZN(n13382) );
  OAI211_X1 U16525 ( .C1(n18851), .C2(n13384), .A(n13383), .B(n13382), .ZN(
        P2_U2873) );
  INV_X1 U16526 ( .A(n14241), .ZN(n19965) );
  OAI222_X1 U16527 ( .A1(n13385), .A2(n14279), .B1(n14272), .B2(n19965), .C1(
        n14270), .C2(n11611), .ZN(P1_U2899) );
  AND2_X1 U16528 ( .A1(n13359), .A2(n13386), .ZN(n13389) );
  OR2_X1 U16529 ( .A1(n13389), .A2(n13388), .ZN(n13483) );
  INV_X1 U16530 ( .A(n14236), .ZN(n19970) );
  OAI222_X1 U16531 ( .A1(n13483), .A2(n14279), .B1(n14272), .B2(n19970), .C1(
        n14270), .C2(n11679), .ZN(P1_U2898) );
  NAND2_X1 U16532 ( .A1(n13391), .A2(n13390), .ZN(n13393) );
  XNOR2_X1 U16533 ( .A(n13393), .B(n13392), .ZN(n13408) );
  NOR2_X1 U16534 ( .A1(n12845), .A2(n15063), .ZN(n13395) );
  INV_X1 U16535 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13574) );
  OAI22_X1 U16536 ( .A1(n13574), .A2(n15953), .B1(n15922), .B2(n13572), .ZN(
        n13394) );
  AOI211_X1 U16537 ( .C1(n18791), .C2(P2_REIP_REG_3__SCAN_IN), .A(n13395), .B(
        n13394), .ZN(n13400) );
  OR2_X1 U16538 ( .A1(n9689), .A2(n13396), .ZN(n13405) );
  NAND3_X1 U16539 ( .A1(n13405), .A2(n15939), .A3(n13398), .ZN(n13399) );
  OAI211_X1 U16540 ( .C1(n13408), .C2(n15946), .A(n13400), .B(n13399), .ZN(
        P2_U3011) );
  OAI22_X1 U16541 ( .A1(n12845), .A2(n15330), .B1(n10292), .B2(n15891), .ZN(
        n13404) );
  AOI21_X1 U16542 ( .B1(n13402), .B2(n13401), .A(n13536), .ZN(n13403) );
  AOI211_X1 U16543 ( .C1(n15982), .C2(n13580), .A(n13404), .B(n13403), .ZN(
        n13407) );
  NAND3_X1 U16544 ( .A1(n13405), .A2(n18977), .A3(n13398), .ZN(n13406) );
  OAI211_X1 U16545 ( .C1(n13408), .C2(n15309), .A(n13407), .B(n13406), .ZN(
        P2_U3043) );
  NAND2_X1 U16546 ( .A1(n19617), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15628) );
  INV_X1 U16547 ( .A(n15342), .ZN(n19691) );
  OAI21_X1 U16548 ( .B1(n15628), .B2(n19691), .A(n16003), .ZN(n13411) );
  NAND2_X1 U16549 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13409), .ZN(n15992) );
  AOI211_X1 U16550 ( .C1(n15996), .C2(n15992), .A(n19617), .B(n10711), .ZN(
        n13410) );
  AOI211_X1 U16551 ( .C1(n15996), .C2(n13411), .A(n18819), .B(n13410), .ZN(
        n13412) );
  INV_X1 U16552 ( .A(n13412), .ZN(P2_U3177) );
  INV_X1 U16553 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13416) );
  OAI22_X1 U16554 ( .A1(n14459), .A2(n13416), .B1(n19921), .B2(n20547), .ZN(
        n13415) );
  NOR2_X1 U16555 ( .A1(n13413), .A2(n19924), .ZN(n13414) );
  AOI211_X1 U16556 ( .C1(n15681), .C2(n13416), .A(n13415), .B(n13414), .ZN(
        n13417) );
  OAI21_X1 U16557 ( .B1(n13418), .B2(n19748), .A(n13417), .ZN(P1_U2998) );
  INV_X1 U16558 ( .A(n13419), .ZN(n13420) );
  NAND2_X1 U16559 ( .A1(n13421), .A2(n13420), .ZN(n13423) );
  OAI21_X1 U16560 ( .B1(n13424), .B2(n13423), .A(n13422), .ZN(n18808) );
  INV_X1 U16561 ( .A(n19277), .ZN(n19696) );
  OAI21_X1 U16562 ( .B1(n19696), .B2(n13580), .A(n13425), .ZN(n13428) );
  XNOR2_X1 U16563 ( .A(n13427), .B(n13426), .ZN(n18804) );
  NAND2_X1 U16564 ( .A1(n13428), .A2(n18804), .ZN(n18886) );
  XOR2_X1 U16565 ( .A(n18808), .B(n18886), .Z(n13432) );
  INV_X1 U16566 ( .A(n18804), .ZN(n13429) );
  AOI22_X1 U16567 ( .A1(n18852), .A2(n13429), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n18881), .ZN(n13431) );
  INV_X1 U16568 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16123) );
  INV_X1 U16569 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U16570 ( .A1(n14848), .A2(n16123), .B1(n17937), .B2(n14847), .ZN(
        n18931) );
  NAND2_X1 U16571 ( .A1(n18883), .A2(n18931), .ZN(n13430) );
  OAI211_X1 U16572 ( .C1(n13432), .C2(n18861), .A(n13431), .B(n13430), .ZN(
        P2_U2915) );
  NAND2_X1 U16573 ( .A1(n19824), .A2(n15693), .ZN(n13436) );
  OAI22_X1 U16574 ( .A1(n14459), .A2(n13433), .B1(n19921), .B2(n13171), .ZN(
        n13434) );
  AOI21_X1 U16575 ( .B1(n19823), .B2(n15681), .A(n13434), .ZN(n13435) );
  OAI211_X1 U16576 ( .C1(n13437), .C2(n19748), .A(n13436), .B(n13435), .ZN(
        P1_U2995) );
  AOI22_X1 U16577 ( .A1(n14848), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14847), .ZN(n18962) );
  OAI21_X1 U16578 ( .B1(n15955), .B2(n13438), .A(n15234), .ZN(n18679) );
  INV_X1 U16579 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n18893) );
  OAI222_X1 U16580 ( .A1(n13439), .A2(n18962), .B1(n18679), .B2(n18890), .C1(
        n18893), .C2(n14858), .ZN(P2_U2904) );
  INV_X1 U16581 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15770) );
  OAI21_X1 U16582 ( .B1(n13951), .B2(n15770), .A(n13938), .ZN(n13440) );
  OAI21_X1 U16583 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n13945), .A(n13440), .ZN(
        n13442) );
  INV_X1 U16584 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19789) );
  NAND2_X1 U16585 ( .A1(n13943), .A2(n19789), .ZN(n13441) );
  NAND2_X1 U16586 ( .A1(n13444), .A2(n13443), .ZN(n13445) );
  NAND2_X1 U16587 ( .A1(n15760), .A2(n13445), .ZN(n19792) );
  OAI222_X1 U16588 ( .A1(n19792), .A2(n14206), .B1(n19789), .B2(n19850), .C1(
        n13483), .C2(n14208), .ZN(P1_U2866) );
  NAND2_X1 U16589 ( .A1(n13454), .A2(n19544), .ZN(n13446) );
  NAND2_X1 U16590 ( .A1(n13264), .A2(n12211), .ZN(n19083) );
  INV_X1 U16591 ( .A(n19083), .ZN(n19085) );
  NAND2_X1 U16592 ( .A1(n19368), .A2(n19085), .ZN(n13453) );
  NAND2_X1 U16593 ( .A1(n13446), .A2(n13453), .ZN(n13449) );
  AND2_X1 U16594 ( .A1(n19277), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19245) );
  NAND2_X1 U16595 ( .A1(n19245), .A2(n19375), .ZN(n13447) );
  NAND2_X1 U16596 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19085), .ZN(
        n13451) );
  NAND2_X1 U16597 ( .A1(n13447), .A2(n13451), .ZN(n13448) );
  MUX2_X1 U16598 ( .A(n13449), .B(n13448), .S(n19688), .Z(n13450) );
  NAND2_X1 U16599 ( .A1(n13450), .A2(n19553), .ZN(n19133) );
  INV_X1 U16600 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13462) );
  INV_X1 U16601 ( .A(n18856), .ZN(n18940) );
  NOR2_X2 U16602 ( .A1(n18940), .A2(n19046), .ZN(n19547) );
  INV_X1 U16603 ( .A(n13451), .ZN(n13452) );
  NAND2_X1 U16604 ( .A1(n13452), .A2(n19688), .ZN(n13456) );
  INV_X1 U16605 ( .A(n13453), .ZN(n19130) );
  OAI21_X1 U16606 ( .B1(n13454), .B2(n19130), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13455) );
  NAND2_X1 U16607 ( .A1(n13456), .A2(n13455), .ZN(n19132) );
  INV_X1 U16608 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16097) );
  INV_X1 U16609 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17917) );
  OAI22_X2 U16610 ( .A1(n16097), .A2(n19039), .B1(n17917), .B2(n19037), .ZN(
        n19555) );
  INV_X1 U16611 ( .A(n19555), .ZN(n13459) );
  INV_X1 U16612 ( .A(n19558), .ZN(n19493) );
  NOR2_X2 U16613 ( .A1(n13457), .A2(n19022), .ZN(n19546) );
  AOI22_X1 U16614 ( .A1(n19493), .A2(n19166), .B1(n19130), .B2(n19546), .ZN(
        n13458) );
  OAI21_X1 U16615 ( .B1(n13459), .B2(n19112), .A(n13458), .ZN(n13460) );
  AOI21_X1 U16616 ( .B1(n19547), .B2(n19132), .A(n13460), .ZN(n13461) );
  OAI21_X1 U16617 ( .B1(n19125), .B2(n13462), .A(n13461), .ZN(P2_U3072) );
  OAI21_X1 U16618 ( .B1(n19822), .B2(n19830), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13468) );
  OAI22_X1 U16619 ( .A1(n19790), .A2(n13464), .B1(n13463), .B2(n19814), .ZN(
        n13466) );
  NOR2_X1 U16620 ( .A1(n19791), .A2(n19909), .ZN(n13465) );
  NOR2_X1 U16621 ( .A1(n13466), .A2(n13465), .ZN(n13467) );
  OAI211_X1 U16622 ( .C1(n19777), .C2(n12944), .A(n13468), .B(n13467), .ZN(
        n13469) );
  AOI21_X1 U16623 ( .B1(n19840), .B2(n13470), .A(n13469), .ZN(n13471) );
  INV_X1 U16624 ( .A(n13471), .ZN(P1_U2840) );
  AOI21_X1 U16625 ( .B1(n13388), .B2(n13472), .A(n13473), .ZN(n13474) );
  OR2_X1 U16626 ( .A1(n9673), .A2(n13474), .ZN(n13676) );
  MUX2_X1 U16627 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n19925), .Z(
        n19887) );
  AOI22_X1 U16628 ( .A1(n14277), .A2(n19887), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14275), .ZN(n13475) );
  OAI21_X1 U16629 ( .B1(n13676), .B2(n14279), .A(n13475), .ZN(P1_U2896) );
  NAND2_X1 U16630 ( .A1(n13476), .A2(n13645), .ZN(n13479) );
  XNOR2_X1 U16631 ( .A(n13647), .B(n13648), .ZN(n13477) );
  NAND2_X1 U16632 ( .A1(n13477), .A2(n13661), .ZN(n13478) );
  NAND2_X1 U16633 ( .A1(n13479), .A2(n13478), .ZN(n13643) );
  XNOR2_X1 U16634 ( .A(n13643), .B(n15770), .ZN(n13641) );
  XNOR2_X1 U16635 ( .A(n13641), .B(n13642), .ZN(n15768) );
  INV_X1 U16636 ( .A(n13483), .ZN(n19797) );
  INV_X2 U16637 ( .A(n19921), .ZN(n15772) );
  AOI22_X1 U16638 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n13484) );
  OAI21_X1 U16639 ( .B1(n15696), .B2(n19800), .A(n13484), .ZN(n13485) );
  AOI21_X1 U16640 ( .B1(n19797), .B2(n15693), .A(n13485), .ZN(n13486) );
  OAI21_X1 U16641 ( .B1(n19748), .B2(n15768), .A(n13486), .ZN(P1_U2993) );
  NAND2_X1 U16642 ( .A1(n19245), .A2(n19308), .ZN(n13488) );
  NOR2_X1 U16643 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19083), .ZN(
        n13495) );
  INV_X1 U16644 ( .A(n13495), .ZN(n13487) );
  NAND2_X1 U16645 ( .A1(n13488), .A2(n13487), .ZN(n13493) );
  NAND2_X1 U16646 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13495), .ZN(
        n19075) );
  NAND2_X1 U16647 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19075), .ZN(n13489) );
  NAND2_X1 U16648 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19075), .ZN(n13491) );
  AND3_X1 U16649 ( .A1(n13498), .A2(n19553), .A3(n13491), .ZN(n13492) );
  NAND2_X1 U16650 ( .A1(n13493), .A2(n13492), .ZN(n19071) );
  INV_X1 U16651 ( .A(n19071), .ZN(n19082) );
  INV_X1 U16652 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13503) );
  INV_X1 U16653 ( .A(n13494), .ZN(n19243) );
  NOR2_X1 U16654 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13495), .ZN(n13496) );
  NOR2_X1 U16655 ( .A1(n19243), .A2(n13496), .ZN(n13497) );
  NAND2_X1 U16656 ( .A1(n13498), .A2(n13497), .ZN(n19076) );
  INV_X1 U16657 ( .A(n19076), .ZN(n19063) );
  INV_X1 U16658 ( .A(n19546), .ZN(n13500) );
  NAND2_X1 U16659 ( .A1(n19308), .A2(n19238), .ZN(n19069) );
  AOI22_X1 U16660 ( .A1(n19078), .A2(n19555), .B1(n19108), .B2(n19493), .ZN(
        n13499) );
  OAI21_X1 U16661 ( .B1(n13500), .B2(n19075), .A(n13499), .ZN(n13501) );
  AOI21_X1 U16662 ( .B1(n19063), .B2(n19547), .A(n13501), .ZN(n13502) );
  OAI21_X1 U16663 ( .B1(n19082), .B2(n13503), .A(n13502), .ZN(P2_U3056) );
  INV_X1 U16664 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19849) );
  NAND2_X1 U16665 ( .A1(n13937), .A2(n19849), .ZN(n13506) );
  INV_X1 U16666 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13668) );
  NAND2_X1 U16667 ( .A1(n13949), .A2(n19849), .ZN(n13504) );
  OAI211_X1 U16668 ( .C1(n13951), .C2(n13668), .A(n13504), .B(n13938), .ZN(
        n13505) );
  NAND2_X1 U16669 ( .A1(n13506), .A2(n13505), .ZN(n15761) );
  INV_X1 U16670 ( .A(n13943), .ZN(n13900) );
  INV_X1 U16671 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13507) );
  OAI21_X1 U16672 ( .B1(n13951), .B2(n13507), .A(n13938), .ZN(n13510) );
  INV_X1 U16673 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13508) );
  NAND2_X1 U16674 ( .A1(n13949), .A2(n13508), .ZN(n13509) );
  NAND2_X1 U16675 ( .A1(n13510), .A2(n13509), .ZN(n13511) );
  OAI21_X1 U16676 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n13900), .A(n13511), .ZN(
        n13512) );
  OR2_X1 U16677 ( .A1(n9648), .A2(n13512), .ZN(n13513) );
  NAND2_X1 U16678 ( .A1(n13562), .A2(n13513), .ZN(n13669) );
  OAI222_X1 U16679 ( .A1(n13669), .A2(n14206), .B1(n19850), .B2(n13508), .C1(
        n13676), .C2(n14208), .ZN(P1_U2864) );
  INV_X1 U16680 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20556) );
  NAND2_X1 U16681 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .ZN(n19807) );
  NOR3_X1 U16682 ( .A1(n20556), .A2(n20554), .A3(n19807), .ZN(n19778) );
  NAND2_X1 U16683 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19778), .ZN(n13517) );
  INV_X1 U16684 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20559) );
  AOI22_X1 U16685 ( .A1(n19834), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n19830), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13514) );
  OAI211_X1 U16686 ( .C1(n19791), .C2(n13669), .A(n13514), .B(n19921), .ZN(
        n13516) );
  AND2_X1 U16687 ( .A1(n19822), .A2(n13673), .ZN(n13515) );
  AOI211_X1 U16688 ( .C1(n13720), .C2(n20559), .A(n13516), .B(n13515), .ZN(
        n13519) );
  NOR3_X1 U16689 ( .A1(n20559), .A2(n13517), .A3(n19802), .ZN(n13722) );
  NOR2_X1 U16690 ( .A1(n13722), .A2(n19777), .ZN(n19769) );
  NAND2_X1 U16691 ( .A1(n19769), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n13518) );
  OAI211_X1 U16692 ( .C1(n13676), .C2(n19771), .A(n13519), .B(n13518), .ZN(
        P1_U2832) );
  NAND2_X1 U16693 ( .A1(n9969), .A2(n13520), .ZN(n13521) );
  XNOR2_X1 U16694 ( .A(n13522), .B(n13521), .ZN(n13529) );
  OAI22_X1 U16695 ( .A1(n11262), .A2(n18833), .B1(n10276), .B2(n18825), .ZN(
        n13525) );
  OAI22_X1 U16696 ( .A1(n18987), .A2(n18823), .B1(n13523), .B2(n18822), .ZN(
        n13524) );
  AOI211_X1 U16697 ( .C1(P2_EBX_REG_2__SCAN_IN), .C2(n18803), .A(n13525), .B(
        n13524), .ZN(n13527) );
  NAND2_X1 U16698 ( .A1(n18983), .A2(n18831), .ZN(n13526) );
  OAI211_X1 U16699 ( .C1(n19139), .C2(n13583), .A(n13527), .B(n13526), .ZN(
        n13528) );
  AOI21_X1 U16700 ( .B1(n13529), .B2(n18819), .A(n13528), .ZN(n13530) );
  INV_X1 U16701 ( .A(n13530), .ZN(P2_U2853) );
  XOR2_X1 U16702 ( .A(n13388), .B(n13472), .Z(n19847) );
  INV_X1 U16703 ( .A(n19847), .ZN(n13532) );
  AOI22_X1 U16704 ( .A1(n14277), .A2(n19977), .B1(P1_EAX_REG_7__SCAN_IN), .B2(
        n14275), .ZN(n13531) );
  OAI21_X1 U16705 ( .B1(n13532), .B2(n14279), .A(n13531), .ZN(P1_U2897) );
  XNOR2_X1 U16706 ( .A(n13533), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13554) );
  XOR2_X1 U16707 ( .A(n13535), .B(n13534), .Z(n13552) );
  NOR2_X1 U16708 ( .A1(n13537), .A2(n13536), .ZN(n13631) );
  INV_X1 U16709 ( .A(n13631), .ZN(n13544) );
  NOR2_X1 U16710 ( .A1(n13539), .A2(n13538), .ZN(n13540) );
  OR2_X1 U16711 ( .A1(n12856), .A2(n13540), .ZN(n18809) );
  NOR2_X1 U16712 ( .A1(n18809), .A2(n15330), .ZN(n13542) );
  OAI22_X1 U16713 ( .A1(n18986), .A2(n18804), .B1(n10613), .B2(n15891), .ZN(
        n13541) );
  AOI211_X1 U16714 ( .C1(n13623), .C2(n20652), .A(n13542), .B(n13541), .ZN(
        n13543) );
  OAI21_X1 U16715 ( .B1(n13544), .B2(n20652), .A(n13543), .ZN(n13545) );
  AOI21_X1 U16716 ( .B1(n13552), .B2(n11303), .A(n13545), .ZN(n13546) );
  OAI21_X1 U16717 ( .B1(n13554), .B2(n15978), .A(n13546), .ZN(P2_U3042) );
  OAI22_X1 U16718 ( .A1(n13547), .A2(n15953), .B1(n10613), .B2(n15891), .ZN(
        n13548) );
  INV_X1 U16719 ( .A(n13548), .ZN(n13550) );
  NAND2_X1 U16720 ( .A1(n15944), .A2(n18814), .ZN(n13549) );
  OAI211_X1 U16721 ( .C1(n18809), .C2(n15063), .A(n13550), .B(n13549), .ZN(
        n13551) );
  AOI21_X1 U16722 ( .B1(n13552), .B2(n10903), .A(n13551), .ZN(n13553) );
  OAI21_X1 U16723 ( .B1(n13554), .B2(n15947), .A(n13553), .ZN(P2_U3010) );
  NOR2_X1 U16724 ( .A1(n9673), .A2(n13555), .ZN(n13556) );
  OR2_X1 U16725 ( .A1(n9684), .A2(n13556), .ZN(n19772) );
  INV_X1 U16726 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13557) );
  NAND2_X1 U16727 ( .A1(n13937), .A2(n13557), .ZN(n13560) );
  INV_X1 U16728 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14282) );
  NAND2_X1 U16729 ( .A1(n13949), .A2(n13557), .ZN(n13558) );
  OAI211_X1 U16730 ( .C1(n13951), .C2(n14282), .A(n13558), .B(n13938), .ZN(
        n13559) );
  NAND2_X1 U16731 ( .A1(n13560), .A2(n13559), .ZN(n13563) );
  INV_X1 U16732 ( .A(n13597), .ZN(n13561) );
  AOI21_X1 U16733 ( .B1(n13563), .B2(n13562), .A(n13561), .ZN(n19765) );
  AOI22_X1 U16734 ( .A1(n19845), .A2(n19765), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14197), .ZN(n13564) );
  OAI21_X1 U16735 ( .B1(n19772), .B2(n14196), .A(n13564), .ZN(P1_U2863) );
  XNOR2_X1 U16736 ( .A(n10007), .B(n13565), .ZN(n13570) );
  AND2_X1 U16737 ( .A1(n13567), .A2(n13566), .ZN(n13568) );
  OR2_X1 U16738 ( .A1(n13568), .A2(n15028), .ZN(n18680) );
  MUX2_X1 U16739 ( .A(n18680), .B(n18673), .S(n18843), .Z(n13569) );
  OAI21_X1 U16740 ( .B1(n13570), .B2(n18844), .A(n13569), .ZN(P2_U2872) );
  NOR2_X1 U16741 ( .A1(n18676), .A2(n13571), .ZN(n13573) );
  XNOR2_X1 U16742 ( .A(n13573), .B(n13572), .ZN(n13585) );
  OAI22_X1 U16743 ( .A1(n13574), .A2(n18833), .B1(n10292), .B2(n18825), .ZN(
        n13579) );
  NOR2_X1 U16744 ( .A1(n12845), .A2(n18796), .ZN(n13578) );
  INV_X1 U16745 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13576) );
  OAI22_X1 U16746 ( .A1(n18828), .A2(n13576), .B1(n13575), .B2(n18822), .ZN(
        n13577) );
  NOR3_X1 U16747 ( .A1(n13579), .A2(n13578), .A3(n13577), .ZN(n13582) );
  NAND2_X1 U16748 ( .A1(n13580), .A2(n18759), .ZN(n13581) );
  OAI211_X1 U16749 ( .C1(n19277), .C2(n13583), .A(n13582), .B(n13581), .ZN(
        n13584) );
  AOI21_X1 U16750 ( .B1(n13585), .B2(n18819), .A(n13584), .ZN(n13586) );
  INV_X1 U16751 ( .A(n13586), .ZN(P2_U2852) );
  OAI21_X1 U16752 ( .B1(n9684), .B2(n13588), .A(n13587), .ZN(n15676) );
  AOI22_X1 U16753 ( .A1(n14277), .A2(n14221), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14275), .ZN(n13589) );
  OAI21_X1 U16754 ( .B1(n15676), .B2(n14279), .A(n13589), .ZN(P1_U2894) );
  INV_X1 U16755 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13591) );
  NAND2_X1 U16756 ( .A1(n13943), .A2(n13591), .ZN(n13595) );
  INV_X1 U16757 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U16758 ( .A1(n13938), .A2(n13590), .ZN(n13593) );
  NAND2_X1 U16759 ( .A1(n13949), .A2(n13591), .ZN(n13592) );
  NAND3_X1 U16760 ( .A1(n13593), .A2(n13977), .A3(n13592), .ZN(n13594) );
  AND2_X1 U16761 ( .A1(n13597), .A2(n13596), .ZN(n13598) );
  OR2_X1 U16762 ( .A1(n13598), .A2(n13726), .ZN(n14700) );
  INV_X1 U16763 ( .A(n14700), .ZN(n15671) );
  AOI22_X1 U16764 ( .A1(n19845), .A2(n15671), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14197), .ZN(n13599) );
  OAI21_X1 U16765 ( .B1(n15676), .B2(n14196), .A(n13599), .ZN(P1_U2862) );
  INV_X1 U16766 ( .A(n14224), .ZN(n13601) );
  OAI222_X1 U16767 ( .A1(n19772), .A2(n14279), .B1(n14272), .B2(n13601), .C1(
        n13600), .C2(n14270), .ZN(P1_U2895) );
  NAND2_X1 U16768 ( .A1(n13603), .A2(n13604), .ZN(n13605) );
  NAND2_X1 U16769 ( .A1(n13602), .A2(n13605), .ZN(n13694) );
  INV_X1 U16770 ( .A(n13606), .ZN(n13607) );
  XNOR2_X1 U16771 ( .A(n15235), .B(n13607), .ZN(n18657) );
  NAND2_X1 U16772 ( .A1(n18657), .A2(n18852), .ZN(n13613) );
  OAI22_X1 U16773 ( .A1(n19007), .A2(n14859), .B1(n14858), .B2(n13608), .ZN(
        n13611) );
  INV_X1 U16774 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13609) );
  NOR2_X1 U16775 ( .A1(n14835), .A2(n13609), .ZN(n13610) );
  AOI211_X1 U16776 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n18859), .A(n13611), .B(
        n13610), .ZN(n13612) );
  OAI211_X1 U16777 ( .C1(n18861), .C2(n13694), .A(n13613), .B(n13612), .ZN(
        P2_U2902) );
  INV_X1 U16778 ( .A(n13614), .ZN(n13618) );
  OAI21_X1 U16779 ( .B1(n13618), .B2(n13616), .A(n13615), .ZN(n13617) );
  OAI21_X1 U16780 ( .B1(n13619), .B2(n13618), .A(n13617), .ZN(n13640) );
  XOR2_X1 U16781 ( .A(n13621), .B(n13620), .Z(n13634) );
  NAND2_X1 U16782 ( .A1(n13634), .A2(n11303), .ZN(n13633) );
  OAI211_X1 U16783 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n13623), .B(n13622), .ZN(n13629) );
  XNOR2_X1 U16784 ( .A(n13625), .B(n13624), .ZN(n18889) );
  INV_X1 U16785 ( .A(n18889), .ZN(n13627) );
  NOR2_X1 U16786 ( .A1(n18970), .A2(n13626), .ZN(n13636) );
  AOI21_X1 U16787 ( .B1(n15982), .B2(n13627), .A(n13636), .ZN(n13628) );
  OAI211_X1 U16788 ( .C1(n15330), .C2(n18795), .A(n13629), .B(n13628), .ZN(
        n13630) );
  AOI21_X1 U16789 ( .B1(n13631), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13630), .ZN(n13632) );
  OAI211_X1 U16790 ( .C1(n13640), .C2(n15978), .A(n13633), .B(n13632), .ZN(
        P2_U3041) );
  NAND2_X1 U16791 ( .A1(n13634), .A2(n10903), .ZN(n13639) );
  INV_X1 U16792 ( .A(n18795), .ZN(n13637) );
  INV_X1 U16793 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18789) );
  OAI22_X1 U16794 ( .A1(n18789), .A2(n15953), .B1(n15922), .B2(n18794), .ZN(
        n13635) );
  AOI211_X1 U16795 ( .C1(n13637), .C2(n15950), .A(n13636), .B(n13635), .ZN(
        n13638) );
  OAI211_X1 U16796 ( .C1(n15947), .C2(n13640), .A(n13639), .B(n13638), .ZN(
        P2_U3009) );
  NAND2_X1 U16797 ( .A1(n13643), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13644) );
  NAND2_X1 U16798 ( .A1(n13646), .A2(n13645), .ZN(n13652) );
  INV_X1 U16799 ( .A(n13647), .ZN(n13649) );
  NAND2_X1 U16800 ( .A1(n13649), .A2(n13648), .ZN(n13659) );
  XNOR2_X1 U16801 ( .A(n13659), .B(n13660), .ZN(n13650) );
  NAND2_X1 U16802 ( .A1(n13650), .A2(n13661), .ZN(n13651) );
  NAND2_X1 U16803 ( .A1(n13652), .A2(n13651), .ZN(n13653) );
  AND2_X1 U16804 ( .A1(n13653), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15687) );
  NOR3_X1 U16805 ( .A1(n13656), .A2(n13655), .A3(n15614), .ZN(n13657) );
  INV_X1 U16806 ( .A(n13659), .ZN(n13662) );
  NAND3_X1 U16807 ( .A1(n13662), .A2(n13661), .A3(n13660), .ZN(n13663) );
  NAND2_X1 U16808 ( .A1(n13658), .A2(n13663), .ZN(n13707) );
  XNOR2_X1 U16809 ( .A(n13707), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13664) );
  XNOR2_X1 U16810 ( .A(n13709), .B(n13664), .ZN(n13679) );
  AOI21_X1 U16811 ( .B1(n13062), .B2(n13666), .A(n13665), .ZN(n15767) );
  OAI21_X1 U16812 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14660), .A(
        n15767), .ZN(n15762) );
  NAND2_X1 U16813 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15771), .ZN(
        n15766) );
  AOI221_X1 U16814 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n13507), .C2(n13668), .A(
        n15766), .ZN(n13671) );
  OAI22_X1 U16815 ( .A1(n19921), .A2(n20559), .B1(n15775), .B2(n13669), .ZN(
        n13670) );
  AOI211_X1 U16816 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n15762), .A(
        n13671), .B(n13670), .ZN(n13672) );
  OAI21_X1 U16817 ( .B1(n13679), .B2(n14704), .A(n13672), .ZN(P1_U3023) );
  AOI22_X1 U16818 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U16819 ( .A1(n15681), .A2(n13673), .ZN(n13674) );
  OAI211_X1 U16820 ( .C1(n13676), .C2(n19924), .A(n13675), .B(n13674), .ZN(
        n13677) );
  INV_X1 U16821 ( .A(n13677), .ZN(n13678) );
  OAI21_X1 U16822 ( .B1(n13679), .B2(n19748), .A(n13678), .ZN(P1_U2991) );
  NAND2_X1 U16823 ( .A1(n13681), .A2(n13680), .ZN(n13682) );
  NAND2_X1 U16824 ( .A1(n14855), .A2(n13682), .ZN(n18649) );
  OAI22_X1 U16825 ( .A1(n19011), .A2(n14859), .B1(n14858), .B2(n13683), .ZN(
        n13686) );
  INV_X1 U16826 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n13684) );
  NOR2_X1 U16827 ( .A1(n14835), .A2(n13684), .ZN(n13685) );
  AOI211_X1 U16828 ( .C1(BUF1_REG_18__SCAN_IN), .C2(n18859), .A(n13686), .B(
        n13685), .ZN(n13690) );
  AOI21_X1 U16829 ( .B1(n13688), .B2(n13602), .A(n13687), .ZN(n15877) );
  NAND2_X1 U16830 ( .A1(n15877), .A2(n18884), .ZN(n13689) );
  OAI211_X1 U16831 ( .C1(n18649), .C2(n18862), .A(n13690), .B(n13689), .ZN(
        P2_U2901) );
  NAND2_X1 U16832 ( .A1(n18843), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13693) );
  AOI21_X1 U16833 ( .B1(n13691), .B2(n9624), .A(n10045), .ZN(n18656) );
  NAND2_X1 U16834 ( .A1(n18656), .A2(n18851), .ZN(n13692) );
  OAI211_X1 U16835 ( .C1(n13694), .C2(n18844), .A(n13693), .B(n13692), .ZN(
        P2_U2870) );
  XNOR2_X1 U16836 ( .A(n13695), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15948) );
  AND2_X1 U16837 ( .A1(n13696), .A2(n15267), .ZN(n15983) );
  INV_X1 U16838 ( .A(n18787), .ZN(n13698) );
  NOR2_X1 U16839 ( .A1(n10618), .A2(n18970), .ZN(n13697) );
  AOI21_X1 U16840 ( .B1(n15982), .B2(n13698), .A(n13697), .ZN(n13700) );
  NAND2_X1 U16841 ( .A1(n18783), .A2(n18982), .ZN(n13699) );
  OAI211_X1 U16842 ( .C1(n13701), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13700), .B(n13699), .ZN(n13702) );
  AOI21_X1 U16843 ( .B1(n15983), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13702), .ZN(n13706) );
  XNOR2_X1 U16844 ( .A(n13703), .B(n13704), .ZN(n15945) );
  OR2_X1 U16845 ( .A1(n15945), .A2(n15309), .ZN(n13705) );
  OAI211_X1 U16846 ( .C1(n15948), .C2(n15978), .A(n13706), .B(n13705), .ZN(
        P2_U3040) );
  NOR2_X1 U16847 ( .A1(n13707), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13708) );
  XNOR2_X1 U16848 ( .A(n9593), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13710) );
  XNOR2_X1 U16849 ( .A(n14281), .B(n13710), .ZN(n15756) );
  INV_X1 U16850 ( .A(n15756), .ZN(n13715) );
  INV_X1 U16851 ( .A(n19772), .ZN(n13713) );
  AOI22_X1 U16852 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13711) );
  OAI21_X1 U16853 ( .B1(n15696), .B2(n19770), .A(n13711), .ZN(n13712) );
  AOI21_X1 U16854 ( .B1(n13713), .B2(n15693), .A(n13712), .ZN(n13714) );
  OAI21_X1 U16855 ( .B1(n13715), .B2(n19748), .A(n13714), .ZN(P1_U2990) );
  INV_X1 U16856 ( .A(n13716), .ZN(n13717) );
  AOI21_X1 U16857 ( .B1(n13719), .B2(n13718), .A(n13717), .ZN(n14498) );
  INV_X1 U16858 ( .A(n14498), .ZN(n13746) );
  NAND2_X1 U16859 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n13721) );
  NOR2_X2 U16860 ( .A1(n19776), .A2(n13721), .ZN(n15659) );
  INV_X1 U16861 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20563) );
  NAND3_X1 U16862 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n13722), .ZN(n15649) );
  NAND2_X1 U16863 ( .A1(n15649), .A2(n19801), .ZN(n15674) );
  MUX2_X1 U16864 ( .A(n13937), .B(n13951), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13724) );
  NOR2_X1 U16865 ( .A1(n13081), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13723) );
  NOR2_X1 U16866 ( .A1(n13724), .A2(n13723), .ZN(n13725) );
  NOR2_X1 U16867 ( .A1(n13726), .A2(n13725), .ZN(n13727) );
  OR2_X1 U16868 ( .A1(n14200), .A2(n13727), .ZN(n13748) );
  INV_X1 U16869 ( .A(n13748), .ZN(n15748) );
  AOI22_X1 U16870 ( .A1(n19832), .A2(n15748), .B1(n19834), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n13728) );
  OAI21_X1 U16871 ( .B1(n20563), .B2(n15674), .A(n13728), .ZN(n13729) );
  AOI211_X1 U16872 ( .C1(n19830), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n13729), .B(n19819), .ZN(n13730) );
  OAI21_X1 U16873 ( .B1(n14496), .B2(n19843), .A(n13730), .ZN(n13731) );
  AOI21_X1 U16874 ( .B1(n15659), .B2(n20563), .A(n13731), .ZN(n13732) );
  OAI21_X1 U16875 ( .B1(n13746), .B2(n19771), .A(n13732), .ZN(P1_U2829) );
  INV_X1 U16876 ( .A(n14217), .ZN(n13733) );
  OAI222_X1 U16877 ( .A1(n13746), .A2(n14279), .B1(n14272), .B2(n13733), .C1(
        n19864), .C2(n14270), .ZN(P1_U2893) );
  INV_X1 U16878 ( .A(n13735), .ZN(n13737) );
  NAND3_X1 U16879 ( .A1(n13716), .A2(n13737), .A3(n13736), .ZN(n13738) );
  AND2_X1 U16880 ( .A1(n13734), .A2(n13738), .ZN(n15665) );
  INV_X1 U16881 ( .A(n15665), .ZN(n13745) );
  MUX2_X1 U16882 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n19925), .Z(
        n19889) );
  AOI22_X1 U16883 ( .A1(n14277), .A2(n19889), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14275), .ZN(n13739) );
  OAI21_X1 U16884 ( .B1(n13745), .B2(n14279), .A(n13739), .ZN(P1_U2892) );
  INV_X1 U16885 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15660) );
  NAND2_X1 U16886 ( .A1(n13943), .A2(n15660), .ZN(n13743) );
  INV_X1 U16887 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15729) );
  NAND2_X1 U16888 ( .A1(n13938), .A2(n15729), .ZN(n13741) );
  NAND2_X1 U16889 ( .A1(n13949), .A2(n15660), .ZN(n13740) );
  NAND3_X1 U16890 ( .A1(n13741), .A2(n13977), .A3(n13740), .ZN(n13742) );
  XNOR2_X1 U16891 ( .A(n14200), .B(n14202), .ZN(n15734) );
  AOI22_X1 U16892 ( .A1(n19845), .A2(n15734), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14197), .ZN(n13744) );
  OAI21_X1 U16893 ( .B1(n13745), .B2(n14196), .A(n13744), .ZN(P1_U2860) );
  INV_X1 U16894 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n13747) );
  OAI222_X1 U16895 ( .A1(n13748), .A2(n14206), .B1(n13747), .B2(n19850), .C1(
        n13746), .C2(n14208), .ZN(P1_U2861) );
  INV_X1 U16896 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18426) );
  INV_X1 U16897 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18520) );
  NAND2_X1 U16898 ( .A1(n18426), .A2(n18520), .ZN(n18530) );
  AOI22_X1 U16899 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13754) );
  AOI22_X1 U16900 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13753) );
  BUF_X2 U16901 ( .A(n16625), .Z(n16825) );
  AOI22_X1 U16902 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13752) );
  AOI22_X1 U16903 ( .A1(n16810), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13751) );
  NAND4_X1 U16904 ( .A1(n13754), .A2(n13753), .A3(n13752), .A4(n13751), .ZN(
        n13764) );
  INV_X2 U16905 ( .A(n10126), .ZN(n16908) );
  AOI22_X1 U16906 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13762) );
  AOI22_X1 U16907 ( .A1(n16894), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U16908 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13760) );
  INV_X1 U16909 ( .A(n15424), .ZN(n13758) );
  AOI22_X1 U16910 ( .A1(n16845), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13759) );
  NAND4_X1 U16911 ( .A1(n13762), .A2(n13761), .A3(n13760), .A4(n13759), .ZN(
        n13763) );
  AOI22_X1 U16912 ( .A1(n16810), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13768) );
  INV_X2 U16913 ( .A(n10112), .ZN(n16799) );
  AOI22_X1 U16914 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13767) );
  AOI22_X1 U16915 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13766) );
  AOI22_X1 U16916 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13765) );
  NAND4_X1 U16917 ( .A1(n13768), .A2(n13767), .A3(n13766), .A4(n13765), .ZN(
        n13774) );
  INV_X2 U16918 ( .A(n10126), .ZN(n15446) );
  AOI22_X1 U16919 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13772) );
  AOI22_X1 U16920 ( .A1(n16894), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U16921 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13770) );
  AOI22_X1 U16922 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13769) );
  NAND4_X1 U16923 ( .A1(n13772), .A2(n13771), .A3(n13770), .A4(n13769), .ZN(
        n13773) );
  AOI22_X1 U16924 ( .A1(n16810), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13778) );
  AOI22_X1 U16925 ( .A1(n9598), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13777) );
  INV_X2 U16926 ( .A(n13827), .ZN(n16871) );
  AOI22_X1 U16927 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13776) );
  AOI22_X1 U16928 ( .A1(n16894), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13775) );
  NAND4_X1 U16929 ( .A1(n13778), .A2(n13777), .A3(n13776), .A4(n13775), .ZN(
        n13784) );
  AOI22_X1 U16930 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13782) );
  BUF_X2 U16931 ( .A(n16625), .Z(n16781) );
  AOI22_X1 U16932 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13781) );
  AOI22_X1 U16933 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13780) );
  AOI22_X1 U16934 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13779) );
  NAND4_X1 U16935 ( .A1(n13782), .A2(n13781), .A3(n13780), .A4(n13779), .ZN(
        n13783) );
  AOI22_X1 U16936 ( .A1(n16888), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13794) );
  AOI22_X1 U16937 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13793) );
  AOI22_X1 U16938 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13785) );
  OAI21_X1 U16939 ( .B1(n10112), .B2(n20659), .A(n13785), .ZN(n13791) );
  AOI22_X1 U16940 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13789) );
  AOI22_X1 U16941 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U16942 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U16943 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13786) );
  NAND4_X1 U16944 ( .A1(n13789), .A2(n13788), .A3(n13787), .A4(n13786), .ZN(
        n13790) );
  AOI211_X1 U16945 ( .C1(n16635), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n13791), .B(n13790), .ZN(n13792) );
  NOR2_X1 U16946 ( .A1(n17036), .A2(n17102), .ZN(n13844) );
  AOI22_X1 U16947 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U16948 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13797) );
  AOI22_X1 U16949 ( .A1(n16894), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15468), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13796) );
  AOI22_X1 U16950 ( .A1(n16810), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16635), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13795) );
  NAND4_X1 U16951 ( .A1(n13798), .A2(n13797), .A3(n13796), .A4(n13795), .ZN(
        n13804) );
  AOI22_X1 U16952 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U16953 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13801) );
  AOI22_X1 U16954 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13800) );
  AOI22_X1 U16955 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13799) );
  NAND4_X1 U16956 ( .A1(n13802), .A2(n13801), .A3(n13800), .A4(n13799), .ZN(
        n13803) );
  AOI22_X1 U16957 ( .A1(n16810), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U16958 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13807) );
  AOI22_X1 U16959 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13806) );
  AOI22_X1 U16960 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13805) );
  AOI22_X1 U16961 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13812) );
  AOI22_X1 U16962 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13811) );
  AOI22_X1 U16963 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U16964 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13809) );
  NAND4_X1 U16965 ( .A1(n15359), .A2(n17933), .A3(n13844), .A4(n13838), .ZN(
        n18359) );
  AOI22_X1 U16966 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16810), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U16967 ( .A1(n16894), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13815) );
  AOI22_X1 U16968 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13814) );
  AOI22_X1 U16969 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13813) );
  NAND4_X1 U16970 ( .A1(n13816), .A2(n13815), .A3(n13814), .A4(n13813), .ZN(
        n13822) );
  AOI22_X1 U16971 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13820) );
  AOI22_X1 U16972 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13819) );
  AOI22_X1 U16973 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13818) );
  AOI22_X1 U16974 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13817) );
  NAND4_X1 U16975 ( .A1(n13820), .A2(n13819), .A3(n13818), .A4(n13817), .ZN(
        n13821) );
  NAND2_X1 U16976 ( .A1(n17927), .A2(n17943), .ZN(n15528) );
  NAND2_X1 U16977 ( .A1(n16953), .A2(n17938), .ZN(n18358) );
  NAND2_X1 U16978 ( .A1(n15528), .A2(n13841), .ZN(n13845) );
  INV_X2 U16979 ( .A(n10112), .ZN(n16887) );
  AOI22_X1 U16980 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U16981 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16810), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13830) );
  AOI22_X1 U16982 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13829) );
  AOI22_X1 U16983 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n16635), .B1(
        n16886), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13828) );
  NAND4_X1 U16984 ( .A1(n13831), .A2(n13830), .A3(n13829), .A4(n13828), .ZN(
        n13837) );
  AOI22_X1 U16985 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13835) );
  AOI22_X1 U16986 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13834) );
  AOI22_X1 U16987 ( .A1(n16888), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U16988 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13832) );
  NAND4_X1 U16989 ( .A1(n13835), .A2(n13834), .A3(n13833), .A4(n13832), .ZN(
        n13836) );
  OAI21_X1 U16990 ( .B1(n17036), .B2(n18379), .A(n15516), .ZN(n13851) );
  INV_X1 U16991 ( .A(n13844), .ZN(n13843) );
  NAND2_X1 U16992 ( .A1(n17916), .A2(n17922), .ZN(n15514) );
  AOI21_X1 U16993 ( .B1(n17927), .B2(n15514), .A(n13838), .ZN(n13842) );
  OAI22_X1 U16994 ( .A1(n17036), .A2(n13839), .B1(n18379), .B2(n17938), .ZN(
        n13840) );
  OAI21_X1 U16995 ( .B1(n17102), .B2(n13841), .A(n13840), .ZN(n13846) );
  AOI211_X1 U16996 ( .C1(n17933), .C2(n13843), .A(n13842), .B(n13846), .ZN(
        n13852) );
  OAI211_X1 U16997 ( .C1(n17933), .C2(n13845), .A(n13851), .B(n13852), .ZN(
        n15519) );
  NAND2_X1 U16998 ( .A1(n17927), .A2(n17933), .ZN(n18357) );
  NAND3_X1 U16999 ( .A1(n13844), .A2(n15358), .A3(n18576), .ZN(n13850) );
  NAND2_X1 U17000 ( .A1(n13848), .A2(n15362), .ZN(n17165) );
  INV_X1 U17001 ( .A(n17165), .ZN(n13849) );
  INV_X1 U17002 ( .A(n13846), .ZN(n13847) );
  NOR2_X1 U17003 ( .A1(n17927), .A2(n18359), .ZN(n13854) );
  NOR2_X1 U17004 ( .A1(n18535), .A2(n18542), .ZN(n18366) );
  AOI21_X1 U17005 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18366), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15380) );
  OR2_X1 U17006 ( .A1(n18400), .A2(n15380), .ZN(n18393) );
  NOR2_X1 U17007 ( .A1(n18530), .A2(n18393), .ZN(n13878) );
  NAND2_X1 U17008 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18426), .ZN(n18428) );
  INV_X1 U17009 ( .A(n13868), .ZN(n13853) );
  OAI211_X1 U17010 ( .C1(n13854), .C2(n13853), .A(n13852), .B(n13851), .ZN(
        n15530) );
  AOI22_X1 U17011 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18385), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18542), .ZN(n13871) );
  XNOR2_X1 U17012 ( .A(n13871), .B(n13869), .ZN(n13866) );
  AND2_X1 U17013 ( .A1(n13871), .A2(n13869), .ZN(n13855) );
  OAI21_X1 U17014 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18535), .A(
        n13856), .ZN(n13857) );
  OAI22_X1 U17015 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18399), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13857), .ZN(n13863) );
  NOR2_X1 U17016 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18399), .ZN(
        n13858) );
  NAND2_X1 U17017 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13857), .ZN(
        n13862) );
  AOI22_X1 U17018 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13863), .B1(
        n13858), .B2(n13862), .ZN(n13870) );
  NAND2_X1 U17019 ( .A1(n13861), .A2(n13860), .ZN(n13859) );
  AND2_X1 U17020 ( .A1(n13862), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13864) );
  OAI22_X1 U17021 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18395), .B1(
        n13864), .B2(n13863), .ZN(n13865) );
  INV_X1 U17022 ( .A(n13865), .ZN(n13873) );
  NAND2_X1 U17023 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18577) );
  NAND2_X1 U17024 ( .A1(n16171), .A2(n18577), .ZN(n13876) );
  INV_X1 U17025 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18449) );
  OR2_X1 U17026 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18441), .ZN(n18585) );
  NAND2_X2 U17027 ( .A1(n18584), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18513) );
  INV_X1 U17028 ( .A(n18574), .ZN(n16193) );
  NAND2_X1 U17029 ( .A1(n16193), .A2(n13867), .ZN(n17101) );
  AOI21_X1 U17030 ( .B1(n18549), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n13869), .ZN(n15521) );
  NAND3_X1 U17031 ( .A1(n13871), .A2(n13870), .A3(n15521), .ZN(n13872) );
  NAND3_X1 U17032 ( .A1(n13873), .A2(n15523), .A3(n13872), .ZN(n18562) );
  INV_X1 U17033 ( .A(n18562), .ZN(n13874) );
  AOI211_X1 U17034 ( .C1(n17165), .C2(n18400), .A(n18403), .B(n18571), .ZN(
        n13875) );
  OAI211_X1 U17035 ( .C1(n13876), .C2(n17101), .A(n15360), .B(n15635), .ZN(
        n13877) );
  INV_X1 U17036 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18425) );
  NAND2_X1 U17037 ( .A1(n18425), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17915) );
  NAND3_X1 U17038 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18518)
         );
  INV_X1 U17039 ( .A(n18518), .ZN(n18433) );
  NAND2_X1 U17040 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18433), .ZN(n15381) );
  OAI211_X1 U17041 ( .C1(n18422), .C2(n18388), .A(n17915), .B(n15381), .ZN(
        n18547) );
  INV_X1 U17042 ( .A(n18547), .ZN(n18550) );
  MUX2_X1 U17043 ( .A(n13878), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18550), .Z(P3_U3284) );
  AOI211_X1 U17044 ( .C1(n13881), .C2(n20429), .A(n20194), .B(n13880), .ZN(
        n13882) );
  AOI21_X1 U17045 ( .B1(n19922), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13882), .ZN(n13883) );
  OAI21_X1 U17046 ( .B1(n13879), .B2(n13884), .A(n13883), .ZN(P1_U3477) );
  INV_X1 U17047 ( .A(n13885), .ZN(n14307) );
  AOI22_X1 U17048 ( .A1(n13081), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13945), .ZN(n13954) );
  AND2_X1 U17049 ( .A1(n13945), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13886) );
  AOI21_X1 U17050 ( .B1(n13081), .B2(P1_EBX_REG_30__SCAN_IN), .A(n13886), .ZN(
        n13979) );
  MUX2_X1 U17051 ( .A(n13927), .B(n13977), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13888) );
  OR2_X1 U17052 ( .A1(n13081), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13887) );
  NAND2_X1 U17053 ( .A1(n13888), .A2(n13887), .ZN(n14201) );
  NOR2_X1 U17054 ( .A1(n14201), .A2(n14202), .ZN(n13889) );
  MUX2_X1 U17055 ( .A(n13937), .B(n13951), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13891) );
  NOR2_X1 U17056 ( .A1(n13081), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13890) );
  NOR2_X1 U17057 ( .A1(n13891), .A2(n13890), .ZN(n14191) );
  INV_X1 U17058 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U17059 ( .A1(n13943), .A2(n14163), .ZN(n13895) );
  INV_X1 U17060 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15723) );
  NAND2_X1 U17061 ( .A1(n13938), .A2(n15723), .ZN(n13893) );
  NAND2_X1 U17062 ( .A1(n13949), .A2(n14163), .ZN(n13892) );
  NAND3_X1 U17063 ( .A1(n13893), .A2(n13977), .A3(n13892), .ZN(n13894) );
  NAND2_X1 U17064 ( .A1(n13895), .A2(n13894), .ZN(n14192) );
  NAND2_X1 U17065 ( .A1(n14191), .A2(n14192), .ZN(n13896) );
  INV_X1 U17066 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15715) );
  NAND2_X1 U17067 ( .A1(n13938), .A2(n15715), .ZN(n13898) );
  INV_X1 U17068 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14147) );
  NAND2_X1 U17069 ( .A1(n13949), .A2(n14147), .ZN(n13897) );
  NAND3_X1 U17070 ( .A1(n13898), .A2(n13977), .A3(n13897), .ZN(n13899) );
  OAI21_X1 U17071 ( .B1(n13900), .B2(P1_EBX_REG_16__SCAN_IN), .A(n13899), .ZN(
        n14149) );
  MUX2_X1 U17072 ( .A(n13927), .B(n13977), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13901) );
  OAI21_X1 U17073 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13081), .A(
        n13901), .ZN(n14138) );
  INV_X1 U17074 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n13902) );
  NAND2_X1 U17075 ( .A1(n13943), .A2(n13902), .ZN(n13906) );
  INV_X1 U17076 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U17077 ( .A1(n13938), .A2(n14390), .ZN(n13904) );
  NAND2_X1 U17078 ( .A1(n13949), .A2(n13902), .ZN(n13903) );
  NAND3_X1 U17079 ( .A1(n13904), .A2(n13977), .A3(n13903), .ZN(n13905) );
  OR2_X2 U17080 ( .A1(n14136), .A2(n14125), .ZN(n14127) );
  INV_X1 U17081 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14184) );
  NAND2_X1 U17082 ( .A1(n13937), .A2(n14184), .ZN(n13910) );
  INV_X1 U17083 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13908) );
  NAND2_X1 U17084 ( .A1(n13949), .A2(n14184), .ZN(n13907) );
  OAI211_X1 U17085 ( .C1(n13951), .C2(n13908), .A(n13907), .B(n13938), .ZN(
        n13909) );
  NAND2_X1 U17086 ( .A1(n13910), .A2(n13909), .ZN(n14111) );
  INV_X1 U17087 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13911) );
  OAI21_X1 U17088 ( .B1(n13951), .B2(n13911), .A(n13938), .ZN(n13912) );
  OAI21_X1 U17089 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n13945), .A(n13912), .ZN(
        n13915) );
  INV_X1 U17090 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n13913) );
  NAND2_X1 U17091 ( .A1(n13943), .A2(n13913), .ZN(n13914) );
  INV_X1 U17092 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14181) );
  NAND2_X1 U17093 ( .A1(n13937), .A2(n14181), .ZN(n13918) );
  INV_X1 U17094 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14634) );
  NAND2_X1 U17095 ( .A1(n13949), .A2(n14181), .ZN(n13916) );
  OAI211_X1 U17096 ( .C1(n13951), .C2(n14634), .A(n13916), .B(n13938), .ZN(
        n13917) );
  AND2_X1 U17097 ( .A1(n13918), .A2(n13917), .ZN(n14086) );
  NAND2_X1 U17098 ( .A1(n14099), .A2(n14086), .ZN(n14088) );
  INV_X1 U17099 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n20755) );
  NAND2_X1 U17100 ( .A1(n13943), .A2(n20755), .ZN(n13922) );
  INV_X1 U17101 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13919) );
  NAND2_X1 U17102 ( .A1(n13938), .A2(n13919), .ZN(n13920) );
  OAI211_X1 U17103 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n13945), .A(n13920), .B(
        n13977), .ZN(n13921) );
  AND2_X1 U17104 ( .A1(n13922), .A2(n13921), .ZN(n14075) );
  INV_X1 U17105 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n13923) );
  NAND2_X1 U17106 ( .A1(n13937), .A2(n13923), .ZN(n13926) );
  INV_X1 U17107 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14601) );
  NAND2_X1 U17108 ( .A1(n13949), .A2(n13923), .ZN(n13924) );
  OAI211_X1 U17109 ( .C1(n13951), .C2(n14601), .A(n13924), .B(n13938), .ZN(
        n13925) );
  NAND2_X1 U17110 ( .A1(n13926), .A2(n13925), .ZN(n14065) );
  MUX2_X1 U17111 ( .A(n13927), .B(n13977), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13929) );
  OR2_X1 U17112 ( .A1(n13081), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13928) );
  NAND2_X1 U17113 ( .A1(n13929), .A2(n13928), .ZN(n14043) );
  INV_X1 U17114 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14179) );
  NAND2_X1 U17115 ( .A1(n13943), .A2(n14179), .ZN(n13932) );
  INV_X1 U17116 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14529) );
  NAND2_X1 U17117 ( .A1(n13938), .A2(n14529), .ZN(n13930) );
  OAI211_X1 U17118 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n13945), .A(n13930), .B(
        n13977), .ZN(n13931) );
  AND2_X1 U17119 ( .A1(n13932), .A2(n13931), .ZN(n14040) );
  NOR2_X1 U17120 ( .A1(n14043), .A2(n14040), .ZN(n13933) );
  INV_X1 U17121 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14584) );
  OAI21_X1 U17122 ( .B1(n13951), .B2(n14584), .A(n13938), .ZN(n13934) );
  OAI21_X1 U17123 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(n13945), .A(n13934), .ZN(
        n13936) );
  INV_X1 U17124 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14177) );
  NAND2_X1 U17125 ( .A1(n13943), .A2(n14177), .ZN(n13935) );
  AND2_X1 U17126 ( .A1(n13936), .A2(n13935), .ZN(n14015) );
  INV_X1 U17127 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14176) );
  NAND2_X1 U17128 ( .A1(n13937), .A2(n14176), .ZN(n13941) );
  INV_X1 U17129 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U17130 ( .A1(n13949), .A2(n14176), .ZN(n13939) );
  OAI211_X1 U17131 ( .C1(n13951), .C2(n14573), .A(n13939), .B(n13938), .ZN(
        n13940) );
  NAND2_X1 U17132 ( .A1(n13941), .A2(n13940), .ZN(n14016) );
  NOR2_X1 U17133 ( .A1(n14015), .A2(n14016), .ZN(n13942) );
  INV_X1 U17134 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14175) );
  NAND2_X1 U17135 ( .A1(n13943), .A2(n14175), .ZN(n13947) );
  INV_X1 U17136 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14562) );
  NAND2_X1 U17137 ( .A1(n13938), .A2(n14562), .ZN(n13944) );
  OAI211_X1 U17138 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n13945), .A(n13944), .B(
        n13977), .ZN(n13946) );
  AND2_X1 U17139 ( .A1(n13947), .A2(n13946), .ZN(n14003) );
  OR2_X1 U17140 ( .A1(n13081), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13950) );
  INV_X1 U17141 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n13948) );
  NAND2_X1 U17142 ( .A1(n13949), .A2(n13948), .ZN(n13952) );
  NAND2_X1 U17143 ( .A1(n13950), .A2(n13952), .ZN(n13976) );
  MUX2_X1 U17144 ( .A(n13976), .B(n13952), .S(n13951), .Z(n13991) );
  MUX2_X1 U17145 ( .A(n13977), .B(n13979), .S(n13993), .Z(n13953) );
  XOR2_X1 U17146 ( .A(n13954), .B(n13953), .Z(n14541) );
  NAND2_X1 U17147 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n13965) );
  INV_X1 U17148 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20568) );
  INV_X1 U17149 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20567) );
  NAND2_X1 U17150 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15650) );
  NOR3_X1 U17151 ( .A1(n20568), .A2(n20567), .A3(n15650), .ZN(n13967) );
  INV_X1 U17152 ( .A(n13967), .ZN(n13955) );
  NOR2_X1 U17153 ( .A1(n13955), .A2(n15649), .ZN(n14109) );
  AND3_X1 U17154 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14110) );
  AND3_X1 U17155 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_19__SCAN_IN), .ZN(n13956) );
  NAND3_X1 U17156 ( .A1(n14109), .A2(n14110), .A3(n13956), .ZN(n13957) );
  NAND2_X1 U17157 ( .A1(n13957), .A2(n19801), .ZN(n14102) );
  INV_X1 U17158 ( .A(n13958), .ZN(n19829) );
  NAND2_X1 U17159 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n13970) );
  INV_X1 U17160 ( .A(n13970), .ZN(n13959) );
  NAND2_X1 U17161 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n13959), .ZN(n13960) );
  NAND2_X1 U17162 ( .A1(n19829), .A2(n13960), .ZN(n13961) );
  NAND2_X1 U17163 ( .A1(n14102), .A2(n13961), .ZN(n14068) );
  AND3_X1 U17164 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_26__SCAN_IN), .ZN(n13971) );
  INV_X1 U17165 ( .A(n13971), .ZN(n13962) );
  AND2_X1 U17166 ( .A1(n19801), .A2(n13962), .ZN(n13963) );
  NOR2_X1 U17167 ( .A1(n14068), .A2(n13963), .ZN(n14029) );
  NAND2_X1 U17168 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n13996) );
  NAND2_X1 U17169 ( .A1(n19801), .A2(n13996), .ZN(n13964) );
  NAND2_X1 U17170 ( .A1(n14029), .A2(n13964), .ZN(n14008) );
  AOI21_X1 U17171 ( .B1(n19801), .B2(n13965), .A(n14008), .ZN(n13982) );
  INV_X1 U17172 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20599) );
  AOI22_X1 U17173 ( .A1(n19834), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13966) );
  OAI21_X1 U17174 ( .B1(n13982), .B2(n20599), .A(n13966), .ZN(n13973) );
  NAND2_X1 U17175 ( .A1(n15659), .A2(n13967), .ZN(n15648) );
  INV_X1 U17176 ( .A(n14110), .ZN(n13968) );
  NOR2_X2 U17177 ( .A1(n15648), .A2(n13968), .ZN(n14117) );
  AND2_X1 U17178 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n13969) );
  NAND2_X1 U17179 ( .A1(n14117), .A2(n13969), .ZN(n14103) );
  INV_X1 U17180 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20577) );
  NAND2_X1 U17182 ( .A1(n14058), .A2(n13971), .ZN(n14009) );
  INV_X1 U17183 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20595) );
  OR3_X1 U17184 ( .A1(n14009), .A2(n13996), .A3(n20595), .ZN(n13984) );
  INV_X1 U17185 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n13983) );
  NOR3_X1 U17186 ( .A1(n13984), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13983), 
        .ZN(n13972) );
  OAI21_X1 U17187 ( .B1(n14307), .B2(n19771), .A(n13974), .ZN(P1_U2809) );
  OAI22_X1 U17188 ( .A1(n13993), .A2(n13977), .B1(n13976), .B2(n9638), .ZN(
        n13978) );
  XOR2_X1 U17189 ( .A(n13979), .B(n13978), .Z(n14547) );
  INV_X1 U17190 ( .A(n14547), .ZN(n13987) );
  INV_X1 U17191 ( .A(n13980), .ZN(n14313) );
  AOI22_X1 U17192 ( .A1(n19834), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13981) );
  OAI21_X1 U17193 ( .B1(n19843), .B2(n14313), .A(n13981), .ZN(n13986) );
  AOI21_X1 U17194 ( .B1(n13984), .B2(n13983), .A(n13982), .ZN(n13985) );
  AOI211_X1 U17195 ( .C1(n13987), .C2(n19832), .A(n13986), .B(n13985), .ZN(
        n13988) );
  OAI21_X1 U17196 ( .B1(n14316), .B2(n19771), .A(n13988), .ZN(P1_U2810) );
  AOI21_X1 U17197 ( .B1(n13990), .B2(n14001), .A(n13989), .ZN(n14173) );
  NAND2_X1 U17198 ( .A1(n14173), .A2(n19796), .ZN(n14000) );
  AND2_X1 U17199 ( .A1(n9638), .A2(n13991), .ZN(n13992) );
  NOR2_X1 U17200 ( .A1(n13993), .A2(n13992), .ZN(n14557) );
  AOI22_X1 U17201 ( .A1(n19834), .A2(P1_EBX_REG_29__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13994) );
  OAI21_X1 U17202 ( .B1(n19843), .B2(n14320), .A(n13994), .ZN(n13995) );
  AOI21_X1 U17203 ( .B1(n14557), .B2(n19832), .A(n13995), .ZN(n13999) );
  NAND2_X1 U17204 ( .A1(n14008), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n13997) );
  NAND4_X1 U17205 ( .A1(n14000), .A2(n13999), .A3(n13998), .A4(n13997), .ZN(
        P1_U2811) );
  OAI21_X1 U17206 ( .B1(n9612), .B2(n14002), .A(n14001), .ZN(n14333) );
  NAND2_X1 U17207 ( .A1(n9656), .A2(n14003), .ZN(n14004) );
  NAND2_X1 U17208 ( .A1(n9638), .A2(n14004), .ZN(n14566) );
  AOI22_X1 U17209 ( .A1(n19834), .A2(P1_EBX_REG_28__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14006) );
  NAND2_X1 U17210 ( .A1(n19822), .A2(n14328), .ZN(n14005) );
  OAI211_X1 U17211 ( .C1(n14566), .C2(n19791), .A(n14006), .B(n14005), .ZN(
        n14007) );
  AOI21_X1 U17212 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14008), .A(n14007), 
        .ZN(n14012) );
  INV_X1 U17213 ( .A(n14009), .ZN(n14025) );
  INV_X1 U17214 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14010) );
  NAND3_X1 U17215 ( .A1(n14025), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14010), 
        .ZN(n14011) );
  OAI211_X1 U17216 ( .C1(n14333), .C2(n19771), .A(n14012), .B(n14011), .ZN(
        P1_U2812) );
  AOI21_X1 U17217 ( .B1(n14014), .B2(n14013), .A(n9612), .ZN(n14341) );
  INV_X1 U17218 ( .A(n14341), .ZN(n14220) );
  INV_X1 U17219 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14024) );
  INV_X1 U17220 ( .A(n14015), .ZN(n14030) );
  NAND2_X1 U17221 ( .A1(n14041), .A2(n14030), .ZN(n14017) );
  NAND2_X1 U17222 ( .A1(n14017), .A2(n14016), .ZN(n14018) );
  NAND2_X1 U17223 ( .A1(n14018), .A2(n9656), .ZN(n14570) );
  INV_X1 U17224 ( .A(n14570), .ZN(n14021) );
  AOI22_X1 U17225 ( .A1(n19834), .A2(P1_EBX_REG_27__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14019) );
  OAI21_X1 U17226 ( .B1(n19843), .B2(n14339), .A(n14019), .ZN(n14020) );
  AOI21_X1 U17227 ( .B1(n14021), .B2(n19832), .A(n14020), .ZN(n14022) );
  OAI21_X1 U17228 ( .B1(n14029), .B2(n14024), .A(n14022), .ZN(n14023) );
  AOI21_X1 U17229 ( .B1(n14025), .B2(n14024), .A(n14023), .ZN(n14026) );
  OAI21_X1 U17230 ( .B1(n14220), .B2(n19771), .A(n14026), .ZN(P1_U2813) );
  OAI21_X1 U17231 ( .B1(n14027), .B2(n14028), .A(n14013), .ZN(n14352) );
  INV_X1 U17232 ( .A(n14029), .ZN(n14034) );
  XNOR2_X1 U17233 ( .A(n14041), .B(n14030), .ZN(n14580) );
  AOI22_X1 U17234 ( .A1(n19834), .A2(P1_EBX_REG_26__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14032) );
  NAND2_X1 U17235 ( .A1(n19822), .A2(n14347), .ZN(n14031) );
  OAI211_X1 U17236 ( .C1(n14580), .C2(n19791), .A(n14032), .B(n14031), .ZN(
        n14033) );
  AOI21_X1 U17237 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n14034), .A(n14033), 
        .ZN(n14036) );
  INV_X1 U17238 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20588) );
  NAND4_X1 U17239 ( .A1(n14058), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .A4(n20588), .ZN(n14035) );
  OAI211_X1 U17240 ( .C1(n14352), .C2(n19771), .A(n14036), .B(n14035), .ZN(
        P1_U2814) );
  AOI21_X1 U17241 ( .B1(n14039), .B2(n14038), .A(n14027), .ZN(n14362) );
  INV_X1 U17242 ( .A(n14362), .ZN(n14227) );
  INV_X1 U17243 ( .A(n14040), .ZN(n14052) );
  NAND2_X1 U17244 ( .A1(n14064), .A2(n14052), .ZN(n14042) );
  AOI21_X1 U17245 ( .B1(n14043), .B2(n14042), .A(n14041), .ZN(n14593) );
  NAND2_X1 U17246 ( .A1(n14593), .A2(n19832), .ZN(n14045) );
  AOI22_X1 U17247 ( .A1(n19834), .A2(P1_EBX_REG_25__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14044) );
  OAI211_X1 U17248 ( .C1(n19843), .C2(n14360), .A(n14045), .B(n14044), .ZN(
        n14046) );
  AOI21_X1 U17249 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n14068), .A(n14046), 
        .ZN(n14049) );
  XOR2_X1 U17250 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .Z(n14047) );
  NAND2_X1 U17251 ( .A1(n14058), .A2(n14047), .ZN(n14048) );
  OAI211_X1 U17252 ( .C1(n14227), .C2(n19771), .A(n14049), .B(n14048), .ZN(
        P1_U2815) );
  OAI21_X1 U17253 ( .B1(n14050), .B2(n14051), .A(n14038), .ZN(n14367) );
  INV_X1 U17254 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20586) );
  XNOR2_X1 U17255 ( .A(n14064), .B(n14052), .ZN(n14600) );
  NAND2_X1 U17256 ( .A1(n14068), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14056) );
  OAI22_X1 U17257 ( .A1(n19782), .A2(n14053), .B1(n19790), .B2(n14179), .ZN(
        n14054) );
  AOI21_X1 U17258 ( .B1(n14368), .B2(n19822), .A(n14054), .ZN(n14055) );
  OAI211_X1 U17259 ( .C1(n14600), .C2(n19791), .A(n14056), .B(n14055), .ZN(
        n14057) );
  AOI21_X1 U17260 ( .B1(n14058), .B2(n20586), .A(n14057), .ZN(n14059) );
  OAI21_X1 U17261 ( .B1(n14367), .B2(n19771), .A(n14059), .ZN(P1_U2816) );
  AOI21_X1 U17262 ( .B1(n14062), .B2(n14061), .A(n14050), .ZN(n14063) );
  INV_X1 U17263 ( .A(n14063), .ZN(n14380) );
  AOI21_X1 U17264 ( .B1(n14065), .B2(n14077), .A(n14064), .ZN(n14611) );
  AOI22_X1 U17265 ( .A1(n19834), .A2(P1_EBX_REG_23__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14066) );
  OAI21_X1 U17266 ( .B1(n19843), .B2(n14377), .A(n14066), .ZN(n14067) );
  AOI21_X1 U17267 ( .B1(n14611), .B2(n19832), .A(n14067), .ZN(n14071) );
  OAI21_X1 U17268 ( .B1(n14069), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14068), 
        .ZN(n14070) );
  OAI211_X1 U17269 ( .C1(n14380), .C2(n19771), .A(n14071), .B(n14070), .ZN(
        P1_U2817) );
  XNOR2_X1 U17270 ( .A(P1_REIP_REG_22__SCAN_IN), .B(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14083) );
  OAI21_X1 U17271 ( .B1(n14072), .B2(n14073), .A(n14061), .ZN(n14389) );
  INV_X1 U17272 ( .A(n14389), .ZN(n14074) );
  NAND2_X1 U17273 ( .A1(n14074), .A2(n19796), .ZN(n14082) );
  INV_X1 U17274 ( .A(n14102), .ZN(n14093) );
  NAND2_X1 U17275 ( .A1(n14088), .A2(n14075), .ZN(n14076) );
  NAND2_X1 U17276 ( .A1(n14077), .A2(n14076), .ZN(n14621) );
  AOI22_X1 U17277 ( .A1(n19834), .A2(P1_EBX_REG_22__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14079) );
  NAND2_X1 U17278 ( .A1(n19822), .A2(n14384), .ZN(n14078) );
  OAI211_X1 U17279 ( .C1(n14621), .C2(n19791), .A(n14079), .B(n14078), .ZN(
        n14080) );
  AOI21_X1 U17280 ( .B1(n14093), .B2(P1_REIP_REG_22__SCAN_IN), .A(n14080), 
        .ZN(n14081) );
  OAI211_X1 U17281 ( .C1(n14096), .C2(n14083), .A(n14082), .B(n14081), .ZN(
        P1_U2818) );
  AOI21_X1 U17282 ( .B1(n14085), .B2(n14084), .A(n14072), .ZN(n14397) );
  NAND2_X1 U17283 ( .A1(n14397), .A2(n19796), .ZN(n14095) );
  OR2_X1 U17284 ( .A1(n14099), .A2(n14086), .ZN(n14087) );
  NAND2_X1 U17285 ( .A1(n14088), .A2(n14087), .ZN(n14628) );
  AOI22_X1 U17286 ( .A1(n19834), .A2(P1_EBX_REG_21__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14091) );
  INV_X1 U17287 ( .A(n14395), .ZN(n14089) );
  NAND2_X1 U17288 ( .A1(n19822), .A2(n14089), .ZN(n14090) );
  OAI211_X1 U17289 ( .C1(n14628), .C2(n19791), .A(n14091), .B(n14090), .ZN(
        n14092) );
  AOI21_X1 U17290 ( .B1(n14093), .B2(P1_REIP_REG_21__SCAN_IN), .A(n14092), 
        .ZN(n14094) );
  OAI211_X1 U17291 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n14096), .A(n14095), 
        .B(n14094), .ZN(P1_U2819) );
  OAI21_X1 U17292 ( .B1(n14097), .B2(n14098), .A(n14084), .ZN(n14401) );
  AOI21_X1 U17293 ( .B1(n14100), .B2(n14113), .A(n14099), .ZN(n14182) );
  INV_X1 U17294 ( .A(n14182), .ZN(n14638) );
  AOI22_X1 U17295 ( .A1(n19834), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14101) );
  OAI21_X1 U17296 ( .B1(n14638), .B2(n19791), .A(n14101), .ZN(n14105) );
  AOI21_X1 U17297 ( .B1(n14103), .B2(n20577), .A(n14102), .ZN(n14104) );
  AOI211_X1 U17298 ( .C1(n19822), .C2(n14402), .A(n14105), .B(n14104), .ZN(
        n14106) );
  OAI21_X1 U17299 ( .B1(n14401), .B2(n19771), .A(n14106), .ZN(P1_U2820) );
  AOI21_X1 U17300 ( .B1(n14108), .B2(n14107), .A(n14097), .ZN(n14418) );
  INV_X1 U17301 ( .A(n14418), .ZN(n14253) );
  OR2_X1 U17302 ( .A1(n14109), .A2(n19777), .ZN(n14161) );
  OAI21_X1 U17303 ( .B1(n19777), .B2(n14110), .A(n14161), .ZN(n14142) );
  NAND2_X1 U17304 ( .A1(n14127), .A2(n14111), .ZN(n14112) );
  NAND2_X1 U17305 ( .A1(n14113), .A2(n14112), .ZN(n14646) );
  OAI22_X1 U17306 ( .A1(n14646), .A2(n19791), .B1(n19782), .B2(n14114), .ZN(
        n14115) );
  AOI211_X1 U17307 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n19834), .A(n19819), .B(
        n14115), .ZN(n14116) );
  OAI21_X1 U17308 ( .B1(n14416), .B2(n19843), .A(n14116), .ZN(n14120) );
  INV_X1 U17309 ( .A(n14117), .ZN(n14131) );
  XNOR2_X1 U17310 ( .A(P1_REIP_REG_18__SCAN_IN), .B(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14118) );
  NOR2_X1 U17311 ( .A1(n14131), .A2(n14118), .ZN(n14119) );
  AOI211_X1 U17312 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(n14142), .A(n14120), 
        .B(n14119), .ZN(n14121) );
  OAI21_X1 U17313 ( .B1(n14253), .B2(n19771), .A(n14121), .ZN(P1_U2821) );
  OAI21_X1 U17314 ( .B1(n14123), .B2(n14124), .A(n14107), .ZN(n14428) );
  NAND2_X1 U17315 ( .A1(n14136), .A2(n14125), .ZN(n14126) );
  NAND2_X1 U17316 ( .A1(n14127), .A2(n14126), .ZN(n15705) );
  AOI22_X1 U17317 ( .A1(n19834), .A2(P1_EBX_REG_18__SCAN_IN), .B1(n19830), 
        .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14128) );
  OAI211_X1 U17318 ( .C1(n19791), .C2(n15705), .A(n14128), .B(n19921), .ZN(
        n14129) );
  AOI21_X1 U17319 ( .B1(n14426), .B2(n19822), .A(n14129), .ZN(n14130) );
  OAI21_X1 U17320 ( .B1(n14131), .B2(P1_REIP_REG_18__SCAN_IN), .A(n14130), 
        .ZN(n14132) );
  AOI21_X1 U17321 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n14142), .A(n14132), 
        .ZN(n14133) );
  OAI21_X1 U17322 ( .B1(n14428), .B2(n19771), .A(n14133), .ZN(P1_U2822) );
  AOI21_X1 U17323 ( .B1(n14135), .B2(n14134), .A(n14123), .ZN(n14440) );
  INV_X1 U17324 ( .A(n14440), .ZN(n14261) );
  INV_X1 U17325 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14140) );
  INV_X1 U17326 ( .A(n14136), .ZN(n14137) );
  AOI21_X1 U17327 ( .B1(n14138), .B2(n14148), .A(n14137), .ZN(n14655) );
  AOI22_X1 U17328 ( .A1(n14655), .A2(n19832), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19830), .ZN(n14139) );
  OAI211_X1 U17329 ( .C1(n19790), .C2(n14140), .A(n14139), .B(n19921), .ZN(
        n14141) );
  AOI21_X1 U17330 ( .B1(n14436), .B2(n19822), .A(n14141), .ZN(n14145) );
  NAND2_X1 U17331 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14154) );
  NOR2_X1 U17332 ( .A1(n15648), .A2(n14154), .ZN(n14143) );
  OAI21_X1 U17333 ( .B1(n14143), .B2(P1_REIP_REG_17__SCAN_IN), .A(n14142), 
        .ZN(n14144) );
  OAI211_X1 U17334 ( .C1(n14261), .C2(n19771), .A(n14145), .B(n14144), .ZN(
        P1_U2823) );
  XNOR2_X1 U17335 ( .A(n9643), .B(n14146), .ZN(n14453) );
  INV_X1 U17336 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20573) );
  INV_X1 U17337 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20571) );
  AOI21_X1 U17338 ( .B1(n20573), .B2(n20571), .A(n15648), .ZN(n14155) );
  OAI21_X1 U17339 ( .B1(n19790), .B2(n14147), .A(n19921), .ZN(n14151) );
  OAI21_X1 U17340 ( .B1(n9674), .B2(n14149), .A(n14148), .ZN(n15708) );
  OAI22_X1 U17341 ( .A1(n19782), .A2(n14442), .B1(n19791), .B2(n15708), .ZN(
        n14150) );
  AOI211_X1 U17342 ( .C1(n14451), .C2(n19822), .A(n14151), .B(n14150), .ZN(
        n14152) );
  OAI21_X1 U17343 ( .B1(n14161), .B2(n20573), .A(n14152), .ZN(n14153) );
  AOI21_X1 U17344 ( .B1(n14155), .B2(n14154), .A(n14153), .ZN(n14156) );
  OAI21_X1 U17345 ( .B1(n14453), .B2(n19771), .A(n14156), .ZN(P1_U2824) );
  OAI21_X1 U17346 ( .B1(n14157), .B2(n14159), .A(n14158), .ZN(n14468) );
  INV_X1 U17347 ( .A(n15650), .ZN(n14160) );
  NAND2_X1 U17348 ( .A1(n15659), .A2(n14160), .ZN(n15653) );
  OAI21_X1 U17349 ( .B1(n20567), .B2(n15653), .A(n20568), .ZN(n14168) );
  INV_X1 U17350 ( .A(n14161), .ZN(n15639) );
  INV_X1 U17351 ( .A(n14162), .ZN(n14470) );
  XNOR2_X1 U17352 ( .A(n14204), .B(n14192), .ZN(n15718) );
  OAI22_X1 U17353 ( .A1(n19782), .A2(n14164), .B1(n14163), .B2(n19790), .ZN(
        n14165) );
  AOI211_X1 U17354 ( .C1(n19832), .C2(n15718), .A(n19819), .B(n14165), .ZN(
        n14166) );
  OAI21_X1 U17355 ( .B1(n14470), .B2(n19843), .A(n14166), .ZN(n14167) );
  AOI21_X1 U17356 ( .B1(n14168), .B2(n15639), .A(n14167), .ZN(n14169) );
  OAI21_X1 U17357 ( .B1(n14468), .B2(n19771), .A(n14169), .ZN(P1_U2826) );
  INV_X1 U17358 ( .A(n14541), .ZN(n14171) );
  INV_X1 U17359 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14170) );
  OAI22_X1 U17360 ( .A1(n14171), .A2(n14206), .B1(n19850), .B2(n14170), .ZN(
        P1_U2841) );
  INV_X1 U17361 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14172) );
  OAI222_X1 U17362 ( .A1(n14206), .A2(n14547), .B1(n14172), .B2(n19850), .C1(
        n14316), .C2(n14208), .ZN(P1_U2842) );
  INV_X1 U17363 ( .A(n14173), .ZN(n14323) );
  AOI22_X1 U17364 ( .A1(n14557), .A2(n19845), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14197), .ZN(n14174) );
  OAI21_X1 U17365 ( .B1(n14323), .B2(n14196), .A(n14174), .ZN(P1_U2843) );
  OAI222_X1 U17366 ( .A1(n14566), .A2(n14206), .B1(n14175), .B2(n19850), .C1(
        n14333), .C2(n14208), .ZN(P1_U2844) );
  OAI222_X1 U17367 ( .A1(n14220), .A2(n14208), .B1(n14176), .B2(n19850), .C1(
        n14570), .C2(n14206), .ZN(P1_U2845) );
  OAI222_X1 U17368 ( .A1(n14208), .A2(n14352), .B1(n14177), .B2(n19850), .C1(
        n14206), .C2(n14580), .ZN(P1_U2846) );
  AOI22_X1 U17369 ( .A1(n14593), .A2(n19845), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14197), .ZN(n14178) );
  OAI21_X1 U17370 ( .B1(n14227), .B2(n14196), .A(n14178), .ZN(P1_U2847) );
  OAI222_X1 U17371 ( .A1(n14367), .A2(n14208), .B1(n14179), .B2(n19850), .C1(
        n14206), .C2(n14600), .ZN(P1_U2848) );
  AOI22_X1 U17372 ( .A1(n14611), .A2(n19845), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14197), .ZN(n14180) );
  OAI21_X1 U17373 ( .B1(n14380), .B2(n14208), .A(n14180), .ZN(P1_U2849) );
  OAI222_X1 U17374 ( .A1(n14621), .A2(n14206), .B1(n20755), .B2(n19850), .C1(
        n14389), .C2(n14208), .ZN(P1_U2850) );
  INV_X1 U17375 ( .A(n14397), .ZN(n14244) );
  OAI222_X1 U17376 ( .A1(n14244), .A2(n14196), .B1(n14181), .B2(n19850), .C1(
        n14628), .C2(n14206), .ZN(P1_U2851) );
  AOI22_X1 U17377 ( .A1(n14182), .A2(n19845), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n14197), .ZN(n14183) );
  OAI21_X1 U17378 ( .B1(n14401), .B2(n14208), .A(n14183), .ZN(P1_U2852) );
  OAI222_X1 U17379 ( .A1(n14253), .A2(n14196), .B1(n14184), .B2(n19850), .C1(
        n14646), .C2(n14206), .ZN(P1_U2853) );
  INV_X1 U17380 ( .A(n15705), .ZN(n14185) );
  AOI22_X1 U17381 ( .A1(n14185), .A2(n19845), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n14197), .ZN(n14186) );
  OAI21_X1 U17382 ( .B1(n14428), .B2(n14196), .A(n14186), .ZN(P1_U2854) );
  AOI22_X1 U17383 ( .A1(n14655), .A2(n19845), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14197), .ZN(n14187) );
  OAI21_X1 U17384 ( .B1(n14261), .B2(n14208), .A(n14187), .ZN(P1_U2855) );
  INV_X1 U17385 ( .A(n15708), .ZN(n14188) );
  AOI22_X1 U17386 ( .A1(n19845), .A2(n14188), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14197), .ZN(n14189) );
  OAI21_X1 U17387 ( .B1(n14453), .B2(n14208), .A(n14189), .ZN(P1_U2856) );
  AOI21_X1 U17388 ( .B1(n14190), .B2(n14158), .A(n9643), .ZN(n15645) );
  INV_X1 U17389 ( .A(n15645), .ZN(n14273) );
  INV_X1 U17390 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14195) );
  INV_X1 U17391 ( .A(n14204), .ZN(n14193) );
  AOI21_X1 U17392 ( .B1(n14193), .B2(n14192), .A(n14191), .ZN(n14194) );
  OR2_X1 U17393 ( .A1(n14194), .A2(n9674), .ZN(n14666) );
  OAI222_X1 U17394 ( .A1(n14273), .A2(n14196), .B1(n14195), .B2(n19850), .C1(
        n14666), .C2(n14206), .ZN(P1_U2857) );
  AOI22_X1 U17395 ( .A1(n19845), .A2(n15718), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14197), .ZN(n14198) );
  OAI21_X1 U17396 ( .B1(n14468), .B2(n14208), .A(n14198), .ZN(P1_U2858) );
  AOI21_X1 U17397 ( .B1(n14199), .B2(n13734), .A(n14157), .ZN(n14480) );
  INV_X1 U17398 ( .A(n14480), .ZN(n15654) );
  INV_X1 U17399 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14207) );
  INV_X1 U17400 ( .A(n14200), .ZN(n14203) );
  OAI21_X1 U17401 ( .B1(n14203), .B2(n14202), .A(n14201), .ZN(n14205) );
  NAND2_X1 U17402 ( .A1(n14205), .A2(n14204), .ZN(n14683) );
  OAI222_X1 U17403 ( .A1(n15654), .A2(n14208), .B1(n14207), .B2(n19850), .C1(
        n14683), .C2(n14206), .ZN(P1_U2859) );
  AOI22_X1 U17404 ( .A1(n14257), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14275), .ZN(n14211) );
  NOR3_X4 U17405 ( .A1(n14275), .A2(n14209), .A3(n11421), .ZN(n14264) );
  MUX2_X1 U17406 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n19925), .Z(
        n19891) );
  AOI22_X1 U17407 ( .A1(n14264), .A2(n19891), .B1(n14268), .B2(DATAI_30_), 
        .ZN(n14210) );
  OAI211_X1 U17408 ( .C1(n14316), .C2(n14279), .A(n14211), .B(n14210), .ZN(
        P1_U2874) );
  AOI22_X1 U17409 ( .A1(n14257), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14275), .ZN(n14213) );
  AOI22_X1 U17410 ( .A1(n14264), .A2(n14276), .B1(n14268), .B2(DATAI_29_), 
        .ZN(n14212) );
  OAI211_X1 U17411 ( .C1(n14323), .C2(n14279), .A(n14213), .B(n14212), .ZN(
        P1_U2875) );
  AOI22_X1 U17412 ( .A1(n14257), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14275), .ZN(n14215) );
  AOI22_X1 U17413 ( .A1(n14264), .A2(n19889), .B1(n14268), .B2(DATAI_28_), 
        .ZN(n14214) );
  OAI211_X1 U17414 ( .C1(n14333), .C2(n14279), .A(n14215), .B(n14214), .ZN(
        P1_U2876) );
  INV_X1 U17415 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19014) );
  OAI22_X1 U17416 ( .A1(n14263), .A2(n19014), .B1(n12811), .B2(n14270), .ZN(
        n14216) );
  INV_X1 U17417 ( .A(n14216), .ZN(n14219) );
  AOI22_X1 U17418 ( .A1(n14264), .A2(n14217), .B1(n14268), .B2(DATAI_27_), 
        .ZN(n14218) );
  OAI211_X1 U17419 ( .C1(n14220), .C2(n14279), .A(n14219), .B(n14218), .ZN(
        P1_U2877) );
  AOI22_X1 U17420 ( .A1(n14257), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14275), .ZN(n14223) );
  AOI22_X1 U17421 ( .A1(n14264), .A2(n14221), .B1(n14268), .B2(DATAI_26_), 
        .ZN(n14222) );
  OAI211_X1 U17422 ( .C1(n14352), .C2(n14279), .A(n14223), .B(n14222), .ZN(
        P1_U2878) );
  AOI22_X1 U17423 ( .A1(n14257), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14275), .ZN(n14226) );
  AOI22_X1 U17424 ( .A1(n14264), .A2(n14224), .B1(n14268), .B2(DATAI_25_), 
        .ZN(n14225) );
  OAI211_X1 U17425 ( .C1(n14227), .C2(n14279), .A(n14226), .B(n14225), .ZN(
        P1_U2879) );
  AOI22_X1 U17426 ( .A1(n14257), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14275), .ZN(n14229) );
  AOI22_X1 U17427 ( .A1(n14264), .A2(n19887), .B1(n14268), .B2(DATAI_24_), 
        .ZN(n14228) );
  OAI211_X1 U17428 ( .C1(n14367), .C2(n14279), .A(n14229), .B(n14228), .ZN(
        P1_U2880) );
  INV_X1 U17429 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n19040) );
  OAI22_X1 U17430 ( .A1(n14263), .A2(n19040), .B1(n14230), .B2(n14270), .ZN(
        n14231) );
  INV_X1 U17431 ( .A(n14231), .ZN(n14233) );
  AOI22_X1 U17432 ( .A1(n14264), .A2(n19977), .B1(n14268), .B2(DATAI_23_), 
        .ZN(n14232) );
  OAI211_X1 U17433 ( .C1(n14380), .C2(n14279), .A(n14233), .B(n14232), .ZN(
        P1_U2881) );
  INV_X1 U17434 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14234) );
  OAI22_X1 U17435 ( .A1(n14263), .A2(n14234), .B1(n12807), .B2(n14270), .ZN(
        n14235) );
  INV_X1 U17436 ( .A(n14235), .ZN(n14238) );
  AOI22_X1 U17437 ( .A1(n14264), .A2(n14236), .B1(n14268), .B2(DATAI_22_), 
        .ZN(n14237) );
  OAI211_X1 U17438 ( .C1(n14389), .C2(n14279), .A(n14238), .B(n14237), .ZN(
        P1_U2882) );
  INV_X1 U17439 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14851) );
  OAI22_X1 U17440 ( .A1(n14263), .A2(n14851), .B1(n14239), .B2(n14270), .ZN(
        n14240) );
  INV_X1 U17441 ( .A(n14240), .ZN(n14243) );
  AOI22_X1 U17442 ( .A1(n14264), .A2(n14241), .B1(n14268), .B2(DATAI_21_), 
        .ZN(n14242) );
  OAI211_X1 U17443 ( .C1(n14244), .C2(n14279), .A(n14243), .B(n14242), .ZN(
        P1_U2883) );
  AOI22_X1 U17444 ( .A1(n14257), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14275), .ZN(n14247) );
  AOI22_X1 U17445 ( .A1(n14264), .A2(n14245), .B1(n14268), .B2(DATAI_20_), 
        .ZN(n14246) );
  OAI211_X1 U17446 ( .C1(n14401), .C2(n14279), .A(n14247), .B(n14246), .ZN(
        P1_U2884) );
  INV_X1 U17447 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16103) );
  OAI22_X1 U17448 ( .A1(n14263), .A2(n16103), .B1(n14248), .B2(n14270), .ZN(
        n14249) );
  INV_X1 U17449 ( .A(n14249), .ZN(n14252) );
  AOI22_X1 U17450 ( .A1(n14264), .A2(n14250), .B1(n14268), .B2(DATAI_19_), 
        .ZN(n14251) );
  OAI211_X1 U17451 ( .C1(n14253), .C2(n14279), .A(n14252), .B(n14251), .ZN(
        P1_U2885) );
  AOI22_X1 U17452 ( .A1(n14257), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14275), .ZN(n14256) );
  AOI22_X1 U17453 ( .A1(n14264), .A2(n14254), .B1(n14268), .B2(DATAI_18_), 
        .ZN(n14255) );
  OAI211_X1 U17454 ( .C1(n14428), .C2(n14279), .A(n14256), .B(n14255), .ZN(
        P1_U2886) );
  AOI22_X1 U17455 ( .A1(n14257), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14275), .ZN(n14260) );
  AOI22_X1 U17456 ( .A1(n14264), .A2(n14258), .B1(n14268), .B2(DATAI_17_), 
        .ZN(n14259) );
  OAI211_X1 U17457 ( .C1(n14261), .C2(n14279), .A(n14260), .B(n14259), .ZN(
        P1_U2887) );
  INV_X1 U17458 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14262) );
  OAI22_X1 U17459 ( .A1(n14263), .A2(n14262), .B1(n12819), .B2(n14270), .ZN(
        n14267) );
  INV_X1 U17460 ( .A(n14264), .ZN(n14265) );
  NOR2_X1 U17461 ( .A1(n14265), .A2(n19938), .ZN(n14266) );
  AOI211_X1 U17462 ( .C1(n14268), .C2(DATAI_16_), .A(n14267), .B(n14266), .ZN(
        n14269) );
  OAI21_X1 U17463 ( .B1(n14453), .B2(n14279), .A(n14269), .ZN(P1_U2888) );
  OAI222_X1 U17464 ( .A1(n14273), .A2(n14279), .B1(n14272), .B2(n14271), .C1(
        n14270), .C2(n19854), .ZN(P1_U2889) );
  AOI22_X1 U17465 ( .A1(n14277), .A2(n19891), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14275), .ZN(n14274) );
  OAI21_X1 U17466 ( .B1(n14468), .B2(n14279), .A(n14274), .ZN(P1_U2890) );
  AOI22_X1 U17467 ( .A1(n14277), .A2(n14276), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14275), .ZN(n14278) );
  OAI21_X1 U17468 ( .B1(n15654), .B2(n14279), .A(n14278), .ZN(P1_U2891) );
  OR2_X1 U17469 ( .A1(n13658), .A2(n14282), .ZN(n14280) );
  NAND2_X1 U17470 ( .A1(n9593), .A2(n14282), .ZN(n14283) );
  XNOR2_X1 U17471 ( .A(n13658), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14476) );
  NAND2_X1 U17472 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14284) );
  NAND2_X1 U17473 ( .A1(n13658), .A2(n14284), .ZN(n14482) );
  NAND2_X1 U17474 ( .A1(n14476), .A2(n14482), .ZN(n14464) );
  NAND2_X1 U17475 ( .A1(n13658), .A2(n15729), .ZN(n14485) );
  NAND2_X1 U17476 ( .A1(n13658), .A2(n15723), .ZN(n14285) );
  NAND2_X1 U17477 ( .A1(n14485), .A2(n14285), .ZN(n14286) );
  INV_X1 U17478 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14668) );
  NOR2_X1 U17479 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14287) );
  OR2_X1 U17480 ( .A1(n13658), .A2(n14287), .ZN(n14289) );
  AND2_X1 U17481 ( .A1(n14454), .A2(n14289), .ZN(n14430) );
  XNOR2_X1 U17482 ( .A(n13658), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14447) );
  NAND2_X1 U17483 ( .A1(n13658), .A2(n14668), .ZN(n14457) );
  NOR2_X1 U17484 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14483) );
  AND2_X1 U17485 ( .A1(n14483), .A2(n15729), .ZN(n14288) );
  OR2_X1 U17486 ( .A1(n13658), .A2(n14288), .ZN(n14429) );
  AND2_X1 U17487 ( .A1(n14289), .A2(n14429), .ZN(n14443) );
  NOR2_X1 U17488 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14290) );
  XNOR2_X1 U17489 ( .A(n9593), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14422) );
  AND2_X1 U17490 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14642) );
  NAND2_X1 U17491 ( .A1(n14642), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14291) );
  NOR2_X1 U17492 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14641) );
  NAND3_X1 U17493 ( .A1(n14641), .A2(n14634), .A3(n14390), .ZN(n14292) );
  INV_X1 U17494 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14357) );
  NAND2_X1 U17495 ( .A1(n14601), .A2(n14357), .ZN(n14324) );
  NAND2_X1 U17496 ( .A1(n14293), .A2(n9593), .ZN(n14354) );
  NAND2_X1 U17497 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14294) );
  NAND3_X1 U17498 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14585) );
  AND2_X1 U17499 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14528) );
  NAND2_X1 U17500 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14297) );
  NOR2_X1 U17501 ( .A1(n14297), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14502) );
  AOI22_X1 U17502 ( .A1(n14492), .A2(n14295), .B1(n14318), .B2(n14502), .ZN(
        n14301) );
  NOR2_X1 U17503 ( .A1(n9593), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14300) );
  NAND2_X1 U17504 ( .A1(n14296), .A2(n14300), .ZN(n14299) );
  OAI211_X1 U17505 ( .C1(n14308), .C2(n14297), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n9593), .ZN(n14298) );
  OAI211_X1 U17506 ( .C1(n14301), .C2(n14300), .A(n14299), .B(n14298), .ZN(
        n14501) );
  INV_X1 U17507 ( .A(n14302), .ZN(n14304) );
  NAND2_X1 U17508 ( .A1(n15772), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14537) );
  NAND2_X1 U17509 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14303) );
  OAI211_X1 U17510 ( .C1(n14304), .C2(n15696), .A(n14537), .B(n14303), .ZN(
        n14305) );
  AOI21_X1 U17511 ( .B1(n14501), .B2(n15692), .A(n14305), .ZN(n14306) );
  OAI21_X1 U17512 ( .B1(n14307), .B2(n19924), .A(n14306), .ZN(P1_U2968) );
  NAND2_X1 U17513 ( .A1(n14309), .A2(n9900), .ZN(n14310) );
  NAND2_X1 U17514 ( .A1(n15772), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14546) );
  NAND2_X1 U17515 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14312) );
  OAI211_X1 U17516 ( .C1(n14313), .C2(n15696), .A(n14546), .B(n14312), .ZN(
        n14314) );
  AOI21_X1 U17517 ( .B1(n14544), .B2(n15692), .A(n14314), .ZN(n14315) );
  XNOR2_X1 U17518 ( .A(n9593), .B(n9900), .ZN(n14317) );
  XNOR2_X1 U17519 ( .A(n14318), .B(n14317), .ZN(n14553) );
  NOR2_X1 U17520 ( .A1(n19921), .A2(n20595), .ZN(n14556) );
  AOI21_X1 U17521 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14556), .ZN(n14319) );
  OAI21_X1 U17522 ( .B1(n15696), .B2(n14320), .A(n14319), .ZN(n14321) );
  AOI21_X1 U17523 ( .B1(n14553), .B2(n15692), .A(n14321), .ZN(n14322) );
  OAI21_X1 U17524 ( .B1(n14323), .B2(n19924), .A(n14322), .ZN(P1_U2970) );
  NOR2_X1 U17525 ( .A1(n9954), .A2(n9899), .ZN(n14344) );
  NOR2_X1 U17526 ( .A1(n14353), .A2(n14344), .ZN(n14327) );
  MUX2_X1 U17527 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14584), .S(
        n9593), .Z(n14326) );
  NOR3_X1 U17528 ( .A1(n14324), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14325) );
  NAND2_X1 U17529 ( .A1(n15681), .A2(n14328), .ZN(n14329) );
  NAND2_X1 U17530 ( .A1(n15772), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14565) );
  OAI211_X1 U17531 ( .C1(n14459), .C2(n14330), .A(n14329), .B(n14565), .ZN(
        n14331) );
  OAI21_X1 U17532 ( .B1(n14333), .B2(n19924), .A(n14332), .ZN(P1_U2971) );
  INV_X1 U17533 ( .A(n14334), .ZN(n14335) );
  MUX2_X1 U17534 ( .A(n14336), .B(n14335), .S(n14492), .Z(n14337) );
  XNOR2_X1 U17535 ( .A(n14337), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14578) );
  AND2_X1 U17536 ( .A1(n15772), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14572) );
  AOI21_X1 U17537 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14572), .ZN(n14338) );
  OAI21_X1 U17538 ( .B1(n15696), .B2(n14339), .A(n14338), .ZN(n14340) );
  AOI21_X1 U17539 ( .B1(n14341), .B2(n15693), .A(n14340), .ZN(n14342) );
  OAI21_X1 U17540 ( .B1(n19748), .B2(n14578), .A(n14342), .ZN(P1_U2972) );
  AOI21_X1 U17541 ( .B1(n9593), .B2(n14375), .A(n14343), .ZN(n14345) );
  NOR2_X1 U17542 ( .A1(n14345), .A2(n14344), .ZN(n14346) );
  XOR2_X1 U17543 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14346), .Z(
        n14579) );
  INV_X1 U17544 ( .A(n14347), .ZN(n14349) );
  NOR2_X1 U17545 ( .A1(n19921), .A2(n20588), .ZN(n14581) );
  AOI21_X1 U17546 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14581), .ZN(n14348) );
  OAI21_X1 U17547 ( .B1(n15696), .B2(n14349), .A(n14348), .ZN(n14350) );
  AOI21_X1 U17548 ( .B1(n14579), .B2(n15692), .A(n14350), .ZN(n14351) );
  OAI21_X1 U17549 ( .B1(n14352), .B2(n19924), .A(n14351), .ZN(P1_U2973) );
  NAND3_X1 U17550 ( .A1(n14353), .A2(n14601), .A3(n14529), .ZN(n14356) );
  AND2_X1 U17551 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14365) );
  NAND2_X1 U17552 ( .A1(n14365), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14355) );
  MUX2_X1 U17553 ( .A(n14356), .B(n14355), .S(n9593), .Z(n14358) );
  XNOR2_X1 U17554 ( .A(n14358), .B(n14357), .ZN(n14599) );
  AND2_X1 U17555 ( .A1(n15772), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14592) );
  AOI21_X1 U17556 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14592), .ZN(n14359) );
  OAI21_X1 U17557 ( .B1(n15696), .B2(n14360), .A(n14359), .ZN(n14361) );
  AOI21_X1 U17558 ( .B1(n14362), .B2(n15693), .A(n14361), .ZN(n14363) );
  OAI21_X1 U17559 ( .B1(n19748), .B2(n14599), .A(n14363), .ZN(P1_U2974) );
  NOR2_X1 U17560 ( .A1(n14365), .A2(n14375), .ZN(n14364) );
  MUX2_X1 U17561 ( .A(n14365), .B(n14364), .S(n14492), .Z(n14366) );
  XNOR2_X1 U17562 ( .A(n14366), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14609) );
  INV_X1 U17563 ( .A(n14367), .ZN(n14372) );
  INV_X1 U17564 ( .A(n14368), .ZN(n14370) );
  AND2_X1 U17565 ( .A1(n15772), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14603) );
  AOI21_X1 U17566 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14603), .ZN(n14369) );
  OAI21_X1 U17567 ( .B1(n15696), .B2(n14370), .A(n14369), .ZN(n14371) );
  AOI21_X1 U17568 ( .B1(n14372), .B2(n15693), .A(n14371), .ZN(n14373) );
  OAI21_X1 U17569 ( .B1(n19748), .B2(n14609), .A(n14373), .ZN(P1_U2975) );
  XNOR2_X1 U17570 ( .A(n9593), .B(n14601), .ZN(n14374) );
  XNOR2_X1 U17571 ( .A(n14375), .B(n14374), .ZN(n14610) );
  INV_X1 U17572 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20583) );
  NOR2_X1 U17573 ( .A1(n19921), .A2(n20583), .ZN(n14614) );
  AOI21_X1 U17574 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n14614), .ZN(n14376) );
  OAI21_X1 U17575 ( .B1(n15696), .B2(n14377), .A(n14376), .ZN(n14378) );
  AOI21_X1 U17576 ( .B1(n14610), .B2(n15692), .A(n14378), .ZN(n14379) );
  OAI21_X1 U17577 ( .B1(n14380), .B2(n19924), .A(n14379), .ZN(P1_U2976) );
  NAND2_X1 U17578 ( .A1(n14382), .A2(n14381), .ZN(n14383) );
  XNOR2_X1 U17579 ( .A(n14383), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14619) );
  NAND2_X1 U17580 ( .A1(n15681), .A2(n14384), .ZN(n14385) );
  NAND2_X1 U17581 ( .A1(n15772), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14620) );
  OAI211_X1 U17582 ( .C1(n14459), .C2(n14386), .A(n14385), .B(n14620), .ZN(
        n14387) );
  AOI21_X1 U17583 ( .B1(n14619), .B2(n15692), .A(n14387), .ZN(n14388) );
  OAI21_X1 U17584 ( .B1(n14389), .B2(n19924), .A(n14388), .ZN(P1_U2977) );
  NOR2_X1 U17585 ( .A1(n9593), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14408) );
  OR2_X1 U17586 ( .A1(n9593), .A2(n14390), .ZN(n14391) );
  NAND2_X1 U17587 ( .A1(n14421), .A2(n14391), .ZN(n14410) );
  OAI22_X1 U17588 ( .A1(n14410), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n14492), .B2(n14421), .ZN(n14392) );
  OAI21_X1 U17589 ( .B1(n14642), .B2(n14408), .A(n14392), .ZN(n14393) );
  XNOR2_X1 U17590 ( .A(n14393), .B(n14634), .ZN(n14637) );
  AND2_X1 U17591 ( .A1(n15772), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14629) );
  AOI21_X1 U17592 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n14629), .ZN(n14394) );
  OAI21_X1 U17593 ( .B1(n15696), .B2(n14395), .A(n14394), .ZN(n14396) );
  AOI21_X1 U17594 ( .B1(n14397), .B2(n15693), .A(n14396), .ZN(n14398) );
  OAI21_X1 U17595 ( .B1(n19748), .B2(n14637), .A(n14398), .ZN(P1_U2978) );
  NAND2_X1 U17596 ( .A1(n9593), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14412) );
  INV_X1 U17597 ( .A(n14410), .ZN(n14399) );
  NAND2_X1 U17598 ( .A1(n14399), .A2(n14408), .ZN(n14413) );
  OAI21_X1 U17599 ( .B1(n14421), .B2(n14412), .A(n14413), .ZN(n14400) );
  XNOR2_X1 U17600 ( .A(n14400), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14645) );
  INV_X1 U17601 ( .A(n14401), .ZN(n14406) );
  INV_X1 U17602 ( .A(n14402), .ZN(n14404) );
  AND2_X1 U17603 ( .A1(n15772), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14640) );
  AOI21_X1 U17604 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14640), .ZN(n14403) );
  OAI21_X1 U17605 ( .B1(n15696), .B2(n14404), .A(n14403), .ZN(n14405) );
  AOI21_X1 U17606 ( .B1(n14406), .B2(n15693), .A(n14405), .ZN(n14407) );
  OAI21_X1 U17607 ( .B1(n14645), .B2(n19748), .A(n14407), .ZN(P1_U2979) );
  INV_X1 U17608 ( .A(n14408), .ZN(n14409) );
  NAND2_X1 U17609 ( .A1(n14409), .A2(n14412), .ZN(n14411) );
  MUX2_X1 U17610 ( .A(n14412), .B(n14411), .S(n14410), .Z(n14414) );
  AND2_X1 U17611 ( .A1(n15772), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14648) );
  AOI21_X1 U17612 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n14648), .ZN(n14415) );
  OAI21_X1 U17613 ( .B1(n15696), .B2(n14416), .A(n14415), .ZN(n14417) );
  AOI21_X1 U17614 ( .B1(n14418), .B2(n15693), .A(n14417), .ZN(n14419) );
  OAI21_X1 U17615 ( .B1(n14653), .B2(n19748), .A(n14419), .ZN(P1_U2980) );
  INV_X1 U17616 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14420) );
  OAI22_X1 U17617 ( .A1(n14459), .A2(n20756), .B1(n14420), .B2(n19921), .ZN(
        n14425) );
  OAI21_X1 U17618 ( .B1(n14423), .B2(n14422), .A(n14421), .ZN(n15700) );
  NOR2_X1 U17619 ( .A1(n15700), .A2(n19748), .ZN(n14424) );
  AOI211_X1 U17620 ( .C1(n15681), .C2(n14426), .A(n14425), .B(n14424), .ZN(
        n14427) );
  OAI21_X1 U17621 ( .B1(n14428), .B2(n19924), .A(n14427), .ZN(P1_U2981) );
  NOR2_X1 U17622 ( .A1(n9593), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14434) );
  NAND2_X1 U17623 ( .A1(n14688), .A2(n14429), .ZN(n14474) );
  INV_X1 U17624 ( .A(n14430), .ZN(n14432) );
  OAI21_X1 U17625 ( .B1(n14474), .B2(n14432), .A(n14431), .ZN(n14433) );
  MUX2_X1 U17626 ( .A(n9593), .B(n14434), .S(n14433), .Z(n14435) );
  XNOR2_X1 U17627 ( .A(n14435), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14665) );
  INV_X1 U17628 ( .A(n14436), .ZN(n14438) );
  AND2_X1 U17629 ( .A1(n15772), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n14654) );
  AOI21_X1 U17630 ( .B1(n15686), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n14654), .ZN(n14437) );
  OAI21_X1 U17631 ( .B1(n15696), .B2(n14438), .A(n14437), .ZN(n14439) );
  AOI21_X1 U17632 ( .B1(n14440), .B2(n15693), .A(n14439), .ZN(n14441) );
  OAI21_X1 U17633 ( .B1(n14665), .B2(n19748), .A(n14441), .ZN(P1_U2982) );
  OAI22_X1 U17634 ( .A1(n14459), .A2(n14442), .B1(n20573), .B2(n19921), .ZN(
        n14450) );
  OAI21_X1 U17635 ( .B1(n14688), .B2(n14444), .A(n14443), .ZN(n14456) );
  INV_X1 U17636 ( .A(n14454), .ZN(n14445) );
  NOR2_X1 U17637 ( .A1(n14456), .A2(n14445), .ZN(n14458) );
  NOR2_X1 U17638 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15707) );
  NOR2_X1 U17639 ( .A1(n14458), .A2(n15707), .ZN(n14448) );
  OAI22_X1 U17640 ( .A1(n14448), .A2(n14447), .B1(n14458), .B2(n14446), .ZN(
        n15709) );
  NOR2_X1 U17641 ( .A1(n15709), .A2(n19748), .ZN(n14449) );
  AOI211_X1 U17642 ( .C1(n15681), .C2(n14451), .A(n14450), .B(n14449), .ZN(
        n14452) );
  OAI21_X1 U17643 ( .B1(n19924), .B2(n14453), .A(n14452), .ZN(P1_U2983) );
  NAND2_X1 U17644 ( .A1(n14454), .A2(n14457), .ZN(n14455) );
  AOI22_X1 U17645 ( .A1(n14458), .A2(n14457), .B1(n14456), .B2(n14455), .ZN(
        n14671) );
  NAND2_X1 U17646 ( .A1(n15645), .A2(n15693), .ZN(n14462) );
  OAI22_X1 U17647 ( .A1(n14459), .A2(n15643), .B1(n20571), .B2(n19921), .ZN(
        n14460) );
  AOI21_X1 U17648 ( .B1(n15681), .B2(n15640), .A(n14460), .ZN(n14461) );
  OAI211_X1 U17649 ( .C1(n14671), .C2(n19748), .A(n14462), .B(n14461), .ZN(
        P1_U2984) );
  INV_X1 U17650 ( .A(n14485), .ZN(n14463) );
  NOR2_X1 U17651 ( .A1(n14464), .A2(n14463), .ZN(n14465) );
  AOI22_X1 U17652 ( .A1(n14474), .A2(n14465), .B1(n9954), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14467) );
  XNOR2_X1 U17653 ( .A(n9593), .B(n15723), .ZN(n14466) );
  XNOR2_X1 U17654 ( .A(n14467), .B(n14466), .ZN(n15717) );
  INV_X1 U17655 ( .A(n14468), .ZN(n14472) );
  AOI22_X1 U17656 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14469) );
  OAI21_X1 U17657 ( .B1(n15696), .B2(n14470), .A(n14469), .ZN(n14471) );
  AOI21_X1 U17658 ( .B1(n14472), .B2(n15693), .A(n14471), .ZN(n14473) );
  OAI21_X1 U17659 ( .B1(n15717), .B2(n19748), .A(n14473), .ZN(P1_U2985) );
  NAND3_X1 U17660 ( .A1(n14474), .A2(n14482), .A3(n14485), .ZN(n14475) );
  XOR2_X1 U17661 ( .A(n14476), .B(n14475), .Z(n14686) );
  INV_X1 U17662 ( .A(n15657), .ZN(n14478) );
  AOI22_X1 U17663 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14477) );
  OAI21_X1 U17664 ( .B1(n15696), .B2(n14478), .A(n14477), .ZN(n14479) );
  AOI21_X1 U17665 ( .B1(n14480), .B2(n15693), .A(n14479), .ZN(n14481) );
  OAI21_X1 U17666 ( .B1(n19748), .B2(n14686), .A(n14481), .ZN(P1_U2986) );
  INV_X1 U17667 ( .A(n14482), .ZN(n14484) );
  OAI22_X1 U17668 ( .A1(n14688), .A2(n14484), .B1(n14483), .B2(n9593), .ZN(
        n14487) );
  OAI21_X1 U17669 ( .B1(n9593), .B2(n15729), .A(n14485), .ZN(n14486) );
  XNOR2_X1 U17670 ( .A(n14487), .B(n14486), .ZN(n15741) );
  INV_X1 U17671 ( .A(n15741), .ZN(n14491) );
  AOI22_X1 U17672 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n14488) );
  OAI21_X1 U17673 ( .B1(n15696), .B2(n15663), .A(n14488), .ZN(n14489) );
  AOI21_X1 U17674 ( .B1(n15665), .B2(n15693), .A(n14489), .ZN(n14490) );
  OAI21_X1 U17675 ( .B1(n14491), .B2(n19748), .A(n14490), .ZN(P1_U2987) );
  NOR3_X1 U17676 ( .A1(n14688), .A2(n9954), .A3(n13590), .ZN(n14691) );
  NOR3_X1 U17677 ( .A1(n14687), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n9593), .ZN(n14493) );
  NOR2_X1 U17678 ( .A1(n14691), .A2(n14493), .ZN(n14494) );
  XNOR2_X1 U17679 ( .A(n14494), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15750) );
  INV_X1 U17680 ( .A(n15750), .ZN(n14500) );
  AOI22_X1 U17681 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n14495) );
  OAI21_X1 U17682 ( .B1(n15696), .B2(n14496), .A(n14495), .ZN(n14497) );
  AOI21_X1 U17683 ( .B1(n14498), .B2(n15693), .A(n14497), .ZN(n14499) );
  OAI21_X1 U17684 ( .B1(n14500), .B2(n19748), .A(n14499), .ZN(P1_U2988) );
  INV_X1 U17685 ( .A(n14501), .ZN(n14543) );
  INV_X1 U17686 ( .A(n14502), .ZN(n14539) );
  INV_X1 U17687 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15746) );
  NAND3_X1 U17688 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14695) );
  NAND2_X1 U17689 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15754) );
  NOR2_X1 U17690 ( .A1(n14695), .A2(n15754), .ZN(n14507) );
  INV_X1 U17691 ( .A(n14507), .ZN(n14503) );
  NOR4_X1 U17692 ( .A1(n14506), .A2(n14505), .A3(n14504), .A4(n14503), .ZN(
        n15739) );
  NAND2_X1 U17693 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15739), .ZN(
        n15731) );
  NOR2_X1 U17694 ( .A1(n15746), .A2(n15731), .ZN(n14677) );
  NAND2_X1 U17695 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14677), .ZN(
        n14657) );
  NAND2_X1 U17696 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14507), .ZN(
        n15745) );
  NOR3_X1 U17697 ( .A1(n15729), .A2(n15737), .A3(n15745), .ZN(n14513) );
  NAND2_X1 U17698 ( .A1(n15736), .A2(n14513), .ZN(n14674) );
  INV_X1 U17699 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14514) );
  NAND2_X1 U17700 ( .A1(n14509), .A2(n14508), .ZN(n15698) );
  INV_X1 U17701 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14661) );
  NAND2_X1 U17702 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15711) );
  NOR2_X1 U17703 ( .A1(n14661), .A2(n15711), .ZN(n14659) );
  NAND2_X1 U17704 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14659), .ZN(
        n15697) );
  INV_X1 U17705 ( .A(n15697), .ZN(n14515) );
  AND2_X1 U17706 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14515), .ZN(
        n14510) );
  NAND2_X1 U17707 ( .A1(n15698), .A2(n14510), .ZN(n14650) );
  INV_X1 U17708 ( .A(n14642), .ZN(n14519) );
  AND2_X1 U17709 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14522) );
  NAND2_X1 U17710 ( .A1(n14635), .A2(n14522), .ZN(n14618) );
  NAND2_X1 U17711 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14525) );
  AND2_X1 U17712 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14532) );
  INV_X1 U17713 ( .A(n14532), .ZN(n14511) );
  NOR2_X1 U17714 ( .A1(n14595), .A2(n14511), .ZN(n14574) );
  NAND2_X1 U17715 ( .A1(n14574), .A2(n14528), .ZN(n14554) );
  INV_X1 U17716 ( .A(n14657), .ZN(n14678) );
  AND3_X1 U17717 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14678), .A3(
        n14515), .ZN(n14512) );
  OR2_X1 U17718 ( .A1(n15740), .A2(n14512), .ZN(n14518) );
  INV_X1 U17719 ( .A(n14513), .ZN(n14681) );
  NOR2_X1 U17720 ( .A1(n14514), .A2(n14681), .ZN(n15724) );
  NAND3_X1 U17721 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15724), .A3(
        n14515), .ZN(n14516) );
  NAND2_X1 U17722 ( .A1(n15736), .A2(n14516), .ZN(n14517) );
  NAND3_X1 U17723 ( .A1(n14518), .A2(n14520), .A3(n14517), .ZN(n14649) );
  OR2_X1 U17724 ( .A1(n14649), .A2(n14519), .ZN(n14521) );
  NAND2_X1 U17725 ( .A1(n14660), .A2(n14520), .ZN(n14696) );
  NAND2_X1 U17726 ( .A1(n14521), .A2(n14696), .ZN(n14632) );
  OR2_X1 U17727 ( .A1(n14660), .A2(n14522), .ZN(n14523) );
  NAND2_X1 U17728 ( .A1(n14632), .A2(n14523), .ZN(n14615) );
  AND2_X1 U17729 ( .A1(n15736), .A2(n14601), .ZN(n14524) );
  INV_X1 U17730 ( .A(n14525), .ZN(n14526) );
  NOR2_X1 U17731 ( .A1(n19914), .A2(n14526), .ZN(n14527) );
  NOR2_X1 U17732 ( .A1(n14606), .A2(n14527), .ZN(n14531) );
  INV_X1 U17733 ( .A(n14531), .ZN(n14535) );
  INV_X1 U17734 ( .A(n14528), .ZN(n14534) );
  INV_X1 U17735 ( .A(n14679), .ZN(n19918) );
  AOI22_X1 U17736 ( .A1(n19918), .A2(n14585), .B1(n15736), .B2(n14529), .ZN(
        n14530) );
  NAND2_X1 U17737 ( .A1(n14583), .A2(n14532), .ZN(n14587) );
  NAND2_X1 U17738 ( .A1(n14583), .A2(n14660), .ZN(n14533) );
  AOI21_X1 U17739 ( .B1(n14534), .B2(n14536), .A(n14575), .ZN(n14560) );
  OAI211_X1 U17740 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14660), .A(
        n14560), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14550) );
  OAI211_X1 U17741 ( .C1(n14536), .C2(n14535), .A(n14550), .B(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14538) );
  OAI211_X1 U17742 ( .C1(n14539), .C2(n14554), .A(n14538), .B(n14537), .ZN(
        n14540) );
  AOI21_X1 U17743 ( .B1(n14541), .B2(n19911), .A(n14540), .ZN(n14542) );
  OAI21_X1 U17744 ( .B1(n14543), .B2(n14704), .A(n14542), .ZN(P1_U3000) );
  INV_X1 U17745 ( .A(n14544), .ZN(n14552) );
  INV_X1 U17746 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14545) );
  OAI21_X1 U17747 ( .B1(n14554), .B2(n9900), .A(n14545), .ZN(n14549) );
  OAI21_X1 U17748 ( .B1(n14547), .B2(n15775), .A(n14546), .ZN(n14548) );
  AOI21_X1 U17749 ( .B1(n14550), .B2(n14549), .A(n14548), .ZN(n14551) );
  OAI21_X1 U17750 ( .B1(n14552), .B2(n14704), .A(n14551), .ZN(P1_U3001) );
  NAND2_X1 U17751 ( .A1(n14553), .A2(n19913), .ZN(n14559) );
  NOR2_X1 U17752 ( .A1(n14554), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14555) );
  AOI211_X1 U17753 ( .C1(n14557), .C2(n19911), .A(n14556), .B(n14555), .ZN(
        n14558) );
  OAI211_X1 U17754 ( .C1(n14560), .C2(n9900), .A(n14559), .B(n14558), .ZN(
        P1_U3002) );
  INV_X1 U17755 ( .A(n14561), .ZN(n14569) );
  XNOR2_X1 U17756 ( .A(n14562), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14563) );
  NAND2_X1 U17757 ( .A1(n14574), .A2(n14563), .ZN(n14564) );
  OAI211_X1 U17758 ( .C1(n14566), .C2(n15775), .A(n14565), .B(n14564), .ZN(
        n14567) );
  AOI21_X1 U17759 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14575), .A(
        n14567), .ZN(n14568) );
  OAI21_X1 U17760 ( .B1(n14569), .B2(n14704), .A(n14568), .ZN(P1_U3003) );
  NOR2_X1 U17761 ( .A1(n14570), .A2(n15775), .ZN(n14571) );
  AOI211_X1 U17762 ( .C1(n14574), .C2(n14573), .A(n14572), .B(n14571), .ZN(
        n14577) );
  NAND2_X1 U17763 ( .A1(n14575), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14576) );
  OAI211_X1 U17764 ( .C1(n14578), .C2(n14704), .A(n14577), .B(n14576), .ZN(
        P1_U3004) );
  INV_X1 U17765 ( .A(n14579), .ZN(n14591) );
  INV_X1 U17766 ( .A(n14580), .ZN(n14582) );
  AOI21_X1 U17767 ( .B1(n14582), .B2(n19911), .A(n14581), .ZN(n14590) );
  INV_X1 U17768 ( .A(n14583), .ZN(n14597) );
  INV_X1 U17769 ( .A(n14595), .ZN(n14588) );
  OAI21_X1 U17770 ( .B1(n14618), .B2(n14585), .A(n14584), .ZN(n14586) );
  OAI211_X1 U17771 ( .C1(n14597), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        n14589) );
  OAI211_X1 U17772 ( .C1(n14591), .C2(n14704), .A(n14590), .B(n14589), .ZN(
        P1_U3005) );
  AOI21_X1 U17773 ( .B1(n14593), .B2(n19911), .A(n14592), .ZN(n14594) );
  OAI21_X1 U17774 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14595), .A(
        n14594), .ZN(n14596) );
  AOI21_X1 U17775 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14597), .A(
        n14596), .ZN(n14598) );
  OAI21_X1 U17776 ( .B1(n14599), .B2(n14704), .A(n14598), .ZN(P1_U3006) );
  INV_X1 U17777 ( .A(n14600), .ZN(n14604) );
  NOR3_X1 U17778 ( .A1(n14618), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14601), .ZN(n14602) );
  AOI211_X1 U17779 ( .C1(n19911), .C2(n14604), .A(n14603), .B(n14602), .ZN(
        n14608) );
  NOR2_X1 U17780 ( .A1(n15730), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14605) );
  OAI21_X1 U17781 ( .B1(n14606), .B2(n14605), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14607) );
  OAI211_X1 U17782 ( .C1(n14609), .C2(n14704), .A(n14608), .B(n14607), .ZN(
        P1_U3007) );
  NAND2_X1 U17783 ( .A1(n14610), .A2(n19913), .ZN(n14617) );
  INV_X1 U17784 ( .A(n14611), .ZN(n14612) );
  NOR2_X1 U17785 ( .A1(n14612), .A2(n15775), .ZN(n14613) );
  AOI211_X1 U17786 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14615), .A(
        n14614), .B(n14613), .ZN(n14616) );
  OAI211_X1 U17787 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14618), .A(
        n14617), .B(n14616), .ZN(P1_U3008) );
  INV_X1 U17788 ( .A(n14635), .ZN(n14627) );
  XNOR2_X1 U17789 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14626) );
  NAND2_X1 U17790 ( .A1(n14619), .A2(n19913), .ZN(n14625) );
  INV_X1 U17791 ( .A(n14632), .ZN(n14623) );
  OAI21_X1 U17792 ( .B1(n14621), .B2(n15775), .A(n14620), .ZN(n14622) );
  AOI21_X1 U17793 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14623), .A(
        n14622), .ZN(n14624) );
  OAI211_X1 U17794 ( .C1(n14627), .C2(n14626), .A(n14625), .B(n14624), .ZN(
        P1_U3009) );
  INV_X1 U17795 ( .A(n14628), .ZN(n14630) );
  AOI21_X1 U17796 ( .B1(n14630), .B2(n19911), .A(n14629), .ZN(n14631) );
  OAI21_X1 U17797 ( .B1(n14634), .B2(n14632), .A(n14631), .ZN(n14633) );
  AOI21_X1 U17798 ( .B1(n14635), .B2(n14634), .A(n14633), .ZN(n14636) );
  OAI21_X1 U17799 ( .B1(n14637), .B2(n14704), .A(n14636), .ZN(P1_U3010) );
  NOR2_X1 U17800 ( .A1(n14638), .A2(n15775), .ZN(n14639) );
  AOI211_X1 U17801 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n14649), .A(
        n14640), .B(n14639), .ZN(n14644) );
  OR3_X1 U17802 ( .A1(n14650), .A2(n14642), .A3(n14641), .ZN(n14643) );
  OAI211_X1 U17803 ( .C1(n14645), .C2(n14704), .A(n14644), .B(n14643), .ZN(
        P1_U3011) );
  NOR2_X1 U17804 ( .A1(n14646), .A2(n15775), .ZN(n14647) );
  AOI211_X1 U17805 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n14649), .A(
        n14648), .B(n14647), .ZN(n14652) );
  OR2_X1 U17806 ( .A1(n14650), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14651) );
  OAI211_X1 U17807 ( .C1(n14653), .C2(n14704), .A(n14652), .B(n14651), .ZN(
        P1_U3012) );
  AOI21_X1 U17808 ( .B1(n14655), .B2(n19911), .A(n14654), .ZN(n14664) );
  AOI21_X1 U17809 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15724), .A(
        n14660), .ZN(n14656) );
  AOI211_X1 U17810 ( .C1(n14658), .C2(n14657), .A(n14656), .B(n15735), .ZN(
        n15716) );
  OAI21_X1 U17811 ( .B1(n14660), .B2(n14659), .A(n15716), .ZN(n15701) );
  NAND2_X1 U17812 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15698), .ZN(
        n15706) );
  OAI21_X1 U17813 ( .B1(n15711), .B2(n15706), .A(n14661), .ZN(n14662) );
  NAND2_X1 U17814 ( .A1(n15701), .A2(n14662), .ZN(n14663) );
  OAI211_X1 U17815 ( .C1(n14665), .C2(n14704), .A(n14664), .B(n14663), .ZN(
        P1_U3014) );
  INV_X1 U17816 ( .A(n14666), .ZN(n15638) );
  NAND2_X1 U17817 ( .A1(n15772), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14667) );
  OAI221_X1 U17818 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15706), 
        .C1(n14668), .C2(n15716), .A(n14667), .ZN(n14669) );
  AOI21_X1 U17819 ( .B1(n15638), .B2(n19911), .A(n14669), .ZN(n14670) );
  OAI21_X1 U17820 ( .B1(n14671), .B2(n14704), .A(n14670), .ZN(P1_U3016) );
  NOR2_X1 U17821 ( .A1(n14678), .A2(n14679), .ZN(n14676) );
  NOR2_X1 U17822 ( .A1(n19921), .A2(n20567), .ZN(n14675) );
  INV_X1 U17823 ( .A(n19914), .ZN(n14672) );
  NAND3_X1 U17824 ( .A1(n14672), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n14677), .ZN(n14673) );
  AOI21_X1 U17825 ( .B1(n14674), .B2(n14673), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15721) );
  AOI211_X1 U17826 ( .C1(n14677), .C2(n14676), .A(n14675), .B(n15721), .ZN(
        n14685) );
  OAI22_X1 U17827 ( .A1(n14679), .A2(n14678), .B1(n19914), .B2(n14677), .ZN(
        n14680) );
  AOI211_X1 U17828 ( .C1(n15736), .C2(n14681), .A(n14680), .B(n15735), .ZN(
        n14682) );
  INV_X1 U17829 ( .A(n14682), .ZN(n15720) );
  INV_X1 U17830 ( .A(n14683), .ZN(n15651) );
  AOI22_X1 U17831 ( .A1(n15720), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n19911), .B2(n15651), .ZN(n14684) );
  OAI211_X1 U17832 ( .C1(n14686), .C2(n14704), .A(n14685), .B(n14684), .ZN(
        P1_U3018) );
  XOR2_X1 U17833 ( .A(n14687), .B(n13590), .Z(n14690) );
  NAND2_X1 U17834 ( .A1(n14688), .A2(n13590), .ZN(n14689) );
  MUX2_X1 U17835 ( .A(n14690), .B(n14689), .S(n9593), .Z(n14693) );
  INV_X1 U17836 ( .A(n14691), .ZN(n14692) );
  NAND2_X1 U17837 ( .A1(n14693), .A2(n14692), .ZN(n15685) );
  INV_X1 U17838 ( .A(n14695), .ZN(n14694) );
  NAND2_X1 U17839 ( .A1(n14694), .A2(n15771), .ZN(n15759) );
  INV_X1 U17840 ( .A(n15759), .ZN(n15747) );
  OAI211_X1 U17841 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15747), .B(n15754), .ZN(n14703) );
  NOR2_X1 U17842 ( .A1(n14695), .A2(n15737), .ZN(n14698) );
  INV_X1 U17843 ( .A(n14696), .ZN(n14697) );
  AOI21_X1 U17844 ( .B1(n14699), .B2(n14698), .A(n14697), .ZN(n15755) );
  INV_X1 U17845 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20561) );
  OAI22_X1 U17846 ( .A1(n19921), .A2(n20561), .B1(n15775), .B2(n14700), .ZN(
        n14701) );
  AOI21_X1 U17847 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15755), .A(
        n14701), .ZN(n14702) );
  OAI211_X1 U17848 ( .C1(n15685), .C2(n14704), .A(n14703), .B(n14702), .ZN(
        P1_U3021) );
  NAND3_X1 U17849 ( .A1(n14705), .A2(n15600), .A3(n15781), .ZN(n15607) );
  NAND2_X1 U17850 ( .A1(n11631), .A2(n14706), .ZN(n14707) );
  OAI211_X1 U17851 ( .C1(n20469), .C2(n20009), .A(n15607), .B(n14707), .ZN(
        n14708) );
  MUX2_X1 U17852 ( .A(n14708), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        n19922), .Z(P1_U3478) );
  INV_X1 U17853 ( .A(n14711), .ZN(n14718) );
  OR2_X1 U17854 ( .A1(n13879), .A2(n14709), .ZN(n14714) );
  AOI22_X1 U17855 ( .A1(n14712), .A2(n11512), .B1(n14711), .B2(n14710), .ZN(
        n14713) );
  NAND2_X1 U17856 ( .A1(n14714), .A2(n14713), .ZN(n15582) );
  NOR2_X1 U17857 ( .A1(n15606), .A2(n14715), .ZN(n14721) );
  INV_X1 U17858 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20697) );
  AOI22_X1 U17859 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n20697), .B2(n12833), .ZN(
        n14720) );
  INV_X1 U17860 ( .A(n14720), .ZN(n14716) );
  AOI22_X1 U17861 ( .A1(n15582), .A2(n14722), .B1(n14721), .B2(n14716), .ZN(
        n14717) );
  OAI21_X1 U17862 ( .B1(n20609), .B2(n14718), .A(n14717), .ZN(n14719) );
  MUX2_X1 U17863 ( .A(n14719), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n20613), .Z(P1_U3473) );
  AOI22_X1 U17864 ( .A1(n14723), .A2(n14722), .B1(n14721), .B2(n14720), .ZN(
        n14724) );
  OAI21_X1 U17865 ( .B1(n20609), .B2(n14725), .A(n14724), .ZN(n14726) );
  MUX2_X1 U17866 ( .A(n14726), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n20613), .Z(P1_U3472) );
  NAND2_X1 U17867 ( .A1(n10918), .A2(n14727), .ZN(n14728) );
  NAND2_X1 U17868 ( .A1(n9637), .A2(n14728), .ZN(n15799) );
  OR2_X1 U17869 ( .A1(n14730), .A2(n14729), .ZN(n14787) );
  NAND3_X1 U17870 ( .A1(n14787), .A2(n14731), .A3(n18848), .ZN(n14733) );
  NAND2_X1 U17871 ( .A1(n18843), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14732) );
  OAI211_X1 U17872 ( .C1(n15799), .C2(n18843), .A(n14733), .B(n14732), .ZN(
        P2_U2858) );
  NOR2_X1 U17873 ( .A1(n14734), .A2(n14735), .ZN(n14737) );
  XNOR2_X1 U17874 ( .A(n14737), .B(n14736), .ZN(n14798) );
  NAND2_X1 U17875 ( .A1(n14798), .A2(n18848), .ZN(n14739) );
  NAND2_X1 U17876 ( .A1(n18843), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14738) );
  OAI211_X1 U17877 ( .C1(n18843), .C2(n15805), .A(n14739), .B(n14738), .ZN(
        P2_U2859) );
  OAI21_X1 U17878 ( .B1(n14742), .B2(n14741), .A(n14740), .ZN(n14810) );
  XNOR2_X1 U17879 ( .A(n14747), .B(n14743), .ZN(n15825) );
  NOR2_X1 U17880 ( .A1(n15825), .A2(n18843), .ZN(n14744) );
  AOI21_X1 U17881 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n18843), .A(n14744), .ZN(
        n14745) );
  OAI21_X1 U17882 ( .B1(n14810), .B2(n18844), .A(n14745), .ZN(P2_U2860) );
  AND2_X1 U17883 ( .A1(n14760), .A2(n14746), .ZN(n14748) );
  OR2_X1 U17884 ( .A1(n14748), .A2(n14747), .ZN(n15106) );
  AOI21_X1 U17885 ( .B1(n14751), .B2(n14750), .A(n14749), .ZN(n14813) );
  NAND2_X1 U17886 ( .A1(n14813), .A2(n18848), .ZN(n14753) );
  NAND2_X1 U17887 ( .A1(n18843), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14752) );
  OAI211_X1 U17888 ( .C1(n15106), .C2(n18843), .A(n14753), .B(n14752), .ZN(
        P2_U2861) );
  OAI21_X1 U17889 ( .B1(n14756), .B2(n14755), .A(n14754), .ZN(n14829) );
  NAND2_X1 U17890 ( .A1(n14757), .A2(n14758), .ZN(n14759) );
  NAND2_X1 U17891 ( .A1(n14760), .A2(n14759), .ZN(n15840) );
  NOR2_X1 U17892 ( .A1(n15840), .A2(n18843), .ZN(n14761) );
  AOI21_X1 U17893 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n18843), .A(n14761), .ZN(
        n14762) );
  OAI21_X1 U17894 ( .B1(n14829), .B2(n18844), .A(n14762), .ZN(P2_U2862) );
  AOI21_X1 U17895 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n14766) );
  XOR2_X1 U17896 ( .A(n14767), .B(n14766), .Z(n14838) );
  OAI21_X1 U17897 ( .B1(n14769), .B2(n14768), .A(n14757), .ZN(n14917) );
  MUX2_X1 U17898 ( .A(n15853), .B(n14917), .S(n18851), .Z(n14770) );
  OAI21_X1 U17899 ( .B1(n14838), .B2(n18844), .A(n14770), .ZN(P2_U2863) );
  NAND2_X1 U17900 ( .A1(n14772), .A2(n14773), .ZN(n14774) );
  AND2_X1 U17901 ( .A1(n14771), .A2(n14774), .ZN(n14853) );
  NAND2_X1 U17902 ( .A1(n14853), .A2(n18848), .ZN(n14777) );
  INV_X1 U17903 ( .A(n15161), .ZN(n14775) );
  NAND2_X1 U17904 ( .A1(n14775), .A2(n18851), .ZN(n14776) );
  OAI211_X1 U17905 ( .C1(n18851), .C2(n10803), .A(n14777), .B(n14776), .ZN(
        P2_U2866) );
  INV_X1 U17906 ( .A(n15871), .ZN(n14778) );
  OAI21_X1 U17907 ( .B1(n13687), .B2(n14779), .A(n14778), .ZN(n14865) );
  NOR2_X1 U17908 ( .A1(n14780), .A2(n14781), .ZN(n14782) );
  OR2_X1 U17909 ( .A1(n14981), .A2(n14782), .ZN(n18640) );
  NOR2_X1 U17910 ( .A1(n18640), .A2(n18843), .ZN(n14783) );
  AOI21_X1 U17911 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n18843), .A(n14783), .ZN(
        n14784) );
  OAI21_X1 U17912 ( .B1(n14865), .B2(n18844), .A(n14784), .ZN(P2_U2868) );
  NOR2_X1 U17913 ( .A1(n14796), .A2(n14785), .ZN(n14786) );
  NAND3_X1 U17914 ( .A1(n14787), .A2(n14731), .A3(n18884), .ZN(n14793) );
  INV_X1 U17915 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n14790) );
  INV_X1 U17916 ( .A(n18953), .ZN(n14788) );
  AOI22_X1 U17917 ( .A1(n18857), .A2(n14788), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n18881), .ZN(n14789) );
  OAI21_X1 U17918 ( .B1(n14835), .B2(n14790), .A(n14789), .ZN(n14791) );
  AOI21_X1 U17919 ( .B1(n18859), .B2(BUF1_REG_29__SCAN_IN), .A(n14791), .ZN(
        n14792) );
  OAI211_X1 U17920 ( .C1(n15803), .C2(n18862), .A(n14793), .B(n14792), .ZN(
        P2_U2890) );
  NOR2_X1 U17921 ( .A1(n14795), .A2(n14794), .ZN(n14797) );
  NOR2_X1 U17922 ( .A1(n14797), .A2(n14796), .ZN(n15806) );
  INV_X1 U17923 ( .A(n15806), .ZN(n15087) );
  NAND2_X1 U17924 ( .A1(n14798), .A2(n18884), .ZN(n14804) );
  INV_X1 U17925 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n14801) );
  INV_X1 U17926 ( .A(n18951), .ZN(n14799) );
  AOI22_X1 U17927 ( .A1(n18857), .A2(n14799), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n18881), .ZN(n14800) );
  OAI21_X1 U17928 ( .B1(n14835), .B2(n14801), .A(n14800), .ZN(n14802) );
  AOI21_X1 U17929 ( .B1(n18859), .B2(BUF1_REG_28__SCAN_IN), .A(n14802), .ZN(
        n14803) );
  OAI211_X1 U17930 ( .C1(n18862), .C2(n15087), .A(n14804), .B(n14803), .ZN(
        P2_U2891) );
  XOR2_X1 U17931 ( .A(n14805), .B(n9636), .Z(n15822) );
  INV_X1 U17932 ( .A(n18859), .ZN(n14860) );
  AOI22_X1 U17933 ( .A1(n18857), .A2(n18871), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n18881), .ZN(n14807) );
  NAND2_X1 U17934 ( .A1(n18858), .A2(BUF2_REG_27__SCAN_IN), .ZN(n14806) );
  OAI211_X1 U17935 ( .C1(n14860), .C2(n19014), .A(n14807), .B(n14806), .ZN(
        n14808) );
  AOI21_X1 U17936 ( .B1(n15822), .B2(n18852), .A(n14808), .ZN(n14809) );
  OAI21_X1 U17937 ( .B1(n14810), .B2(n18861), .A(n14809), .ZN(P2_U2892) );
  NAND2_X1 U17938 ( .A1(n14825), .A2(n14811), .ZN(n14812) );
  AND2_X1 U17939 ( .A1(n9636), .A2(n14812), .ZN(n15827) );
  INV_X1 U17940 ( .A(n15827), .ZN(n14819) );
  NAND2_X1 U17941 ( .A1(n14813), .A2(n18884), .ZN(n14818) );
  INV_X1 U17942 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n14815) );
  AOI22_X1 U17943 ( .A1(n18857), .A2(n18874), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n18881), .ZN(n14814) );
  OAI21_X1 U17944 ( .B1(n14835), .B2(n14815), .A(n14814), .ZN(n14816) );
  AOI21_X1 U17945 ( .B1(n18859), .B2(BUF1_REG_26__SCAN_IN), .A(n14816), .ZN(
        n14817) );
  OAI211_X1 U17946 ( .C1(n14819), .C2(n18862), .A(n14818), .B(n14817), .ZN(
        P2_U2893) );
  NAND2_X1 U17947 ( .A1(n18858), .A2(BUF2_REG_25__SCAN_IN), .ZN(n14822) );
  INV_X1 U17948 ( .A(n18949), .ZN(n14820) );
  AOI22_X1 U17949 ( .A1(n18857), .A2(n14820), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n18881), .ZN(n14821) );
  NAND2_X1 U17950 ( .A1(n14822), .A2(n14821), .ZN(n14827) );
  OR2_X1 U17951 ( .A1(n14830), .A2(n14823), .ZN(n14824) );
  NAND2_X1 U17952 ( .A1(n14825), .A2(n14824), .ZN(n15848) );
  NOR2_X1 U17953 ( .A1(n15848), .A2(n18862), .ZN(n14826) );
  AOI211_X1 U17954 ( .C1(BUF1_REG_25__SCAN_IN), .C2(n18859), .A(n14827), .B(
        n14826), .ZN(n14828) );
  OAI21_X1 U17955 ( .B1(n14829), .B2(n18861), .A(n14828), .ZN(P2_U2894) );
  AOI21_X1 U17956 ( .B1(n14832), .B2(n14831), .A(n14830), .ZN(n15859) );
  AOI22_X1 U17957 ( .A1(n18857), .A2(n18878), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n18881), .ZN(n14834) );
  NAND2_X1 U17958 ( .A1(n18859), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14833) );
  OAI211_X1 U17959 ( .C1(n14835), .C2(n17917), .A(n14834), .B(n14833), .ZN(
        n14836) );
  AOI21_X1 U17960 ( .B1(n15859), .B2(n18852), .A(n14836), .ZN(n14837) );
  OAI21_X1 U17961 ( .B1(n14838), .B2(n18861), .A(n14837), .ZN(P2_U2895) );
  OAI22_X1 U17962 ( .A1(n19047), .A2(n14859), .B1(n14858), .B2(n14839), .ZN(
        n14841) );
  NOR2_X1 U17963 ( .A1(n14860), .A2(n19040), .ZN(n14840) );
  AOI211_X1 U17964 ( .C1(n18858), .C2(BUF2_REG_23__SCAN_IN), .A(n14841), .B(
        n14840), .ZN(n14846) );
  AOI21_X1 U17965 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(n15863) );
  NAND2_X1 U17966 ( .A1(n15863), .A2(n18884), .ZN(n14845) );
  OAI211_X1 U17967 ( .C1(n15140), .C2(n18862), .A(n14846), .B(n14845), .ZN(
        P2_U2896) );
  AOI22_X1 U17968 ( .A1(n14848), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14847), .ZN(n19029) );
  INV_X1 U17969 ( .A(n19029), .ZN(n18882) );
  AOI22_X1 U17970 ( .A1(n18857), .A2(n18882), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n18881), .ZN(n14850) );
  NAND2_X1 U17971 ( .A1(n18858), .A2(BUF2_REG_21__SCAN_IN), .ZN(n14849) );
  OAI211_X1 U17972 ( .C1(n14860), .C2(n14851), .A(n14850), .B(n14849), .ZN(
        n14852) );
  AOI21_X1 U17973 ( .B1(n14853), .B2(n18884), .A(n14852), .ZN(n14854) );
  OAI21_X1 U17974 ( .B1(n15168), .B2(n18862), .A(n14854), .ZN(P2_U2898) );
  XOR2_X1 U17975 ( .A(n14856), .B(n14855), .Z(n18638) );
  NAND2_X1 U17976 ( .A1(n18638), .A2(n18852), .ZN(n14864) );
  OAI22_X1 U17977 ( .A1(n19017), .A2(n14859), .B1(n14858), .B2(n14857), .ZN(
        n14862) );
  NOR2_X1 U17978 ( .A1(n14860), .A2(n16103), .ZN(n14861) );
  AOI211_X1 U17979 ( .C1(n18858), .C2(BUF2_REG_19__SCAN_IN), .A(n14862), .B(
        n14861), .ZN(n14863) );
  OAI211_X1 U17980 ( .C1(n18861), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        P2_U2900) );
  INV_X1 U17981 ( .A(n15788), .ZN(n14869) );
  INV_X1 U17982 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14867) );
  OAI21_X1 U17983 ( .B1(n15953), .B2(n14867), .A(n14866), .ZN(n14868) );
  AOI21_X1 U17984 ( .B1(n15944), .B2(n14869), .A(n14868), .ZN(n14870) );
  OAI21_X1 U17985 ( .B1(n14871), .B2(n15063), .A(n14870), .ZN(n14872) );
  OAI21_X1 U17986 ( .B1(n14875), .B2(n15946), .A(n14874), .ZN(P2_U2984) );
  NOR2_X1 U17987 ( .A1(n14888), .A2(n20769), .ZN(n14877) );
  OAI21_X1 U17988 ( .B1(n14877), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14876), .ZN(n15081) );
  INV_X1 U17989 ( .A(n14878), .ZN(n14879) );
  NOR2_X1 U17990 ( .A1(n14880), .A2(n14879), .ZN(n14881) );
  XNOR2_X1 U17991 ( .A(n14882), .B(n14881), .ZN(n15078) );
  NOR2_X1 U17992 ( .A1(n15891), .A2(n20752), .ZN(n15068) );
  AOI21_X1 U17993 ( .B1(n15915), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15068), .ZN(n14884) );
  NAND2_X1 U17994 ( .A1(n15944), .A2(n15794), .ZN(n14883) );
  OAI211_X1 U17995 ( .C1(n15799), .C2(n15063), .A(n14884), .B(n14883), .ZN(
        n14885) );
  AOI21_X1 U17996 ( .B1(n15078), .B2(n10903), .A(n14885), .ZN(n14886) );
  OAI21_X1 U17997 ( .B1(n15081), .B2(n15947), .A(n14886), .ZN(P2_U2985) );
  XNOR2_X1 U17998 ( .A(n14887), .B(n15097), .ZN(n15102) );
  INV_X1 U17999 ( .A(n14888), .ZN(n14889) );
  AOI21_X1 U18000 ( .B1(n15097), .B2(n14902), .A(n14889), .ZN(n15100) );
  OR2_X1 U18001 ( .A1(n15891), .A2(n19674), .ZN(n15092) );
  OAI21_X1 U18002 ( .B1(n15953), .B2(n14890), .A(n15092), .ZN(n14891) );
  AOI21_X1 U18003 ( .B1(n15944), .B2(n15819), .A(n14891), .ZN(n14892) );
  OAI21_X1 U18004 ( .B1(n15825), .B2(n15063), .A(n14892), .ZN(n14893) );
  AOI21_X1 U18005 ( .B1(n15100), .B2(n15939), .A(n14893), .ZN(n14894) );
  OAI21_X1 U18006 ( .B1(n15102), .B2(n15946), .A(n14894), .ZN(P2_U2987) );
  AOI21_X1 U18007 ( .B1(n9896), .B2(n14906), .A(n14895), .ZN(n14897) );
  XNOR2_X1 U18008 ( .A(n14897), .B(n14896), .ZN(n15115) );
  INV_X1 U18009 ( .A(n15106), .ZN(n15828) );
  NAND2_X1 U18010 ( .A1(n15944), .A2(n15831), .ZN(n14899) );
  OR2_X1 U18011 ( .A1(n15891), .A2(n14898), .ZN(n15105) );
  OAI211_X1 U18012 ( .C1(n14900), .C2(n15953), .A(n14899), .B(n15105), .ZN(
        n14904) );
  OAI21_X1 U18013 ( .B1(n14901), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14902), .ZN(n15103) );
  NOR2_X1 U18014 ( .A1(n15103), .A2(n15947), .ZN(n14903) );
  OAI21_X1 U18015 ( .B1(n15946), .B2(n15115), .A(n14905), .ZN(P2_U2988) );
  NAND2_X1 U18016 ( .A1(n14907), .A2(n14906), .ZN(n14908) );
  XNOR2_X1 U18017 ( .A(n9896), .B(n14908), .ZN(n15126) );
  AOI21_X1 U18018 ( .B1(n15118), .B2(n14909), .A(n14901), .ZN(n15124) );
  OR2_X1 U18019 ( .A1(n15891), .A2(n19669), .ZN(n15116) );
  OAI21_X1 U18020 ( .B1(n15953), .B2(n9985), .A(n15116), .ZN(n14910) );
  AOI21_X1 U18021 ( .B1(n15944), .B2(n15842), .A(n14910), .ZN(n14911) );
  OAI21_X1 U18022 ( .B1(n15840), .B2(n15063), .A(n14911), .ZN(n14912) );
  AOI21_X1 U18023 ( .B1(n15124), .B2(n15939), .A(n14912), .ZN(n14913) );
  OAI21_X1 U18024 ( .B1(n15946), .B2(n15126), .A(n14913), .ZN(P2_U2989) );
  XNOR2_X1 U18025 ( .A(n14914), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14915) );
  XNOR2_X1 U18026 ( .A(n14916), .B(n14915), .ZN(n15135) );
  INV_X1 U18027 ( .A(n14917), .ZN(n15849) );
  NOR2_X1 U18028 ( .A1(n15891), .A2(n19667), .ZN(n15127) );
  AOI21_X1 U18029 ( .B1(n15915), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15127), .ZN(n14918) );
  OAI21_X1 U18030 ( .B1(n15922), .B2(n14919), .A(n14918), .ZN(n14921) );
  OAI21_X1 U18031 ( .B1(n9611), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14909), .ZN(n15131) );
  NOR2_X1 U18032 ( .A1(n15131), .A2(n15947), .ZN(n14920) );
  AOI211_X1 U18033 ( .C1(n15849), .C2(n15950), .A(n14921), .B(n14920), .ZN(
        n14922) );
  OAI21_X1 U18034 ( .B1(n15135), .B2(n15946), .A(n14922), .ZN(P2_U2990) );
  XNOR2_X1 U18035 ( .A(n14924), .B(n14923), .ZN(n15145) );
  INV_X1 U18036 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14925) );
  NAND2_X1 U18037 ( .A1(n9642), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14933) );
  AOI21_X1 U18038 ( .B1(n14925), .B2(n14933), .A(n9611), .ZN(n15136) );
  NAND2_X1 U18039 ( .A1(n15136), .A2(n15939), .ZN(n14932) );
  NAND2_X1 U18040 ( .A1(n15944), .A2(n14926), .ZN(n14927) );
  NAND2_X1 U18041 ( .A1(n18791), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15138) );
  OAI211_X1 U18042 ( .C1(n14928), .C2(n15953), .A(n14927), .B(n15138), .ZN(
        n14929) );
  AOI21_X1 U18043 ( .B1(n14930), .B2(n15950), .A(n14929), .ZN(n14931) );
  OAI211_X1 U18044 ( .C1(n15145), .C2(n15946), .A(n14932), .B(n14931), .ZN(
        P2_U2991) );
  OAI21_X1 U18045 ( .B1(n9642), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n14933), .ZN(n15158) );
  NAND2_X1 U18046 ( .A1(n14935), .A2(n14934), .ZN(n14936) );
  XNOR2_X1 U18047 ( .A(n14937), .B(n14936), .ZN(n15155) );
  NAND2_X1 U18048 ( .A1(n14939), .A2(n14938), .ZN(n14940) );
  AND2_X1 U18049 ( .A1(n14941), .A2(n14940), .ZN(n15570) );
  INV_X1 U18050 ( .A(n15570), .ZN(n15869) );
  NOR2_X1 U18051 ( .A1(n15891), .A2(n14942), .ZN(n15149) );
  NOR2_X1 U18052 ( .A1(n15922), .A2(n14943), .ZN(n14944) );
  AOI211_X1 U18053 ( .C1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n15915), .A(
        n15149), .B(n14944), .ZN(n14945) );
  OAI21_X1 U18054 ( .B1(n15869), .B2(n15063), .A(n14945), .ZN(n14946) );
  AOI21_X1 U18055 ( .B1(n15155), .B2(n10903), .A(n14946), .ZN(n14947) );
  OAI21_X1 U18056 ( .B1(n15158), .B2(n15947), .A(n14947), .ZN(P2_U2992) );
  XNOR2_X1 U18057 ( .A(n14950), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15053) );
  INV_X1 U18058 ( .A(n14951), .ZN(n14952) );
  INV_X1 U18059 ( .A(n15894), .ZN(n14953) );
  INV_X1 U18060 ( .A(n15039), .ZN(n14955) );
  INV_X1 U18061 ( .A(n14956), .ZN(n15026) );
  NOR2_X1 U18062 ( .A1(n14959), .A2(n10865), .ZN(n15001) );
  NOR2_X1 U18063 ( .A1(n14961), .A2(n10865), .ZN(n14975) );
  OAI21_X1 U18064 ( .B1(n14963), .B2(n10865), .A(n14962), .ZN(n14964) );
  XNOR2_X1 U18065 ( .A(n14965), .B(n14964), .ZN(n15172) );
  AOI21_X1 U18066 ( .B1(n14967), .B2(n14966), .A(n9642), .ZN(n15170) );
  NAND2_X1 U18067 ( .A1(n18791), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15160) );
  OAI21_X1 U18068 ( .B1(n15953), .B2(n14968), .A(n15160), .ZN(n14969) );
  AOI21_X1 U18069 ( .B1(n15944), .B2(n14970), .A(n14969), .ZN(n14971) );
  OAI21_X1 U18070 ( .B1(n15161), .B2(n15063), .A(n14971), .ZN(n14972) );
  AOI21_X1 U18071 ( .B1(n15170), .B2(n15939), .A(n14972), .ZN(n14973) );
  OAI21_X1 U18072 ( .B1(n15172), .B2(n15946), .A(n14973), .ZN(P2_U2993) );
  NOR2_X1 U18073 ( .A1(n14975), .A2(n10088), .ZN(n14976) );
  XNOR2_X1 U18074 ( .A(n14977), .B(n14976), .ZN(n15188) );
  INV_X1 U18075 ( .A(n14966), .ZN(n14979) );
  AOI21_X1 U18076 ( .B1(n15183), .B2(n14978), .A(n14979), .ZN(n15186) );
  OR2_X1 U18077 ( .A1(n14981), .A2(n14980), .ZN(n14982) );
  AND2_X1 U18078 ( .A1(n14983), .A2(n14982), .ZN(n18621) );
  NAND2_X1 U18079 ( .A1(n18621), .A2(n15950), .ZN(n14985) );
  NOR2_X1 U18080 ( .A1(n15891), .A2(n19661), .ZN(n15181) );
  AOI21_X1 U18081 ( .B1(n15915), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15181), .ZN(n14984) );
  OAI211_X1 U18082 ( .C1(n15922), .C2(n14986), .A(n14985), .B(n14984), .ZN(
        n14987) );
  AOI21_X1 U18083 ( .B1(n15186), .B2(n15939), .A(n14987), .ZN(n14988) );
  OAI21_X1 U18084 ( .B1(n15188), .B2(n15946), .A(n14988), .ZN(P2_U2994) );
  NAND2_X1 U18085 ( .A1(n14990), .A2(n14989), .ZN(n14993) );
  INV_X1 U18086 ( .A(n14991), .ZN(n15000) );
  XOR2_X1 U18087 ( .A(n14993), .B(n14992), .Z(n15200) );
  INV_X1 U18088 ( .A(n14994), .ZN(n15011) );
  INV_X1 U18089 ( .A(n14978), .ZN(n14995) );
  AOI21_X1 U18090 ( .B1(n15195), .B2(n15011), .A(n14995), .ZN(n15198) );
  NOR2_X1 U18091 ( .A1(n18970), .A2(n19660), .ZN(n15191) );
  AOI21_X1 U18092 ( .B1(n15915), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15191), .ZN(n14997) );
  NAND2_X1 U18093 ( .A1(n15944), .A2(n18632), .ZN(n14996) );
  OAI211_X1 U18094 ( .C1(n18640), .C2(n15063), .A(n14997), .B(n14996), .ZN(
        n14998) );
  AOI21_X1 U18095 ( .B1(n15198), .B2(n15939), .A(n14998), .ZN(n14999) );
  OAI21_X1 U18096 ( .B1(n15200), .B2(n15946), .A(n14999), .ZN(P2_U2995) );
  NOR2_X1 U18097 ( .A1(n15001), .A2(n15000), .ZN(n15002) );
  XNOR2_X1 U18098 ( .A(n15015), .B(n15002), .ZN(n15216) );
  AND2_X1 U18099 ( .A1(n15004), .A2(n15003), .ZN(n15005) );
  NOR2_X1 U18100 ( .A1(n15891), .A2(n19658), .ZN(n15207) );
  AOI21_X1 U18101 ( .B1(n15915), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15207), .ZN(n15006) );
  OAI21_X1 U18102 ( .B1(n15922), .B2(n15007), .A(n15006), .ZN(n15013) );
  OAI21_X1 U18103 ( .B1(n15220), .B2(n15009), .A(n15209), .ZN(n15010) );
  NAND2_X1 U18104 ( .A1(n15011), .A2(n15010), .ZN(n15211) );
  NOR2_X1 U18105 ( .A1(n15211), .A2(n15947), .ZN(n15012) );
  AOI211_X1 U18106 ( .C1(n15950), .C2(n10111), .A(n15013), .B(n15012), .ZN(
        n15014) );
  OAI21_X1 U18107 ( .B1(n15216), .B2(n15946), .A(n15014), .ZN(P2_U2996) );
  INV_X1 U18108 ( .A(n15015), .ZN(n15019) );
  AOI22_X1 U18109 ( .A1(n15019), .A2(n15018), .B1(n15017), .B2(n15016), .ZN(
        n15231) );
  XNOR2_X1 U18110 ( .A(n15220), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15023) );
  NAND2_X1 U18111 ( .A1(n18656), .A2(n15950), .ZN(n15021) );
  NOR2_X1 U18112 ( .A1(n18970), .A2(n19656), .ZN(n15224) );
  AOI21_X1 U18113 ( .B1(n15915), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15224), .ZN(n15020) );
  OAI211_X1 U18114 ( .C1(n15922), .C2(n18661), .A(n15021), .B(n15020), .ZN(
        n15022) );
  AOI21_X1 U18115 ( .B1(n15023), .B2(n15939), .A(n15022), .ZN(n15024) );
  OAI21_X1 U18116 ( .B1(n15231), .B2(n15946), .A(n15024), .ZN(P2_U2997) );
  XNOR2_X1 U18117 ( .A(n15025), .B(n15026), .ZN(n15244) );
  OR2_X1 U18118 ( .A1(n15028), .A2(n15027), .ZN(n15029) );
  AND2_X1 U18119 ( .A1(n9624), .A2(n15029), .ZN(n18841) );
  NAND2_X1 U18120 ( .A1(n15944), .A2(n18664), .ZN(n15030) );
  NAND2_X1 U18121 ( .A1(n18791), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15238) );
  OAI211_X1 U18122 ( .C1(n15031), .C2(n15953), .A(n15030), .B(n15238), .ZN(
        n15036) );
  INV_X1 U18123 ( .A(n15220), .ZN(n15223) );
  AOI21_X1 U18124 ( .B1(n15033), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15034) );
  NOR3_X1 U18125 ( .A1(n15223), .A2(n15034), .A3(n15947), .ZN(n15035) );
  AOI211_X1 U18126 ( .C1(n15950), .C2(n18841), .A(n15036), .B(n15035), .ZN(
        n15037) );
  OAI21_X1 U18127 ( .B1(n15244), .B2(n15946), .A(n15037), .ZN(P2_U2998) );
  NAND2_X1 U18128 ( .A1(n15039), .A2(n15038), .ZN(n15041) );
  XOR2_X1 U18129 ( .A(n15041), .B(n15040), .Z(n15256) );
  XNOR2_X1 U18130 ( .A(n15033), .B(n15250), .ZN(n15254) );
  OAI22_X1 U18131 ( .A1(n15953), .A2(n18685), .B1(n15042), .B2(n15891), .ZN(
        n15043) );
  AOI21_X1 U18132 ( .B1(n15944), .B2(n15044), .A(n15043), .ZN(n15045) );
  OAI21_X1 U18133 ( .B1(n15063), .B2(n18680), .A(n15045), .ZN(n15046) );
  AOI21_X1 U18134 ( .B1(n15254), .B2(n15939), .A(n15046), .ZN(n15047) );
  OAI21_X1 U18135 ( .B1(n15256), .B2(n15946), .A(n15047), .ZN(P2_U2999) );
  INV_X1 U18136 ( .A(n15313), .ZN(n15049) );
  INV_X1 U18137 ( .A(n15293), .ZN(n15312) );
  INV_X1 U18138 ( .A(n15266), .ZN(n15285) );
  NOR2_X1 U18139 ( .A1(n15312), .A2(n15285), .ZN(n15278) );
  NAND2_X1 U18140 ( .A1(n15313), .A2(n15050), .ZN(n15262) );
  OAI21_X1 U18141 ( .B1(n15278), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15262), .ZN(n15977) );
  NAND2_X1 U18142 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18791), .ZN(n15969) );
  INV_X1 U18143 ( .A(n15969), .ZN(n15052) );
  INV_X1 U18144 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20739) );
  OAI22_X1 U18145 ( .A1(n20739), .A2(n15953), .B1(n15922), .B2(n18710), .ZN(
        n15051) );
  AOI211_X1 U18146 ( .C1(n18715), .C2(n15950), .A(n15052), .B(n15051), .ZN(
        n15056) );
  XNOR2_X1 U18147 ( .A(n15054), .B(n15053), .ZN(n15974) );
  NAND2_X1 U18148 ( .A1(n15974), .A2(n10903), .ZN(n15055) );
  OAI211_X1 U18149 ( .C1(n15977), .C2(n15947), .A(n15056), .B(n15055), .ZN(
        P2_U3002) );
  XNOR2_X1 U18150 ( .A(n15058), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15059) );
  XNOR2_X1 U18151 ( .A(n15057), .B(n15059), .ZN(n15335) );
  NAND2_X1 U18152 ( .A1(n10099), .A2(n15933), .ZN(n15060) );
  OAI22_X1 U18153 ( .A1(n10622), .A2(n15891), .B1(n15922), .B2(n18766), .ZN(
        n15061) );
  AOI21_X1 U18154 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n15915), .A(
        n15061), .ZN(n15062) );
  OAI21_X1 U18155 ( .B1(n15063), .B2(n18769), .A(n15062), .ZN(n15064) );
  AOI21_X1 U18156 ( .B1(n15333), .B2(n10903), .A(n15064), .ZN(n15065) );
  OAI21_X1 U18157 ( .B1(n15335), .B2(n15947), .A(n15065), .ZN(P2_U3007) );
  INV_X1 U18158 ( .A(n15803), .ZN(n15077) );
  NAND2_X1 U18159 ( .A1(n15203), .A2(n15097), .ZN(n15066) );
  NAND2_X1 U18160 ( .A1(n15098), .A2(n15066), .ZN(n15085) );
  NAND2_X1 U18161 ( .A1(n20769), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15067) );
  NOR2_X1 U18162 ( .A1(n15070), .A2(n15067), .ZN(n15083) );
  OAI21_X1 U18163 ( .B1(n15085), .B2(n15083), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15075) );
  INV_X1 U18164 ( .A(n15799), .ZN(n15069) );
  AOI21_X1 U18165 ( .B1(n15069), .B2(n18982), .A(n15068), .ZN(n15074) );
  INV_X1 U18166 ( .A(n15070), .ZN(n15094) );
  NAND3_X1 U18167 ( .A1(n15094), .A2(n15072), .A3(n15071), .ZN(n15073) );
  NAND3_X1 U18168 ( .A1(n15075), .A2(n15074), .A3(n15073), .ZN(n15076) );
  AOI21_X1 U18169 ( .B1(n15077), .B2(n15982), .A(n15076), .ZN(n15080) );
  NAND2_X1 U18170 ( .A1(n15078), .A2(n11303), .ZN(n15079) );
  OAI211_X1 U18171 ( .C1(n15081), .C2(n15978), .A(n15080), .B(n15079), .ZN(
        P2_U3017) );
  OAI21_X1 U18172 ( .B1(n15805), .B2(n15330), .A(n15082), .ZN(n15084) );
  OAI21_X1 U18173 ( .B1(n15087), .B2(n18986), .A(n15086), .ZN(n15088) );
  OAI21_X1 U18174 ( .B1(n15091), .B2(n15309), .A(n15090), .ZN(P2_U3018) );
  NAND2_X1 U18175 ( .A1(n15822), .A2(n15982), .ZN(n15096) );
  OAI21_X1 U18176 ( .B1(n15825), .B2(n15330), .A(n15092), .ZN(n15093) );
  AOI21_X1 U18177 ( .B1(n15094), .B2(n15097), .A(n15093), .ZN(n15095) );
  OAI211_X1 U18178 ( .C1(n15098), .C2(n15097), .A(n15096), .B(n15095), .ZN(
        n15099) );
  AOI21_X1 U18179 ( .B1(n15100), .B2(n18977), .A(n15099), .ZN(n15101) );
  OAI21_X1 U18180 ( .B1(n15102), .B2(n15309), .A(n15101), .ZN(P2_U3019) );
  INV_X1 U18181 ( .A(n15103), .ZN(n15113) );
  NAND2_X1 U18182 ( .A1(n15827), .A2(n15982), .ZN(n15111) );
  INV_X1 U18183 ( .A(n15104), .ZN(n15119) );
  XNOR2_X1 U18184 ( .A(n15118), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15108) );
  OAI21_X1 U18185 ( .B1(n15106), .B2(n15330), .A(n15105), .ZN(n15107) );
  AOI21_X1 U18186 ( .B1(n15119), .B2(n15108), .A(n15107), .ZN(n15110) );
  INV_X1 U18187 ( .A(n15130), .ZN(n15120) );
  NAND3_X1 U18188 ( .A1(n15120), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15267), .ZN(n15109) );
  NAND3_X1 U18189 ( .A1(n15111), .A2(n15110), .A3(n15109), .ZN(n15112) );
  AOI21_X1 U18190 ( .B1(n15113), .B2(n18977), .A(n15112), .ZN(n15114) );
  OAI21_X1 U18191 ( .B1(n15309), .B2(n15115), .A(n15114), .ZN(P2_U3020) );
  OAI21_X1 U18192 ( .B1(n15840), .B2(n15330), .A(n15116), .ZN(n15117) );
  AOI21_X1 U18193 ( .B1(n15119), .B2(n15118), .A(n15117), .ZN(n15122) );
  NAND3_X1 U18194 ( .A1(n15120), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15267), .ZN(n15121) );
  OAI211_X1 U18195 ( .C1(n15848), .C2(n18986), .A(n15122), .B(n15121), .ZN(
        n15123) );
  AOI21_X1 U18196 ( .B1(n15124), .B2(n18977), .A(n15123), .ZN(n15125) );
  OAI21_X1 U18197 ( .B1(n15309), .B2(n15126), .A(n15125), .ZN(P2_U3021) );
  AOI21_X1 U18198 ( .B1(n15148), .B2(n9825), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15129) );
  AOI21_X1 U18199 ( .B1(n15849), .B2(n18982), .A(n15127), .ZN(n15128) );
  OAI21_X1 U18200 ( .B1(n15130), .B2(n15129), .A(n15128), .ZN(n15133) );
  NOR2_X1 U18201 ( .A1(n15131), .A2(n15978), .ZN(n15132) );
  AOI211_X1 U18202 ( .C1(n15982), .C2(n15859), .A(n15133), .B(n15132), .ZN(
        n15134) );
  NAND2_X1 U18203 ( .A1(n15136), .A2(n18977), .ZN(n15144) );
  OAI211_X1 U18204 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15148), .B(n15137), .ZN(
        n15139) );
  OAI211_X1 U18205 ( .C1(n15865), .C2(n15330), .A(n15139), .B(n15138), .ZN(
        n15142) );
  NOR2_X1 U18206 ( .A1(n15140), .A2(n18986), .ZN(n15141) );
  AOI211_X1 U18207 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15150), .A(
        n15142), .B(n15141), .ZN(n15143) );
  OAI211_X1 U18208 ( .C1(n15145), .C2(n15309), .A(n15144), .B(n15143), .ZN(
        P2_U3023) );
  AOI21_X1 U18209 ( .B1(n15147), .B2(n9675), .A(n15146), .ZN(n15882) );
  INV_X1 U18210 ( .A(n15148), .ZN(n15153) );
  AOI21_X1 U18211 ( .B1(n15570), .B2(n18982), .A(n15149), .ZN(n15152) );
  NAND2_X1 U18212 ( .A1(n15150), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15151) );
  OAI211_X1 U18213 ( .C1(n15153), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15152), .B(n15151), .ZN(n15154) );
  AOI21_X1 U18214 ( .B1(n15882), .B2(n15982), .A(n15154), .ZN(n15157) );
  NAND2_X1 U18215 ( .A1(n15155), .A2(n11303), .ZN(n15156) );
  OAI211_X1 U18216 ( .C1(n15158), .C2(n15978), .A(n15157), .B(n15156), .ZN(
        P2_U3024) );
  OAI21_X1 U18217 ( .B1(n15221), .B2(n15159), .A(n15319), .ZN(n15166) );
  OAI21_X1 U18218 ( .B1(n15161), .B2(n15330), .A(n15160), .ZN(n15165) );
  INV_X1 U18219 ( .A(n15162), .ZN(n15201) );
  NOR2_X1 U18220 ( .A1(n15959), .A2(n15201), .ZN(n15245) );
  NAND2_X1 U18221 ( .A1(n15245), .A2(n15163), .ZN(n15189) );
  NOR3_X1 U18222 ( .A1(n15189), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15178), .ZN(n15164) );
  AOI211_X1 U18223 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15166), .A(
        n15165), .B(n15164), .ZN(n15167) );
  OAI21_X1 U18224 ( .B1(n15168), .B2(n18986), .A(n15167), .ZN(n15169) );
  AOI21_X1 U18225 ( .B1(n15170), .B2(n18977), .A(n15169), .ZN(n15171) );
  OAI21_X1 U18226 ( .B1(n15172), .B2(n15309), .A(n15171), .ZN(P2_U3025) );
  NOR2_X1 U18227 ( .A1(n15174), .A2(n15173), .ZN(n15175) );
  OR2_X1 U18228 ( .A1(n15176), .A2(n15175), .ZN(n18619) );
  NOR2_X1 U18229 ( .A1(n18619), .A2(n18986), .ZN(n15185) );
  OAI21_X1 U18230 ( .B1(n15268), .B2(n15177), .A(n15267), .ZN(n15196) );
  OAI21_X1 U18231 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15178), .ZN(n15179) );
  NOR2_X1 U18232 ( .A1(n15189), .A2(n15179), .ZN(n15180) );
  AOI211_X1 U18233 ( .C1(n18621), .C2(n18982), .A(n15181), .B(n15180), .ZN(
        n15182) );
  OAI21_X1 U18234 ( .B1(n15183), .B2(n15196), .A(n15182), .ZN(n15184) );
  AOI211_X1 U18235 ( .C1(n15186), .C2(n18977), .A(n15185), .B(n15184), .ZN(
        n15187) );
  OAI21_X1 U18236 ( .B1(n15188), .B2(n15309), .A(n15187), .ZN(P2_U3026) );
  NAND2_X1 U18237 ( .A1(n18638), .A2(n15982), .ZN(n15194) );
  INV_X1 U18238 ( .A(n18640), .ZN(n15192) );
  NOR2_X1 U18239 ( .A1(n15189), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15190) );
  AOI211_X1 U18240 ( .C1(n15192), .C2(n18982), .A(n15191), .B(n15190), .ZN(
        n15193) );
  OAI211_X1 U18241 ( .C1(n15196), .C2(n15195), .A(n15194), .B(n15193), .ZN(
        n15197) );
  AOI21_X1 U18242 ( .B1(n15198), .B2(n18977), .A(n15197), .ZN(n15199) );
  OAI21_X1 U18243 ( .B1(n15200), .B2(n15309), .A(n15199), .ZN(P2_U3027) );
  INV_X1 U18244 ( .A(n18649), .ZN(n15214) );
  OAI21_X1 U18245 ( .B1(n15268), .B2(n15201), .A(n15267), .ZN(n15251) );
  INV_X1 U18246 ( .A(n15251), .ZN(n15202) );
  AOI21_X1 U18247 ( .B1(n15203), .B2(n15204), .A(n15202), .ZN(n15210) );
  INV_X1 U18248 ( .A(n15245), .ZN(n15205) );
  NOR3_X1 U18249 ( .A1(n15205), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15204), .ZN(n15206) );
  AOI211_X1 U18250 ( .C1(n10111), .C2(n18982), .A(n15207), .B(n15206), .ZN(
        n15208) );
  OAI21_X1 U18251 ( .B1(n15210), .B2(n15209), .A(n15208), .ZN(n15213) );
  NOR2_X1 U18252 ( .A1(n15211), .A2(n15978), .ZN(n15212) );
  AOI211_X1 U18253 ( .C1(n15982), .C2(n15214), .A(n15213), .B(n15212), .ZN(
        n15215) );
  OAI21_X1 U18254 ( .B1(n15216), .B2(n15309), .A(n15215), .ZN(P2_U3028) );
  OR2_X1 U18255 ( .A1(n18977), .A2(n18973), .ZN(n15219) );
  NAND2_X1 U18256 ( .A1(n18964), .A2(n15250), .ZN(n15217) );
  NAND2_X1 U18257 ( .A1(n15251), .A2(n15217), .ZN(n15218) );
  AOI21_X1 U18258 ( .B1(n15220), .B2(n15219), .A(n15218), .ZN(n15232) );
  OAI21_X1 U18259 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15221), .A(
        n15232), .ZN(n15229) );
  AOI22_X1 U18260 ( .A1(n15223), .A2(n18977), .B1(n15222), .B2(n15245), .ZN(
        n15227) );
  AOI21_X1 U18261 ( .B1(n18656), .B2(n18982), .A(n15224), .ZN(n15226) );
  NAND2_X1 U18262 ( .A1(n18657), .A2(n15982), .ZN(n15225) );
  OAI211_X1 U18263 ( .C1(n15227), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15226), .B(n15225), .ZN(n15228) );
  AOI21_X1 U18264 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15229), .A(
        n15228), .ZN(n15230) );
  OAI21_X1 U18265 ( .B1(n15231), .B2(n15309), .A(n15230), .ZN(P2_U3029) );
  INV_X1 U18266 ( .A(n15232), .ZN(n15242) );
  AND2_X1 U18267 ( .A1(n15234), .A2(n15233), .ZN(n15236) );
  OR2_X1 U18268 ( .A1(n15236), .A2(n15235), .ZN(n18863) );
  NAND2_X1 U18269 ( .A1(n18982), .A2(n18841), .ZN(n15237) );
  OAI211_X1 U18270 ( .C1(n18863), .C2(n18986), .A(n15238), .B(n15237), .ZN(
        n15241) );
  AOI21_X1 U18271 ( .B1(n15033), .B2(n18977), .A(n15245), .ZN(n15239) );
  NOR3_X1 U18272 ( .A1(n15239), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15250), .ZN(n15240) );
  AOI211_X1 U18273 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15242), .A(
        n15241), .B(n15240), .ZN(n15243) );
  OAI21_X1 U18274 ( .B1(n15244), .B2(n15309), .A(n15243), .ZN(P2_U3030) );
  NOR2_X1 U18275 ( .A1(n18679), .A2(n18986), .ZN(n15253) );
  NAND2_X1 U18276 ( .A1(n15245), .A2(n15250), .ZN(n15249) );
  INV_X1 U18277 ( .A(n18680), .ZN(n15247) );
  NOR2_X1 U18278 ( .A1(n15042), .A2(n15891), .ZN(n15246) );
  AOI21_X1 U18279 ( .B1(n18982), .B2(n15247), .A(n15246), .ZN(n15248) );
  OAI211_X1 U18280 ( .C1(n15251), .C2(n15250), .A(n15249), .B(n15248), .ZN(
        n15252) );
  AOI211_X1 U18281 ( .C1(n15254), .C2(n18977), .A(n15253), .B(n15252), .ZN(
        n15255) );
  OAI21_X1 U18282 ( .B1(n15256), .B2(n15309), .A(n15255), .ZN(P2_U3031) );
  INV_X1 U18283 ( .A(n15257), .ZN(n15261) );
  AOI21_X1 U18284 ( .B1(n15892), .B2(n15259), .A(n15258), .ZN(n15260) );
  AOI21_X1 U18285 ( .B1(n15261), .B2(n15892), .A(n15260), .ZN(n15906) );
  INV_X1 U18286 ( .A(n15906), .ZN(n15277) );
  NAND2_X1 U18287 ( .A1(n15262), .A2(n10817), .ZN(n15264) );
  INV_X1 U18288 ( .A(n15958), .ZN(n15263) );
  NAND2_X1 U18289 ( .A1(n15313), .A2(n15263), .ZN(n15897) );
  NOR2_X1 U18290 ( .A1(n15318), .A2(n15959), .ZN(n15302) );
  NAND2_X1 U18291 ( .A1(n15266), .A2(n15302), .ZN(n15265) );
  NOR2_X1 U18292 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15265), .ZN(
        n15964) );
  NAND3_X1 U18293 ( .A1(n15266), .A2(n15302), .A3(n15972), .ZN(n15970) );
  OAI21_X1 U18294 ( .B1(n15269), .B2(n15268), .A(n15267), .ZN(n15971) );
  NAND2_X1 U18295 ( .A1(n15970), .A2(n15971), .ZN(n15963) );
  INV_X1 U18296 ( .A(n15963), .ZN(n15272) );
  INV_X1 U18297 ( .A(n18703), .ZN(n15904) );
  NOR2_X1 U18298 ( .A1(n10602), .A2(n18970), .ZN(n15270) );
  AOI21_X1 U18299 ( .B1(n18982), .B2(n15904), .A(n15270), .ZN(n15271) );
  OAI21_X1 U18300 ( .B1(n15272), .B2(n10817), .A(n15271), .ZN(n15273) );
  AOI21_X1 U18301 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15964), .A(
        n15273), .ZN(n15274) );
  OAI21_X1 U18302 ( .B1(n18702), .B2(n18986), .A(n15274), .ZN(n15275) );
  AOI21_X1 U18303 ( .B1(n15905), .B2(n18977), .A(n15275), .ZN(n15276) );
  OAI21_X1 U18304 ( .B1(n15277), .B2(n15309), .A(n15276), .ZN(P2_U3033) );
  NAND2_X1 U18305 ( .A1(n15293), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15292) );
  AOI21_X1 U18306 ( .B1(n15292), .B2(n15280), .A(n15278), .ZN(n15909) );
  INV_X1 U18307 ( .A(n15909), .ZN(n15291) );
  XNOR2_X1 U18308 ( .A(n15281), .B(n15280), .ZN(n15282) );
  XNOR2_X1 U18309 ( .A(n15279), .B(n15282), .ZN(n15911) );
  OAI21_X1 U18310 ( .B1(n9693), .B2(n15284), .A(n15283), .ZN(n18873) );
  NOR2_X1 U18311 ( .A1(n18873), .A2(n18986), .ZN(n15289) );
  OAI211_X1 U18312 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n15302), .B(n15285), .ZN(
        n15287) );
  OAI21_X1 U18313 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15959), .A(
        n15319), .ZN(n15301) );
  AOI22_X1 U18314 ( .A1(n18791), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15301), .ZN(n15286) );
  OAI211_X1 U18315 ( .C1(n15330), .C2(n18724), .A(n15287), .B(n15286), .ZN(
        n15288) );
  AOI211_X1 U18316 ( .C1(n15911), .C2(n11303), .A(n15289), .B(n15288), .ZN(
        n15290) );
  OAI21_X1 U18317 ( .B1(n15291), .B2(n15978), .A(n15290), .ZN(P2_U3035) );
  OAI21_X1 U18318 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15292), .ZN(n15917) );
  INV_X1 U18319 ( .A(n15294), .ZN(n15314) );
  OR2_X1 U18320 ( .A1(n15295), .A2(n15314), .ZN(n15299) );
  AND2_X1 U18321 ( .A1(n15297), .A2(n15296), .ZN(n15298) );
  XNOR2_X1 U18322 ( .A(n15299), .B(n15298), .ZN(n15916) );
  NOR2_X1 U18323 ( .A1(n10631), .A2(n15891), .ZN(n15300) );
  AOI221_X1 U18324 ( .B1(n15302), .B2(n10786), .C1(n15301), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15300), .ZN(n15308) );
  XNOR2_X1 U18325 ( .A(n15304), .B(n15303), .ZN(n18876) );
  INV_X1 U18326 ( .A(n18736), .ZN(n15305) );
  OAI22_X1 U18327 ( .A1(n18876), .A2(n18986), .B1(n15330), .B2(n15305), .ZN(
        n15306) );
  INV_X1 U18328 ( .A(n15306), .ZN(n15307) );
  OAI211_X1 U18329 ( .C1(n15916), .C2(n15309), .A(n15308), .B(n15307), .ZN(
        n15310) );
  INV_X1 U18330 ( .A(n15310), .ZN(n15311) );
  OAI21_X1 U18331 ( .B1(n15917), .B2(n15978), .A(n15311), .ZN(P2_U3036) );
  OAI21_X1 U18332 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15313), .A(
        n15312), .ZN(n15924) );
  NOR2_X1 U18333 ( .A1(n15315), .A2(n15314), .ZN(n15316) );
  XNOR2_X1 U18334 ( .A(n15317), .B(n15316), .ZN(n15925) );
  NOR2_X1 U18335 ( .A1(n15319), .A2(n15318), .ZN(n15325) );
  NOR2_X1 U18336 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15959), .ZN(
        n15322) );
  NOR2_X1 U18337 ( .A1(n18970), .A2(n15320), .ZN(n15321) );
  AOI211_X1 U18338 ( .C1(n18747), .C2(n18982), .A(n15322), .B(n15321), .ZN(
        n15323) );
  OAI21_X1 U18339 ( .B1(n18750), .B2(n18986), .A(n15323), .ZN(n15324) );
  AOI211_X1 U18340 ( .C1(n15925), .C2(n11303), .A(n15325), .B(n15324), .ZN(
        n15326) );
  OAI21_X1 U18341 ( .B1(n15924), .B2(n15978), .A(n15326), .ZN(P2_U3037) );
  NOR2_X1 U18342 ( .A1(n10622), .A2(n18970), .ZN(n15327) );
  AOI221_X1 U18343 ( .B1(n15983), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n15987), .C2(n15328), .A(n15327), .ZN(n15329) );
  INV_X1 U18344 ( .A(n15329), .ZN(n15332) );
  OAI22_X1 U18345 ( .A1(n18769), .A2(n15330), .B1(n18986), .B2(n18770), .ZN(
        n15331) );
  AOI211_X1 U18346 ( .C1(n15333), .C2(n11303), .A(n15332), .B(n15331), .ZN(
        n15334) );
  OAI21_X1 U18347 ( .B1(n15335), .B2(n15978), .A(n15334), .ZN(P2_U3039) );
  OAI22_X1 U18348 ( .A1(n9969), .A2(n15336), .B1(n18837), .B2(n18676), .ZN(
        n15341) );
  OAI222_X1 U18349 ( .A1(n15995), .A2(n12204), .B1(n19691), .B2(n15337), .C1(
        n10711), .C2(n15341), .ZN(n15338) );
  MUX2_X1 U18350 ( .A(n15338), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15356), .Z(P2_U3601) );
  INV_X1 U18351 ( .A(n15995), .ZN(n15345) );
  OAI21_X1 U18352 ( .B1(n9969), .B2(n15340), .A(n15339), .ZN(n15351) );
  INV_X1 U18353 ( .A(n15351), .ZN(n15344) );
  AND2_X1 U18354 ( .A1(n15341), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15350) );
  AOI222_X1 U18355 ( .A1(n19709), .A2(n15345), .B1(n15344), .B2(n15350), .C1(
        n15343), .C2(n15342), .ZN(n15347) );
  NAND2_X1 U18356 ( .A1(n15356), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15346) );
  OAI21_X1 U18357 ( .B1(n15347), .B2(n15356), .A(n15346), .ZN(P2_U3600) );
  OAI22_X1 U18358 ( .A1(n19139), .A2(n15995), .B1(n15348), .B2(n19691), .ZN(
        n15349) );
  AOI21_X1 U18359 ( .B1(n15351), .B2(n15350), .A(n15349), .ZN(n15353) );
  MUX2_X1 U18360 ( .A(n15353), .B(n15352), .S(n15356), .Z(n15354) );
  INV_X1 U18361 ( .A(n15354), .ZN(P2_U3599) );
  OAI22_X1 U18362 ( .A1(n19277), .A2(n15995), .B1(n15355), .B2(n19691), .ZN(
        n15357) );
  MUX2_X1 U18363 ( .A(n15357), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15356), .Z(P2_U3596) );
  INV_X1 U18364 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16578) );
  INV_X1 U18365 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16750) );
  INV_X1 U18366 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16807) );
  INV_X1 U18367 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16837) );
  INV_X1 U18368 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16462) );
  INV_X1 U18369 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16486) );
  NAND3_X1 U18370 ( .A1(n15359), .A2(n15358), .A3(n17036), .ZN(n15361) );
  NAND2_X1 U18371 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16933) );
  NOR2_X1 U18372 ( .A1(n16948), .A2(n16933), .ZN(n15363) );
  NAND4_X1 U18373 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .A4(n15363), .ZN(n16930) );
  NAND3_X1 U18374 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n16780), .ZN(n16736) );
  NAND3_X1 U18375 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(P3_EBX_REG_23__SCAN_IN), .ZN(n15364) );
  NAND3_X1 U18376 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(P3_EBX_REG_26__SCAN_IN), .ZN(n16684) );
  NOR3_X1 U18377 ( .A1(n16736), .A2(n15364), .A3(n16684), .ZN(n15365) );
  NAND4_X1 U18378 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n15365), .ZN(n16577) );
  NOR2_X1 U18379 ( .A1(n16578), .A2(n16577), .ZN(n16679) );
  NAND2_X1 U18380 ( .A1(n16941), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n15367) );
  NAND2_X1 U18381 ( .A1(n16679), .A2(n17036), .ZN(n15366) );
  OAI22_X1 U18382 ( .A1(n16679), .A2(n15367), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n15366), .ZN(P3_U2672) );
  AOI22_X1 U18383 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15371) );
  AOI22_X1 U18384 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16894), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15370) );
  AOI22_X1 U18385 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16635), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U18386 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15368) );
  NAND4_X1 U18387 ( .A1(n15371), .A2(n15370), .A3(n15369), .A4(n15368), .ZN(
        n15377) );
  AOI22_X1 U18388 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15375) );
  AOI22_X1 U18389 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15374) );
  AOI22_X1 U18390 ( .A1(n16810), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15373) );
  AOI22_X1 U18391 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15372) );
  NAND4_X1 U18392 ( .A1(n15375), .A2(n15374), .A3(n15373), .A4(n15372), .ZN(
        n15376) );
  NOR2_X1 U18393 ( .A1(n15377), .A2(n15376), .ZN(n17043) );
  AOI21_X1 U18394 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16865), .A(n16927), .ZN(
        n16836) );
  NOR2_X1 U18395 ( .A1(n17959), .A2(n15378), .ZN(n16853) );
  AOI22_X1 U18396 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16836), .B1(n16853), 
        .B2(n16835), .ZN(n15379) );
  OAI21_X1 U18397 ( .B1(n17043), .B2(n16941), .A(n15379), .ZN(P3_U2690) );
  NOR2_X1 U18398 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18520), .ZN(
        n17905) );
  INV_X1 U18399 ( .A(n17905), .ZN(n17966) );
  NAND2_X1 U18400 ( .A1(n15380), .A2(n10126), .ZN(n17903) );
  INV_X1 U18401 ( .A(n17903), .ZN(n15382) );
  NAND2_X1 U18402 ( .A1(n18426), .A2(n18415), .ZN(n18411) );
  NAND2_X1 U18403 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17902) );
  NOR2_X1 U18404 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18520), .ZN(
        n18543) );
  AOI21_X1 U18405 ( .B1(n18411), .B2(n17902), .A(n18543), .ZN(n17914) );
  INV_X1 U18406 ( .A(n18264), .ZN(n18119) );
  OAI211_X1 U18407 ( .C1(n18518), .C2(n15382), .A(n18119), .B(n15381), .ZN(
        n17910) );
  NAND2_X1 U18408 ( .A1(n17966), .A2(n17910), .ZN(n15385) );
  INV_X1 U18409 ( .A(n15385), .ZN(n15384) );
  INV_X1 U18410 ( .A(n18118), .ZN(n18261) );
  NAND2_X1 U18411 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17534) );
  INV_X1 U18412 ( .A(n17534), .ZN(n17474) );
  NAND2_X1 U18413 ( .A1(n18520), .A2(n17902), .ZN(n18568) );
  OAI22_X1 U18414 ( .A1(n17474), .A2(n18568), .B1(n18166), .B2(n18520), .ZN(
        n15387) );
  NAND3_X1 U18415 ( .A1(n18385), .A2(n17910), .A3(n15387), .ZN(n15383) );
  OAI221_X1 U18416 ( .B1(n18385), .B2(n15384), .C1(n18385), .C2(n18261), .A(
        n15383), .ZN(P3_U2864) );
  NAND2_X1 U18417 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18071) );
  NOR2_X1 U18418 ( .A1(n17474), .A2(n18568), .ZN(n15386) );
  AOI221_X1 U18419 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18071), .C1(n15386), 
        .C2(n18071), .A(n15385), .ZN(n17909) );
  OAI221_X1 U18420 ( .B1(n18118), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18118), .C2(n15387), .A(n17910), .ZN(n17907) );
  AOI22_X1 U18421 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17909), .B1(
        n17907), .B2(n18390), .ZN(P3_U2865) );
  INV_X1 U18422 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17588) );
  INV_X1 U18423 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U18424 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15391) );
  AOI22_X1 U18425 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15390) );
  AOI22_X1 U18426 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U18427 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15388) );
  NAND4_X1 U18428 ( .A1(n15391), .A2(n15390), .A3(n15389), .A4(n15388), .ZN(
        n15397) );
  AOI22_X1 U18429 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15395) );
  AOI22_X1 U18430 ( .A1(n16810), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15394) );
  AOI22_X1 U18431 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15393) );
  AOI22_X1 U18432 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15392) );
  NAND4_X1 U18433 ( .A1(n15395), .A2(n15394), .A3(n15393), .A4(n15392), .ZN(
        n15396) );
  AOI22_X1 U18434 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15401) );
  AOI22_X1 U18435 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15400) );
  AOI22_X1 U18436 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15399) );
  AOI22_X1 U18437 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15398) );
  NAND4_X1 U18438 ( .A1(n15401), .A2(n15400), .A3(n15399), .A4(n15398), .ZN(
        n15407) );
  AOI22_X1 U18439 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15405) );
  AOI22_X1 U18440 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U18441 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15403) );
  INV_X2 U18442 ( .A(n13758), .ZN(n16845) );
  AOI22_X1 U18443 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15402) );
  NAND4_X1 U18444 ( .A1(n15405), .A2(n15404), .A3(n15403), .A4(n15402), .ZN(
        n15406) );
  AOI22_X1 U18445 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15411) );
  AOI22_X1 U18446 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15410) );
  AOI22_X1 U18447 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15409) );
  AOI22_X1 U18448 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16894), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15408) );
  NAND4_X1 U18449 ( .A1(n15411), .A2(n15410), .A3(n15409), .A4(n15408), .ZN(
        n15417) );
  AOI22_X1 U18450 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15415) );
  AOI22_X1 U18451 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U18452 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U18453 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15412) );
  NAND4_X1 U18454 ( .A1(n15415), .A2(n15414), .A3(n15413), .A4(n15412), .ZN(
        n15416) );
  INV_X1 U18455 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20735) );
  AOI22_X1 U18456 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n16889), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n15418), .ZN(n15419) );
  OAI21_X1 U18457 ( .B1(n20735), .B2(n9639), .A(n15419), .ZN(n15420) );
  INV_X1 U18458 ( .A(n15420), .ZN(n15431) );
  AOI22_X1 U18459 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16781), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n16870), .ZN(n15421) );
  INV_X1 U18460 ( .A(n15421), .ZN(n15422) );
  AOI22_X1 U18461 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16894), .B1(
        n16635), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15429) );
  AOI22_X1 U18462 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U18463 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15435), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15427) );
  AOI22_X1 U18464 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n16886), .ZN(n15426) );
  AOI22_X1 U18465 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n16845), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15425) );
  AOI22_X1 U18466 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15444) );
  INV_X1 U18467 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n20722) );
  AOI22_X1 U18468 ( .A1(n15432), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15434) );
  OAI211_X1 U18469 ( .C1(n9596), .C2(n20722), .A(n15434), .B(n15433), .ZN(
        n15442) );
  AOI22_X1 U18471 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15440) );
  AOI22_X1 U18472 ( .A1(n15436), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15438) );
  AOI22_X1 U18473 ( .A1(n16894), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15468), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15437) );
  NAND4_X1 U18474 ( .A1(n15440), .A2(n15439), .A3(n15438), .A4(n15437), .ZN(
        n15441) );
  AOI211_X1 U18475 ( .C1(n9605), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n15442), .B(n15441), .ZN(n15443) );
  NAND2_X1 U18476 ( .A1(n17092), .A2(n15546), .ZN(n15484) );
  NOR2_X2 U18477 ( .A1(n17082), .A2(n15484), .ZN(n15487) );
  AOI22_X1 U18478 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16810), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U18479 ( .A1(n16888), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15454) );
  INV_X1 U18480 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n20698) );
  AOI22_X1 U18481 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15445) );
  OAI21_X1 U18482 ( .B1(n13827), .B2(n20698), .A(n15445), .ZN(n15452) );
  AOI22_X1 U18483 ( .A1(n15446), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15450) );
  AOI22_X1 U18484 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15449) );
  AOI22_X1 U18485 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U18486 ( .A1(n16845), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15447) );
  NAND4_X1 U18487 ( .A1(n15450), .A2(n15449), .A3(n15448), .A4(n15447), .ZN(
        n15451) );
  AOI211_X1 U18488 ( .C1(n16825), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n15452), .B(n15451), .ZN(n15453) );
  NAND3_X1 U18489 ( .A1(n15455), .A2(n15454), .A3(n15453), .ZN(n15537) );
  NAND2_X1 U18490 ( .A1(n15487), .A2(n15537), .ZN(n15490) );
  AOI22_X1 U18491 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15465) );
  AOI22_X1 U18492 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15464) );
  INV_X1 U18493 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17954) );
  AOI22_X1 U18494 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15456) );
  OAI21_X1 U18495 ( .B1(n9644), .B2(n17954), .A(n15456), .ZN(n15462) );
  AOI22_X1 U18496 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15460) );
  AOI22_X1 U18497 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U18498 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16894), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15458) );
  AOI22_X1 U18499 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15457) );
  NAND4_X1 U18500 ( .A1(n15460), .A2(n15459), .A3(n15458), .A4(n15457), .ZN(
        n15461) );
  AOI211_X1 U18501 ( .C1(n16905), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n15462), .B(n15461), .ZN(n15463) );
  NAND3_X1 U18502 ( .A1(n15465), .A2(n15464), .A3(n15463), .ZN(n15538) );
  INV_X1 U18503 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17782) );
  NOR2_X1 U18504 ( .A1(n17800), .A2(n17782), .ZN(n17767) );
  NAND2_X1 U18505 ( .A1(n17767), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17753) );
  NOR2_X1 U18506 ( .A1(n17753), .A2(n17758), .ZN(n17410) );
  NAND2_X1 U18507 ( .A1(n17410), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17731) );
  INV_X1 U18508 ( .A(n17731), .ZN(n17725) );
  NAND2_X1 U18509 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17725), .ZN(
        n17712) );
  AOI21_X1 U18510 ( .B1(n17068), .B2(n16072), .A(n17312), .ZN(n15498) );
  INV_X1 U18511 ( .A(n15538), .ZN(n17071) );
  XNOR2_X1 U18512 ( .A(n17071), .B(n15466), .ZN(n15495) );
  NAND2_X1 U18513 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15495), .ZN(
        n15496) );
  NAND2_X1 U18514 ( .A1(n15536), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15480) );
  AOI22_X1 U18515 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16894), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U18516 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U18517 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U18518 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15469) );
  NAND4_X1 U18519 ( .A1(n15472), .A2(n15471), .A3(n15470), .A4(n15469), .ZN(
        n15479) );
  AOI22_X1 U18520 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U18521 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15476) );
  AOI22_X1 U18522 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15475) );
  AOI22_X1 U18523 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15474) );
  NAND4_X1 U18524 ( .A1(n15477), .A2(n15476), .A3(n15475), .A4(n15474), .ZN(
        n15478) );
  NOR2_X1 U18525 ( .A1(n15479), .A2(n15478), .ZN(n17572) );
  INV_X1 U18526 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18546) );
  NOR2_X1 U18527 ( .A1(n17572), .A2(n18546), .ZN(n17571) );
  NAND2_X1 U18528 ( .A1(n15480), .A2(n17562), .ZN(n17554) );
  INV_X1 U18529 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17879) );
  XOR2_X1 U18530 ( .A(n17082), .B(n15484), .Z(n17543) );
  INV_X1 U18531 ( .A(n15537), .ZN(n17078) );
  XNOR2_X1 U18532 ( .A(n17078), .B(n15487), .ZN(n15488) );
  XNOR2_X1 U18533 ( .A(n20762), .B(n15488), .ZN(n17527) );
  NAND2_X1 U18534 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15488), .ZN(
        n15489) );
  XOR2_X1 U18535 ( .A(n17075), .B(n15490), .Z(n15493) );
  INV_X1 U18536 ( .A(n15493), .ZN(n15491) );
  NAND2_X1 U18537 ( .A1(n15493), .A2(n15492), .ZN(n15494) );
  INV_X1 U18538 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17836) );
  XNOR2_X1 U18539 ( .A(n17836), .B(n15495), .ZN(n17505) );
  NAND2_X1 U18540 ( .A1(n15498), .A2(n15497), .ZN(n15499) );
  INV_X1 U18541 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17442) );
  INV_X1 U18542 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20690) );
  NAND2_X1 U18543 ( .A1(n17404), .A2(n20690), .ZN(n17389) );
  INV_X1 U18544 ( .A(n15500), .ZN(n15501) );
  NOR2_X2 U18545 ( .A1(n15501), .A2(n17710), .ZN(n17369) );
  INV_X1 U18546 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17685) );
  NOR2_X1 U18547 ( .A1(n17704), .A2(n17685), .ZN(n17680) );
  NAND2_X1 U18548 ( .A1(n17680), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17635) );
  INV_X1 U18549 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17318) );
  NAND2_X1 U18550 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17651) );
  NOR2_X1 U18551 ( .A1(n17318), .A2(n17651), .ZN(n17642) );
  NAND2_X1 U18552 ( .A1(n17642), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15506) );
  NOR2_X1 U18553 ( .A1(n17635), .A2(n15506), .ZN(n17627) );
  NAND2_X1 U18554 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17627), .ZN(
        n17614) );
  INV_X1 U18555 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17357) );
  NAND2_X1 U18556 ( .A1(n17357), .A2(n17483), .ZN(n17352) );
  NOR2_X1 U18557 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17352), .ZN(
        n15502) );
  INV_X1 U18558 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17331) );
  NAND2_X1 U18559 ( .A1(n15502), .A2(n17331), .ZN(n17313) );
  NOR2_X1 U18560 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17313), .ZN(
        n17295) );
  INV_X1 U18561 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20685) );
  INV_X1 U18562 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17643) );
  NAND3_X1 U18563 ( .A1(n17295), .A2(n20685), .A3(n17643), .ZN(n15503) );
  INV_X1 U18564 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17620) );
  MUX2_X1 U18565 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17266), .S(
        n17483), .Z(n15508) );
  INV_X1 U18566 ( .A(n17680), .ZN(n17682) );
  NOR2_X1 U18567 ( .A1(n17369), .A2(n17682), .ZN(n17311) );
  NOR2_X2 U18568 ( .A1(n17327), .A2(n17311), .ZN(n17353) );
  NAND2_X1 U18569 ( .A1(n15509), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15507) );
  INV_X1 U18570 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17253) );
  NAND2_X1 U18571 ( .A1(n17312), .A2(n15509), .ZN(n17265) );
  NOR2_X1 U18572 ( .A1(n17599), .A2(n17253), .ZN(n17579) );
  INV_X1 U18573 ( .A(n16071), .ZN(n17232) );
  NAND2_X1 U18574 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17312), .ZN(
        n15511) );
  NOR2_X1 U18575 ( .A1(n15616), .A2(n15617), .ZN(n15512) );
  INV_X1 U18576 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16037) );
  XNOR2_X1 U18577 ( .A(n15512), .B(n16037), .ZN(n16052) );
  INV_X1 U18578 ( .A(n15514), .ZN(n15515) );
  NOR2_X1 U18579 ( .A1(n15516), .A2(n15515), .ZN(n18588) );
  NOR2_X1 U18580 ( .A1(n18576), .A2(n15518), .ZN(n15520) );
  AOI21_X1 U18581 ( .B1(n15520), .B2(n18401), .A(n15519), .ZN(n18356) );
  XNOR2_X1 U18582 ( .A(n18576), .B(n17927), .ZN(n15525) );
  INV_X1 U18583 ( .A(n15521), .ZN(n15522) );
  OAI21_X1 U18584 ( .B1(n15523), .B2(n15522), .A(n16171), .ZN(n18560) );
  INV_X1 U18585 ( .A(n18560), .ZN(n15524) );
  NAND4_X1 U18586 ( .A1(n15524), .A2(n17927), .A3(n17922), .A4(n17950), .ZN(
        n15527) );
  AOI21_X1 U18587 ( .B1(n15525), .B2(n18574), .A(n18571), .ZN(n16175) );
  NAND3_X1 U18588 ( .A1(n16171), .A2(n16175), .A3(n15528), .ZN(n15526) );
  OAI211_X1 U18589 ( .C1(n18562), .C2(n15528), .A(n15527), .B(n15526), .ZN(
        n15529) );
  NAND2_X1 U18590 ( .A1(n18415), .A2(n18545), .ZN(n18587) );
  OR2_X2 U18591 ( .A1(n18587), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n17894) );
  NAND2_X1 U18592 ( .A1(n17894), .A2(n17886), .ZN(n17880) );
  NOR3_X1 U18593 ( .A1(n17601), .A2(n17599), .A3(n17253), .ZN(n16067) );
  NAND2_X1 U18594 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17802) );
  NOR2_X1 U18595 ( .A1(n17811), .A2(n17802), .ZN(n17687) );
  INV_X1 U18596 ( .A(n17687), .ZN(n15531) );
  INV_X1 U18597 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17840) );
  NOR3_X1 U18598 ( .A1(n17840), .A2(n15483), .A3(n20762), .ZN(n15532) );
  NOR2_X1 U18599 ( .A1(n17879), .A2(n15467), .ZN(n17847) );
  NAND2_X1 U18600 ( .A1(n15532), .A2(n17847), .ZN(n17804) );
  NOR2_X1 U18601 ( .A1(n15531), .A2(n17804), .ZN(n17724) );
  NAND2_X1 U18602 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17724), .ZN(
        n17790) );
  NOR2_X1 U18603 ( .A1(n17689), .A2(n17790), .ZN(n17700) );
  NAND3_X1 U18604 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16067), .A3(
        n17700), .ZN(n15534) );
  NAND2_X1 U18605 ( .A1(n17370), .A2(n17724), .ZN(n17678) );
  INV_X1 U18606 ( .A(n17678), .ZN(n15565) );
  AOI21_X1 U18607 ( .B1(n16067), .B2(n15565), .A(n18380), .ZN(n15533) );
  AOI21_X1 U18608 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17869) );
  INV_X1 U18609 ( .A(n15532), .ZN(n17686) );
  NOR2_X1 U18610 ( .A1(n17869), .A2(n17686), .ZN(n17806) );
  NAND2_X1 U18611 ( .A1(n17806), .A2(n17687), .ZN(n17726) );
  NOR2_X1 U18612 ( .A1(n17689), .A2(n17726), .ZN(n17679) );
  AOI21_X1 U18613 ( .B1(n17679), .B2(n16067), .A(n18374), .ZN(n17581) );
  AOI211_X1 U18614 ( .C1(n18378), .C2(n15534), .A(n15533), .B(n17581), .ZN(
        n15619) );
  INV_X1 U18615 ( .A(n15619), .ZN(n15535) );
  AOI211_X1 U18616 ( .C1(n17780), .C2(n17588), .A(n17888), .B(n15535), .ZN(
        n16076) );
  NAND2_X1 U18617 ( .A1(n17068), .A2(n17834), .ZN(n17740) );
  INV_X1 U18618 ( .A(n17740), .ZN(n17816) );
  NAND2_X1 U18619 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16048) );
  NOR2_X1 U18620 ( .A1(n16048), .A2(n16037), .ZN(n16005) );
  NAND2_X1 U18621 ( .A1(n17579), .A2(n17264), .ZN(n17225) );
  INV_X1 U18622 ( .A(n17225), .ZN(n17584) );
  NAND2_X1 U18623 ( .A1(n16005), .A2(n17584), .ZN(n16028) );
  NOR2_X1 U18624 ( .A1(n17572), .A2(n15536), .ZN(n15547) );
  NOR2_X1 U18625 ( .A1(n15547), .A2(n15546), .ZN(n15544) );
  NOR2_X1 U18626 ( .A1(n15544), .A2(n17082), .ZN(n15543) );
  NAND2_X1 U18627 ( .A1(n15543), .A2(n15537), .ZN(n15541) );
  NOR2_X1 U18628 ( .A1(n17075), .A2(n15541), .ZN(n15540) );
  NAND2_X1 U18629 ( .A1(n15540), .A2(n15538), .ZN(n15539) );
  NOR2_X1 U18630 ( .A1(n17068), .A2(n15539), .ZN(n15562) );
  INV_X1 U18631 ( .A(n17068), .ZN(n16074) );
  XNOR2_X1 U18632 ( .A(n15539), .B(n16074), .ZN(n17496) );
  XNOR2_X1 U18633 ( .A(n15540), .B(n17071), .ZN(n15555) );
  XOR2_X1 U18634 ( .A(n15541), .B(n17075), .Z(n15542) );
  NAND2_X1 U18635 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15542), .ZN(
        n15554) );
  XNOR2_X1 U18636 ( .A(n17840), .B(n15542), .ZN(n17519) );
  XNOR2_X1 U18637 ( .A(n15543), .B(n17078), .ZN(n17529) );
  XOR2_X1 U18638 ( .A(n17082), .B(n15544), .Z(n15545) );
  NAND2_X1 U18639 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15545), .ZN(
        n15552) );
  XNOR2_X1 U18640 ( .A(n15483), .B(n15545), .ZN(n17541) );
  INV_X1 U18641 ( .A(n15546), .ZN(n17087) );
  XNOR2_X1 U18642 ( .A(n15547), .B(n17087), .ZN(n15550) );
  OR2_X1 U18643 ( .A1(n17879), .A2(n15550), .ZN(n15551) );
  INV_X1 U18644 ( .A(n17572), .ZN(n15636) );
  AOI21_X1 U18645 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17092), .A(
        n15636), .ZN(n15549) );
  NOR2_X1 U18646 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17092), .ZN(
        n15548) );
  AOI221_X1 U18647 ( .B1(n15636), .B2(n17092), .C1(n15549), .C2(n18546), .A(
        n15548), .ZN(n17552) );
  XNOR2_X1 U18648 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15550), .ZN(
        n17551) );
  NAND2_X1 U18649 ( .A1(n17552), .A2(n17551), .ZN(n17550) );
  NAND2_X1 U18650 ( .A1(n15551), .A2(n17550), .ZN(n17540) );
  NAND2_X1 U18651 ( .A1(n17541), .A2(n17540), .ZN(n17539) );
  NAND2_X1 U18652 ( .A1(n15552), .A2(n17539), .ZN(n17530) );
  NAND2_X1 U18653 ( .A1(n17529), .A2(n17530), .ZN(n17528) );
  NOR2_X1 U18654 ( .A1(n17529), .A2(n17530), .ZN(n15553) );
  AOI21_X1 U18655 ( .B1(n20762), .B2(n17528), .A(n15553), .ZN(n17518) );
  NAND2_X1 U18656 ( .A1(n17519), .A2(n17518), .ZN(n17517) );
  NAND2_X1 U18657 ( .A1(n15554), .A2(n17517), .ZN(n15556) );
  NAND2_X1 U18658 ( .A1(n15555), .A2(n15556), .ZN(n15557) );
  XOR2_X1 U18659 ( .A(n15556), .B(n15555), .Z(n17502) );
  NAND2_X1 U18660 ( .A1(n17502), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17501) );
  NAND2_X1 U18661 ( .A1(n15557), .A2(n17501), .ZN(n17495) );
  NOR2_X1 U18662 ( .A1(n17496), .A2(n17495), .ZN(n17494) );
  INV_X1 U18663 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17807) );
  NOR2_X1 U18664 ( .A1(n17494), .A2(n17807), .ZN(n15558) );
  NAND2_X1 U18665 ( .A1(n15562), .A2(n15558), .ZN(n15563) );
  INV_X1 U18666 ( .A(n15558), .ZN(n15561) );
  NAND2_X1 U18667 ( .A1(n17496), .A2(n17495), .ZN(n15560) );
  NAND2_X1 U18668 ( .A1(n15562), .A2(n15561), .ZN(n15559) );
  OAI211_X1 U18669 ( .C1(n15562), .C2(n15561), .A(n15560), .B(n15559), .ZN(
        n17471) );
  NAND2_X1 U18670 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17471), .ZN(
        n17470) );
  NAND2_X1 U18671 ( .A1(n17255), .A2(n17579), .ZN(n17582) );
  INV_X1 U18672 ( .A(n16005), .ZN(n16053) );
  NOR2_X1 U18673 ( .A1(n17582), .A2(n16053), .ZN(n16029) );
  INV_X1 U18674 ( .A(n16029), .ZN(n16049) );
  AOI22_X1 U18675 ( .A1(n17816), .A2(n16028), .B1(n17885), .B2(n16049), .ZN(
        n15621) );
  NOR2_X1 U18676 ( .A1(n17703), .A2(n17886), .ZN(n16055) );
  INV_X1 U18677 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16068) );
  NAND2_X1 U18678 ( .A1(n16055), .A2(n16068), .ZN(n15564) );
  OAI211_X1 U18679 ( .C1(n17896), .C2(n16076), .A(n15621), .B(n15564), .ZN(
        n15568) );
  INV_X1 U18680 ( .A(n18378), .ZN(n17773) );
  OAI21_X1 U18681 ( .B1(n17773), .B2(n18546), .A(n18380), .ZN(n17864) );
  AOI22_X1 U18682 ( .A1(n18404), .A2(n17679), .B1(n15565), .B2(n17864), .ZN(
        n17600) );
  NAND2_X1 U18683 ( .A1(n17892), .A2(n16067), .ZN(n17585) );
  NOR2_X1 U18684 ( .A1(n17600), .A2(n17585), .ZN(n16059) );
  OAI22_X1 U18685 ( .A1(n17582), .A2(n17900), .B1(n17225), .B2(n17740), .ZN(
        n15566) );
  NOR2_X1 U18686 ( .A1(n16059), .A2(n15566), .ZN(n15624) );
  OAI21_X1 U18687 ( .B1(n16048), .B2(n15624), .A(n16037), .ZN(n15567) );
  OAI21_X1 U18688 ( .B1(n16037), .B2(n15568), .A(n15567), .ZN(n15569) );
  NAND2_X1 U18689 ( .A1(n17896), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16043) );
  OAI211_X1 U18690 ( .C1(n16052), .C2(n17788), .A(n15569), .B(n16043), .ZN(
        P3_U2833) );
  AOI22_X1 U18691 ( .A1(n15570), .A2(n18831), .B1(n15882), .B2(n18759), .ZN(
        n15579) );
  AOI211_X1 U18692 ( .C1(n15573), .C2(n15572), .A(n15571), .B(n18811), .ZN(
        n15577) );
  AOI22_X1 U18693 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18802), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18807), .ZN(n15574) );
  OAI21_X1 U18694 ( .B1(n15575), .B2(n18822), .A(n15574), .ZN(n15576) );
  AOI211_X1 U18695 ( .C1(P2_EBX_REG_22__SCAN_IN), .C2(n18803), .A(n15577), .B(
        n15576), .ZN(n15578) );
  NAND2_X1 U18696 ( .A1(n15579), .A2(n15578), .ZN(P2_U2833) );
  NOR3_X1 U18697 ( .A1(n15581), .A2(n15580), .A3(n20397), .ZN(n15583) );
  NAND2_X1 U18698 ( .A1(n15583), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15587) );
  INV_X1 U18699 ( .A(n15582), .ZN(n15584) );
  OAI22_X1 U18700 ( .A1(n15585), .A2(n15584), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15583), .ZN(n15586) );
  NAND2_X1 U18701 ( .A1(n15587), .A2(n15586), .ZN(n15590) );
  INV_X1 U18702 ( .A(n15588), .ZN(n15589) );
  AOI222_X1 U18703 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15590), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15589), .C1(n15590), 
        .C2(n15589), .ZN(n15591) );
  AOI222_X1 U18704 ( .A1(n20276), .A2(n15592), .B1(n20276), .B2(n15591), .C1(
        n15592), .C2(n15591), .ZN(n15601) );
  AOI21_X1 U18705 ( .B1(n19749), .B2(n15594), .A(n15593), .ZN(n15596) );
  NOR4_X1 U18706 ( .A1(n15598), .A2(n15597), .A3(n15596), .A4(n15595), .ZN(
        n15599) );
  OAI211_X1 U18707 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15601), .A(
        n15600), .B(n15599), .ZN(n15610) );
  NAND2_X1 U18708 ( .A1(n15603), .A2(n15602), .ZN(n15604) );
  AOI21_X1 U18709 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATE2_REG_1__SCAN_IN), .A(n11609), .ZN(n20529) );
  NAND2_X1 U18710 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20623), .ZN(n15777) );
  OAI211_X1 U18711 ( .C1(n15605), .C2(n15604), .A(n20529), .B(n15777), .ZN(
        n15780) );
  AOI221_X1 U18712 ( .B1(n15614), .B2(n15606), .C1(n15610), .C2(n15606), .A(
        n15780), .ZN(n15615) );
  NOR2_X1 U18713 ( .A1(n20626), .A2(n20609), .ZN(n15613) );
  INV_X1 U18714 ( .A(n15777), .ZN(n15608) );
  OAI21_X1 U18715 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20631), .A(n11609), 
        .ZN(n15778) );
  NOR2_X1 U18716 ( .A1(n15615), .A2(n15614), .ZN(n15783) );
  OAI211_X1 U18717 ( .C1(n15608), .C2(n15778), .A(n15783), .B(n15607), .ZN(
        n15609) );
  AOI21_X1 U18718 ( .B1(n15611), .B2(n15610), .A(n15609), .ZN(n15612) );
  AOI221_X1 U18719 ( .B1(n15615), .B2(n15614), .C1(n15613), .C2(n15614), .A(
        n15612), .ZN(P1_U3161) );
  INV_X1 U18720 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16054) );
  NAND2_X1 U18721 ( .A1(n16005), .A2(n16054), .ZN(n16034) );
  NAND2_X1 U18722 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15616), .ZN(
        n16017) );
  NAND2_X1 U18723 ( .A1(n15617), .A2(n16037), .ZN(n16015) );
  NAND2_X1 U18724 ( .A1(n16017), .A2(n16015), .ZN(n15618) );
  XNOR2_X1 U18725 ( .A(n15618), .B(n16054), .ZN(n16030) );
  OAI21_X1 U18726 ( .B1(n15619), .B2(n17886), .A(n17880), .ZN(n15620) );
  AOI21_X1 U18727 ( .B1(n16055), .B2(n16053), .A(n15620), .ZN(n16056) );
  AOI21_X1 U18728 ( .B1(n16056), .B2(n15621), .A(n16054), .ZN(n15622) );
  AOI21_X1 U18729 ( .B1(n17814), .B2(n16030), .A(n15622), .ZN(n15623) );
  NAND2_X1 U18730 ( .A1(n17896), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16024) );
  OAI211_X1 U18731 ( .C1(n15624), .C2(n16034), .A(n15623), .B(n16024), .ZN(
        P3_U2832) );
  NAND2_X1 U18732 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20537) );
  INV_X1 U18733 ( .A(n20537), .ZN(n15625) );
  INV_X1 U18734 ( .A(HOLD), .ZN(n19627) );
  NOR2_X1 U18735 ( .A1(n20532), .A2(n19627), .ZN(n20531) );
  NAND2_X1 U18736 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n20534) );
  OAI21_X1 U18737 ( .B1(n15625), .B2(n20531), .A(n20534), .ZN(n15626) );
  OAI211_X1 U18738 ( .C1(n20623), .C2(n20532), .A(n15627), .B(n15626), .ZN(
        P1_U3195) );
  INV_X1 U18739 ( .A(n19882), .ZN(n19862) );
  INV_X1 U18740 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16165) );
  NOR2_X1 U18741 ( .A1(n19862), .A2(n16165), .ZN(P1_U2905) );
  OR2_X1 U18742 ( .A1(n15628), .A2(n10711), .ZN(n15630) );
  AND2_X1 U18743 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19705) );
  AOI21_X1 U18744 ( .B1(n19705), .B2(n18596), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15629) );
  AOI21_X1 U18745 ( .B1(n15630), .B2(n15629), .A(n15632), .ZN(P2_U3178) );
  INV_X1 U18746 ( .A(n15631), .ZN(n19729) );
  INV_X1 U18747 ( .A(n19721), .ZN(n19718) );
  NOR2_X1 U18748 ( .A1(n20684), .A2(n19718), .ZN(P2_U3047) );
  NAND3_X1 U18749 ( .A1(n17916), .A2(n18576), .A3(n15633), .ZN(n15634) );
  NAND2_X1 U18750 ( .A1(n17036), .A2(n16950), .ZN(n17095) );
  NAND2_X2 U18751 ( .A1(n16950), .A2(n17959), .ZN(n17086) );
  AOI22_X1 U18752 ( .A1(n17094), .A2(BUF2_REG_0__SCAN_IN), .B1(n17093), .B2(
        n15636), .ZN(n15637) );
  OAI221_X1 U18753 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17095), .C1(n17163), 
        .C2(n16950), .A(n15637), .ZN(P3_U2735) );
  AOI22_X1 U18754 ( .A1(n15639), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n19832), 
        .B2(n15638), .ZN(n15647) );
  NAND2_X1 U18755 ( .A1(n19822), .A2(n15640), .ZN(n15642) );
  AOI21_X1 U18756 ( .B1(n19834), .B2(P1_EBX_REG_15__SCAN_IN), .A(n19819), .ZN(
        n15641) );
  OAI211_X1 U18757 ( .C1(n15643), .C2(n19782), .A(n15642), .B(n15641), .ZN(
        n15644) );
  AOI21_X1 U18758 ( .B1(n15645), .B2(n19796), .A(n15644), .ZN(n15646) );
  OAI211_X1 U18759 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15648), .A(n15647), 
        .B(n15646), .ZN(P1_U2825) );
  OAI21_X1 U18760 ( .B1(n15650), .B2(n15649), .A(n19801), .ZN(n15669) );
  AOI22_X1 U18761 ( .A1(n19832), .A2(n15651), .B1(n19834), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15652) );
  OAI211_X1 U18762 ( .C1(n19782), .C2(n11775), .A(n15652), .B(n19921), .ZN(
        n15656) );
  OAI22_X1 U18763 ( .A1(n15654), .A2(n19771), .B1(P1_REIP_REG_13__SCAN_IN), 
        .B2(n15653), .ZN(n15655) );
  AOI211_X1 U18764 ( .C1(n15657), .C2(n19822), .A(n15656), .B(n15655), .ZN(
        n15658) );
  OAI21_X1 U18765 ( .B1(n15669), .B2(n20567), .A(n15658), .ZN(P1_U2827) );
  AOI21_X1 U18766 ( .B1(n15659), .B2(P1_REIP_REG_11__SCAN_IN), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15668) );
  INV_X1 U18767 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15661) );
  OAI22_X1 U18768 ( .A1(n19782), .A2(n15661), .B1(n15660), .B2(n19790), .ZN(
        n15662) );
  AOI211_X1 U18769 ( .C1(n19832), .C2(n15734), .A(n19819), .B(n15662), .ZN(
        n15667) );
  NOR2_X1 U18770 ( .A1(n19843), .A2(n15663), .ZN(n15664) );
  AOI21_X1 U18771 ( .B1(n15665), .B2(n19796), .A(n15664), .ZN(n15666) );
  OAI211_X1 U18772 ( .C1(n15669), .C2(n15668), .A(n15667), .B(n15666), .ZN(
        P1_U2828) );
  NAND2_X1 U18773 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20561), .ZN(n15679) );
  OAI21_X1 U18774 ( .B1(n19790), .B2(n13591), .A(n19921), .ZN(n15670) );
  INV_X1 U18775 ( .A(n15670), .ZN(n15673) );
  AOI22_X1 U18776 ( .A1(n19832), .A2(n15671), .B1(n19830), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15672) );
  OAI211_X1 U18777 ( .C1(n15674), .C2(n20561), .A(n15673), .B(n15672), .ZN(
        n15675) );
  INV_X1 U18778 ( .A(n15675), .ZN(n15678) );
  INV_X1 U18779 ( .A(n15676), .ZN(n15682) );
  AOI22_X1 U18780 ( .A1(n15682), .A2(n19796), .B1(n19822), .B2(n15680), .ZN(
        n15677) );
  OAI211_X1 U18781 ( .C1(n19776), .C2(n15679), .A(n15678), .B(n15677), .ZN(
        P1_U2830) );
  AOI22_X1 U18782 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15684) );
  AOI22_X1 U18783 ( .A1(n15682), .A2(n15693), .B1(n15681), .B2(n15680), .ZN(
        n15683) );
  OAI211_X1 U18784 ( .C1(n19748), .C2(n15685), .A(n15684), .B(n15683), .ZN(
        P1_U2989) );
  AOI22_X1 U18785 ( .A1(n15686), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n15772), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15695) );
  INV_X1 U18786 ( .A(n15687), .ZN(n15689) );
  NAND2_X1 U18787 ( .A1(n15689), .A2(n15688), .ZN(n15690) );
  XNOR2_X1 U18788 ( .A(n15691), .B(n15690), .ZN(n15763) );
  AOI22_X1 U18789 ( .A1(n19847), .A2(n15693), .B1(n15763), .B2(n15692), .ZN(
        n15694) );
  OAI211_X1 U18790 ( .C1(n15696), .C2(n19787), .A(n15695), .B(n15694), .ZN(
        P1_U2992) );
  NOR2_X1 U18791 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15697), .ZN(
        n15699) );
  AOI22_X1 U18792 ( .A1(n15772), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n15699), 
        .B2(n15698), .ZN(n15704) );
  INV_X1 U18793 ( .A(n15700), .ZN(n15702) );
  AOI22_X1 U18794 ( .A1(n15702), .A2(n19913), .B1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15701), .ZN(n15703) );
  OAI211_X1 U18795 ( .C1(n15775), .C2(n15705), .A(n15704), .B(n15703), .ZN(
        P1_U3013) );
  NOR2_X1 U18796 ( .A1(n15707), .A2(n15706), .ZN(n15712) );
  OAI22_X1 U18797 ( .A1(n15709), .A2(n14704), .B1(n15775), .B2(n15708), .ZN(
        n15710) );
  AOI21_X1 U18798 ( .B1(n15712), .B2(n15711), .A(n15710), .ZN(n15714) );
  NAND2_X1 U18799 ( .A1(n15772), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15713) );
  OAI211_X1 U18800 ( .C1(n15716), .C2(n15715), .A(n15714), .B(n15713), .ZN(
        P1_U3015) );
  INV_X1 U18801 ( .A(n15717), .ZN(n15719) );
  AOI22_X1 U18802 ( .A1(n15719), .A2(n19913), .B1(n19911), .B2(n15718), .ZN(
        n15728) );
  NAND2_X1 U18803 ( .A1(n15772), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15727) );
  OAI21_X1 U18804 ( .B1(n15721), .B2(n15720), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15726) );
  NAND3_X1 U18805 ( .A1(n15724), .A2(n15723), .A3(n15722), .ZN(n15725) );
  NAND4_X1 U18806 ( .A1(n15728), .A2(n15727), .A3(n15726), .A4(n15725), .ZN(
        P1_U3017) );
  NAND2_X1 U18807 ( .A1(n15771), .A2(n15729), .ZN(n15744) );
  AND2_X1 U18808 ( .A1(n15772), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15733) );
  NOR3_X1 U18809 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15731), .A3(
        n15730), .ZN(n15732) );
  AOI211_X1 U18810 ( .C1(n19911), .C2(n15734), .A(n15733), .B(n15732), .ZN(
        n15743) );
  AOI221_X1 U18811 ( .B1(n15737), .B2(n15736), .C1(n15745), .C2(n15736), .A(
        n15735), .ZN(n15738) );
  OAI21_X1 U18812 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(n15749) );
  AOI22_X1 U18813 ( .A1(n15741), .A2(n19913), .B1(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15749), .ZN(n15742) );
  OAI211_X1 U18814 ( .C1(n15745), .C2(n15744), .A(n15743), .B(n15742), .ZN(
        P1_U3019) );
  NAND2_X1 U18815 ( .A1(n15747), .A2(n15746), .ZN(n15753) );
  AOI22_X1 U18816 ( .A1(n15772), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n19911), 
        .B2(n15748), .ZN(n15752) );
  AOI22_X1 U18817 ( .A1(n15750), .A2(n19913), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15749), .ZN(n15751) );
  OAI211_X1 U18818 ( .C1(n15754), .C2(n15753), .A(n15752), .B(n15751), .ZN(
        P1_U3020) );
  AOI22_X1 U18819 ( .A1(n15772), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n19911), 
        .B2(n19765), .ZN(n15758) );
  AOI22_X1 U18820 ( .A1(n15756), .A2(n19913), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15755), .ZN(n15757) );
  OAI211_X1 U18821 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15759), .A(
        n15758), .B(n15757), .ZN(P1_U3022) );
  AOI21_X1 U18822 ( .B1(n15761), .B2(n15760), .A(n9648), .ZN(n19844) );
  AOI22_X1 U18823 ( .A1(n15772), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n19911), 
        .B2(n19844), .ZN(n15765) );
  AOI22_X1 U18824 ( .A1(n15763), .A2(n19913), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15762), .ZN(n15764) );
  OAI211_X1 U18825 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n15766), .A(
        n15765), .B(n15764), .ZN(P1_U3024) );
  OAI22_X1 U18826 ( .A1(n15768), .A2(n14704), .B1(n15767), .B2(n15770), .ZN(
        n15769) );
  AOI21_X1 U18827 ( .B1(n15771), .B2(n15770), .A(n15769), .ZN(n15774) );
  NAND2_X1 U18828 ( .A1(n15772), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n15773) );
  OAI211_X1 U18829 ( .C1(n15775), .C2(n19792), .A(n15774), .B(n15773), .ZN(
        P1_U3025) );
  NAND2_X1 U18830 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11609), .ZN(n19744) );
  OAI21_X1 U18831 ( .B1(n15777), .B2(n19744), .A(n15776), .ZN(n20528) );
  AOI21_X1 U18832 ( .B1(n15783), .B2(n15778), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n15779) );
  AOI221_X1 U18833 ( .B1(n15781), .B2(n15780), .C1(n20528), .C2(n15780), .A(
        n15779), .ZN(P1_U3162) );
  OAI21_X1 U18834 ( .B1(n15783), .B2(n20357), .A(n15782), .ZN(P1_U3466) );
  AOI22_X1 U18835 ( .A1(n15784), .A2(n18775), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n18807), .ZN(n15792) );
  AOI22_X1 U18836 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18802), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n15785), .ZN(n15791) );
  INV_X1 U18837 ( .A(n15862), .ZN(n15787) );
  AOI22_X1 U18838 ( .A1(n18759), .A2(n18853), .B1(n18831), .B2(n15787), .ZN(
        n15790) );
  NAND4_X1 U18839 ( .A1(n18819), .A2(n15793), .A3(n15788), .A4(n9969), .ZN(
        n15789) );
  NAND4_X1 U18840 ( .A1(n15792), .A2(n15791), .A3(n15790), .A4(n15789), .ZN(
        P2_U2824) );
  AOI21_X1 U18841 ( .B1(n15795), .B2(n15794), .A(n15793), .ZN(n15801) );
  AOI22_X1 U18842 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n18807), .B1(n15796), 
        .B2(n18775), .ZN(n15798) );
  AOI22_X1 U18843 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n18803), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18802), .ZN(n15797) );
  OAI211_X1 U18844 ( .C1(n15799), .C2(n18796), .A(n15798), .B(n15797), .ZN(
        n15800) );
  AOI21_X1 U18845 ( .B1(n18819), .B2(n15801), .A(n15800), .ZN(n15802) );
  OAI21_X1 U18846 ( .B1(n15803), .B2(n18823), .A(n15802), .ZN(P2_U2826) );
  AOI22_X1 U18847 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n18807), .B1(n15804), 
        .B2(n18775), .ZN(n15814) );
  AOI22_X1 U18848 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18802), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n18803), .ZN(n15813) );
  INV_X1 U18849 ( .A(n15805), .ZN(n15807) );
  AOI22_X1 U18850 ( .A1(n15807), .A2(n18831), .B1(n15806), .B2(n18759), .ZN(
        n15812) );
  AOI21_X1 U18851 ( .B1(n15809), .B2(n9669), .A(n15808), .ZN(n15810) );
  NAND2_X1 U18852 ( .A1(n18819), .A2(n15810), .ZN(n15811) );
  NAND4_X1 U18853 ( .A1(n15814), .A2(n15813), .A3(n15812), .A4(n15811), .ZN(
        P2_U2827) );
  AOI22_X1 U18854 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18802), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n18807), .ZN(n15815) );
  OAI21_X1 U18855 ( .B1(n15816), .B2(n18822), .A(n15815), .ZN(n15817) );
  AOI21_X1 U18856 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n18803), .A(n15817), .ZN(
        n15824) );
  AOI21_X1 U18857 ( .B1(n15820), .B2(n15819), .A(n15818), .ZN(n15821) );
  AOI22_X1 U18858 ( .A1(n15822), .A2(n18759), .B1(n18819), .B2(n15821), .ZN(
        n15823) );
  OAI211_X1 U18859 ( .C1(n15825), .C2(n18796), .A(n15824), .B(n15823), .ZN(
        P2_U2828) );
  AOI22_X1 U18860 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18802), .B1(
        n15826), .B2(n18775), .ZN(n15836) );
  AOI22_X1 U18861 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18803), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18807), .ZN(n15835) );
  AOI22_X1 U18862 ( .A1(n15828), .A2(n18831), .B1(n15827), .B2(n18759), .ZN(
        n15834) );
  AOI21_X1 U18863 ( .B1(n15831), .B2(n15830), .A(n15829), .ZN(n15832) );
  NAND2_X1 U18864 ( .A1(n18819), .A2(n15832), .ZN(n15833) );
  NAND4_X1 U18865 ( .A1(n15836), .A2(n15835), .A3(n15834), .A4(n15833), .ZN(
        P2_U2829) );
  AOI211_X1 U18866 ( .C1(P2_EBX_REG_25__SCAN_IN), .C2(n15852), .A(n15837), .B(
        n18822), .ZN(n15839) );
  OAI22_X1 U18867 ( .A1(n9985), .A2(n18833), .B1(n19669), .B2(n18825), .ZN(
        n15838) );
  AOI211_X1 U18868 ( .C1(P2_EBX_REG_25__SCAN_IN), .C2(n18803), .A(n15839), .B(
        n15838), .ZN(n15847) );
  INV_X1 U18869 ( .A(n15840), .ZN(n15845) );
  AOI21_X1 U18870 ( .B1(n15843), .B2(n15842), .A(n15841), .ZN(n15844) );
  AOI22_X1 U18871 ( .A1(n15845), .A2(n18831), .B1(n18819), .B2(n15844), .ZN(
        n15846) );
  OAI211_X1 U18872 ( .C1(n15848), .C2(n18823), .A(n15847), .B(n15846), .ZN(
        P2_U2830) );
  AOI211_X1 U18873 ( .C1(n15851), .C2(n9980), .A(n15850), .B(n18811), .ZN(
        n15858) );
  AOI22_X1 U18874 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18802), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n18803), .ZN(n15856) );
  OAI211_X1 U18875 ( .C1(n15854), .C2(n15853), .A(n15852), .B(n18775), .ZN(
        n15855) );
  OAI211_X1 U18876 ( .C1(n18825), .C2(n19667), .A(n15856), .B(n15855), .ZN(
        n15857) );
  AOI211_X1 U18877 ( .C1(n18759), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        n15860) );
  OAI21_X1 U18878 ( .B1(n14917), .B2(n18796), .A(n15860), .ZN(P2_U2831) );
  AOI22_X1 U18879 ( .A1(n18851), .A2(n15862), .B1(n15861), .B2(n18843), .ZN(
        P2_U2856) );
  AOI22_X1 U18880 ( .A1(n15863), .A2(n18848), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n18843), .ZN(n15864) );
  OAI21_X1 U18881 ( .B1(n18843), .B2(n15865), .A(n15864), .ZN(P2_U2864) );
  AND2_X1 U18882 ( .A1(n14771), .A2(n15866), .ZN(n15867) );
  NOR2_X1 U18883 ( .A1(n12351), .A2(n15867), .ZN(n15881) );
  AOI22_X1 U18884 ( .A1(n15881), .A2(n18848), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n18843), .ZN(n15868) );
  OAI21_X1 U18885 ( .B1(n18843), .B2(n15869), .A(n15868), .ZN(P2_U2865) );
  INV_X1 U18886 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15876) );
  OR2_X1 U18887 ( .A1(n15871), .A2(n15870), .ZN(n15872) );
  NAND2_X1 U18888 ( .A1(n14772), .A2(n15872), .ZN(n15886) );
  INV_X1 U18889 ( .A(n18621), .ZN(n15873) );
  OAI22_X1 U18890 ( .A1(n15886), .A2(n18844), .B1(n15873), .B2(n18843), .ZN(
        n15874) );
  INV_X1 U18891 ( .A(n15874), .ZN(n15875) );
  OAI21_X1 U18892 ( .B1(n18851), .B2(n15876), .A(n15875), .ZN(P2_U2867) );
  AOI22_X1 U18893 ( .A1(n15877), .A2(n18848), .B1(n18851), .B2(n10111), .ZN(
        n15878) );
  OAI21_X1 U18894 ( .B1(n18851), .B2(n15879), .A(n15878), .ZN(P2_U2869) );
  INV_X1 U18895 ( .A(n19034), .ZN(n15880) );
  AOI22_X1 U18896 ( .A1(n18857), .A2(n15880), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n18881), .ZN(n15885) );
  AOI22_X1 U18897 ( .A1(n18859), .A2(BUF1_REG_22__SCAN_IN), .B1(n18858), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n15884) );
  AOI22_X1 U18898 ( .A1(n15882), .A2(n18852), .B1(n18884), .B2(n15881), .ZN(
        n15883) );
  NAND3_X1 U18899 ( .A1(n15885), .A2(n15884), .A3(n15883), .ZN(P2_U2897) );
  AOI22_X1 U18900 ( .A1(n18857), .A2(n18931), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n18881), .ZN(n15890) );
  AOI22_X1 U18901 ( .A1(n18859), .A2(BUF1_REG_20__SCAN_IN), .B1(n18858), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15889) );
  OAI22_X1 U18902 ( .A1(n18619), .A2(n18862), .B1(n18861), .B2(n15886), .ZN(
        n15887) );
  INV_X1 U18903 ( .A(n15887), .ZN(n15888) );
  NAND3_X1 U18904 ( .A1(n15890), .A2(n15889), .A3(n15888), .ZN(P2_U2899) );
  AOI22_X1 U18905 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n15915), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18791), .ZN(n15902) );
  NAND2_X1 U18906 ( .A1(n15257), .A2(n15892), .ZN(n15896) );
  NAND2_X1 U18907 ( .A1(n15894), .A2(n15893), .ZN(n15895) );
  XNOR2_X1 U18908 ( .A(n15896), .B(n15895), .ZN(n15962) );
  AOI21_X1 U18909 ( .B1(n15898), .B2(n15897), .A(n15033), .ZN(n15961) );
  AOI22_X1 U18910 ( .A1(n15962), .A2(n10903), .B1(n15939), .B2(n15961), .ZN(
        n15899) );
  INV_X1 U18911 ( .A(n15899), .ZN(n15900) );
  AOI21_X1 U18912 ( .B1(n15950), .B2(n18692), .A(n15900), .ZN(n15901) );
  OAI211_X1 U18913 ( .C1(n15922), .C2(n18688), .A(n15902), .B(n15901), .ZN(
        P2_U3000) );
  AOI22_X1 U18914 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n18791), .B1(n15944), 
        .B2(n15903), .ZN(n15908) );
  AOI222_X1 U18915 ( .A1(n15906), .A2(n10903), .B1(n15939), .B2(n15905), .C1(
        n15950), .C2(n15904), .ZN(n15907) );
  OAI211_X1 U18916 ( .C1(n18697), .C2(n15953), .A(n15908), .B(n15907), .ZN(
        P2_U3001) );
  AOI22_X1 U18917 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18791), .B1(n15944), 
        .B2(n18720), .ZN(n15913) );
  INV_X1 U18918 ( .A(n18724), .ZN(n15910) );
  AOI222_X1 U18919 ( .A1(n15911), .A2(n10903), .B1(n15950), .B2(n15910), .C1(
        n15939), .C2(n15909), .ZN(n15912) );
  OAI211_X1 U18920 ( .C1(n15914), .C2(n15953), .A(n15913), .B(n15912), .ZN(
        P2_U3003) );
  AOI22_X1 U18921 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n15915), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18791), .ZN(n15920) );
  OAI22_X1 U18922 ( .A1(n15917), .A2(n15947), .B1(n15916), .B2(n15946), .ZN(
        n15918) );
  AOI21_X1 U18923 ( .B1(n15950), .B2(n18736), .A(n15918), .ZN(n15919) );
  OAI211_X1 U18924 ( .C1(n15922), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        P2_U3004) );
  AOI22_X1 U18925 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18791), .B1(n15944), 
        .B2(n15923), .ZN(n15928) );
  INV_X1 U18926 ( .A(n15924), .ZN(n15926) );
  AOI222_X1 U18927 ( .A1(n15926), .A2(n15939), .B1(n10903), .B2(n15925), .C1(
        n15950), .C2(n18747), .ZN(n15927) );
  OAI211_X1 U18928 ( .C1(n18741), .C2(n15953), .A(n15928), .B(n15927), .ZN(
        P2_U3005) );
  AOI22_X1 U18929 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18791), .B1(n15944), 
        .B2(n18753), .ZN(n15943) );
  INV_X1 U18930 ( .A(n15929), .ZN(n18758) );
  XOR2_X1 U18931 ( .A(n15930), .B(n15931), .Z(n15984) );
  INV_X1 U18932 ( .A(n15934), .ZN(n15936) );
  NOR2_X1 U18933 ( .A1(n15936), .A2(n15935), .ZN(n15937) );
  XNOR2_X1 U18934 ( .A(n15938), .B(n15937), .ZN(n15985) );
  AOI22_X1 U18935 ( .A1(n15984), .A2(n15939), .B1(n10903), .B2(n15985), .ZN(
        n15940) );
  INV_X1 U18936 ( .A(n15940), .ZN(n15941) );
  AOI21_X1 U18937 ( .B1(n15950), .B2(n18758), .A(n15941), .ZN(n15942) );
  OAI211_X1 U18938 ( .C1(n18756), .C2(n15953), .A(n15943), .B(n15942), .ZN(
        P2_U3006) );
  AOI22_X1 U18939 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n18791), .B1(n15944), 
        .B2(n18782), .ZN(n15952) );
  OAI22_X1 U18940 ( .A1(n15948), .A2(n15947), .B1(n15946), .B2(n15945), .ZN(
        n15949) );
  AOI21_X1 U18941 ( .B1(n15950), .B2(n18783), .A(n15949), .ZN(n15951) );
  OAI211_X1 U18942 ( .C1(n15954), .C2(n15953), .A(n15952), .B(n15951), .ZN(
        P2_U3008) );
  AOI21_X1 U18943 ( .B1(n15957), .B2(n15956), .A(n15955), .ZN(n18868) );
  NOR3_X1 U18944 ( .A1(n15959), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15958), .ZN(n15960) );
  AOI21_X1 U18945 ( .B1(n18868), .B2(n15982), .A(n15960), .ZN(n15968) );
  AOI222_X1 U18946 ( .A1(n15962), .A2(n11303), .B1(n18982), .B2(n18692), .C1(
        n18977), .C2(n15961), .ZN(n15967) );
  NAND2_X1 U18947 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18791), .ZN(n15966) );
  OAI21_X1 U18948 ( .B1(n15964), .B2(n15963), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15965) );
  NAND4_X1 U18949 ( .A1(n15968), .A2(n15967), .A3(n15966), .A4(n15965), .ZN(
        P2_U3032) );
  OAI211_X1 U18950 ( .C1(n15972), .C2(n15971), .A(n15970), .B(n15969), .ZN(
        n15973) );
  AOI21_X1 U18951 ( .B1(n15982), .B2(n18714), .A(n15973), .ZN(n15976) );
  AOI22_X1 U18952 ( .A1(n15974), .A2(n11303), .B1(n18982), .B2(n18715), .ZN(
        n15975) );
  OAI211_X1 U18953 ( .C1(n15978), .C2(n15977), .A(n15976), .B(n15975), .ZN(
        P2_U3034) );
  AOI21_X1 U18954 ( .B1(n15981), .B2(n15980), .A(n15979), .ZN(n18877) );
  AOI22_X1 U18955 ( .A1(n15983), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n15982), .B2(n18877), .ZN(n15991) );
  AOI222_X1 U18956 ( .A1(n15985), .A2(n11303), .B1(n18982), .B2(n18758), .C1(
        n15984), .C2(n18977), .ZN(n15990) );
  NAND2_X1 U18957 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18791), .ZN(n15989) );
  OAI211_X1 U18958 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n15987), .B(n15986), .ZN(n15988) );
  NAND4_X1 U18959 ( .A1(n15991), .A2(n15990), .A3(n15989), .A4(n15988), .ZN(
        P2_U3038) );
  OAI22_X1 U18960 ( .A1(n19729), .A2(n15993), .B1(n15992), .B2(n19617), .ZN(
        n16000) );
  NOR2_X1 U18961 ( .A1(n15996), .A2(n19617), .ZN(n15998) );
  AOI21_X1 U18962 ( .B1(n15995), .B2(n18596), .A(n15994), .ZN(n15997) );
  OAI22_X1 U18963 ( .A1(n15998), .A2(n15997), .B1(n18596), .B2(n15996), .ZN(
        n15999) );
  NOR3_X1 U18964 ( .A1(n16001), .A2(n16000), .A3(n15999), .ZN(n16002) );
  OAI21_X1 U18965 ( .B1(n16004), .B2(n16003), .A(n16002), .ZN(P2_U3176) );
  NAND3_X1 U18966 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17584), .A3(
        n16005), .ZN(n16006) );
  XOR2_X1 U18967 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16006), .Z(
        n16065) );
  NAND2_X1 U18968 ( .A1(n17068), .A2(n16014), .ZN(n17421) );
  INV_X1 U18969 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16231) );
  NAND2_X1 U18970 ( .A1(n17535), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17516) );
  NAND4_X1 U18971 ( .A1(n17477), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17397) );
  INV_X1 U18972 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17428) );
  NAND2_X1 U18973 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17376) );
  NAND2_X1 U18974 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17335) );
  NAND2_X1 U18975 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17302) );
  NAND2_X1 U18976 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17259) );
  NAND2_X1 U18977 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17219) );
  NAND2_X1 U18978 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16039), .ZN(
        n16008) );
  INV_X1 U18979 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18510) );
  NOR2_X1 U18980 ( .A1(n18510), .A2(n17894), .ZN(n16057) );
  NAND2_X1 U18981 ( .A1(n16038), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16010) );
  INV_X1 U18982 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17566) );
  NOR2_X1 U18983 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18415), .ZN(n16009) );
  OAI21_X1 U18984 ( .B1(n17566), .B2(n17359), .A(n17958), .ZN(n17374) );
  INV_X1 U18985 ( .A(n17374), .ZN(n17334) );
  OR2_X1 U18986 ( .A1(n16010), .A2(n17334), .ZN(n16026) );
  INV_X1 U18987 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16217) );
  XOR2_X1 U18988 ( .A(n16217), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16011) );
  NOR2_X1 U18989 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17359), .ZN(
        n16041) );
  INV_X1 U18990 ( .A(n16040), .ZN(n16198) );
  NAND2_X1 U18991 ( .A1(n18299), .A2(n16010), .ZN(n16044) );
  OAI211_X1 U18992 ( .C1(n16198), .C2(n17574), .A(n17573), .B(n16044), .ZN(
        n16047) );
  NOR2_X1 U18993 ( .A1(n16041), .A2(n16047), .ZN(n16025) );
  OAI22_X1 U18994 ( .A1(n16026), .A2(n16011), .B1(n16025), .B2(n16217), .ZN(
        n16012) );
  AOI211_X1 U18995 ( .C1(n9610), .C2(n16478), .A(n16057), .B(n16012), .ZN(
        n16023) );
  NOR2_X2 U18996 ( .A1(n17922), .A2(n16177), .ZN(n17565) );
  NAND2_X1 U18997 ( .A1(n16029), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16013) );
  XNOR2_X1 U18998 ( .A(n16013), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16062) );
  INV_X1 U18999 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18529) );
  OAI221_X1 U19000 ( .B1(n18529), .B2(n16054), .C1(n16017), .C2(n16054), .A(
        n16018), .ZN(n16016) );
  AOI22_X1 U19001 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17483), .B1(
        n17312), .B2(n18529), .ZN(n16022) );
  NAND2_X1 U19002 ( .A1(n16018), .A2(n16017), .ZN(n16020) );
  NOR2_X1 U19003 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16054), .ZN(
        n16019) );
  OAI22_X1 U19004 ( .A1(n16020), .A2(n16019), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18529), .ZN(n16021) );
  AOI22_X1 U19005 ( .A1(n17565), .A2(n17768), .B1(n17485), .B2(n17771), .ZN(
        n17469) );
  NAND2_X1 U19006 ( .A1(n16067), .A2(n17382), .ZN(n17239) );
  XOR2_X1 U19007 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16039), .Z(
        n16220) );
  INV_X1 U19008 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16221) );
  OAI221_X1 U19009 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16026), .C1(
        n16221), .C2(n16025), .A(n16024), .ZN(n16027) );
  AOI21_X1 U19010 ( .B1(n9610), .B2(n16220), .A(n16027), .ZN(n16033) );
  NAND2_X1 U19011 ( .A1(n17485), .A2(n16028), .ZN(n16035) );
  OAI21_X1 U19012 ( .B1(n16029), .B2(n17578), .A(n16035), .ZN(n16031) );
  AOI22_X1 U19013 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16031), .B1(
        n17484), .B2(n16030), .ZN(n16032) );
  OAI211_X1 U19014 ( .C1(n16034), .C2(n17239), .A(n16033), .B(n16032), .ZN(
        P3_U2800) );
  NOR2_X1 U19015 ( .A1(n16048), .A2(n17225), .ZN(n16075) );
  INV_X1 U19016 ( .A(n16075), .ZN(n16036) );
  AOI21_X1 U19017 ( .B1(n16037), .B2(n16036), .A(n16035), .ZN(n16046) );
  AOI21_X1 U19018 ( .B1(n16231), .B2(n16040), .A(n16039), .ZN(n16230) );
  OAI21_X1 U19019 ( .B1(n16041), .B2(n9610), .A(n16230), .ZN(n16042) );
  OAI211_X1 U19020 ( .C1(n16044), .C2(n9859), .A(n16043), .B(n16042), .ZN(
        n16045) );
  AOI211_X1 U19021 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16047), .A(
        n16046), .B(n16045), .ZN(n16051) );
  NOR2_X1 U19022 ( .A1(n17582), .A2(n16048), .ZN(n16077) );
  OAI211_X1 U19023 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16077), .A(
        n17565), .B(n16049), .ZN(n16050) );
  OAI211_X1 U19024 ( .C1(n16052), .C2(n17458), .A(n16051), .B(n16050), .ZN(
        P3_U2801) );
  NOR3_X1 U19025 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16054), .A3(
        n16053), .ZN(n16060) );
  INV_X1 U19026 ( .A(n16055), .ZN(n17881) );
  AOI221_X1 U19027 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16056), 
        .C1(n17881), .C2(n16056), .A(n18529), .ZN(n16058) );
  AOI211_X1 U19028 ( .C1(n16060), .C2(n16059), .A(n16058), .B(n16057), .ZN(
        n16064) );
  AOI22_X1 U19029 ( .A1(n16062), .A2(n17885), .B1(n16061), .B2(n17814), .ZN(
        n16063) );
  OAI211_X1 U19030 ( .C1(n16065), .C2(n17740), .A(n16064), .B(n16063), .ZN(
        P3_U2831) );
  OR4_X1 U19031 ( .A1(n17588), .A2(n17483), .A3(n16066), .A4(n17898), .ZN(
        n16082) );
  INV_X1 U19032 ( .A(n17769), .ZN(n18563) );
  NAND2_X1 U19033 ( .A1(n18561), .A2(n17068), .ZN(n17770) );
  INV_X1 U19034 ( .A(n17770), .ZN(n17637) );
  AOI22_X1 U19035 ( .A1(n17768), .A2(n18563), .B1(n17771), .B2(n17637), .ZN(
        n17688) );
  OAI21_X1 U19036 ( .B1(n17689), .B2(n17688), .A(n17600), .ZN(n17628) );
  INV_X1 U19037 ( .A(n17628), .ZN(n17586) );
  NOR2_X1 U19038 ( .A1(n17586), .A2(n17886), .ZN(n17613) );
  AND3_X1 U19039 ( .A1(n16068), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16067), .ZN(n17224) );
  AOI22_X1 U19040 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17312), .B1(
        n17483), .B2(n16068), .ZN(n17228) );
  NOR3_X1 U19041 ( .A1(n17228), .A2(n17788), .A3(n16069), .ZN(n16070) );
  INV_X1 U19042 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18506) );
  NOR2_X1 U19043 ( .A1(n17894), .A2(n18506), .ZN(n17223) );
  AOI211_X1 U19044 ( .C1(n17613), .C2(n17224), .A(n16070), .B(n17223), .ZN(
        n16081) );
  OAI21_X1 U19045 ( .B1(n16071), .B2(n17483), .A(n16069), .ZN(n17227) );
  NAND2_X1 U19046 ( .A1(n17228), .A2(n17227), .ZN(n17226) );
  OAI21_X1 U19047 ( .B1(n17232), .B2(n16072), .A(n17226), .ZN(n16073) );
  AOI221_X1 U19048 ( .B1(n17068), .B2(n16075), .C1(n16074), .C2(n16073), .A(
        n18405), .ZN(n16079) );
  OAI21_X1 U19049 ( .B1(n16077), .B2(n17769), .A(n16076), .ZN(n16078) );
  OAI211_X1 U19050 ( .C1(n16079), .C2(n16078), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17894), .ZN(n16080) );
  OAI211_X1 U19051 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16082), .A(
        n16081), .B(n16080), .ZN(P3_U2834) );
  NOR3_X1 U19052 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16084) );
  NOR4_X1 U19053 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16083) );
  NAND4_X1 U19054 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16084), .A3(n16083), .A4(
        U215), .ZN(U213) );
  INV_X1 U19055 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18891) );
  INV_X2 U19056 ( .A(U214), .ZN(n16128) );
  NOR2_X1 U19057 ( .A1(n16128), .A2(n16085), .ZN(n16126) );
  OAI222_X1 U19058 ( .A1(U212), .A2(n18891), .B1(n16131), .B2(n16086), .C1(
        U214), .C2(n16165), .ZN(U216) );
  INV_X1 U19059 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19032) );
  INV_X1 U19060 ( .A(U212), .ZN(n16129) );
  AOI22_X1 U19061 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16128), .ZN(n16087) );
  OAI21_X1 U19062 ( .B1(n19032), .B2(n16131), .A(n16087), .ZN(U217) );
  INV_X1 U19063 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n19027) );
  AOI22_X1 U19064 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16128), .ZN(n16088) );
  OAI21_X1 U19065 ( .B1(n19027), .B2(n16131), .A(n16088), .ZN(U218) );
  INV_X1 U19066 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16090) );
  AOI22_X1 U19067 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16128), .ZN(n16089) );
  OAI21_X1 U19068 ( .B1(n16090), .B2(n16131), .A(n16089), .ZN(U219) );
  AOI22_X1 U19069 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16128), .ZN(n16091) );
  OAI21_X1 U19070 ( .B1(n19014), .B2(n16131), .A(n16091), .ZN(U220) );
  INV_X1 U19071 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16093) );
  AOI22_X1 U19072 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16128), .ZN(n16092) );
  OAI21_X1 U19073 ( .B1(n16093), .B2(n16131), .A(n16092), .ZN(U221) );
  INV_X1 U19074 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16095) );
  AOI22_X1 U19075 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16128), .ZN(n16094) );
  OAI21_X1 U19076 ( .B1(n16095), .B2(n16131), .A(n16094), .ZN(U222) );
  AOI22_X1 U19077 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16128), .ZN(n16096) );
  OAI21_X1 U19078 ( .B1(n16097), .B2(n16131), .A(n16096), .ZN(U223) );
  INV_X1 U19079 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n16098) );
  OAI222_X1 U19080 ( .A1(U214), .A2(n16098), .B1(n16131), .B2(n19040), .C1(
        U212), .C2(n16154), .ZN(U224) );
  AOI22_X1 U19081 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16128), .ZN(n16099) );
  OAI21_X1 U19082 ( .B1(n14234), .B2(n16131), .A(n16099), .ZN(U225) );
  AOI22_X1 U19083 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16128), .ZN(n16100) );
  OAI21_X1 U19084 ( .B1(n14851), .B2(n16131), .A(n16100), .ZN(U226) );
  INV_X1 U19085 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n19021) );
  AOI22_X1 U19086 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16128), .ZN(n16101) );
  OAI21_X1 U19087 ( .B1(n19021), .B2(n16131), .A(n16101), .ZN(U227) );
  AOI22_X1 U19088 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16128), .ZN(n16102) );
  OAI21_X1 U19089 ( .B1(n16103), .B2(n16131), .A(n16102), .ZN(U228) );
  INV_X1 U19090 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16105) );
  AOI22_X1 U19091 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16128), .ZN(n16104) );
  OAI21_X1 U19092 ( .B1(n16105), .B2(n16131), .A(n16104), .ZN(U229) );
  AOI222_X1 U19093 ( .A1(n16128), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n16126), 
        .B2(BUF1_REG_17__SCAN_IN), .C1(n16129), .C2(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n16106) );
  INV_X1 U19094 ( .A(n16106), .ZN(U230) );
  AOI22_X1 U19095 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16128), .ZN(n16107) );
  OAI21_X1 U19096 ( .B1(n14262), .B2(n16131), .A(n16107), .ZN(U231) );
  INV_X1 U19097 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n20688) );
  AOI22_X1 U19098 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16126), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16129), .ZN(n16108) );
  OAI21_X1 U19099 ( .B1(n20688), .B2(U214), .A(n16108), .ZN(U232) );
  INV_X1 U19100 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n20771) );
  AOI22_X1 U19101 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16126), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16128), .ZN(n16109) );
  OAI21_X1 U19102 ( .B1(n20771), .B2(U212), .A(n16109), .ZN(U233) );
  INV_X1 U19103 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16145) );
  AOI22_X1 U19104 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16126), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16128), .ZN(n16110) );
  OAI21_X1 U19105 ( .B1(n16145), .B2(U212), .A(n16110), .ZN(U234) );
  INV_X1 U19106 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n20753) );
  AOI22_X1 U19107 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16126), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16129), .ZN(n16111) );
  OAI21_X1 U19108 ( .B1(n20753), .B2(U214), .A(n16111), .ZN(U235) );
  AOI22_X1 U19109 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16128), .ZN(n16112) );
  OAI21_X1 U19110 ( .B1(n16113), .B2(n16131), .A(n16112), .ZN(U236) );
  AOI22_X1 U19111 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16128), .ZN(n16114) );
  OAI21_X1 U19112 ( .B1(n20765), .B2(n16131), .A(n16114), .ZN(U237) );
  INV_X1 U19113 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16141) );
  AOI22_X1 U19114 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16126), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16128), .ZN(n16115) );
  OAI21_X1 U19115 ( .B1(n16141), .B2(U212), .A(n16115), .ZN(U238) );
  AOI22_X1 U19116 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16128), .ZN(n16116) );
  OAI21_X1 U19117 ( .B1(n16117), .B2(n16131), .A(n16116), .ZN(U239) );
  INV_X1 U19118 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n20671) );
  AOI22_X1 U19119 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16126), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16128), .ZN(n16118) );
  OAI21_X1 U19120 ( .B1(n20671), .B2(U212), .A(n16118), .ZN(U240) );
  INV_X1 U19121 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16120) );
  AOI22_X1 U19122 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16128), .ZN(n16119) );
  OAI21_X1 U19123 ( .B1(n16120), .B2(n16131), .A(n16119), .ZN(U241) );
  INV_X1 U19124 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16138) );
  AOI22_X1 U19125 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16126), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16128), .ZN(n16121) );
  OAI21_X1 U19126 ( .B1(n16138), .B2(U212), .A(n16121), .ZN(U242) );
  AOI22_X1 U19127 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16128), .ZN(n16122) );
  OAI21_X1 U19128 ( .B1(n16123), .B2(n16131), .A(n16122), .ZN(U243) );
  INV_X1 U19129 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16136) );
  AOI22_X1 U19130 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16126), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16128), .ZN(n16124) );
  OAI21_X1 U19131 ( .B1(n16136), .B2(U212), .A(n16124), .ZN(U244) );
  INV_X1 U19132 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16135) );
  AOI22_X1 U19133 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16126), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16128), .ZN(n16125) );
  OAI21_X1 U19134 ( .B1(n16135), .B2(U212), .A(n16125), .ZN(U245) );
  INV_X1 U19135 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16134) );
  AOI22_X1 U19136 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16126), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16128), .ZN(n16127) );
  OAI21_X1 U19137 ( .B1(n16134), .B2(U212), .A(n16127), .ZN(U246) );
  AOI22_X1 U19138 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16129), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16128), .ZN(n16130) );
  OAI21_X1 U19139 ( .B1(n16132), .B2(n16131), .A(n16130), .ZN(U247) );
  INV_X1 U19140 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16133) );
  AOI22_X1 U19141 ( .A1(n16163), .A2(n16133), .B1(n17913), .B2(U215), .ZN(U251) );
  INV_X1 U19142 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n17921) );
  AOI22_X1 U19143 ( .A1(n16163), .A2(n16134), .B1(n17921), .B2(U215), .ZN(U252) );
  INV_X1 U19144 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n17926) );
  AOI22_X1 U19145 ( .A1(n16163), .A2(n16135), .B1(n17926), .B2(U215), .ZN(U253) );
  INV_X1 U19146 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n17931) );
  AOI22_X1 U19147 ( .A1(n16163), .A2(n16136), .B1(n17931), .B2(U215), .ZN(U254) );
  INV_X1 U19148 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16137) );
  AOI22_X1 U19149 ( .A1(n16163), .A2(n16137), .B1(n17937), .B2(U215), .ZN(U255) );
  INV_X1 U19150 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n17942) );
  AOI22_X1 U19151 ( .A1(n16163), .A2(n16138), .B1(n17942), .B2(U215), .ZN(U256) );
  INV_X1 U19152 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16139) );
  INV_X1 U19153 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n17949) );
  AOI22_X1 U19154 ( .A1(n16163), .A2(n16139), .B1(n17949), .B2(U215), .ZN(U257) );
  INV_X1 U19155 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n17955) );
  AOI22_X1 U19156 ( .A1(n16163), .A2(n20671), .B1(n17955), .B2(U215), .ZN(U258) );
  INV_X1 U19157 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16140) );
  INV_X1 U19158 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U19159 ( .A1(n16163), .A2(n16140), .B1(n17195), .B2(U215), .ZN(U259) );
  INV_X1 U19160 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U19161 ( .A1(n16156), .A2(n16141), .B1(n17198), .B2(U215), .ZN(U260) );
  INV_X1 U19162 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16142) );
  INV_X1 U19163 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U19164 ( .A1(n16156), .A2(n16142), .B1(n17200), .B2(U215), .ZN(U261) );
  INV_X1 U19165 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16143) );
  INV_X1 U19166 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U19167 ( .A1(n16163), .A2(n16143), .B1(n17202), .B2(U215), .ZN(U262) );
  INV_X1 U19168 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16144) );
  INV_X1 U19169 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U19170 ( .A1(n16163), .A2(n16144), .B1(n17204), .B2(U215), .ZN(U263) );
  INV_X1 U19171 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U19172 ( .A1(n16163), .A2(n16145), .B1(n17208), .B2(U215), .ZN(U264) );
  INV_X1 U19173 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n16146) );
  AOI22_X1 U19174 ( .A1(n16156), .A2(n20771), .B1(n16146), .B2(U215), .ZN(U265) );
  OAI22_X1 U19175 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16163), .ZN(n16147) );
  INV_X1 U19176 ( .A(n16147), .ZN(U266) );
  OAI22_X1 U19177 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16163), .ZN(n16148) );
  INV_X1 U19178 ( .A(n16148), .ZN(U267) );
  AOI22_X1 U19179 ( .A1(n16163), .A2(n20726), .B1(n13609), .B2(U215), .ZN(U268) );
  OAI22_X1 U19180 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16156), .ZN(n16149) );
  INV_X1 U19181 ( .A(n16149), .ZN(U269) );
  OAI22_X1 U19182 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16156), .ZN(n16150) );
  INV_X1 U19183 ( .A(n16150), .ZN(U270) );
  INV_X1 U19184 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n16151) );
  INV_X1 U19185 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19020) );
  AOI22_X1 U19186 ( .A1(n16156), .A2(n16151), .B1(n19020), .B2(U215), .ZN(U271) );
  INV_X1 U19187 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16152) );
  INV_X1 U19188 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n17944) );
  AOI22_X1 U19189 ( .A1(n16163), .A2(n16152), .B1(n17944), .B2(U215), .ZN(U272) );
  OAI22_X1 U19190 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16156), .ZN(n16153) );
  INV_X1 U19191 ( .A(n16153), .ZN(U273) );
  INV_X1 U19192 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19038) );
  AOI22_X1 U19193 ( .A1(n16156), .A2(n16154), .B1(n19038), .B2(U215), .ZN(U274) );
  INV_X1 U19194 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16155) );
  AOI22_X1 U19195 ( .A1(n16156), .A2(n16155), .B1(n17917), .B2(U215), .ZN(U275) );
  OAI22_X1 U19196 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16156), .ZN(n16157) );
  INV_X1 U19197 ( .A(n16157), .ZN(U276) );
  OAI22_X1 U19198 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16163), .ZN(n16158) );
  INV_X1 U19199 ( .A(n16158), .ZN(U277) );
  INV_X1 U19200 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16159) );
  INV_X1 U19201 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19015) );
  AOI22_X1 U19202 ( .A1(n16163), .A2(n16159), .B1(n19015), .B2(U215), .ZN(U278) );
  OAI22_X1 U19203 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16163), .ZN(n16160) );
  INV_X1 U19204 ( .A(n16160), .ZN(U279) );
  INV_X1 U19205 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16161) );
  AOI22_X1 U19206 ( .A1(n16163), .A2(n16161), .B1(n14790), .B2(U215), .ZN(U280) );
  INV_X1 U19207 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16162) );
  AOI22_X1 U19208 ( .A1(n16163), .A2(n16162), .B1(n12527), .B2(U215), .ZN(U281) );
  INV_X1 U19209 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17957) );
  AOI22_X1 U19210 ( .A1(n16163), .A2(n18891), .B1(n17957), .B2(U215), .ZN(U282) );
  INV_X1 U19211 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16164) );
  AOI222_X1 U19212 ( .A1(n18891), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16165), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16164), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16166) );
  INV_X2 U19213 ( .A(n16168), .ZN(n16167) );
  INV_X1 U19214 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18470) );
  INV_X1 U19215 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U19216 ( .A1(n16167), .A2(n18470), .B1(n19650), .B2(n16168), .ZN(
        U347) );
  INV_X1 U19217 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18468) );
  INV_X1 U19218 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19649) );
  AOI22_X1 U19219 ( .A1(n16166), .A2(n18468), .B1(n19649), .B2(n16168), .ZN(
        U348) );
  INV_X1 U19220 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18466) );
  INV_X1 U19221 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19648) );
  AOI22_X1 U19222 ( .A1(n16167), .A2(n18466), .B1(n19648), .B2(n16168), .ZN(
        U349) );
  INV_X1 U19223 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18464) );
  INV_X1 U19224 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19647) );
  AOI22_X1 U19225 ( .A1(n16167), .A2(n18464), .B1(n19647), .B2(n16168), .ZN(
        U350) );
  INV_X1 U19226 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18462) );
  INV_X1 U19227 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19646) );
  AOI22_X1 U19228 ( .A1(n16167), .A2(n18462), .B1(n19646), .B2(n16168), .ZN(
        U351) );
  INV_X1 U19229 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18461) );
  INV_X1 U19230 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19645) );
  AOI22_X1 U19231 ( .A1(n16167), .A2(n18461), .B1(n19645), .B2(n16168), .ZN(
        U352) );
  INV_X1 U19232 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18459) );
  INV_X1 U19233 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19644) );
  AOI22_X1 U19234 ( .A1(n16167), .A2(n18459), .B1(n19644), .B2(n16168), .ZN(
        U353) );
  INV_X1 U19235 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18457) );
  AOI22_X1 U19236 ( .A1(n16167), .A2(n18457), .B1(n19643), .B2(n16168), .ZN(
        U354) );
  INV_X1 U19237 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18511) );
  INV_X1 U19238 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19680) );
  AOI22_X1 U19239 ( .A1(n16167), .A2(n18511), .B1(n19680), .B2(n16168), .ZN(
        U355) );
  INV_X1 U19240 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18508) );
  INV_X1 U19241 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19677) );
  AOI22_X1 U19242 ( .A1(n16167), .A2(n18508), .B1(n19677), .B2(n16168), .ZN(
        U356) );
  INV_X1 U19243 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18505) );
  INV_X1 U19244 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19676) );
  AOI22_X1 U19245 ( .A1(n16167), .A2(n18505), .B1(n19676), .B2(n16168), .ZN(
        U357) );
  INV_X1 U19246 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18504) );
  INV_X1 U19247 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19673) );
  AOI22_X1 U19248 ( .A1(n16167), .A2(n18504), .B1(n19673), .B2(n16168), .ZN(
        U358) );
  INV_X1 U19249 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18502) );
  INV_X1 U19250 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19671) );
  AOI22_X1 U19251 ( .A1(n16167), .A2(n18502), .B1(n19671), .B2(n16168), .ZN(
        U359) );
  INV_X1 U19252 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18500) );
  INV_X1 U19253 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19670) );
  AOI22_X1 U19254 ( .A1(n16167), .A2(n18500), .B1(n19670), .B2(n16168), .ZN(
        U360) );
  INV_X1 U19255 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18497) );
  INV_X1 U19256 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19668) );
  AOI22_X1 U19257 ( .A1(n16167), .A2(n18497), .B1(n19668), .B2(n16168), .ZN(
        U361) );
  INV_X1 U19258 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18494) );
  INV_X1 U19259 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19666) );
  AOI22_X1 U19260 ( .A1(n16167), .A2(n18494), .B1(n19666), .B2(n16168), .ZN(
        U362) );
  INV_X1 U19261 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18493) );
  INV_X1 U19262 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19664) );
  AOI22_X1 U19263 ( .A1(n16167), .A2(n18493), .B1(n19664), .B2(n16168), .ZN(
        U363) );
  INV_X1 U19264 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18490) );
  INV_X1 U19265 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19663) );
  AOI22_X1 U19266 ( .A1(n16167), .A2(n18490), .B1(n19663), .B2(n16168), .ZN(
        U364) );
  INV_X1 U19267 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18455) );
  INV_X1 U19268 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19642) );
  AOI22_X1 U19269 ( .A1(n16167), .A2(n18455), .B1(n19642), .B2(n16168), .ZN(
        U365) );
  INV_X1 U19270 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18489) );
  INV_X1 U19271 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U19272 ( .A1(n16167), .A2(n18489), .B1(n19662), .B2(n16168), .ZN(
        U366) );
  INV_X1 U19273 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18487) );
  INV_X1 U19274 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20704) );
  AOI22_X1 U19275 ( .A1(n16167), .A2(n18487), .B1(n20704), .B2(n16168), .ZN(
        U367) );
  INV_X1 U19276 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18485) );
  INV_X1 U19277 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19659) );
  AOI22_X1 U19278 ( .A1(n16167), .A2(n18485), .B1(n19659), .B2(n16168), .ZN(
        U368) );
  INV_X1 U19279 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18483) );
  INV_X1 U19280 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19657) );
  AOI22_X1 U19281 ( .A1(n16167), .A2(n18483), .B1(n19657), .B2(n16168), .ZN(
        U369) );
  INV_X1 U19282 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18481) );
  INV_X1 U19283 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19655) );
  AOI22_X1 U19284 ( .A1(n16167), .A2(n18481), .B1(n19655), .B2(n16168), .ZN(
        U370) );
  INV_X1 U19285 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18479) );
  INV_X1 U19286 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19654) );
  AOI22_X1 U19287 ( .A1(n16166), .A2(n18479), .B1(n19654), .B2(n16168), .ZN(
        U371) );
  INV_X1 U19288 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18476) );
  INV_X1 U19289 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19653) );
  AOI22_X1 U19290 ( .A1(n16167), .A2(n18476), .B1(n19653), .B2(n16168), .ZN(
        U372) );
  INV_X1 U19291 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18475) );
  INV_X1 U19292 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19652) );
  AOI22_X1 U19293 ( .A1(n16167), .A2(n18475), .B1(n19652), .B2(n16168), .ZN(
        U373) );
  INV_X1 U19294 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18473) );
  INV_X1 U19295 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20705) );
  AOI22_X1 U19296 ( .A1(n16167), .A2(n18473), .B1(n20705), .B2(n16168), .ZN(
        U374) );
  INV_X1 U19297 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20733) );
  INV_X1 U19298 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19651) );
  AOI22_X1 U19299 ( .A1(n16166), .A2(n20733), .B1(n19651), .B2(n16168), .ZN(
        U375) );
  INV_X1 U19300 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18453) );
  INV_X1 U19301 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19641) );
  AOI22_X1 U19302 ( .A1(n16166), .A2(n18453), .B1(n19641), .B2(n16168), .ZN(
        U376) );
  INV_X1 U19303 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16170) );
  NAND3_X1 U19304 ( .A1(n18452), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n16169) );
  NAND2_X1 U19305 ( .A1(n18449), .A2(n18441), .ZN(n18437) );
  NAND2_X1 U19306 ( .A1(n16169), .A2(n18437), .ZN(n18517) );
  OAI21_X1 U19307 ( .B1(n18449), .B2(n16170), .A(n18436), .ZN(P3_U2633) );
  OAI21_X1 U19308 ( .B1(n16176), .B2(n17164), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16172) );
  OAI21_X1 U19309 ( .B1(n18587), .B2(n18425), .A(n16172), .ZN(P3_U2634) );
  AOI21_X1 U19310 ( .B1(n18449), .B2(n18452), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16173) );
  AOI22_X1 U19311 ( .A1(n18584), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16173), 
        .B2(n18585), .ZN(P3_U2635) );
  NOR2_X1 U19312 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n16174) );
  OAI21_X1 U19313 ( .B1(n16174), .B2(BS16), .A(n18517), .ZN(n18516) );
  OAI21_X1 U19314 ( .B1(n18517), .B2(n18575), .A(n18516), .ZN(P3_U2636) );
  NOR3_X1 U19315 ( .A1(n16176), .A2(n16175), .A3(n18403), .ZN(n18392) );
  NOR2_X1 U19316 ( .A1(n18392), .A2(n18422), .ZN(n18566) );
  INV_X1 U19317 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17904) );
  OAI21_X1 U19318 ( .B1(n18566), .B2(n17904), .A(n16177), .ZN(P3_U2637) );
  NOR4_X1 U19319 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_19__SCAN_IN), .A3(P3_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_21__SCAN_IN), .ZN(n16181) );
  NOR4_X1 U19320 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16180) );
  NOR4_X1 U19321 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16179) );
  NOR4_X1 U19322 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16178) );
  NAND4_X1 U19323 ( .A1(n16181), .A2(n16180), .A3(n16179), .A4(n16178), .ZN(
        n16187) );
  NOR4_X1 U19324 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16185) );
  AOI211_X1 U19325 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_26__SCAN_IN), .B(
        P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n16184) );
  NOR4_X1 U19326 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n16183) );
  NOR4_X1 U19327 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n16182) );
  NAND4_X1 U19328 ( .A1(n16185), .A2(n16184), .A3(n16183), .A4(n16182), .ZN(
        n16186) );
  NOR2_X1 U19329 ( .A1(n16187), .A2(n16186), .ZN(n16190) );
  NOR2_X1 U19330 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18552) );
  INV_X1 U19331 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n16188) );
  NAND3_X1 U19332 ( .A1(n16190), .A2(n18552), .A3(n16188), .ZN(n16191) );
  INV_X1 U19333 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18551) );
  NAND2_X1 U19334 ( .A1(n16190), .A2(n18551), .ZN(n18553) );
  OAI21_X1 U19335 ( .B1(n16190), .B2(P3_BYTEENABLE_REG_1__SCAN_IN), .A(n18553), 
        .ZN(n16189) );
  NAND2_X1 U19336 ( .A1(n16191), .A2(n16189), .ZN(P3_U2638) );
  INV_X1 U19337 ( .A(n16190), .ZN(n18559) );
  NAND2_X1 U19338 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n18559), .ZN(n16192) );
  OAI211_X1 U19339 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(n18553), .A(n16192), 
        .B(n16191), .ZN(P3_U2639) );
  NAND2_X1 U19340 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18415), .ZN(n18419) );
  INV_X2 U19341 ( .A(n17894), .ZN(n17896) );
  NOR3_X1 U19342 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18435) );
  NOR2_X1 U19343 ( .A1(n17896), .A2(n18432), .ZN(n16523) );
  OAI211_X1 U19344 ( .C1(n17922), .C2(n16193), .A(n18577), .B(n18575), .ZN(
        n18414) );
  INV_X1 U19345 ( .A(n18414), .ZN(n16194) );
  NAND2_X1 U19346 ( .A1(n18573), .A2(n17102), .ZN(n16197) );
  AOI211_X4 U19347 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17922), .A(n16194), .B(
        n16197), .ZN(n16559) );
  INV_X1 U19348 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18512) );
  INV_X1 U19349 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18503) );
  NOR2_X1 U19350 ( .A1(n18506), .A2(n18503), .ZN(n16240) );
  INV_X1 U19351 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18499) );
  INV_X1 U19352 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18495) );
  INV_X1 U19353 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18477) );
  INV_X1 U19354 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18472) );
  INV_X1 U19355 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18469) );
  INV_X1 U19356 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18465) );
  INV_X1 U19357 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18463) );
  INV_X1 U19358 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18460) );
  INV_X1 U19359 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18456) );
  NAND2_X1 U19360 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16552) );
  NOR2_X1 U19361 ( .A1(n18456), .A2(n16552), .ZN(n16519) );
  NAND2_X1 U19362 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16519), .ZN(n16475) );
  NOR2_X1 U19363 ( .A1(n18460), .A2(n16475), .ZN(n16474) );
  NAND2_X1 U19364 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16474), .ZN(n16463) );
  NOR3_X1 U19365 ( .A1(n18465), .A2(n18463), .A3(n16463), .ZN(n16444) );
  NAND2_X1 U19366 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16444), .ZN(n16440) );
  NOR2_X1 U19367 ( .A1(n18469), .A2(n16440), .ZN(n16425) );
  NAND2_X1 U19368 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16425), .ZN(n16408) );
  NOR2_X1 U19369 ( .A1(n18472), .A2(n16408), .ZN(n16410) );
  NAND2_X1 U19370 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16410), .ZN(n16396) );
  NOR2_X1 U19371 ( .A1(n18477), .A2(n16396), .ZN(n16311) );
  INV_X1 U19372 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18491) );
  INV_X1 U19373 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18484) );
  NAND3_X1 U19374 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16336) );
  NOR2_X1 U19375 ( .A1(n18484), .A2(n16336), .ZN(n16326) );
  NAND3_X1 U19376 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(n16326), .ZN(n16313) );
  NOR2_X1 U19377 ( .A1(n18491), .A2(n16313), .ZN(n16303) );
  NAND3_X1 U19378 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16311), .A3(n16303), 
        .ZN(n16294) );
  NOR2_X1 U19379 ( .A1(n18495), .A2(n16294), .ZN(n16289) );
  NAND2_X1 U19380 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16289), .ZN(n16281) );
  NOR2_X1 U19381 ( .A1(n18499), .A2(n16281), .ZN(n16262) );
  NAND2_X1 U19382 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16262), .ZN(n16210) );
  NOR2_X1 U19383 ( .A1(n16517), .A2(n16210), .ZN(n16255) );
  NAND3_X1 U19384 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16240), .A3(n16255), 
        .ZN(n16212) );
  NOR3_X1 U19385 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18512), .A3(n16212), 
        .ZN(n16195) );
  AOI21_X1 U19386 ( .B1(n16559), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16195), .ZN(
        n16216) );
  NAND2_X1 U19387 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17922), .ZN(n16196) );
  AOI211_X4 U19388 ( .C1(n18575), .C2(n18577), .A(n16197), .B(n16196), .ZN(
        n16562) );
  NOR3_X1 U19389 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16542) );
  INV_X1 U19390 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16934) );
  NAND2_X1 U19391 ( .A1(n16542), .A2(n16934), .ZN(n16537) );
  NOR2_X1 U19392 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16537), .ZN(n16511) );
  NAND2_X1 U19393 ( .A1(n16511), .A2(n16508), .ZN(n16507) );
  NAND2_X1 U19394 ( .A1(n16489), .A2(n16486), .ZN(n16485) );
  NAND2_X1 U19395 ( .A1(n16467), .A2(n16462), .ZN(n16453) );
  NAND2_X1 U19396 ( .A1(n16445), .A2(n16433), .ZN(n16432) );
  NAND2_X1 U19397 ( .A1(n16415), .A2(n16835), .ZN(n16409) );
  INV_X1 U19398 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16388) );
  NAND2_X1 U19399 ( .A1(n16391), .A2(n16388), .ZN(n16387) );
  INV_X1 U19400 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16362) );
  NAND2_X1 U19401 ( .A1(n16374), .A2(n16362), .ZN(n16361) );
  INV_X1 U19402 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16341) );
  NAND2_X1 U19403 ( .A1(n16348), .A2(n16341), .ZN(n16340) );
  INV_X1 U19404 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16737) );
  NAND2_X1 U19405 ( .A1(n16327), .A2(n16737), .ZN(n16322) );
  INV_X1 U19406 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16302) );
  NAND2_X1 U19407 ( .A1(n16306), .A2(n16302), .ZN(n16299) );
  INV_X1 U19408 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16278) );
  NAND2_X1 U19409 ( .A1(n16286), .A2(n16278), .ZN(n16277) );
  INV_X1 U19410 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16257) );
  NAND2_X1 U19411 ( .A1(n16263), .A2(n16257), .ZN(n16256) );
  NOR2_X1 U19412 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16256), .ZN(n16242) );
  INV_X1 U19413 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16687) );
  NAND2_X1 U19414 ( .A1(n16242), .A2(n16687), .ZN(n16218) );
  NOR2_X1 U19415 ( .A1(n16569), .A2(n16218), .ZN(n16225) );
  INV_X1 U19416 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16249) );
  NOR2_X1 U19417 ( .A1(n17566), .A2(n17218), .ZN(n16200) );
  NAND2_X1 U19418 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16200), .ZN(
        n16199) );
  AOI21_X1 U19419 ( .B1(n16249), .B2(n16199), .A(n16198), .ZN(n17217) );
  OAI21_X1 U19420 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16200), .A(
        n16199), .ZN(n17234) );
  INV_X1 U19421 ( .A(n17234), .ZN(n16252) );
  INV_X1 U19422 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17261) );
  INV_X1 U19423 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16205) );
  NAND2_X1 U19424 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17321), .ZN(
        n16337) );
  NAND2_X1 U19425 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17292), .ZN(
        n16208) );
  NOR2_X1 U19426 ( .A1(n17302), .A2(n16208), .ZN(n17256) );
  INV_X1 U19427 ( .A(n17256), .ZN(n16204) );
  NOR2_X1 U19428 ( .A1(n16205), .A2(n16204), .ZN(n16203) );
  NAND2_X1 U19429 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16203), .ZN(
        n16202) );
  NOR2_X1 U19430 ( .A1(n17261), .A2(n16202), .ZN(n17215) );
  INV_X1 U19431 ( .A(n17215), .ZN(n16201) );
  AOI21_X1 U19432 ( .B1(n9858), .B2(n16201), .A(n16200), .ZN(n17248) );
  AOI21_X1 U19433 ( .B1(n17261), .B2(n16202), .A(n17215), .ZN(n17263) );
  OAI21_X1 U19434 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16203), .A(
        n16202), .ZN(n17270) );
  INV_X1 U19435 ( .A(n17270), .ZN(n16285) );
  AOI21_X1 U19436 ( .B1(n16205), .B2(n16204), .A(n16203), .ZN(n17285) );
  INV_X1 U19437 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16307) );
  INV_X1 U19438 ( .A(n16208), .ZN(n16207) );
  NAND2_X1 U19439 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16207), .ZN(
        n16206) );
  AOI21_X1 U19440 ( .B1(n16307), .B2(n16206), .A(n17256), .ZN(n17294) );
  OAI21_X1 U19441 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16207), .A(
        n16206), .ZN(n17306) );
  OAI21_X1 U19442 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17292), .A(
        n16208), .ZN(n16209) );
  INV_X1 U19443 ( .A(n16209), .ZN(n17326) );
  INV_X2 U19444 ( .A(n16478), .ZN(n16529) );
  NOR2_X1 U19445 ( .A1(n17566), .A2(n17372), .ZN(n17373) );
  NAND2_X1 U19446 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17373), .ZN(
        n16381) );
  OAI21_X1 U19447 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16381), .A(
        n16478), .ZN(n16371) );
  OAI21_X1 U19448 ( .B1(n17292), .B2(n16529), .A(n16371), .ZN(n16329) );
  NOR2_X1 U19449 ( .A1(n17326), .A2(n16329), .ZN(n16328) );
  OR2_X1 U19450 ( .A1(n16328), .A2(n16529), .ZN(n16317) );
  NOR2_X1 U19451 ( .A1(n17285), .A2(n16296), .ZN(n16295) );
  NOR2_X1 U19452 ( .A1(n16295), .A2(n16529), .ZN(n16284) );
  NOR2_X1 U19453 ( .A1(n16285), .A2(n16284), .ZN(n16283) );
  NOR2_X1 U19454 ( .A1(n16283), .A2(n16529), .ZN(n16273) );
  NOR2_X1 U19455 ( .A1(n17263), .A2(n16273), .ZN(n16272) );
  NOR2_X1 U19456 ( .A1(n16250), .A2(n16529), .ZN(n16244) );
  NOR2_X1 U19457 ( .A1(n17217), .A2(n16244), .ZN(n16243) );
  NOR2_X1 U19458 ( .A1(n16243), .A2(n16529), .ZN(n16229) );
  NAND2_X1 U19459 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16240), .ZN(n16211) );
  INV_X1 U19460 ( .A(n16473), .ZN(n16572) );
  AND2_X1 U19461 ( .A1(n16561), .A2(n16210), .ZN(n16261) );
  NOR2_X1 U19462 ( .A1(n16572), .A2(n16261), .ZN(n16260) );
  INV_X1 U19463 ( .A(n16260), .ZN(n16268) );
  AOI21_X1 U19464 ( .B1(n16561), .B2(n16211), .A(n16268), .ZN(n16239) );
  NOR2_X1 U19465 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16212), .ZN(n16223) );
  INV_X1 U19466 ( .A(n16223), .ZN(n16213) );
  AOI21_X1 U19467 ( .B1(n16239), .B2(n16213), .A(n18510), .ZN(n16214) );
  OAI211_X1 U19468 ( .C1(n16217), .C2(n16549), .A(n16216), .B(n16215), .ZN(
        P3_U2640) );
  NAND2_X1 U19469 ( .A1(n16562), .A2(n16218), .ZN(n16235) );
  XOR2_X1 U19470 ( .A(n16220), .B(n16219), .Z(n16224) );
  OAI22_X1 U19471 ( .A1(n16239), .A2(n18512), .B1(n16221), .B2(n16549), .ZN(
        n16222) );
  AOI211_X1 U19472 ( .C1(n16224), .C2(n18432), .A(n16223), .B(n16222), .ZN(
        n16227) );
  OAI21_X1 U19473 ( .B1(n16559), .B2(n16225), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16226) );
  OAI211_X1 U19474 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16235), .A(n16227), .B(
        n16226), .ZN(P3_U2641) );
  INV_X1 U19475 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18507) );
  AOI211_X1 U19476 ( .C1(n16230), .C2(n16229), .A(n16228), .B(n16531), .ZN(
        n16234) );
  NAND2_X1 U19477 ( .A1(n16240), .A2(n16255), .ZN(n16232) );
  OAI22_X1 U19478 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16232), .B1(n16231), 
        .B2(n16549), .ZN(n16233) );
  AOI211_X1 U19479 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16559), .A(n16234), .B(
        n16233), .ZN(n16238) );
  INV_X1 U19480 ( .A(n16235), .ZN(n16236) );
  OAI21_X1 U19481 ( .B1(n16242), .B2(n16687), .A(n16236), .ZN(n16237) );
  OAI211_X1 U19482 ( .C1(n16239), .C2(n18507), .A(n16238), .B(n16237), .ZN(
        P3_U2642) );
  AOI21_X1 U19483 ( .B1(n18506), .B2(n18503), .A(n16240), .ZN(n16241) );
  AOI22_X1 U19484 ( .A1(n16559), .A2(P3_EBX_REG_28__SCAN_IN), .B1(n16255), 
        .B2(n16241), .ZN(n16248) );
  AOI211_X1 U19485 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16256), .A(n16242), .B(
        n16569), .ZN(n16246) );
  AOI211_X1 U19486 ( .C1(n17217), .C2(n16244), .A(n16243), .B(n16531), .ZN(
        n16245) );
  AOI211_X1 U19487 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16268), .A(n16246), 
        .B(n16245), .ZN(n16247) );
  OAI211_X1 U19488 ( .C1(n16249), .C2(n16549), .A(n16248), .B(n16247), .ZN(
        P3_U2643) );
  AOI211_X1 U19489 ( .C1(n16252), .C2(n16251), .A(n16250), .B(n16531), .ZN(
        n16254) );
  INV_X1 U19490 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17237) );
  OAI22_X1 U19491 ( .A1(n17237), .A2(n16549), .B1(n16570), .B2(n16257), .ZN(
        n16253) );
  AOI211_X1 U19492 ( .C1(n16255), .C2(n18503), .A(n16254), .B(n16253), .ZN(
        n16259) );
  OAI211_X1 U19493 ( .C1(n16263), .C2(n16257), .A(n16562), .B(n16256), .ZN(
        n16258) );
  OAI211_X1 U19494 ( .C1(n16260), .C2(n18503), .A(n16259), .B(n16258), .ZN(
        P3_U2644) );
  AOI22_X1 U19495 ( .A1(n16559), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16262), 
        .B2(n16261), .ZN(n16270) );
  AOI211_X1 U19496 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16277), .A(n16263), .B(
        n16569), .ZN(n16267) );
  AOI211_X1 U19497 ( .C1(n17248), .C2(n16265), .A(n16264), .B(n16531), .ZN(
        n16266) );
  AOI211_X1 U19498 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16268), .A(n16267), 
        .B(n16266), .ZN(n16269) );
  OAI211_X1 U19499 ( .C1(n9858), .C2(n16549), .A(n16270), .B(n16269), .ZN(
        P3_U2645) );
  NAND2_X1 U19500 ( .A1(n16561), .A2(n18499), .ZN(n16282) );
  INV_X1 U19501 ( .A(n16289), .ZN(n16271) );
  AOI21_X1 U19502 ( .B1(n16561), .B2(n16271), .A(n16572), .ZN(n16293) );
  OAI21_X1 U19503 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16517), .A(n16293), 
        .ZN(n16276) );
  AOI211_X1 U19504 ( .C1(n17263), .C2(n16273), .A(n16272), .B(n16531), .ZN(
        n16275) );
  OAI22_X1 U19505 ( .A1(n17261), .A2(n16549), .B1(n16570), .B2(n16278), .ZN(
        n16274) );
  AOI211_X1 U19506 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16276), .A(n16275), 
        .B(n16274), .ZN(n16280) );
  OAI211_X1 U19507 ( .C1(n16286), .C2(n16278), .A(n16562), .B(n16277), .ZN(
        n16279) );
  OAI211_X1 U19508 ( .C1(n16282), .C2(n16281), .A(n16280), .B(n16279), .ZN(
        P3_U2646) );
  INV_X1 U19509 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18496) );
  AOI22_X1 U19510 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16564), .B1(
        n16559), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16292) );
  NOR2_X1 U19511 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16517), .ZN(n16290) );
  AOI211_X1 U19512 ( .C1(n16285), .C2(n16284), .A(n16283), .B(n16531), .ZN(
        n16288) );
  AOI211_X1 U19513 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16299), .A(n16286), .B(
        n16569), .ZN(n16287) );
  AOI211_X1 U19514 ( .C1(n16290), .C2(n16289), .A(n16288), .B(n16287), .ZN(
        n16291) );
  OAI211_X1 U19515 ( .C1(n18496), .C2(n16293), .A(n16292), .B(n16291), .ZN(
        P3_U2647) );
  AOI221_X1 U19516 ( .B1(n16517), .B2(n18495), .C1(n16294), .C2(n18495), .A(
        n16293), .ZN(n16298) );
  AOI211_X1 U19517 ( .C1(n17285), .C2(n16296), .A(n16295), .B(n16531), .ZN(
        n16297) );
  AOI211_X1 U19518 ( .C1(n16564), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16298), .B(n16297), .ZN(n16301) );
  OAI211_X1 U19519 ( .C1(n16306), .C2(n16302), .A(n16562), .B(n16299), .ZN(
        n16300) );
  OAI211_X1 U19520 ( .C1(n16302), .C2(n16570), .A(n16301), .B(n16300), .ZN(
        P3_U2648) );
  NOR3_X1 U19521 ( .A1(n16517), .A2(n18477), .A3(n16396), .ZN(n16325) );
  NAND2_X1 U19522 ( .A1(n16303), .A2(n16325), .ZN(n16316) );
  AOI211_X1 U19523 ( .C1(n17294), .C2(n16305), .A(n16304), .B(n16531), .ZN(
        n16310) );
  AOI211_X1 U19524 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16322), .A(n16306), .B(
        n16569), .ZN(n16309) );
  INV_X1 U19525 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16680) );
  OAI22_X1 U19526 ( .A1(n16307), .A2(n16549), .B1(n16570), .B2(n16680), .ZN(
        n16308) );
  NOR3_X1 U19527 ( .A1(n16310), .A2(n16309), .A3(n16308), .ZN(n16315) );
  NAND2_X1 U19528 ( .A1(n16311), .A2(n16473), .ZN(n16397) );
  NAND2_X1 U19529 ( .A1(n16473), .A2(n16517), .ZN(n16575) );
  OAI21_X1 U19530 ( .B1(n16313), .B2(n16397), .A(n16575), .ZN(n16312) );
  INV_X1 U19531 ( .A(n16312), .ZN(n16332) );
  INV_X1 U19532 ( .A(n16325), .ZN(n16380) );
  NOR3_X1 U19533 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16313), .A3(n16380), 
        .ZN(n16321) );
  OAI21_X1 U19534 ( .B1(n16332), .B2(n16321), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16314) );
  OAI211_X1 U19535 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16316), .A(n16315), 
        .B(n16314), .ZN(P3_U2649) );
  OAI21_X1 U19536 ( .B1(n17306), .B2(n16317), .A(n18432), .ZN(n16318) );
  INV_X1 U19537 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17309) );
  OAI22_X1 U19538 ( .A1(n16319), .A2(n16318), .B1(n17309), .B2(n16549), .ZN(
        n16320) );
  AOI211_X1 U19539 ( .C1(n16332), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16321), 
        .B(n16320), .ZN(n16324) );
  OAI211_X1 U19540 ( .C1(n16327), .C2(n16737), .A(n16562), .B(n16322), .ZN(
        n16323) );
  OAI211_X1 U19541 ( .C1(n16737), .C2(n16570), .A(n16324), .B(n16323), .ZN(
        P3_U2650) );
  NAND2_X1 U19542 ( .A1(n16326), .A2(n16325), .ZN(n16347) );
  INV_X1 U19543 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18488) );
  NAND2_X1 U19544 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18488), .ZN(n16335) );
  AOI22_X1 U19545 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16564), .B1(
        n16559), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16334) );
  AOI211_X1 U19546 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16340), .A(n16327), .B(
        n16569), .ZN(n16331) );
  AOI211_X1 U19547 ( .C1(n17326), .C2(n16329), .A(n16328), .B(n16531), .ZN(
        n16330) );
  AOI211_X1 U19548 ( .C1(n16332), .C2(P3_REIP_REG_20__SCAN_IN), .A(n16331), 
        .B(n16330), .ZN(n16333) );
  OAI211_X1 U19549 ( .C1(n16347), .C2(n16335), .A(n16334), .B(n16333), .ZN(
        P3_U2651) );
  AOI22_X1 U19550 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16564), .B1(
        n16559), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16346) );
  OAI21_X1 U19551 ( .B1(n16336), .B2(n16397), .A(n16575), .ZN(n16357) );
  INV_X1 U19552 ( .A(n16357), .ZN(n16360) );
  NOR3_X1 U19553 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16336), .A3(n16380), 
        .ZN(n16354) );
  INV_X1 U19554 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16363) );
  NAND2_X1 U19555 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17358), .ZN(
        n16369) );
  NOR2_X1 U19556 ( .A1(n16363), .A2(n16369), .ZN(n17332) );
  NAND2_X1 U19557 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17332), .ZN(
        n16349) );
  INV_X1 U19558 ( .A(n16349), .ZN(n16338) );
  OAI21_X1 U19559 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16338), .A(
        n16337), .ZN(n17337) );
  OAI21_X1 U19560 ( .B1(n16338), .B2(n16529), .A(n16371), .ZN(n16339) );
  XOR2_X1 U19561 ( .A(n17337), .B(n16339), .Z(n16343) );
  OAI211_X1 U19562 ( .C1(n16348), .C2(n16341), .A(n16562), .B(n16340), .ZN(
        n16342) );
  OAI211_X1 U19563 ( .C1(n16343), .C2(n16531), .A(n17894), .B(n16342), .ZN(
        n16344) );
  AOI221_X1 U19564 ( .B1(n16360), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n16354), 
        .C2(P3_REIP_REG_19__SCAN_IN), .A(n16344), .ZN(n16345) );
  OAI211_X1 U19565 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16347), .A(n16346), 
        .B(n16345), .ZN(P3_U2652) );
  AOI22_X1 U19566 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16564), .B1(
        n16559), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16356) );
  AOI211_X1 U19567 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16361), .A(n16348), .B(
        n16569), .ZN(n16353) );
  OAI21_X1 U19568 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17332), .A(
        n16349), .ZN(n17347) );
  INV_X1 U19569 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16571) );
  NAND2_X1 U19570 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16571), .ZN(
        n16514) );
  OAI21_X1 U19571 ( .B1(n17333), .B2(n16514), .A(n16478), .ZN(n16351) );
  OAI21_X1 U19572 ( .B1(n17347), .B2(n16351), .A(n18432), .ZN(n16350) );
  AOI21_X1 U19573 ( .B1(n17347), .B2(n16351), .A(n16350), .ZN(n16352) );
  NOR4_X1 U19574 ( .A1(n17896), .A2(n16354), .A3(n16353), .A4(n16352), .ZN(
        n16355) );
  OAI211_X1 U19575 ( .C1(n18484), .C2(n16357), .A(n16356), .B(n16355), .ZN(
        P3_U2653) );
  INV_X1 U19576 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18480) );
  INV_X1 U19577 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18478) );
  NOR4_X1 U19578 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18480), .A3(n18478), 
        .A4(n16380), .ZN(n16359) );
  OAI22_X1 U19579 ( .A1(n16363), .A2(n16549), .B1(n16570), .B2(n16362), .ZN(
        n16358) );
  AOI211_X1 U19580 ( .C1(n16360), .C2(P3_REIP_REG_17__SCAN_IN), .A(n16359), 
        .B(n16358), .ZN(n16368) );
  OAI211_X1 U19581 ( .C1(n16374), .C2(n16362), .A(n16562), .B(n16361), .ZN(
        n16367) );
  AOI21_X1 U19582 ( .B1(n16363), .B2(n16369), .A(n17332), .ZN(n17360) );
  INV_X1 U19583 ( .A(n16514), .ZN(n16546) );
  AOI21_X1 U19584 ( .B1(n17358), .B2(n16546), .A(n16529), .ZN(n16365) );
  AOI21_X1 U19585 ( .B1(n17360), .B2(n16365), .A(n16531), .ZN(n16364) );
  OAI21_X1 U19586 ( .B1(n17360), .B2(n16365), .A(n16364), .ZN(n16366) );
  NAND4_X1 U19587 ( .A1(n16368), .A2(n17894), .A3(n16367), .A4(n16366), .ZN(
        P3_U2654) );
  OAI21_X1 U19588 ( .B1(n18478), .B2(n16397), .A(n16575), .ZN(n16379) );
  INV_X1 U19589 ( .A(n16371), .ZN(n16382) );
  INV_X1 U19590 ( .A(n16381), .ZN(n16370) );
  OAI21_X1 U19591 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16370), .A(
        n16369), .ZN(n17379) );
  INV_X1 U19592 ( .A(n17379), .ZN(n16372) );
  AOI221_X1 U19593 ( .B1(n16382), .B2(n16372), .C1(n16371), .C2(n17379), .A(
        n16531), .ZN(n16373) );
  AOI211_X1 U19594 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n16564), .A(
        n17896), .B(n16373), .ZN(n16378) );
  NOR3_X1 U19595 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18478), .A3(n16380), 
        .ZN(n16376) );
  AOI211_X1 U19596 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16387), .A(n16374), .B(
        n16569), .ZN(n16375) );
  AOI211_X1 U19597 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16559), .A(n16376), .B(
        n16375), .ZN(n16377) );
  OAI211_X1 U19598 ( .C1(n16379), .C2(n18480), .A(n16378), .B(n16377), .ZN(
        P3_U2655) );
  INV_X1 U19599 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17387) );
  AOI21_X1 U19600 ( .B1(n18478), .B2(n16380), .A(n16379), .ZN(n16386) );
  OAI21_X1 U19601 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17373), .A(
        n16381), .ZN(n17384) );
  NOR2_X1 U19602 ( .A1(n16529), .A2(n16571), .ZN(n16563) );
  NOR2_X1 U19603 ( .A1(n16563), .A2(n16531), .ZN(n16556) );
  OAI21_X1 U19604 ( .B1(n17373), .B2(n16529), .A(n16556), .ZN(n16384) );
  NAND3_X1 U19605 ( .A1(n16382), .A2(n18432), .A3(n17384), .ZN(n16383) );
  OAI211_X1 U19606 ( .C1(n17384), .C2(n16384), .A(n17894), .B(n16383), .ZN(
        n16385) );
  AOI211_X1 U19607 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16559), .A(n16386), .B(
        n16385), .ZN(n16390) );
  OAI211_X1 U19608 ( .C1(n16391), .C2(n16388), .A(n16562), .B(n16387), .ZN(
        n16389) );
  OAI211_X1 U19609 ( .C1(n16549), .C2(n17387), .A(n16390), .B(n16389), .ZN(
        P3_U2656) );
  AOI211_X1 U19610 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16409), .A(n16391), .B(
        n16569), .ZN(n16392) );
  AOI21_X1 U19611 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16559), .A(n16392), .ZN(
        n16401) );
  INV_X1 U19612 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16393) );
  NAND3_X1 U19613 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17509), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16476) );
  NOR2_X1 U19614 ( .A1(n17397), .A2(n16476), .ZN(n17414) );
  NAND2_X1 U19615 ( .A1(n17413), .A2(n17414), .ZN(n16404) );
  AOI21_X1 U19616 ( .B1(n16393), .B2(n16404), .A(n17373), .ZN(n17401) );
  OAI21_X1 U19617 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16404), .A(
        n16478), .ZN(n16394) );
  XNOR2_X1 U19618 ( .A(n17401), .B(n16394), .ZN(n16395) );
  AOI22_X1 U19619 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16564), .B1(
        n18432), .B2(n16395), .ZN(n16400) );
  NOR2_X1 U19620 ( .A1(n16517), .A2(n16396), .ZN(n16398) );
  OAI211_X1 U19621 ( .C1(n16398), .C2(P3_REIP_REG_14__SCAN_IN), .A(n16575), 
        .B(n16397), .ZN(n16399) );
  NAND4_X1 U19622 ( .A1(n16401), .A2(n16400), .A3(n16399), .A4(n17894), .ZN(
        P3_U2657) );
  INV_X1 U19623 ( .A(n17414), .ZN(n16428) );
  NOR2_X1 U19624 ( .A1(n17428), .A2(n16428), .ZN(n16417) );
  OAI21_X1 U19625 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16417), .A(
        n16404), .ZN(n17417) );
  INV_X1 U19626 ( .A(n16556), .ZN(n16402) );
  AOI211_X1 U19627 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16478), .A(
        n17417), .B(n16402), .ZN(n16407) );
  NOR2_X1 U19628 ( .A1(n16529), .A2(n16531), .ZN(n16403) );
  OAI211_X1 U19629 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n16404), .A(
        n16403), .B(n17417), .ZN(n16405) );
  OAI211_X1 U19630 ( .C1(n16570), .C2(n16835), .A(n17894), .B(n16405), .ZN(
        n16406) );
  AOI211_X1 U19631 ( .C1(n16564), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16407), .B(n16406), .ZN(n16414) );
  INV_X1 U19632 ( .A(n16408), .ZN(n16421) );
  OAI21_X1 U19633 ( .B1(n16421), .B2(n16517), .A(n16473), .ZN(n16426) );
  NOR2_X1 U19634 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16517), .ZN(n16420) );
  OAI21_X1 U19635 ( .B1(n16426), .B2(n16420), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16413) );
  OAI211_X1 U19636 ( .C1(n16415), .C2(n16835), .A(n16562), .B(n16409), .ZN(
        n16412) );
  INV_X1 U19637 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18474) );
  NAND3_X1 U19638 ( .A1(n16561), .A2(n16410), .A3(n18474), .ZN(n16411) );
  NAND4_X1 U19639 ( .A1(n16414), .A2(n16413), .A3(n16412), .A4(n16411), .ZN(
        P3_U2658) );
  AOI211_X1 U19640 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16432), .A(n16415), .B(
        n16569), .ZN(n16416) );
  AOI21_X1 U19641 ( .B1(n16564), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16416), .ZN(n16424) );
  AOI21_X1 U19642 ( .B1(n17428), .B2(n16428), .A(n16417), .ZN(n17431) );
  OAI21_X1 U19643 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16428), .A(
        n16478), .ZN(n16418) );
  XNOR2_X1 U19644 ( .A(n17431), .B(n16418), .ZN(n16419) );
  AOI22_X1 U19645 ( .A1(n16559), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n18432), 
        .B2(n16419), .ZN(n16423) );
  AOI22_X1 U19646 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16426), .B1(n16421), 
        .B2(n16420), .ZN(n16422) );
  NAND4_X1 U19647 ( .A1(n16424), .A2(n16423), .A3(n16422), .A4(n17894), .ZN(
        P3_U2659) );
  AOI21_X1 U19648 ( .B1(n16561), .B2(n16425), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16437) );
  INV_X1 U19649 ( .A(n16426), .ZN(n16436) );
  NOR2_X1 U19650 ( .A1(n17473), .A2(n17492), .ZN(n17472) );
  NAND2_X1 U19651 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17472), .ZN(
        n16477) );
  NOR2_X1 U19652 ( .A1(n17475), .A2(n16477), .ZN(n16464) );
  NAND2_X1 U19653 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16464), .ZN(
        n16450) );
  NOR2_X1 U19654 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16450), .ZN(
        n16427) );
  AOI21_X1 U19655 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16427), .A(
        n16529), .ZN(n16429) );
  INV_X1 U19656 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17450) );
  NOR2_X1 U19657 ( .A1(n17450), .A2(n16450), .ZN(n16438) );
  OAI21_X1 U19658 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16438), .A(
        n16428), .ZN(n17436) );
  XOR2_X1 U19659 ( .A(n16429), .B(n17436), .Z(n16430) );
  OAI22_X1 U19660 ( .A1(n16570), .A2(n16433), .B1(n16531), .B2(n16430), .ZN(
        n16431) );
  AOI211_X1 U19661 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n16564), .A(
        n17896), .B(n16431), .ZN(n16435) );
  OAI211_X1 U19662 ( .C1(n16445), .C2(n16433), .A(n16562), .B(n16432), .ZN(
        n16434) );
  OAI211_X1 U19663 ( .C1(n16437), .C2(n16436), .A(n16435), .B(n16434), .ZN(
        P3_U2660) );
  AOI21_X1 U19664 ( .B1(n17450), .B2(n16450), .A(n16438), .ZN(n17453) );
  INV_X1 U19665 ( .A(n16450), .ZN(n16439) );
  AOI21_X1 U19666 ( .B1(n16571), .B2(n16439), .A(n16529), .ZN(n16451) );
  XOR2_X1 U19667 ( .A(n17453), .B(n16451), .Z(n16442) );
  NOR3_X1 U19668 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16517), .A3(n16440), 
        .ZN(n16441) );
  AOI211_X1 U19669 ( .C1(n18432), .C2(n16442), .A(n17896), .B(n16441), .ZN(
        n16449) );
  OAI21_X1 U19670 ( .B1(n16517), .B2(n16444), .A(n16473), .ZN(n16443) );
  INV_X1 U19671 ( .A(n16443), .ZN(n16471) );
  INV_X1 U19672 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18467) );
  NAND3_X1 U19673 ( .A1(n16561), .A2(n16444), .A3(n18467), .ZN(n16460) );
  AOI21_X1 U19674 ( .B1(n16471), .B2(n16460), .A(n18469), .ZN(n16447) );
  AOI211_X1 U19675 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16453), .A(n16445), .B(
        n16569), .ZN(n16446) );
  AOI211_X1 U19676 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16559), .A(n16447), .B(
        n16446), .ZN(n16448) );
  OAI211_X1 U19677 ( .C1(n17450), .C2(n16549), .A(n16449), .B(n16448), .ZN(
        P3_U2661) );
  OAI21_X1 U19678 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16464), .A(
        n16450), .ZN(n17462) );
  INV_X1 U19679 ( .A(n17462), .ZN(n16459) );
  NOR2_X1 U19680 ( .A1(n16478), .A2(n16531), .ZN(n16543) );
  NOR3_X1 U19681 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17473), .A3(
        n16514), .ZN(n16452) );
  AOI22_X1 U19682 ( .A1(n17477), .A2(n16452), .B1(n16451), .B2(n17462), .ZN(
        n16455) );
  OAI211_X1 U19683 ( .C1(n16467), .C2(n16462), .A(n16562), .B(n16453), .ZN(
        n16454) );
  OAI211_X1 U19684 ( .C1(n16455), .C2(n16531), .A(n17894), .B(n16454), .ZN(
        n16458) );
  INV_X1 U19685 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16456) );
  OAI22_X1 U19686 ( .A1(n16456), .A2(n16549), .B1(n18467), .B2(n16471), .ZN(
        n16457) );
  AOI211_X1 U19687 ( .C1(n16459), .C2(n16543), .A(n16458), .B(n16457), .ZN(
        n16461) );
  OAI211_X1 U19688 ( .C1(n16462), .C2(n16570), .A(n16461), .B(n16460), .ZN(
        P3_U2662) );
  NOR2_X1 U19689 ( .A1(n16517), .A2(n16463), .ZN(n16484) );
  AOI21_X1 U19690 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16484), .A(
        P3_REIP_REG_8__SCAN_IN), .ZN(n16472) );
  AOI21_X1 U19691 ( .B1(n17475), .B2(n16477), .A(n16464), .ZN(n17479) );
  AOI21_X1 U19692 ( .B1(n17472), .B2(n16546), .A(n16529), .ZN(n16480) );
  OAI21_X1 U19693 ( .B1(n17479), .B2(n16480), .A(n18432), .ZN(n16465) );
  AOI21_X1 U19694 ( .B1(n17479), .B2(n16480), .A(n16465), .ZN(n16466) );
  AOI211_X1 U19695 ( .C1(n16559), .C2(P3_EBX_REG_8__SCAN_IN), .A(n17896), .B(
        n16466), .ZN(n16470) );
  AOI211_X1 U19696 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16485), .A(n16467), .B(
        n16569), .ZN(n16468) );
  AOI21_X1 U19697 ( .B1(n16564), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16468), .ZN(n16469) );
  OAI211_X1 U19698 ( .C1(n16472), .C2(n16471), .A(n16470), .B(n16469), .ZN(
        P3_U2663) );
  OAI21_X1 U19699 ( .B1(n16517), .B2(n16474), .A(n16473), .ZN(n16506) );
  INV_X1 U19700 ( .A(n16506), .ZN(n16495) );
  NOR2_X1 U19701 ( .A1(n16517), .A2(n16475), .ZN(n16505) );
  INV_X1 U19702 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20750) );
  NAND3_X1 U19703 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16505), .A3(n20750), 
        .ZN(n16498) );
  NAND2_X1 U19704 ( .A1(n16495), .A2(n16498), .ZN(n16483) );
  INV_X1 U19705 ( .A(n16476), .ZN(n16490) );
  OAI21_X1 U19706 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16490), .A(
        n16477), .ZN(n16479) );
  INV_X1 U19707 ( .A(n16479), .ZN(n17498) );
  OAI21_X1 U19708 ( .B1(n17473), .B2(n16514), .A(n16478), .ZN(n16491) );
  OAI221_X1 U19709 ( .B1(n17498), .B2(n16480), .C1(n16479), .C2(n16491), .A(
        n18432), .ZN(n16481) );
  OAI211_X1 U19710 ( .C1(n16570), .C2(n16486), .A(n17894), .B(n16481), .ZN(
        n16482) );
  AOI221_X1 U19711 ( .B1(n16484), .B2(n18463), .C1(n16483), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n16482), .ZN(n16488) );
  OAI211_X1 U19712 ( .C1(n16489), .C2(n16486), .A(n16562), .B(n16485), .ZN(
        n16487) );
  OAI211_X1 U19713 ( .C1(n16549), .C2(n17492), .A(n16488), .B(n16487), .ZN(
        P3_U2664) );
  AOI211_X1 U19714 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16507), .A(n16489), .B(
        n16569), .ZN(n16497) );
  NAND2_X1 U19715 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17509), .ZN(
        n16500) );
  AOI21_X1 U19716 ( .B1(n9872), .B2(n16500), .A(n16490), .ZN(n17510) );
  NOR3_X1 U19717 ( .A1(n17510), .A2(n16531), .A3(n16491), .ZN(n16492) );
  AOI211_X1 U19718 ( .C1(n16559), .C2(P3_EBX_REG_6__SCAN_IN), .A(n17896), .B(
        n16492), .ZN(n16494) );
  OAI211_X1 U19719 ( .C1(n9872), .C2(n16529), .A(n17510), .B(n16556), .ZN(
        n16493) );
  OAI211_X1 U19720 ( .C1(n16495), .C2(n20750), .A(n16494), .B(n16493), .ZN(
        n16496) );
  AOI211_X1 U19721 ( .C1(n16564), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16497), .B(n16496), .ZN(n16499) );
  NAND2_X1 U19722 ( .A1(n16499), .A2(n16498), .ZN(P3_U2665) );
  NOR2_X1 U19723 ( .A1(n17566), .A2(n17516), .ZN(n16512) );
  OAI21_X1 U19724 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16512), .A(
        n16500), .ZN(n17520) );
  INV_X1 U19725 ( .A(n17520), .ZN(n16502) );
  AOI21_X1 U19726 ( .B1(n16571), .B2(n16512), .A(n16529), .ZN(n16501) );
  INV_X1 U19727 ( .A(n16501), .ZN(n16515) );
  AOI221_X1 U19728 ( .B1(n16502), .B2(n16515), .C1(n17520), .C2(n16501), .A(
        n17896), .ZN(n16503) );
  OAI22_X1 U19729 ( .A1(n16523), .A2(n16503), .B1(n16570), .B2(n16508), .ZN(
        n16504) );
  AOI221_X1 U19730 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n16506), .C1(n16505), 
        .C2(n16506), .A(n16504), .ZN(n16510) );
  OAI211_X1 U19731 ( .C1(n16511), .C2(n16508), .A(n16562), .B(n16507), .ZN(
        n16509) );
  OAI211_X1 U19732 ( .C1(n16549), .C2(n17515), .A(n16510), .B(n16509), .ZN(
        P3_U2666) );
  NOR2_X1 U19733 ( .A1(n16519), .A2(n16517), .ZN(n16532) );
  NOR2_X1 U19734 ( .A1(n16572), .A2(n16532), .ZN(n16534) );
  INV_X1 U19735 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18458) );
  AOI211_X1 U19736 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16537), .A(n16511), .B(
        n16569), .ZN(n16525) );
  INV_X1 U19737 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16513) );
  NAND2_X1 U19738 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17535), .ZN(
        n16527) );
  AOI21_X1 U19739 ( .B1(n16513), .B2(n16527), .A(n16512), .ZN(n17536) );
  NAND2_X1 U19740 ( .A1(n17535), .A2(n16513), .ZN(n17532) );
  OAI22_X1 U19741 ( .A1(n17536), .A2(n16515), .B1(n16514), .B2(n17532), .ZN(
        n16516) );
  AOI211_X1 U19742 ( .C1(n17536), .C2(n16529), .A(n17896), .B(n16516), .ZN(
        n16522) );
  NOR2_X1 U19743 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16517), .ZN(n16518) );
  AOI22_X1 U19744 ( .A1(n16559), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n16519), .B2(
        n16518), .ZN(n16521) );
  NOR2_X1 U19745 ( .A1(n17102), .A2(n18589), .ZN(n16558) );
  OAI21_X1 U19746 ( .B1(n16635), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16558), .ZN(n16520) );
  OAI211_X1 U19747 ( .C1(n16523), .C2(n16522), .A(n16521), .B(n16520), .ZN(
        n16524) );
  AOI211_X1 U19748 ( .C1(n16564), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16525), .B(n16524), .ZN(n16526) );
  OAI21_X1 U19749 ( .B1(n16534), .B2(n18458), .A(n16526), .ZN(P3_U2667) );
  NAND2_X1 U19750 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18366), .ZN(
        n18363) );
  INV_X1 U19751 ( .A(n18363), .ZN(n16541) );
  OAI21_X1 U19752 ( .B1(n16541), .B2(n18528), .A(n13827), .ZN(n18525) );
  NOR2_X1 U19753 ( .A1(n17566), .A2(n17560), .ZN(n16528) );
  OAI21_X1 U19754 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16528), .A(
        n16527), .ZN(n17545) );
  AOI21_X1 U19755 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16546), .A(
        n16529), .ZN(n16545) );
  XOR2_X1 U19756 ( .A(n17545), .B(n16545), .Z(n16530) );
  OAI22_X1 U19757 ( .A1(n16570), .A2(n16934), .B1(n16531), .B2(n16530), .ZN(
        n16536) );
  INV_X1 U19758 ( .A(n16532), .ZN(n16533) );
  OAI22_X1 U19759 ( .A1(n16534), .A2(n18456), .B1(n16552), .B2(n16533), .ZN(
        n16535) );
  AOI211_X1 U19760 ( .C1(n16558), .C2(n18525), .A(n16536), .B(n16535), .ZN(
        n16539) );
  OAI211_X1 U19761 ( .C1(n16542), .C2(n16934), .A(n16562), .B(n16537), .ZN(
        n16538) );
  OAI211_X1 U19762 ( .C1(n16549), .C2(n16540), .A(n16539), .B(n16538), .ZN(
        P3_U2668) );
  INV_X1 U19763 ( .A(n16558), .ZN(n18591) );
  AOI21_X1 U19764 ( .B1(n18535), .B2(n18371), .A(n16541), .ZN(n18533) );
  INV_X1 U19765 ( .A(n18533), .ZN(n16555) );
  OR2_X1 U19766 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n16560) );
  AOI211_X1 U19767 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16560), .A(n16542), .B(
        n16569), .ZN(n16551) );
  AOI22_X1 U19768 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17560), .B1(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17566), .ZN(n17556) );
  INV_X1 U19769 ( .A(n17556), .ZN(n16544) );
  AOI22_X1 U19770 ( .A1(n16572), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n16544), 
        .B2(n16543), .ZN(n16548) );
  OAI211_X1 U19771 ( .C1(n16546), .C2(n17556), .A(n18432), .B(n16545), .ZN(
        n16547) );
  OAI211_X1 U19772 ( .C1(n16549), .C2(n17560), .A(n16548), .B(n16547), .ZN(
        n16550) );
  AOI211_X1 U19773 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16559), .A(n16551), .B(
        n16550), .ZN(n16554) );
  OAI211_X1 U19774 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16561), .B(n16552), .ZN(n16553) );
  OAI211_X1 U19775 ( .C1(n18591), .C2(n16555), .A(n16554), .B(n16553), .ZN(
        P3_U2669) );
  AOI22_X1 U19776 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16572), .B1(n16556), 
        .B2(n17566), .ZN(n16568) );
  NAND2_X1 U19777 ( .A1(n18371), .A2(n16557), .ZN(n18382) );
  INV_X1 U19778 ( .A(n18382), .ZN(n18539) );
  AOI22_X1 U19779 ( .A1(n16559), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n18539), .B2(
        n16558), .ZN(n16567) );
  AND2_X1 U19780 ( .A1(n16560), .A2(n16933), .ZN(n16944) );
  AOI22_X1 U19781 ( .A1(n16562), .A2(n16944), .B1(n16561), .B2(n18551), .ZN(
        n16566) );
  OAI221_X1 U19782 ( .B1(n16564), .B2(n16563), .C1(n16564), .C2(n18432), .A(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16565) );
  NAND4_X1 U19783 ( .A1(n16568), .A2(n16567), .A3(n16566), .A4(n16565), .ZN(
        P3_U2670) );
  INV_X1 U19784 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n16946) );
  AOI21_X1 U19785 ( .B1(n16570), .B2(n16569), .A(n16946), .ZN(n16574) );
  NOR3_X1 U19786 ( .A1(n18545), .A2(n16572), .A3(n16571), .ZN(n16573) );
  AOI211_X1 U19787 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n16575), .A(n16574), .B(
        n16573), .ZN(n16576) );
  OAI21_X1 U19788 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18591), .A(
        n16576), .ZN(P3_U2671) );
  NAND2_X1 U19789 ( .A1(n16578), .A2(n16577), .ZN(n16579) );
  NAND2_X1 U19790 ( .A1(n16579), .A2(n16941), .ZN(n16678) );
  AOI22_X1 U19791 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16583) );
  AOI22_X1 U19792 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16582) );
  AOI22_X1 U19793 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16581) );
  AOI22_X1 U19794 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16580) );
  NAND4_X1 U19795 ( .A1(n16583), .A2(n16582), .A3(n16581), .A4(n16580), .ZN(
        n16589) );
  AOI22_X1 U19796 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16587) );
  AOI22_X1 U19797 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16586) );
  AOI22_X1 U19798 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16585) );
  AOI22_X1 U19799 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16584) );
  NAND4_X1 U19800 ( .A1(n16587), .A2(n16586), .A3(n16585), .A4(n16584), .ZN(
        n16588) );
  NOR2_X1 U19801 ( .A1(n16589), .A2(n16588), .ZN(n16683) );
  AOI22_X1 U19802 ( .A1(n16886), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16593) );
  AOI22_X1 U19803 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16592) );
  AOI22_X1 U19804 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16591) );
  AOI22_X1 U19805 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16590) );
  NAND4_X1 U19806 ( .A1(n16593), .A2(n16592), .A3(n16591), .A4(n16590), .ZN(
        n16599) );
  AOI22_X1 U19807 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16597) );
  AOI22_X1 U19808 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16596) );
  AOI22_X1 U19809 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16595) );
  AOI22_X1 U19810 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16594) );
  NAND4_X1 U19811 ( .A1(n16597), .A2(n16596), .A3(n16595), .A4(n16594), .ZN(
        n16598) );
  NOR2_X1 U19812 ( .A1(n16599), .A2(n16598), .ZN(n16692) );
  AOI22_X1 U19813 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16603) );
  AOI22_X1 U19814 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16602) );
  AOI22_X1 U19815 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16601) );
  AOI22_X1 U19816 ( .A1(n16886), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16600) );
  NAND4_X1 U19817 ( .A1(n16603), .A2(n16602), .A3(n16601), .A4(n16600), .ZN(
        n16609) );
  AOI22_X1 U19818 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16607) );
  AOI22_X1 U19819 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16606) );
  AOI22_X1 U19820 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16605) );
  AOI22_X1 U19821 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16604) );
  NAND4_X1 U19822 ( .A1(n16607), .A2(n16606), .A3(n16605), .A4(n16604), .ZN(
        n16608) );
  NOR2_X1 U19823 ( .A1(n16609), .A2(n16608), .ZN(n16700) );
  AOI22_X1 U19824 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16614) );
  AOI22_X1 U19825 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16613) );
  AOI22_X1 U19826 ( .A1(n16886), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16612) );
  AOI22_X1 U19827 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16610), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16611) );
  NAND4_X1 U19828 ( .A1(n16614), .A2(n16613), .A3(n16612), .A4(n16611), .ZN(
        n16620) );
  AOI22_X1 U19829 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16618) );
  AOI22_X1 U19830 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16617) );
  AOI22_X1 U19831 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16616) );
  AOI22_X1 U19832 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16615) );
  NAND4_X1 U19833 ( .A1(n16618), .A2(n16617), .A3(n16616), .A4(n16615), .ZN(
        n16619) );
  NOR2_X1 U19834 ( .A1(n16620), .A2(n16619), .ZN(n16710) );
  AOI22_X1 U19835 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16624) );
  AOI22_X1 U19836 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16623) );
  AOI22_X1 U19837 ( .A1(n16887), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16622) );
  AOI22_X1 U19838 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16621) );
  NAND4_X1 U19839 ( .A1(n16624), .A2(n16623), .A3(n16622), .A4(n16621), .ZN(
        n16631) );
  AOI22_X1 U19840 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16629) );
  AOI22_X1 U19841 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16628) );
  AOI22_X1 U19842 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16627) );
  AOI22_X1 U19843 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16626) );
  NAND4_X1 U19844 ( .A1(n16629), .A2(n16628), .A3(n16627), .A4(n16626), .ZN(
        n16630) );
  NOR2_X1 U19845 ( .A1(n16631), .A2(n16630), .ZN(n16709) );
  NOR2_X1 U19846 ( .A1(n16710), .A2(n16709), .ZN(n16705) );
  AOI22_X1 U19847 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16643) );
  INV_X1 U19848 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16634) );
  AOI22_X1 U19849 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n9598), .ZN(n16633) );
  AOI22_X1 U19850 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n16781), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n15473), .ZN(n16632) );
  OAI211_X1 U19851 ( .C1(n16634), .C2(n9596), .A(n16633), .B(n16632), .ZN(
        n16641) );
  AOI22_X1 U19852 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16639) );
  AOI22_X1 U19853 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16638) );
  AOI22_X1 U19854 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n16799), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n16888), .ZN(n16637) );
  AOI22_X1 U19855 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16635), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16636) );
  NAND4_X1 U19856 ( .A1(n16639), .A2(n16638), .A3(n16637), .A4(n16636), .ZN(
        n16640) );
  AOI211_X1 U19857 ( .C1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .C2(n9605), .A(
        n16641), .B(n16640), .ZN(n16642) );
  NAND2_X1 U19858 ( .A1(n16643), .A2(n16642), .ZN(n16704) );
  NAND2_X1 U19859 ( .A1(n16705), .A2(n16704), .ZN(n16703) );
  NOR2_X1 U19860 ( .A1(n16700), .A2(n16703), .ZN(n16698) );
  AOI22_X1 U19861 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16654) );
  INV_X1 U19862 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16646) );
  AOI22_X1 U19863 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16905), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16645) );
  AOI22_X1 U19864 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16644) );
  OAI211_X1 U19865 ( .C1(n9594), .C2(n16646), .A(n16645), .B(n16644), .ZN(
        n16652) );
  AOI22_X1 U19866 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16650) );
  AOI22_X1 U19867 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16649) );
  AOI22_X1 U19868 ( .A1(n16886), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16648) );
  AOI22_X1 U19869 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16647) );
  NAND4_X1 U19870 ( .A1(n16650), .A2(n16649), .A3(n16648), .A4(n16647), .ZN(
        n16651) );
  AOI211_X1 U19871 ( .C1(n9607), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n16652), .B(n16651), .ZN(n16653) );
  NAND2_X1 U19872 ( .A1(n16654), .A2(n16653), .ZN(n16697) );
  NAND2_X1 U19873 ( .A1(n16698), .A2(n16697), .ZN(n16696) );
  NOR2_X1 U19874 ( .A1(n16692), .A2(n16696), .ZN(n16968) );
  AOI22_X1 U19875 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16666) );
  INV_X1 U19876 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16657) );
  AOI22_X1 U19877 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16656) );
  AOI22_X1 U19878 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16655) );
  OAI211_X1 U19879 ( .C1(n9594), .C2(n16657), .A(n16656), .B(n16655), .ZN(
        n16664) );
  AOI22_X1 U19880 ( .A1(n16886), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16662) );
  AOI22_X1 U19881 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16661) );
  AOI22_X1 U19882 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16660) );
  AOI22_X1 U19883 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16659) );
  NAND4_X1 U19884 ( .A1(n16662), .A2(n16661), .A3(n16660), .A4(n16659), .ZN(
        n16663) );
  AOI211_X1 U19885 ( .C1(n9605), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n16664), .B(n16663), .ZN(n16665) );
  NAND2_X1 U19886 ( .A1(n16666), .A2(n16665), .ZN(n16967) );
  NAND2_X1 U19887 ( .A1(n16968), .A2(n16967), .ZN(n16966) );
  NOR2_X1 U19888 ( .A1(n16683), .A2(n16966), .ZN(n16682) );
  AOI22_X1 U19889 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16670) );
  AOI22_X1 U19890 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16669) );
  AOI22_X1 U19891 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16668) );
  AOI22_X1 U19892 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16667) );
  NAND4_X1 U19893 ( .A1(n16670), .A2(n16669), .A3(n16668), .A4(n16667), .ZN(
        n16676) );
  AOI22_X1 U19894 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16674) );
  AOI22_X1 U19895 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16673) );
  AOI22_X1 U19896 ( .A1(n16888), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16672) );
  AOI22_X1 U19897 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16671) );
  NAND4_X1 U19898 ( .A1(n16674), .A2(n16673), .A3(n16672), .A4(n16671), .ZN(
        n16675) );
  NOR2_X1 U19899 ( .A1(n16676), .A2(n16675), .ZN(n16677) );
  XOR2_X1 U19900 ( .A(n16682), .B(n16677), .Z(n16957) );
  OAI22_X1 U19901 ( .A1(n16679), .A2(n16678), .B1(n16957), .B2(n16941), .ZN(
        P3_U2673) );
  NOR2_X1 U19902 ( .A1(n17959), .A2(n16948), .ZN(n16947) );
  NAND2_X1 U19903 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16681) );
  NAND2_X1 U19904 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16702), .ZN(n16695) );
  AOI21_X1 U19905 ( .B1(n16683), .B2(n16966), .A(n16682), .ZN(n16961) );
  NOR2_X1 U19906 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16684), .ZN(n16685) );
  AOI22_X1 U19907 ( .A1(n16927), .A2(n16961), .B1(n16702), .B2(n16685), .ZN(
        n16686) );
  OAI21_X1 U19908 ( .B1(n16689), .B2(n16687), .A(n16686), .ZN(P3_U2674) );
  NAND2_X1 U19909 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n9709), .ZN(n16691) );
  INV_X1 U19910 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16690) );
  OAI211_X1 U19911 ( .C1(n16968), .C2(n16967), .A(n16927), .B(n16966), .ZN(
        n16688) );
  AOI21_X1 U19912 ( .B1(n16692), .B2(n16696), .A(n16968), .ZN(n16973) );
  AOI22_X1 U19913 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16693), .B1(n16927), 
        .B2(n16973), .ZN(n16694) );
  OAI21_X1 U19914 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16695), .A(n16694), .ZN(
        P3_U2676) );
  AOI21_X1 U19915 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16941), .A(n16702), .ZN(
        n16699) );
  OAI21_X1 U19916 ( .B1(n16698), .B2(n16697), .A(n16696), .ZN(n16981) );
  OAI22_X1 U19917 ( .A1(n9709), .A2(n16699), .B1(n16941), .B2(n16981), .ZN(
        P3_U2677) );
  AOI21_X1 U19918 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16941), .A(n16707), .ZN(
        n16701) );
  XNOR2_X1 U19919 ( .A(n16700), .B(n16703), .ZN(n16986) );
  OAI22_X1 U19920 ( .A1(n16702), .A2(n16701), .B1(n16941), .B2(n16986), .ZN(
        P3_U2678) );
  AOI21_X1 U19921 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16941), .A(n16712), .ZN(
        n16706) );
  OAI21_X1 U19922 ( .B1(n16705), .B2(n16704), .A(n16703), .ZN(n16991) );
  OAI22_X1 U19923 ( .A1(n16707), .A2(n16706), .B1(n16941), .B2(n16991), .ZN(
        P3_U2679) );
  AOI21_X1 U19924 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16941), .A(n16708), .ZN(
        n16711) );
  XNOR2_X1 U19925 ( .A(n16710), .B(n16709), .ZN(n16996) );
  OAI22_X1 U19926 ( .A1(n16712), .A2(n16711), .B1(n16941), .B2(n16996), .ZN(
        P3_U2680) );
  AOI22_X1 U19927 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16722) );
  AOI22_X1 U19928 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16721) );
  AOI22_X1 U19929 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16720) );
  NOR2_X1 U19930 ( .A1(n10126), .A2(n17954), .ZN(n16718) );
  AOI22_X1 U19931 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16716) );
  AOI22_X1 U19932 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16715) );
  AOI22_X1 U19933 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16714) );
  AOI22_X1 U19934 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16713) );
  NAND4_X1 U19935 ( .A1(n16716), .A2(n16715), .A3(n16714), .A4(n16713), .ZN(
        n16717) );
  AOI211_X1 U19936 ( .C1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .C2(n9609), .A(
        n16718), .B(n16717), .ZN(n16719) );
  NAND4_X1 U19937 ( .A1(n16722), .A2(n16721), .A3(n16720), .A4(n16719), .ZN(
        n16997) );
  INV_X1 U19938 ( .A(n16997), .ZN(n16724) );
  NAND3_X1 U19939 ( .A1(n16725), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n16941), 
        .ZN(n16723) );
  OAI221_X1 U19940 ( .B1(n16725), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n16941), 
        .C2(n16724), .A(n16723), .ZN(P3_U2681) );
  AOI22_X1 U19941 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16729) );
  AOI22_X1 U19942 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16728) );
  AOI22_X1 U19943 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16727) );
  AOI22_X1 U19944 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16726) );
  NAND4_X1 U19945 ( .A1(n16729), .A2(n16728), .A3(n16727), .A4(n16726), .ZN(
        n16735) );
  AOI22_X1 U19946 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16733) );
  AOI22_X1 U19947 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16732) );
  AOI22_X1 U19948 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16731) );
  AOI22_X1 U19949 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16730) );
  NAND4_X1 U19950 ( .A1(n16733), .A2(n16732), .A3(n16731), .A4(n16730), .ZN(
        n16734) );
  NOR2_X1 U19951 ( .A1(n16735), .A2(n16734), .ZN(n17003) );
  AND2_X1 U19952 ( .A1(n16941), .A2(n16736), .ZN(n16751) );
  AOI22_X1 U19953 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16751), .B1(n16738), 
        .B2(n16737), .ZN(n16739) );
  OAI21_X1 U19954 ( .B1(n17003), .B2(n16941), .A(n16739), .ZN(P3_U2682) );
  AOI22_X1 U19955 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16749) );
  AOI22_X1 U19956 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16886), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16748) );
  AOI22_X1 U19957 ( .A1(n16845), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16747) );
  AND2_X1 U19958 ( .A1(n9609), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16745) );
  AOI22_X1 U19959 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16743) );
  AOI22_X1 U19960 ( .A1(n16888), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16742) );
  AOI22_X1 U19961 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16741) );
  AOI22_X1 U19962 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16740) );
  NAND4_X1 U19963 ( .A1(n16743), .A2(n16742), .A3(n16741), .A4(n16740), .ZN(
        n16744) );
  AOI211_X1 U19964 ( .C1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .C2(n16908), .A(
        n16745), .B(n16744), .ZN(n16746) );
  NAND4_X1 U19965 ( .A1(n16749), .A2(n16748), .A3(n16747), .A4(n16746), .ZN(
        n17007) );
  INV_X1 U19966 ( .A(n17007), .ZN(n16753) );
  NOR3_X1 U19967 ( .A1(n17959), .A2(n16750), .A3(n16792), .ZN(n16765) );
  OAI221_X1 U19968 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(P3_EBX_REG_19__SCAN_IN), 
        .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16765), .A(n16751), .ZN(n16752) );
  OAI21_X1 U19969 ( .B1(n16753), .B2(n16941), .A(n16752), .ZN(P3_U2683) );
  AOI22_X1 U19970 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16757) );
  AOI22_X1 U19971 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16756) );
  AOI22_X1 U19972 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16755) );
  AOI22_X1 U19973 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16754) );
  NAND4_X1 U19974 ( .A1(n16757), .A2(n16756), .A3(n16755), .A4(n16754), .ZN(
        n16763) );
  AOI22_X1 U19975 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16761) );
  AOI22_X1 U19976 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16760) );
  AOI22_X1 U19977 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16759) );
  AOI22_X1 U19978 ( .A1(n16845), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16758) );
  NAND4_X1 U19979 ( .A1(n16761), .A2(n16760), .A3(n16759), .A4(n16758), .ZN(
        n16762) );
  NOR2_X1 U19980 ( .A1(n16763), .A2(n16762), .ZN(n17015) );
  OAI21_X1 U19981 ( .B1(n16927), .B2(n16780), .A(P3_EBX_REG_19__SCAN_IN), .ZN(
        n16764) );
  OAI21_X1 U19982 ( .B1(n16765), .B2(P3_EBX_REG_19__SCAN_IN), .A(n16764), .ZN(
        n16766) );
  OAI21_X1 U19983 ( .B1(n17015), .B2(n16941), .A(n16766), .ZN(P3_U2684) );
  NOR2_X1 U19984 ( .A1(n17959), .A2(n16792), .ZN(n16767) );
  AOI21_X1 U19985 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16941), .A(n16767), .ZN(
        n16779) );
  AOI22_X1 U19986 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16771) );
  AOI22_X1 U19987 ( .A1(n16886), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16770) );
  AOI22_X1 U19988 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16810), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16769) );
  AOI22_X1 U19989 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16768) );
  NAND4_X1 U19990 ( .A1(n16771), .A2(n16770), .A3(n16769), .A4(n16768), .ZN(
        n16778) );
  AOI22_X1 U19991 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16776) );
  AOI22_X1 U19992 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16775) );
  AOI22_X1 U19993 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16772), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U19994 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16773) );
  NAND4_X1 U19995 ( .A1(n16776), .A2(n16775), .A3(n16774), .A4(n16773), .ZN(
        n16777) );
  NOR2_X1 U19996 ( .A1(n16778), .A2(n16777), .ZN(n17019) );
  OAI22_X1 U19997 ( .A1(n16780), .A2(n16779), .B1(n17019), .B2(n16941), .ZN(
        P3_U2685) );
  AOI22_X1 U19998 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16888), .B1(
        n16781), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16785) );
  AOI22_X1 U19999 ( .A1(n16870), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n16889), .ZN(n16784) );
  AOI22_X1 U20000 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16894), .B1(
        n16886), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16783) );
  AOI22_X1 U20001 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n16869), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9598), .ZN(n16782) );
  NAND4_X1 U20002 ( .A1(n16785), .A2(n16784), .A3(n16783), .A4(n16782), .ZN(
        n16791) );
  AOI22_X1 U20003 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16789) );
  AOI22_X1 U20004 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16788) );
  AOI22_X1 U20005 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16635), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16787) );
  AOI22_X1 U20006 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9606), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n16845), .ZN(n16786) );
  NAND4_X1 U20007 ( .A1(n16789), .A2(n16788), .A3(n16787), .A4(n16786), .ZN(
        n16790) );
  NOR2_X1 U20008 ( .A1(n16791), .A2(n16790), .ZN(n17025) );
  OAI21_X1 U20009 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16793), .A(n16792), .ZN(
        n16794) );
  AOI22_X1 U20010 ( .A1(n16927), .A2(n17025), .B1(n16794), .B2(n16941), .ZN(
        P3_U2686) );
  AOI22_X1 U20011 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16798) );
  AOI22_X1 U20012 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16797) );
  AOI22_X1 U20013 ( .A1(n16781), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16796) );
  AOI22_X1 U20014 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16795) );
  NAND4_X1 U20015 ( .A1(n16798), .A2(n16797), .A3(n16796), .A4(n16795), .ZN(
        n16805) );
  AOI22_X1 U20016 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16803) );
  AOI22_X1 U20017 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16802) );
  AOI22_X1 U20018 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U20019 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16800) );
  NAND4_X1 U20020 ( .A1(n16803), .A2(n16802), .A3(n16801), .A4(n16800), .ZN(
        n16804) );
  NOR2_X1 U20021 ( .A1(n16805), .A2(n16804), .ZN(n17031) );
  INV_X1 U20022 ( .A(n16821), .ZN(n16806) );
  OAI33_X1 U20023 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17959), .A3(n16821), 
        .B1(n16807), .B2(n16927), .B3(n16806), .ZN(n16808) );
  INV_X1 U20024 ( .A(n16808), .ZN(n16809) );
  OAI21_X1 U20025 ( .B1(n17031), .B2(n16941), .A(n16809), .ZN(P3_U2687) );
  AOI22_X1 U20026 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16814) );
  AOI22_X1 U20027 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16813) );
  AOI22_X1 U20028 ( .A1(n16909), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15473), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16812) );
  AOI22_X1 U20029 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16810), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16811) );
  NAND4_X1 U20030 ( .A1(n16814), .A2(n16813), .A3(n16812), .A4(n16811), .ZN(
        n16820) );
  AOI22_X1 U20031 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16818) );
  AOI22_X1 U20032 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16817) );
  AOI22_X1 U20033 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16816) );
  AOI22_X1 U20034 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16815) );
  NAND4_X1 U20035 ( .A1(n16818), .A2(n16817), .A3(n16816), .A4(n16815), .ZN(
        n16819) );
  NOR2_X1 U20036 ( .A1(n16820), .A2(n16819), .ZN(n17035) );
  OAI211_X1 U20037 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16822), .A(n16821), .B(
        n16941), .ZN(n16823) );
  OAI21_X1 U20038 ( .B1(n17035), .B2(n16941), .A(n16823), .ZN(P3_U2688) );
  AOI22_X1 U20039 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U20040 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16886), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16833) );
  AOI22_X1 U20041 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16824) );
  OAI21_X1 U20042 ( .B1(n9639), .B2(n17954), .A(n16824), .ZN(n16831) );
  AOI22_X1 U20043 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U20044 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U20045 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16827) );
  AOI22_X1 U20046 ( .A1(n16845), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16826) );
  NAND4_X1 U20047 ( .A1(n16829), .A2(n16828), .A3(n16827), .A4(n16826), .ZN(
        n16830) );
  AOI211_X1 U20048 ( .C1(n16658), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16831), .B(n16830), .ZN(n16832) );
  NAND3_X1 U20049 ( .A1(n16834), .A2(n16833), .A3(n16832), .ZN(n17038) );
  INV_X1 U20050 ( .A(n17038), .ZN(n16840) );
  OAI221_X1 U20051 ( .B1(n16836), .B2(n16947), .C1(n16836), .C2(n16835), .A(
        P3_EBX_REG_14__SCAN_IN), .ZN(n16839) );
  NAND3_X1 U20052 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16853), .A3(n16837), 
        .ZN(n16838) );
  OAI211_X1 U20053 ( .C1(n16840), .C2(n16941), .A(n16839), .B(n16838), .ZN(
        P3_U2689) );
  AOI22_X1 U20054 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16844) );
  AOI22_X1 U20055 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16843) );
  AOI22_X1 U20056 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16842) );
  AOI22_X1 U20057 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16841) );
  NAND4_X1 U20058 ( .A1(n16844), .A2(n16843), .A3(n16842), .A4(n16841), .ZN(
        n16851) );
  AOI22_X1 U20059 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9608), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16849) );
  AOI22_X1 U20060 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U20061 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16847) );
  AOI22_X1 U20062 ( .A1(n16845), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16846) );
  NAND4_X1 U20063 ( .A1(n16849), .A2(n16848), .A3(n16847), .A4(n16846), .ZN(
        n16850) );
  NOR2_X1 U20064 ( .A1(n16851), .A2(n16850), .ZN(n17047) );
  NOR3_X1 U20065 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16927), .A3(n16865), .ZN(
        n16852) );
  AOI211_X1 U20066 ( .C1(n17047), .C2(n16927), .A(n16853), .B(n16852), .ZN(
        P3_U2691) );
  AOI22_X1 U20067 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16857) );
  AOI22_X1 U20068 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16856) );
  AOI22_X1 U20069 ( .A1(n9598), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16855) );
  AOI22_X1 U20070 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16854) );
  NAND4_X1 U20071 ( .A1(n16857), .A2(n16856), .A3(n16855), .A4(n16854), .ZN(
        n16863) );
  AOI22_X1 U20072 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20073 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16860) );
  AOI22_X1 U20074 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20075 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16858) );
  NAND4_X1 U20076 ( .A1(n16861), .A2(n16860), .A3(n16859), .A4(n16858), .ZN(
        n16862) );
  NOR2_X1 U20077 ( .A1(n16863), .A2(n16862), .ZN(n17050) );
  INV_X1 U20078 ( .A(n16864), .ZN(n16867) );
  NOR2_X1 U20079 ( .A1(n16927), .A2(n16865), .ZN(n16866) );
  OAI21_X1 U20080 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n16867), .A(n16866), .ZN(
        n16868) );
  OAI21_X1 U20081 ( .B1(n17050), .B2(n16941), .A(n16868), .ZN(P3_U2692) );
  AOI22_X1 U20082 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16876) );
  AOI22_X1 U20083 ( .A1(n16658), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16889), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U20084 ( .A1(n16871), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16870), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16874) );
  AOI22_X1 U20085 ( .A1(n16799), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16873) );
  NAND4_X1 U20086 ( .A1(n16876), .A2(n16875), .A3(n16874), .A4(n16873), .ZN(
        n16882) );
  AOI22_X1 U20087 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20088 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16635), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20089 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16878) );
  AOI22_X1 U20090 ( .A1(n16845), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16877) );
  NAND4_X1 U20091 ( .A1(n16880), .A2(n16879), .A3(n16878), .A4(n16877), .ZN(
        n16881) );
  NOR2_X1 U20092 ( .A1(n16882), .A2(n16881), .ZN(n17057) );
  NOR2_X1 U20093 ( .A1(n16927), .A2(n16884), .ZN(n16903) );
  NOR2_X1 U20094 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17959), .ZN(n16883) );
  AOI22_X1 U20095 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16903), .B1(n16884), 
        .B2(n16883), .ZN(n16885) );
  OAI21_X1 U20096 ( .B1(n17057), .B2(n16941), .A(n16885), .ZN(P3_U2693) );
  AOI22_X1 U20097 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16886), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20098 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n16869), .B1(
        n16887), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16892) );
  AOI22_X1 U20099 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n15473), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16888), .ZN(n16891) );
  AOI22_X1 U20100 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16658), .B1(
        n16825), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16890) );
  NAND4_X1 U20101 ( .A1(n16893), .A2(n16892), .A3(n16891), .A4(n16890), .ZN(
        n16901) );
  AOI22_X1 U20102 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20103 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16894), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20104 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n16909), .B1(
        n16635), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16897) );
  AOI22_X1 U20105 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16895), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16896) );
  NAND4_X1 U20106 ( .A1(n16899), .A2(n16898), .A3(n16897), .A4(n16896), .ZN(
        n16900) );
  NOR2_X1 U20107 ( .A1(n16901), .A2(n16900), .ZN(n17058) );
  INV_X1 U20108 ( .A(n16902), .ZN(n16921) );
  OAI21_X1 U20109 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16921), .A(n16903), .ZN(
        n16904) );
  OAI21_X1 U20110 ( .B1(n17058), .B2(n16941), .A(n16904), .ZN(P3_U2694) );
  AOI22_X1 U20111 ( .A1(n17036), .A2(n16925), .B1(P3_EBX_REG_8__SCAN_IN), .B2(
        n16941), .ZN(n16920) );
  AOI22_X1 U20112 ( .A1(n16825), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16888), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20113 ( .A1(n16905), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16799), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16917) );
  INV_X1 U20114 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20678) );
  AOI22_X1 U20115 ( .A1(n16869), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9598), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16906) );
  OAI21_X1 U20116 ( .B1(n16907), .B2(n20678), .A(n16906), .ZN(n16915) );
  AOI22_X1 U20117 ( .A1(n16908), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9609), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20118 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16909), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20119 ( .A1(n16635), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16871), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U20120 ( .A1(n16895), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16910) );
  NAND4_X1 U20121 ( .A1(n16913), .A2(n16912), .A3(n16911), .A4(n16910), .ZN(
        n16914) );
  AOI211_X1 U20122 ( .C1(n16658), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n16915), .B(n16914), .ZN(n16916) );
  NAND3_X1 U20123 ( .A1(n16918), .A2(n16917), .A3(n16916), .ZN(n17061) );
  INV_X1 U20124 ( .A(n17061), .ZN(n16919) );
  OAI22_X1 U20125 ( .A1(n16921), .A2(n16920), .B1(n16919), .B2(n16941), .ZN(
        P3_U2695) );
  INV_X1 U20126 ( .A(n16922), .ZN(n16923) );
  OAI21_X1 U20127 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n16923), .A(n16941), .ZN(
        n16924) );
  INV_X1 U20128 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17964) );
  OAI22_X1 U20129 ( .A1(n16925), .A2(n16924), .B1(n17964), .B2(n16941), .ZN(
        P3_U2696) );
  NAND2_X1 U20130 ( .A1(n17036), .A2(n16926), .ZN(n16929) );
  NOR2_X1 U20131 ( .A1(n16927), .A2(n16926), .ZN(n16931) );
  AOI22_X1 U20132 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n16927), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n16931), .ZN(n16928) );
  OAI21_X1 U20133 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n16929), .A(n16928), .ZN(
        P3_U2697) );
  INV_X1 U20134 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17948) );
  INV_X1 U20135 ( .A(n16930), .ZN(n16936) );
  OAI21_X1 U20136 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n16936), .A(n16931), .ZN(
        n16932) );
  OAI21_X1 U20137 ( .B1(n16941), .B2(n17948), .A(n16932), .ZN(P3_U2698) );
  INV_X1 U20138 ( .A(n16933), .ZN(n16940) );
  NAND3_X1 U20139 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n16940), .A3(n16947), .ZN(
        n16937) );
  NOR2_X1 U20140 ( .A1(n16934), .A2(n16937), .ZN(n16939) );
  AOI21_X1 U20141 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n16941), .A(n16939), .ZN(
        n16935) );
  INV_X1 U20142 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17941) );
  OAI22_X1 U20143 ( .A1(n16936), .A2(n16935), .B1(n17941), .B2(n16941), .ZN(
        P3_U2699) );
  INV_X1 U20144 ( .A(n16937), .ZN(n16943) );
  AOI21_X1 U20145 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n16941), .A(n16943), .ZN(
        n16938) );
  INV_X1 U20146 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17936) );
  OAI22_X1 U20147 ( .A1(n16939), .A2(n16938), .B1(n17936), .B2(n16941), .ZN(
        P3_U2700) );
  AOI22_X1 U20148 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n16941), .B1(n16940), .B2(
        n16947), .ZN(n16942) );
  INV_X1 U20149 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17930) );
  OAI22_X1 U20150 ( .A1(n16943), .A2(n16942), .B1(n17930), .B2(n16941), .ZN(
        P3_U2701) );
  INV_X1 U20151 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17925) );
  AOI22_X1 U20152 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n16948), .B1(n16947), .B2(
        n16944), .ZN(n16945) );
  OAI21_X1 U20153 ( .B1(n17925), .B2(n16941), .A(n16945), .ZN(P3_U2702) );
  INV_X1 U20154 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17920) );
  AOI22_X1 U20155 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16948), .B1(n16947), .B2(
        n16946), .ZN(n16949) );
  OAI21_X1 U20156 ( .B1(n17920), .B2(n16941), .A(n16949), .ZN(P3_U2703) );
  INV_X1 U20157 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17109) );
  INV_X1 U20158 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17113) );
  INV_X1 U20159 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17214) );
  NAND2_X1 U20160 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .ZN(n17067) );
  INV_X1 U20161 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17138) );
  INV_X1 U20162 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17140) );
  INV_X1 U20163 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17142) );
  NAND2_X1 U20164 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .ZN(n17037) );
  NOR4_X1 U20165 ( .A1(n17138), .A2(n17140), .A3(n17142), .A4(n17037), .ZN(
        n16951) );
  NAND4_X1 U20166 ( .A1(n17062), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n16951), .ZN(n17039) );
  INV_X1 U20167 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17119) );
  INV_X1 U20168 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17121) );
  NAND4_X1 U20169 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n16952)
         );
  NAND2_X1 U20170 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n16993), .ZN(n16992) );
  INV_X1 U20171 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17184) );
  OR2_X1 U20172 ( .A1(n16962), .A2(n17184), .ZN(n16956) );
  NOR2_X2 U20173 ( .A1(n16953), .A2(n17086), .ZN(n17026) );
  OAI21_X1 U20174 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17095), .A(n16960), .ZN(
        n16954) );
  AOI22_X1 U20175 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17026), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n16954), .ZN(n16955) );
  OAI21_X1 U20176 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n16956), .A(n16955), .ZN(
        P3_U2704) );
  NOR2_X2 U20177 ( .A1(n17943), .A2(n17086), .ZN(n17027) );
  INV_X1 U20178 ( .A(n17026), .ZN(n17002) );
  OAI22_X1 U20179 ( .A1(n16957), .A2(n17088), .B1(n12527), .B2(n17002), .ZN(
        n16958) );
  AOI21_X1 U20180 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17027), .A(n16958), .ZN(
        n16959) );
  OAI221_X1 U20181 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n16962), .C1(n17184), 
        .C2(n16960), .A(n16959), .ZN(P3_U2705) );
  AOI22_X1 U20182 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17027), .B1(n17093), .B2(
        n16961), .ZN(n16965) );
  OAI211_X1 U20183 ( .C1(n16963), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17086), .B(
        n16962), .ZN(n16964) );
  OAI211_X1 U20184 ( .C1(n17002), .C2(n14790), .A(n16965), .B(n16964), .ZN(
        P3_U2706) );
  OAI21_X1 U20185 ( .B1(n16968), .B2(n16967), .A(n16966), .ZN(n16972) );
  AOI22_X1 U20186 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17026), .ZN(n16971) );
  OAI211_X1 U20187 ( .C1(n16974), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17086), .B(
        n16969), .ZN(n16970) );
  OAI211_X1 U20188 ( .C1(n16972), .C2(n17088), .A(n16971), .B(n16970), .ZN(
        P3_U2707) );
  AOI22_X1 U20189 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17027), .B1(n17093), .B2(
        n16973), .ZN(n16977) );
  AOI211_X1 U20190 ( .C1(n17109), .C2(n16978), .A(n16974), .B(n17063), .ZN(
        n16975) );
  INV_X1 U20191 ( .A(n16975), .ZN(n16976) );
  OAI211_X1 U20192 ( .C1(n17002), .C2(n19015), .A(n16977), .B(n16976), .ZN(
        P3_U2708) );
  AOI22_X1 U20193 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17026), .ZN(n16980) );
  OAI211_X1 U20194 ( .C1(n16982), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17086), .B(
        n16978), .ZN(n16979) );
  OAI211_X1 U20195 ( .C1(n16981), .C2(n17088), .A(n16980), .B(n16979), .ZN(
        P3_U2709) );
  AOI22_X1 U20196 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17026), .ZN(n16985) );
  AOI211_X1 U20197 ( .C1(n17113), .C2(n16987), .A(n16982), .B(n17063), .ZN(
        n16983) );
  INV_X1 U20198 ( .A(n16983), .ZN(n16984) );
  OAI211_X1 U20199 ( .C1(n16986), .C2(n17088), .A(n16985), .B(n16984), .ZN(
        P3_U2710) );
  AOI22_X1 U20200 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17026), .ZN(n16990) );
  OAI211_X1 U20201 ( .C1(n16988), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17086), .B(
        n16987), .ZN(n16989) );
  OAI211_X1 U20202 ( .C1(n16991), .C2(n17088), .A(n16990), .B(n16989), .ZN(
        P3_U2711) );
  AOI22_X1 U20203 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17026), .ZN(n16995) );
  OAI211_X1 U20204 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n16993), .A(n17086), .B(
        n16992), .ZN(n16994) );
  OAI211_X1 U20205 ( .C1(n16996), .C2(n17088), .A(n16995), .B(n16994), .ZN(
        P3_U2712) );
  INV_X1 U20206 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17125) );
  INV_X1 U20207 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17169) );
  NAND2_X1 U20208 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17020), .ZN(n17016) );
  NAND2_X1 U20209 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17011), .ZN(n17006) );
  NAND2_X1 U20210 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17119), .ZN(n17001) );
  AOI22_X1 U20211 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17026), .B1(n17093), .B2(
        n16997), .ZN(n17000) );
  NAND2_X1 U20212 ( .A1(n17086), .A2(n17006), .ZN(n17010) );
  OAI21_X1 U20213 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17095), .A(n17010), .ZN(
        n16998) );
  AOI22_X1 U20214 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17027), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n16998), .ZN(n16999) );
  OAI211_X1 U20215 ( .C1(n17006), .C2(n17001), .A(n17000), .B(n16999), .ZN(
        P3_U2713) );
  OAI22_X1 U20216 ( .A1(n17003), .A2(n17088), .B1(n17944), .B2(n17002), .ZN(
        n17004) );
  AOI21_X1 U20217 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17027), .A(n17004), .ZN(
        n17005) );
  OAI221_X1 U20218 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17006), .C1(n17121), 
        .C2(n17010), .A(n17005), .ZN(P3_U2714) );
  INV_X1 U20219 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U20220 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17026), .B1(n17093), .B2(
        n17007), .ZN(n17009) );
  AOI22_X1 U20221 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17027), .B1(n17011), .B2(
        n17123), .ZN(n17008) );
  OAI211_X1 U20222 ( .C1(n17123), .C2(n17010), .A(n17009), .B(n17008), .ZN(
        P3_U2715) );
  AOI22_X1 U20223 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17026), .ZN(n17014) );
  AOI211_X1 U20224 ( .C1(n17125), .C2(n17016), .A(n17011), .B(n17063), .ZN(
        n17012) );
  INV_X1 U20225 ( .A(n17012), .ZN(n17013) );
  OAI211_X1 U20226 ( .C1(n17015), .C2(n17088), .A(n17014), .B(n17013), .ZN(
        P3_U2716) );
  AOI22_X1 U20227 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17026), .ZN(n17018) );
  OAI211_X1 U20228 ( .C1(n17020), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17086), .B(
        n17016), .ZN(n17017) );
  OAI211_X1 U20229 ( .C1(n17019), .C2(n17088), .A(n17018), .B(n17017), .ZN(
        P3_U2717) );
  AOI22_X1 U20230 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17026), .ZN(n17024) );
  INV_X1 U20231 ( .A(n17028), .ZN(n17022) );
  INV_X1 U20232 ( .A(n17020), .ZN(n17021) );
  OAI211_X1 U20233 ( .C1(n17022), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17086), .B(
        n17021), .ZN(n17023) );
  OAI211_X1 U20234 ( .C1(n17025), .C2(n17088), .A(n17024), .B(n17023), .ZN(
        P3_U2718) );
  AOI22_X1 U20235 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17027), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17026), .ZN(n17030) );
  OAI211_X1 U20236 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17032), .A(n17086), .B(
        n17028), .ZN(n17029) );
  OAI211_X1 U20237 ( .C1(n17031), .C2(n17088), .A(n17030), .B(n17029), .ZN(
        P3_U2719) );
  AOI21_X1 U20238 ( .B1(n17214), .B2(n17039), .A(n17032), .ZN(n17033) );
  AOI22_X1 U20239 ( .A1(n17094), .A2(BUF2_REG_15__SCAN_IN), .B1(n17033), .B2(
        n17086), .ZN(n17034) );
  OAI21_X1 U20240 ( .B1(n17035), .B2(n17088), .A(n17034), .ZN(P3_U2720) );
  NAND2_X1 U20241 ( .A1(n17036), .A2(n17062), .ZN(n17066) );
  NOR2_X1 U20242 ( .A1(n17037), .A2(n17066), .ZN(n17060) );
  INV_X1 U20243 ( .A(n17060), .ZN(n17054) );
  NOR2_X1 U20244 ( .A1(n17142), .A2(n17054), .ZN(n17053) );
  NAND2_X1 U20245 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17053), .ZN(n17046) );
  NOR2_X1 U20246 ( .A1(n17138), .A2(n17046), .ZN(n17049) );
  NAND2_X1 U20247 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17049), .ZN(n17042) );
  AOI22_X1 U20248 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17094), .B1(n17093), .B2(
        n17038), .ZN(n17041) );
  NAND3_X1 U20249 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17086), .A3(n17039), 
        .ZN(n17040) );
  OAI211_X1 U20250 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17042), .A(n17041), .B(
        n17040), .ZN(P3_U2721) );
  INV_X1 U20251 ( .A(n17042), .ZN(n17045) );
  AOI21_X1 U20252 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17086), .A(n17049), .ZN(
        n17044) );
  OAI222_X1 U20253 ( .A1(n17091), .A2(n17208), .B1(n17045), .B2(n17044), .C1(
        n17088), .C2(n17043), .ZN(P3_U2722) );
  INV_X1 U20254 ( .A(n17046), .ZN(n17052) );
  AOI21_X1 U20255 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17086), .A(n17052), .ZN(
        n17048) );
  OAI222_X1 U20256 ( .A1(n17091), .A2(n17204), .B1(n17049), .B2(n17048), .C1(
        n17088), .C2(n17047), .ZN(P3_U2723) );
  AOI21_X1 U20257 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17086), .A(n17053), .ZN(
        n17051) );
  OAI222_X1 U20258 ( .A1(n17091), .A2(n17202), .B1(n17052), .B2(n17051), .C1(
        n17088), .C2(n17050), .ZN(P3_U2724) );
  AOI21_X1 U20259 ( .B1(n17142), .B2(n17054), .A(n17053), .ZN(n17055) );
  AOI22_X1 U20260 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17094), .B1(n17055), .B2(
        n17086), .ZN(n17056) );
  OAI21_X1 U20261 ( .B1(n17057), .B2(n17088), .A(n17056), .ZN(P3_U2725) );
  INV_X1 U20262 ( .A(n17066), .ZN(n17070) );
  AOI22_X1 U20263 ( .A1(n17070), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17086), .ZN(n17059) );
  OAI222_X1 U20264 ( .A1(n17091), .A2(n17198), .B1(n17060), .B2(n17059), .C1(
        n17088), .C2(n17058), .ZN(P3_U2726) );
  AOI22_X1 U20265 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17094), .B1(n17093), .B2(
        n17061), .ZN(n17065) );
  INV_X1 U20266 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17146) );
  OR3_X1 U20267 ( .A1(n17146), .A2(n17063), .A3(n17062), .ZN(n17064) );
  OAI211_X1 U20268 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n17066), .A(n17065), .B(
        n17064), .ZN(P3_U2727) );
  INV_X1 U20269 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17156) );
  INV_X1 U20270 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17187) );
  NOR3_X1 U20271 ( .A1(n17187), .A2(n17163), .A3(n17095), .ZN(n17085) );
  NAND2_X1 U20272 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17085), .ZN(n17081) );
  NOR2_X1 U20273 ( .A1(n17156), .A2(n17081), .ZN(n17084) );
  NAND2_X1 U20274 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17084), .ZN(n17074) );
  NOR2_X1 U20275 ( .A1(n17067), .A2(n17074), .ZN(n17073) );
  AOI21_X1 U20276 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17086), .A(n17073), .ZN(
        n17069) );
  OAI222_X1 U20277 ( .A1(n17091), .A2(n17955), .B1(n17070), .B2(n17069), .C1(
        n17088), .C2(n17068), .ZN(P3_U2728) );
  INV_X1 U20278 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20708) );
  NOR2_X1 U20279 ( .A1(n20708), .A2(n17074), .ZN(n17077) );
  AOI21_X1 U20280 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17086), .A(n17077), .ZN(
        n17072) );
  OAI222_X1 U20281 ( .A1(n17949), .A2(n17091), .B1(n17073), .B2(n17072), .C1(
        n17088), .C2(n17071), .ZN(P3_U2729) );
  INV_X1 U20282 ( .A(n17074), .ZN(n17080) );
  AOI21_X1 U20283 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17086), .A(n17080), .ZN(
        n17076) );
  OAI222_X1 U20284 ( .A1(n17942), .A2(n17091), .B1(n17077), .B2(n17076), .C1(
        n17088), .C2(n17075), .ZN(P3_U2730) );
  AOI21_X1 U20285 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17086), .A(n17084), .ZN(
        n17079) );
  OAI222_X1 U20286 ( .A1(n17937), .A2(n17091), .B1(n17080), .B2(n17079), .C1(
        n17088), .C2(n17078), .ZN(P3_U2731) );
  INV_X1 U20287 ( .A(n17081), .ZN(n17090) );
  AOI21_X1 U20288 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17086), .A(n17090), .ZN(
        n17083) );
  OAI222_X1 U20289 ( .A1(n17931), .A2(n17091), .B1(n17084), .B2(n17083), .C1(
        n17088), .C2(n17082), .ZN(P3_U2732) );
  AOI21_X1 U20290 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17086), .A(n17085), .ZN(
        n17089) );
  OAI222_X1 U20291 ( .A1(n17926), .A2(n17091), .B1(n17090), .B2(n17089), .C1(
        n17088), .C2(n17087), .ZN(P3_U2733) );
  AOI22_X1 U20292 ( .A1(n17094), .A2(BUF2_REG_1__SCAN_IN), .B1(n17093), .B2(
        n17092), .ZN(n17100) );
  NOR2_X1 U20293 ( .A1(n17163), .A2(n17095), .ZN(n17098) );
  NOR2_X1 U20294 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17095), .ZN(n17097) );
  OAI22_X1 U20295 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17098), .B1(n17097), .B2(
        n17096), .ZN(n17099) );
  NAND2_X1 U20296 ( .A1(n17100), .A2(n17099), .ZN(P3_U2734) );
  NOR2_X4 U20297 ( .A1(n17160), .A2(n17132), .ZN(n17149) );
  AND2_X1 U20298 ( .A1(n17149), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20299 ( .A1(n17132), .A2(n17102), .ZN(n17130) );
  AOI22_X1 U20300 ( .A1(n17160), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17103) );
  OAI21_X1 U20301 ( .B1(n17184), .B2(n17130), .A(n17103), .ZN(P3_U2737) );
  INV_X1 U20302 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20303 ( .A1(n17160), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17104) );
  OAI21_X1 U20304 ( .B1(n17105), .B2(n17130), .A(n17104), .ZN(P3_U2738) );
  INV_X1 U20305 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U20306 ( .A1(n17160), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17106) );
  OAI21_X1 U20307 ( .B1(n17107), .B2(n17130), .A(n17106), .ZN(P3_U2739) );
  AOI22_X1 U20308 ( .A1(n17160), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17108) );
  OAI21_X1 U20309 ( .B1(n17109), .B2(n17130), .A(n17108), .ZN(P3_U2740) );
  INV_X1 U20310 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17111) );
  INV_X2 U20311 ( .A(n18570), .ZN(n17160) );
  AOI22_X1 U20312 ( .A1(n17160), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17110) );
  OAI21_X1 U20313 ( .B1(n17111), .B2(n17130), .A(n17110), .ZN(P3_U2741) );
  AOI22_X1 U20314 ( .A1(n17160), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17112) );
  OAI21_X1 U20315 ( .B1(n17113), .B2(n17130), .A(n17112), .ZN(P3_U2742) );
  INV_X1 U20316 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20317 ( .A1(n17160), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17114) );
  OAI21_X1 U20318 ( .B1(n17115), .B2(n17130), .A(n17114), .ZN(P3_U2743) );
  INV_X1 U20319 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20320 ( .A1(n17160), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17116) );
  OAI21_X1 U20321 ( .B1(n17117), .B2(n17130), .A(n17116), .ZN(P3_U2744) );
  AOI22_X1 U20322 ( .A1(n17160), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17118) );
  OAI21_X1 U20323 ( .B1(n17119), .B2(n17130), .A(n17118), .ZN(P3_U2745) );
  AOI22_X1 U20324 ( .A1(n17160), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17120) );
  OAI21_X1 U20325 ( .B1(n17121), .B2(n17130), .A(n17120), .ZN(P3_U2746) );
  AOI22_X1 U20326 ( .A1(P3_DATAO_REG_20__SCAN_IN), .A2(n17149), .B1(n17160), 
        .B2(P3_UWORD_REG_4__SCAN_IN), .ZN(n17122) );
  OAI21_X1 U20327 ( .B1(n17123), .B2(n17130), .A(n17122), .ZN(P3_U2747) );
  AOI22_X1 U20328 ( .A1(n17160), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17124) );
  OAI21_X1 U20329 ( .B1(n17125), .B2(n17130), .A(n17124), .ZN(P3_U2748) );
  INV_X1 U20330 ( .A(P3_UWORD_REG_2__SCAN_IN), .ZN(n20768) );
  INV_X1 U20331 ( .A(n17130), .ZN(n17126) );
  AOI22_X1 U20332 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17126), .B1(n17149), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17127) );
  OAI21_X1 U20333 ( .B1(n20768), .B2(n18570), .A(n17127), .ZN(P3_U2749) );
  AOI22_X1 U20334 ( .A1(n17160), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17128) );
  OAI21_X1 U20335 ( .B1(n17169), .B2(n17130), .A(n17128), .ZN(P3_U2750) );
  INV_X1 U20336 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20337 ( .A1(n17160), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17129) );
  OAI21_X1 U20338 ( .B1(n17131), .B2(n17130), .A(n17129), .ZN(P3_U2751) );
  AOI22_X1 U20339 ( .A1(n17160), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17133) );
  OAI21_X1 U20340 ( .B1(n17214), .B2(n17162), .A(n17133), .ZN(P3_U2752) );
  INV_X1 U20341 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20342 ( .A1(n17160), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17134) );
  OAI21_X1 U20343 ( .B1(n17210), .B2(n17162), .A(n17134), .ZN(P3_U2753) );
  INV_X1 U20344 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20345 ( .A1(n17160), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17135) );
  OAI21_X1 U20346 ( .B1(n17136), .B2(n17162), .A(n17135), .ZN(P3_U2754) );
  AOI22_X1 U20347 ( .A1(n17160), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17137) );
  OAI21_X1 U20348 ( .B1(n17138), .B2(n17162), .A(n17137), .ZN(P3_U2755) );
  AOI22_X1 U20349 ( .A1(n17160), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17139) );
  OAI21_X1 U20350 ( .B1(n17140), .B2(n17162), .A(n17139), .ZN(P3_U2756) );
  AOI22_X1 U20351 ( .A1(n17160), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17141) );
  OAI21_X1 U20352 ( .B1(n17142), .B2(n17162), .A(n17141), .ZN(P3_U2757) );
  INV_X1 U20353 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20354 ( .A1(n17160), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17143) );
  OAI21_X1 U20355 ( .B1(n17144), .B2(n17162), .A(n17143), .ZN(P3_U2758) );
  AOI22_X1 U20356 ( .A1(n17160), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17145) );
  OAI21_X1 U20357 ( .B1(n17146), .B2(n17162), .A(n17145), .ZN(P3_U2759) );
  INV_X1 U20358 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20359 ( .A1(n17160), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17147) );
  OAI21_X1 U20360 ( .B1(n17148), .B2(n17162), .A(n17147), .ZN(P3_U2760) );
  INV_X1 U20361 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20362 ( .A1(n17160), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17150) );
  OAI21_X1 U20363 ( .B1(n17151), .B2(n17162), .A(n17150), .ZN(P3_U2761) );
  AOI22_X1 U20364 ( .A1(n17160), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17152) );
  OAI21_X1 U20365 ( .B1(n20708), .B2(n17162), .A(n17152), .ZN(P3_U2762) );
  INV_X1 U20366 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20367 ( .A1(n17160), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17153) );
  OAI21_X1 U20368 ( .B1(n17154), .B2(n17162), .A(n17153), .ZN(P3_U2763) );
  AOI22_X1 U20369 ( .A1(n17160), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17155) );
  OAI21_X1 U20370 ( .B1(n17156), .B2(n17162), .A(n17155), .ZN(P3_U2764) );
  INV_X1 U20371 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20372 ( .A1(n17160), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17157) );
  OAI21_X1 U20373 ( .B1(n17158), .B2(n17162), .A(n17157), .ZN(P3_U2765) );
  AOI22_X1 U20374 ( .A1(P3_LWORD_REG_1__SCAN_IN), .A2(n17160), .B1(n17149), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17159) );
  OAI21_X1 U20375 ( .B1(n17187), .B2(n17162), .A(n17159), .ZN(P3_U2766) );
  AOI22_X1 U20376 ( .A1(n17160), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17149), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17161) );
  OAI21_X1 U20377 ( .B1(n17163), .B2(n17162), .A(n17161), .ZN(P3_U2767) );
  NAND2_X2 U20378 ( .A1(n17166), .A2(n17922), .ZN(n17207) );
  AOI22_X1 U20379 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17205), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17196), .ZN(n17167) );
  OAI21_X1 U20380 ( .B1(n17913), .B2(n17207), .A(n17167), .ZN(P3_U2768) );
  AOI22_X1 U20381 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17211), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17196), .ZN(n17168) );
  OAI21_X1 U20382 ( .B1(n17169), .B2(n17213), .A(n17168), .ZN(P3_U2769) );
  AOI22_X1 U20383 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17205), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17196), .ZN(n17170) );
  OAI21_X1 U20384 ( .B1(n17926), .B2(n17207), .A(n17170), .ZN(P3_U2770) );
  AOI22_X1 U20385 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17205), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17196), .ZN(n17171) );
  OAI21_X1 U20386 ( .B1(n17931), .B2(n17207), .A(n17171), .ZN(P3_U2771) );
  AOI22_X1 U20387 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17179), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17196), .ZN(n17172) );
  OAI21_X1 U20388 ( .B1(n17937), .B2(n17207), .A(n17172), .ZN(P3_U2772) );
  AOI22_X1 U20389 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17179), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17196), .ZN(n17173) );
  OAI21_X1 U20390 ( .B1(n17942), .B2(n17207), .A(n17173), .ZN(P3_U2773) );
  AOI22_X1 U20391 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17179), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17196), .ZN(n17174) );
  OAI21_X1 U20392 ( .B1(n17949), .B2(n17207), .A(n17174), .ZN(P3_U2774) );
  AOI22_X1 U20393 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17179), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17196), .ZN(n17175) );
  OAI21_X1 U20394 ( .B1(n17955), .B2(n17207), .A(n17175), .ZN(P3_U2775) );
  AOI22_X1 U20395 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17179), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17196), .ZN(n17176) );
  OAI21_X1 U20396 ( .B1(n17195), .B2(n17207), .A(n17176), .ZN(P3_U2776) );
  AOI22_X1 U20397 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17179), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17196), .ZN(n17177) );
  OAI21_X1 U20398 ( .B1(n17198), .B2(n17207), .A(n17177), .ZN(P3_U2777) );
  AOI22_X1 U20399 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17179), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17196), .ZN(n17178) );
  OAI21_X1 U20400 ( .B1(n17200), .B2(n17207), .A(n17178), .ZN(P3_U2778) );
  AOI22_X1 U20401 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17179), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17196), .ZN(n17180) );
  OAI21_X1 U20402 ( .B1(n17202), .B2(n17207), .A(n17180), .ZN(P3_U2779) );
  AOI22_X1 U20403 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17205), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17196), .ZN(n17181) );
  OAI21_X1 U20404 ( .B1(n17204), .B2(n17207), .A(n17181), .ZN(P3_U2780) );
  AOI22_X1 U20405 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17205), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17196), .ZN(n17182) );
  OAI21_X1 U20406 ( .B1(n17208), .B2(n17207), .A(n17182), .ZN(P3_U2781) );
  AOI22_X1 U20407 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17211), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17196), .ZN(n17183) );
  OAI21_X1 U20408 ( .B1(n17184), .B2(n17213), .A(n17183), .ZN(P3_U2782) );
  AOI22_X1 U20409 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17196), .ZN(n17185) );
  OAI21_X1 U20410 ( .B1(n17913), .B2(n17207), .A(n17185), .ZN(P3_U2783) );
  AOI22_X1 U20411 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17211), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17196), .ZN(n17186) );
  OAI21_X1 U20412 ( .B1(n17187), .B2(n17213), .A(n17186), .ZN(P3_U2784) );
  AOI22_X1 U20413 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17196), .ZN(n17188) );
  OAI21_X1 U20414 ( .B1(n17926), .B2(n17207), .A(n17188), .ZN(P3_U2785) );
  AOI22_X1 U20415 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17196), .ZN(n17189) );
  OAI21_X1 U20416 ( .B1(n17931), .B2(n17207), .A(n17189), .ZN(P3_U2786) );
  AOI22_X1 U20417 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17196), .ZN(n17190) );
  OAI21_X1 U20418 ( .B1(n17937), .B2(n17207), .A(n17190), .ZN(P3_U2787) );
  AOI22_X1 U20419 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17196), .ZN(n17191) );
  OAI21_X1 U20420 ( .B1(n17942), .B2(n17207), .A(n17191), .ZN(P3_U2788) );
  AOI22_X1 U20421 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17196), .ZN(n17192) );
  OAI21_X1 U20422 ( .B1(n17949), .B2(n17207), .A(n17192), .ZN(P3_U2789) );
  AOI22_X1 U20423 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17196), .ZN(n17193) );
  OAI21_X1 U20424 ( .B1(n17955), .B2(n17207), .A(n17193), .ZN(P3_U2790) );
  AOI22_X1 U20425 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17196), .ZN(n17194) );
  OAI21_X1 U20426 ( .B1(n17195), .B2(n17207), .A(n17194), .ZN(P3_U2791) );
  AOI22_X1 U20427 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17196), .ZN(n17197) );
  OAI21_X1 U20428 ( .B1(n17198), .B2(n17207), .A(n17197), .ZN(P3_U2792) );
  AOI22_X1 U20429 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17196), .ZN(n17199) );
  OAI21_X1 U20430 ( .B1(n17200), .B2(n17207), .A(n17199), .ZN(P3_U2793) );
  AOI22_X1 U20431 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17196), .ZN(n17201) );
  OAI21_X1 U20432 ( .B1(n17202), .B2(n17207), .A(n17201), .ZN(P3_U2794) );
  AOI22_X1 U20433 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17196), .ZN(n17203) );
  OAI21_X1 U20434 ( .B1(n17204), .B2(n17207), .A(n17203), .ZN(P3_U2795) );
  AOI22_X1 U20435 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17205), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17196), .ZN(n17206) );
  OAI21_X1 U20436 ( .B1(n17208), .B2(n17207), .A(n17206), .ZN(P3_U2796) );
  AOI22_X1 U20437 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17211), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17196), .ZN(n17209) );
  OAI21_X1 U20438 ( .B1(n17210), .B2(n17213), .A(n17209), .ZN(P3_U2797) );
  AOI22_X1 U20439 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17211), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17196), .ZN(n17212) );
  OAI21_X1 U20440 ( .B1(n17214), .B2(n17213), .A(n17212), .ZN(P3_U2798) );
  OAI21_X1 U20441 ( .B1(n17215), .B2(n17574), .A(n17573), .ZN(n17216) );
  AOI21_X1 U20442 ( .B1(n17474), .B2(n17218), .A(n17216), .ZN(n17246) );
  OAI21_X1 U20443 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17359), .A(
        n17246), .ZN(n17236) );
  AOI22_X1 U20444 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17236), .B1(
        n9610), .B2(n17217), .ZN(n17221) );
  NOR2_X1 U20445 ( .A1(n17334), .A2(n17218), .ZN(n17238) );
  OAI211_X1 U20446 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17238), .B(n17219), .ZN(n17220) );
  NAND2_X1 U20447 ( .A1(n17221), .A2(n17220), .ZN(n17222) );
  AOI211_X1 U20448 ( .C1(n17224), .C2(n17382), .A(n17223), .B(n17222), .ZN(
        n17231) );
  NAND2_X1 U20449 ( .A1(n17578), .A2(n17421), .ZN(n17320) );
  AOI22_X1 U20450 ( .A1(n17565), .A2(n17582), .B1(n17485), .B2(n17225), .ZN(
        n17254) );
  NAND2_X1 U20451 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17254), .ZN(
        n17240) );
  NAND3_X1 U20452 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17320), .A3(
        n17240), .ZN(n17230) );
  OAI211_X1 U20453 ( .C1(n17228), .C2(n17227), .A(n17484), .B(n17226), .ZN(
        n17229) );
  NAND3_X1 U20454 ( .A1(n17231), .A2(n17230), .A3(n17229), .ZN(P3_U2802) );
  NAND2_X1 U20455 ( .A1(n16069), .A2(n17232), .ZN(n17233) );
  XNOR2_X1 U20456 ( .A(n17312), .B(n17233), .ZN(n17591) );
  OAI22_X1 U20457 ( .A1(n17894), .A2(n18503), .B1(n9591), .B2(n17234), .ZN(
        n17235) );
  AOI221_X1 U20458 ( .B1(n17238), .B2(n17237), .C1(n17236), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17235), .ZN(n17243) );
  INV_X1 U20459 ( .A(n17239), .ZN(n17241) );
  OAI21_X1 U20460 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17241), .A(
        n17240), .ZN(n17242) );
  OAI211_X1 U20461 ( .C1(n17591), .C2(n17458), .A(n17243), .B(n17242), .ZN(
        P3_U2803) );
  AOI21_X1 U20462 ( .B1(n17244), .B2(n18299), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17245) );
  INV_X1 U20463 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18501) );
  OAI22_X1 U20464 ( .A1(n17246), .A2(n17245), .B1(n17894), .B2(n18501), .ZN(
        n17247) );
  AOI221_X1 U20465 ( .B1(n9610), .B2(n17248), .C1(n17325), .C2(n17248), .A(
        n17247), .ZN(n17252) );
  OAI21_X1 U20466 ( .B1(n17250), .B2(n17253), .A(n17249), .ZN(n17593) );
  NOR3_X1 U20467 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17599), .A3(
        n17601), .ZN(n17592) );
  AOI22_X1 U20468 ( .A1(n17484), .A2(n17593), .B1(n17382), .B2(n17592), .ZN(
        n17251) );
  OAI211_X1 U20469 ( .C1(n17254), .C2(n17253), .A(n17252), .B(n17251), .ZN(
        P3_U2804) );
  XNOR2_X1 U20470 ( .A(n17255), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17612) );
  INV_X1 U20471 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17273) );
  OAI21_X1 U20472 ( .B1(n17256), .B2(n17574), .A(n17573), .ZN(n17257) );
  AOI21_X1 U20473 ( .B1(n18299), .B2(n17258), .A(n17257), .ZN(n17283) );
  OAI21_X1 U20474 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17359), .A(
        n17283), .ZN(n17272) );
  NOR2_X1 U20475 ( .A1(n17334), .A2(n17258), .ZN(n17274) );
  AOI22_X1 U20476 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17272), .B1(
        n17274), .B2(n17259), .ZN(n17260) );
  AOI21_X1 U20477 ( .B1(n17273), .B2(n17261), .A(n17260), .ZN(n17262) );
  NOR2_X1 U20478 ( .A1(n17894), .A2(n18499), .ZN(n17607) );
  AOI211_X1 U20479 ( .C1(n9610), .C2(n17263), .A(n17262), .B(n17607), .ZN(
        n17269) );
  XNOR2_X1 U20480 ( .A(n17599), .B(n17264), .ZN(n17609) );
  OAI21_X1 U20481 ( .B1(n17312), .B2(n17266), .A(n17265), .ZN(n17267) );
  XNOR2_X1 U20482 ( .A(n17267), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17608) );
  AOI22_X1 U20483 ( .A1(n17485), .A2(n17609), .B1(n17484), .B2(n17608), .ZN(
        n17268) );
  OAI211_X1 U20484 ( .C1(n17578), .C2(n17612), .A(n17269), .B(n17268), .ZN(
        P3_U2805) );
  INV_X1 U20485 ( .A(n17382), .ZN(n17315) );
  OR2_X1 U20486 ( .A1(n17614), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17626) );
  OAI22_X1 U20487 ( .A1(n17894), .A2(n18496), .B1(n9591), .B2(n17270), .ZN(
        n17271) );
  AOI221_X1 U20488 ( .B1(n17274), .B2(n17273), .C1(n17272), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17271), .ZN(n17277) );
  OAI21_X1 U20489 ( .B1(n17614), .B2(n17636), .A(n17485), .ZN(n17286) );
  OAI21_X1 U20490 ( .B1(n17638), .B2(n17614), .A(n17565), .ZN(n17287) );
  NAND2_X1 U20491 ( .A1(n17286), .A2(n17287), .ZN(n17289) );
  AOI22_X1 U20492 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17289), .B1(
        n17484), .B2(n17623), .ZN(n17276) );
  OAI211_X1 U20493 ( .C1(n17315), .C2(n17626), .A(n17277), .B(n17276), .ZN(
        P3_U2806) );
  OAI22_X1 U20494 ( .A1(n17312), .A2(n17643), .B1(n17278), .B2(n17295), .ZN(
        n17279) );
  NOR2_X1 U20495 ( .A1(n17279), .A2(n17327), .ZN(n17280) );
  XNOR2_X1 U20496 ( .A(n17280), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17633) );
  AOI21_X1 U20497 ( .B1(n18299), .B2(n17281), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17282) );
  OAI22_X1 U20498 ( .A1(n17283), .A2(n17282), .B1(n17894), .B2(n18495), .ZN(
        n17284) );
  AOI221_X1 U20499 ( .B1(n9610), .B2(n17285), .C1(n17325), .C2(n17285), .A(
        n17284), .ZN(n17291) );
  OAI22_X1 U20500 ( .A1(n17638), .A2(n17287), .B1(n17636), .B2(n17286), .ZN(
        n17288) );
  AOI22_X1 U20501 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17289), .B1(
        n17627), .B2(n17288), .ZN(n17290) );
  OAI211_X1 U20502 ( .C1(n17458), .C2(n17633), .A(n17291), .B(n17290), .ZN(
        P3_U2807) );
  OAI21_X1 U20503 ( .B1(n17292), .B2(n17574), .A(n17573), .ZN(n17293) );
  AOI21_X1 U20504 ( .B1(n17474), .B2(n17301), .A(n17293), .ZN(n17323) );
  OAI21_X1 U20505 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17359), .A(
        n17323), .ZN(n17308) );
  AOI22_X1 U20506 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17308), .B1(
        n9610), .B2(n17294), .ZN(n17305) );
  INV_X1 U20507 ( .A(n17295), .ZN(n17296) );
  INV_X1 U20508 ( .A(n17635), .ZN(n17652) );
  NAND2_X1 U20509 ( .A1(n17652), .A2(n17642), .ZN(n17641) );
  AOI221_X1 U20510 ( .B1(n17369), .B2(n17296), .C1(n17641), .C2(n17296), .A(
        n17327), .ZN(n17297) );
  XNOR2_X1 U20511 ( .A(n17297), .B(n17643), .ZN(n17646) );
  NOR2_X1 U20512 ( .A1(n17315), .A2(n17641), .ZN(n17299) );
  INV_X1 U20513 ( .A(n17638), .ZN(n17717) );
  OAI22_X1 U20514 ( .A1(n17717), .A2(n17578), .B1(n17710), .B2(n17421), .ZN(
        n17381) );
  AOI21_X1 U20515 ( .B1(n17320), .B2(n17641), .A(n17381), .ZN(n17319) );
  INV_X1 U20516 ( .A(n17319), .ZN(n17298) );
  MUX2_X1 U20517 ( .A(n17299), .B(n17298), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17300) );
  AOI21_X1 U20518 ( .B1(n17484), .B2(n17646), .A(n17300), .ZN(n17304) );
  NAND2_X1 U20519 ( .A1(n17896), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17647) );
  NOR2_X1 U20520 ( .A1(n17334), .A2(n17301), .ZN(n17310) );
  OAI211_X1 U20521 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17310), .B(n17302), .ZN(n17303) );
  NAND4_X1 U20522 ( .A1(n17305), .A2(n17304), .A3(n17647), .A4(n17303), .ZN(
        P3_U2808) );
  OAI22_X1 U20523 ( .A1(n17894), .A2(n18491), .B1(n9591), .B2(n17306), .ZN(
        n17307) );
  AOI221_X1 U20524 ( .B1(n17310), .B2(n17309), .C1(n17308), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17307), .ZN(n17317) );
  NAND3_X1 U20525 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17312), .A3(
        n17311), .ZN(n17339) );
  INV_X1 U20526 ( .A(n17353), .ZN(n17340) );
  OAI22_X1 U20527 ( .A1(n17651), .A2(n17339), .B1(n17340), .B2(n17313), .ZN(
        n17314) );
  XNOR2_X1 U20528 ( .A(n17318), .B(n17314), .ZN(n17659) );
  NOR2_X1 U20529 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17651), .ZN(
        n17658) );
  NOR2_X1 U20530 ( .A1(n17635), .A2(n17315), .ZN(n17342) );
  AOI22_X1 U20531 ( .A1(n17484), .A2(n17659), .B1(n17658), .B2(n17342), .ZN(
        n17316) );
  OAI211_X1 U20532 ( .C1(n17319), .C2(n17318), .A(n17317), .B(n17316), .ZN(
        P3_U2809) );
  NAND2_X1 U20533 ( .A1(n17652), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17666) );
  AOI21_X1 U20534 ( .B1(n17320), .B2(n17666), .A(n17381), .ZN(n17346) );
  INV_X1 U20535 ( .A(n17359), .ZN(n17325) );
  AOI21_X1 U20536 ( .B1(n17321), .B2(n18299), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17322) );
  OAI22_X1 U20537 ( .A1(n17323), .A2(n17322), .B1(n17894), .B2(n18488), .ZN(
        n17324) );
  AOI221_X1 U20538 ( .B1(n9610), .B2(n17326), .C1(n17325), .C2(n17326), .A(
        n17324), .ZN(n17330) );
  INV_X1 U20539 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17345) );
  AOI221_X1 U20540 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17339), 
        .C1(n17345), .C2(n17352), .A(n17327), .ZN(n17328) );
  XNOR2_X1 U20541 ( .A(n17328), .B(n17331), .ZN(n17663) );
  NOR2_X1 U20542 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17345), .ZN(
        n17662) );
  AOI22_X1 U20543 ( .A1(n17484), .A2(n17663), .B1(n17342), .B2(n17662), .ZN(
        n17329) );
  OAI211_X1 U20544 ( .C1(n17346), .C2(n17331), .A(n17330), .B(n17329), .ZN(
        P3_U2810) );
  AOI21_X1 U20545 ( .B1(n17474), .B2(n17333), .A(n17559), .ZN(n17367) );
  OAI21_X1 U20546 ( .B1(n17332), .B2(n17574), .A(n17367), .ZN(n17349) );
  NOR2_X1 U20547 ( .A1(n17334), .A2(n17333), .ZN(n17351) );
  OAI211_X1 U20548 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17351), .B(n17335), .ZN(n17336) );
  NAND2_X1 U20549 ( .A1(n17896), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17675) );
  OAI211_X1 U20550 ( .C1(n9591), .C2(n17337), .A(n17336), .B(n17675), .ZN(
        n17338) );
  AOI21_X1 U20551 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17349), .A(
        n17338), .ZN(n17344) );
  OAI21_X1 U20552 ( .B1(n17340), .B2(n17352), .A(n17339), .ZN(n17341) );
  XNOR2_X1 U20553 ( .A(n17341), .B(n17345), .ZN(n17673) );
  AOI22_X1 U20554 ( .A1(n17484), .A2(n17673), .B1(n17342), .B2(n17345), .ZN(
        n17343) );
  OAI211_X1 U20555 ( .C1(n17346), .C2(n17345), .A(n17344), .B(n17343), .ZN(
        P3_U2811) );
  AOI21_X1 U20556 ( .B1(n17382), .B2(n17682), .A(n17381), .ZN(n17363) );
  INV_X1 U20557 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17350) );
  OAI22_X1 U20558 ( .A1(n17894), .A2(n18484), .B1(n9591), .B2(n17347), .ZN(
        n17348) );
  AOI221_X1 U20559 ( .B1(n17351), .B2(n17350), .C1(n17349), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17348), .ZN(n17356) );
  OAI21_X1 U20560 ( .B1(n17357), .B2(n17483), .A(n17352), .ZN(n17354) );
  XNOR2_X1 U20561 ( .A(n17354), .B(n17353), .ZN(n17691) );
  NOR2_X1 U20562 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17682), .ZN(
        n17690) );
  AOI22_X1 U20563 ( .A1(n17484), .A2(n17691), .B1(n17382), .B2(n17690), .ZN(
        n17355) );
  OAI211_X1 U20564 ( .C1(n17363), .C2(n17357), .A(n17356), .B(n17355), .ZN(
        P3_U2812) );
  AOI21_X1 U20565 ( .B1(n17358), .B2(n18299), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U20566 ( .A1(n17896), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17360), 
        .B2(n17567), .ZN(n17366) );
  NOR2_X1 U20567 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17704), .ZN(
        n17694) );
  AOI21_X1 U20568 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17362), .A(
        n17361), .ZN(n17698) );
  OAI22_X1 U20569 ( .A1(n17363), .A2(n17685), .B1(n17698), .B2(n17458), .ZN(
        n17364) );
  AOI21_X1 U20570 ( .B1(n17382), .B2(n17694), .A(n17364), .ZN(n17365) );
  OAI211_X1 U20571 ( .C1(n17368), .C2(n17367), .A(n17366), .B(n17365), .ZN(
        P3_U2813) );
  NOR2_X1 U20572 ( .A1(n17483), .A2(n17481), .ZN(n17459) );
  AOI22_X1 U20573 ( .A1(n17370), .A2(n17459), .B1(n17369), .B2(n17483), .ZN(
        n17371) );
  XNOR2_X1 U20574 ( .A(n17371), .B(n17704), .ZN(n17709) );
  AOI21_X1 U20575 ( .B1(n17474), .B2(n17372), .A(n17559), .ZN(n17399) );
  OAI21_X1 U20576 ( .B1(n17373), .B2(n17574), .A(n17399), .ZN(n17386) );
  AOI22_X1 U20577 ( .A1(n17896), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17386), .ZN(n17378) );
  NAND2_X1 U20578 ( .A1(n17413), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17375) );
  NAND2_X1 U20579 ( .A1(n17415), .A2(n17374), .ZN(n17429) );
  NOR2_X1 U20580 ( .A1(n17375), .A2(n17429), .ZN(n17388) );
  OAI211_X1 U20581 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17388), .B(n17376), .ZN(n17377) );
  OAI211_X1 U20582 ( .C1(n17379), .C2(n9591), .A(n17378), .B(n17377), .ZN(
        n17380) );
  AOI221_X1 U20583 ( .B1(n17382), .B2(n17704), .C1(n17381), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17380), .ZN(n17383) );
  OAI21_X1 U20584 ( .B1(n17709), .B2(n17458), .A(n17383), .ZN(P3_U2814) );
  INV_X1 U20585 ( .A(n17768), .ZN(n17440) );
  NOR3_X1 U20586 ( .A1(n17440), .A2(n20690), .A3(n17731), .ZN(n17402) );
  NOR2_X1 U20587 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17402), .ZN(
        n17716) );
  NAND2_X1 U20588 ( .A1(n17565), .A2(n17638), .ZN(n17394) );
  OAI22_X1 U20589 ( .A1(n17894), .A2(n18478), .B1(n9591), .B2(n17384), .ZN(
        n17385) );
  AOI221_X1 U20590 ( .B1(n17388), .B2(n17387), .C1(n17386), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17385), .ZN(n17393) );
  NAND2_X1 U20591 ( .A1(n17410), .A2(n17459), .ZN(n17406) );
  NOR2_X1 U20592 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17758), .ZN(
        n17422) );
  AOI221_X1 U20593 ( .B1(n20690), .B2(n17389), .C1(n17406), .C2(n17389), .A(
        n17422), .ZN(n17390) );
  XNOR2_X1 U20594 ( .A(n17390), .B(n17718), .ZN(n17721) );
  NOR2_X1 U20595 ( .A1(n17710), .A2(n17421), .ZN(n17391) );
  NAND2_X1 U20596 ( .A1(n17718), .A2(n17395), .ZN(n17714) );
  AOI22_X1 U20597 ( .A1(n17484), .A2(n17721), .B1(n17391), .B2(n17714), .ZN(
        n17392) );
  OAI211_X1 U20598 ( .C1(n17716), .C2(n17394), .A(n17393), .B(n17392), .ZN(
        P3_U2815) );
  OAI21_X1 U20599 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17396), .A(
        n17395), .ZN(n17739) );
  NOR3_X1 U20600 ( .A1(n17958), .A2(n17473), .A3(n17397), .ZN(n17438) );
  AOI21_X1 U20601 ( .B1(n17413), .B2(n17438), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17398) );
  OAI22_X1 U20602 ( .A1(n17399), .A2(n17398), .B1(n17894), .B2(n18477), .ZN(
        n17400) );
  AOI21_X1 U20603 ( .B1(n17401), .B2(n17567), .A(n17400), .ZN(n17409) );
  NAND2_X1 U20604 ( .A1(n17725), .A2(n17768), .ZN(n17403) );
  AOI21_X1 U20605 ( .B1(n20690), .B2(n17403), .A(n17402), .ZN(n17736) );
  INV_X1 U20606 ( .A(n17404), .ZN(n17405) );
  AOI21_X1 U20607 ( .B1(n17406), .B2(n17405), .A(n17422), .ZN(n17407) );
  XNOR2_X1 U20608 ( .A(n17407), .B(n20690), .ZN(n17735) );
  AOI22_X1 U20609 ( .A1(n17565), .A2(n17736), .B1(n17484), .B2(n17735), .ZN(
        n17408) );
  OAI211_X1 U20610 ( .C1(n17421), .C2(n17739), .A(n17409), .B(n17408), .ZN(
        P3_U2816) );
  INV_X1 U20611 ( .A(n17410), .ZN(n17741) );
  NOR2_X1 U20612 ( .A1(n17741), .A2(n17481), .ZN(n17743) );
  AOI21_X1 U20613 ( .B1(n17758), .B2(n17483), .A(n17743), .ZN(n17411) );
  AOI21_X1 U20614 ( .B1(n17483), .B2(n17425), .A(n17411), .ZN(n17412) );
  XNOR2_X1 U20615 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17412), .ZN(
        n17752) );
  AOI211_X1 U20616 ( .C1(n17428), .C2(n17418), .A(n17413), .B(n17429), .ZN(
        n17420) );
  OAI22_X1 U20617 ( .A1(n17415), .A2(n17534), .B1(n17414), .B2(n17574), .ZN(
        n17416) );
  NOR2_X1 U20618 ( .A1(n17559), .A2(n17416), .ZN(n17427) );
  OAI22_X1 U20619 ( .A1(n17427), .A2(n17418), .B1(n9591), .B2(n17417), .ZN(
        n17419) );
  AOI211_X1 U20620 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17896), .A(n17420), 
        .B(n17419), .ZN(n17424) );
  NOR2_X1 U20621 ( .A1(n17741), .A2(n17440), .ZN(n17744) );
  OAI22_X1 U20622 ( .A1(n17743), .A2(n17421), .B1(n17744), .B2(n17578), .ZN(
        n17433) );
  NOR2_X1 U20623 ( .A1(n17469), .A2(n17753), .ZN(n17432) );
  AOI22_X1 U20624 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17433), .B1(
        n17422), .B2(n17432), .ZN(n17423) );
  OAI211_X1 U20625 ( .C1(n17458), .C2(n17752), .A(n17424), .B(n17423), .ZN(
        P3_U2817) );
  NAND2_X1 U20626 ( .A1(n17767), .A2(n17459), .ZN(n17441) );
  OAI21_X1 U20627 ( .B1(n17442), .B2(n17441), .A(n17425), .ZN(n17426) );
  XOR2_X1 U20628 ( .A(n17426), .B(n17758), .Z(n17757) );
  NAND2_X1 U20629 ( .A1(n17896), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17761) );
  OAI221_X1 U20630 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17429), .C1(
        n17428), .C2(n17427), .A(n17761), .ZN(n17430) );
  AOI21_X1 U20631 ( .B1(n9610), .B2(n17431), .A(n17430), .ZN(n17435) );
  AOI22_X1 U20632 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17433), .B1(
        n17432), .B2(n17758), .ZN(n17434) );
  OAI211_X1 U20633 ( .C1(n17757), .C2(n17458), .A(n17435), .B(n17434), .ZN(
        P3_U2818) );
  NAND2_X1 U20634 ( .A1(n17767), .A2(n17442), .ZN(n17777) );
  NOR2_X1 U20635 ( .A1(n17958), .A2(n17473), .ZN(n17493) );
  NAND3_X1 U20636 ( .A1(n17477), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17493), .ZN(n17461) );
  NOR2_X1 U20637 ( .A1(n17450), .A2(n17461), .ZN(n17449) );
  AOI21_X1 U20638 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17568), .A(
        n17449), .ZN(n17437) );
  OAI22_X1 U20639 ( .A1(n17438), .A2(n17437), .B1(n17557), .B2(n17436), .ZN(
        n17439) );
  AOI21_X1 U20640 ( .B1(n17896), .B2(P3_REIP_REG_11__SCAN_IN), .A(n17439), 
        .ZN(n17445) );
  AOI22_X1 U20641 ( .A1(n17565), .A2(n17440), .B1(n17485), .B2(n17481), .ZN(
        n17468) );
  OAI21_X1 U20642 ( .B1(n17767), .B2(n17469), .A(n17468), .ZN(n17454) );
  OAI21_X1 U20643 ( .B1(n17446), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17441), .ZN(n17443) );
  XNOR2_X1 U20644 ( .A(n17443), .B(n17442), .ZN(n17763) );
  AOI22_X1 U20645 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17454), .B1(
        n17484), .B2(n17763), .ZN(n17444) );
  OAI211_X1 U20646 ( .C1(n17469), .C2(n17777), .A(n17445), .B(n17444), .ZN(
        P3_U2819) );
  INV_X1 U20647 ( .A(n17459), .ZN(n17447) );
  OAI21_X1 U20648 ( .B1(n17800), .B2(n17447), .A(n17446), .ZN(n17448) );
  XNOR2_X1 U20649 ( .A(n17448), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17789) );
  INV_X1 U20650 ( .A(n17568), .ZN(n17508) );
  AOI211_X1 U20651 ( .C1(n17461), .C2(n17450), .A(n17508), .B(n17449), .ZN(
        n17452) );
  NOR2_X1 U20652 ( .A1(n17894), .A2(n18469), .ZN(n17451) );
  AOI211_X1 U20653 ( .C1(n17453), .C2(n17567), .A(n17452), .B(n17451), .ZN(
        n17457) );
  INV_X1 U20654 ( .A(n17469), .ZN(n17455) );
  OAI221_X1 U20655 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17455), .A(n17454), .ZN(
        n17456) );
  OAI211_X1 U20656 ( .C1(n17789), .C2(n17458), .A(n17457), .B(n17456), .ZN(
        P3_U2820) );
  NOR2_X1 U20657 ( .A1(n17459), .A2(n9682), .ZN(n17460) );
  XNOR2_X1 U20658 ( .A(n17460), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17797) );
  NOR2_X1 U20659 ( .A1(n17894), .A2(n18467), .ZN(n17466) );
  INV_X1 U20660 ( .A(n17461), .ZN(n17464) );
  AOI22_X1 U20661 ( .A1(n17477), .A2(n17493), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17568), .ZN(n17463) );
  OAI22_X1 U20662 ( .A1(n17464), .A2(n17463), .B1(n17557), .B2(n17462), .ZN(
        n17465) );
  AOI211_X1 U20663 ( .C1(n17484), .C2(n17797), .A(n17466), .B(n17465), .ZN(
        n17467) );
  OAI221_X1 U20664 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17469), .C1(
        n17800), .C2(n17468), .A(n17467), .ZN(P3_U2821) );
  OAI21_X1 U20665 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17471), .A(
        n17470), .ZN(n17819) );
  NOR2_X1 U20666 ( .A1(n17894), .A2(n18465), .ZN(n17809) );
  OAI21_X1 U20667 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17472), .A(
        n18299), .ZN(n17476) );
  AOI21_X1 U20668 ( .B1(n17474), .B2(n17473), .A(n17559), .ZN(n17490) );
  OAI22_X1 U20669 ( .A1(n17477), .A2(n17476), .B1(n17490), .B2(n17475), .ZN(
        n17478) );
  AOI211_X1 U20670 ( .C1(n17479), .C2(n17567), .A(n17809), .B(n17478), .ZN(
        n17487) );
  NAND2_X1 U20671 ( .A1(n17481), .A2(n17480), .ZN(n17482) );
  INV_X1 U20672 ( .A(n17482), .ZN(n17815) );
  XNOR2_X1 U20673 ( .A(n17483), .B(n17482), .ZN(n17813) );
  AOI22_X1 U20674 ( .A1(n17485), .A2(n17815), .B1(n17484), .B2(n17813), .ZN(
        n17486) );
  OAI211_X1 U20675 ( .C1(n17578), .C2(n17819), .A(n17487), .B(n17486), .ZN(
        P3_U2822) );
  OAI21_X1 U20676 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17489), .A(
        n17488), .ZN(n17828) );
  INV_X1 U20677 ( .A(n17490), .ZN(n17491) );
  NOR2_X1 U20678 ( .A1(n17894), .A2(n18463), .ZN(n17820) );
  AOI221_X1 U20679 ( .B1(n17493), .B2(n17492), .C1(n17491), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17820), .ZN(n17500) );
  AOI21_X1 U20680 ( .B1(n17496), .B2(n17495), .A(n17494), .ZN(n17497) );
  XNOR2_X1 U20681 ( .A(n17497), .B(n17807), .ZN(n17824) );
  AOI22_X1 U20682 ( .A1(n17565), .A2(n17824), .B1(n17498), .B2(n17567), .ZN(
        n17499) );
  OAI211_X1 U20683 ( .C1(n17577), .C2(n17828), .A(n17500), .B(n17499), .ZN(
        P3_U2823) );
  OAI21_X1 U20684 ( .B1(n17502), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17501), .ZN(n17831) );
  NAND2_X1 U20685 ( .A1(n18299), .A2(n17509), .ZN(n17506) );
  OAI21_X1 U20686 ( .B1(n17505), .B2(n17504), .A(n17503), .ZN(n17830) );
  OAI22_X1 U20687 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17506), .B1(
        n17577), .B2(n17830), .ZN(n17507) );
  AOI21_X1 U20688 ( .B1(n17896), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17507), .ZN(
        n17512) );
  AOI21_X1 U20689 ( .B1(n17509), .B2(n18299), .A(n17508), .ZN(n17523) );
  AOI22_X1 U20690 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17523), .B1(
        n17510), .B2(n17567), .ZN(n17511) );
  OAI211_X1 U20691 ( .C1(n17578), .C2(n17831), .A(n17512), .B(n17511), .ZN(
        P3_U2824) );
  OAI21_X1 U20692 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17514), .A(
        n17513), .ZN(n17838) );
  OAI21_X1 U20693 ( .B1(n17559), .B2(n17516), .A(n17515), .ZN(n17522) );
  OAI21_X1 U20694 ( .B1(n17519), .B2(n17518), .A(n17517), .ZN(n17845) );
  OAI22_X1 U20695 ( .A1(n17557), .A2(n17520), .B1(n17578), .B2(n17845), .ZN(
        n17521) );
  AOI21_X1 U20696 ( .B1(n17523), .B2(n17522), .A(n17521), .ZN(n17524) );
  NAND2_X1 U20697 ( .A1(n17896), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n17843) );
  OAI211_X1 U20698 ( .C1(n17577), .C2(n17838), .A(n17524), .B(n17843), .ZN(
        P3_U2825) );
  OAI21_X1 U20699 ( .B1(n17527), .B2(n17526), .A(n17525), .ZN(n17855) );
  OAI21_X1 U20700 ( .B1(n17530), .B2(n17529), .A(n17528), .ZN(n17531) );
  XNOR2_X1 U20701 ( .A(n17531), .B(n20762), .ZN(n17850) );
  OAI22_X1 U20702 ( .A1(n17578), .A2(n17850), .B1(n17958), .B2(n17532), .ZN(
        n17533) );
  AOI21_X1 U20703 ( .B1(n17896), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17533), .ZN(
        n17538) );
  OAI21_X1 U20704 ( .B1(n17535), .B2(n17534), .A(n17573), .ZN(n17548) );
  AOI22_X1 U20705 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17548), .B1(
        n17536), .B2(n17567), .ZN(n17537) );
  OAI211_X1 U20706 ( .C1(n17577), .C2(n17855), .A(n17538), .B(n17537), .ZN(
        P3_U2826) );
  OAI21_X1 U20707 ( .B1(n17541), .B2(n17540), .A(n17539), .ZN(n17858) );
  NOR2_X1 U20708 ( .A1(n17559), .A2(n17560), .ZN(n17547) );
  OAI21_X1 U20709 ( .B1(n17544), .B2(n17543), .A(n17542), .ZN(n17859) );
  OAI22_X1 U20710 ( .A1(n17557), .A2(n17545), .B1(n17577), .B2(n17859), .ZN(
        n17546) );
  AOI221_X1 U20711 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17548), .C1(
        n17547), .C2(n17548), .A(n17546), .ZN(n17549) );
  NAND2_X1 U20712 ( .A1(n17896), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n17862) );
  OAI211_X1 U20713 ( .C1(n17578), .C2(n17858), .A(n17549), .B(n17862), .ZN(
        P3_U2827) );
  OAI21_X1 U20714 ( .B1(n17552), .B2(n17551), .A(n17550), .ZN(n17873) );
  OAI21_X1 U20715 ( .B1(n17555), .B2(n17554), .A(n17553), .ZN(n17874) );
  OAI22_X1 U20716 ( .A1(n17557), .A2(n17556), .B1(n17577), .B2(n17874), .ZN(
        n17558) );
  AOI221_X1 U20717 ( .B1(n18299), .B2(n17560), .C1(n17559), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17558), .ZN(n17561) );
  NAND2_X1 U20718 ( .A1(n17896), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n17877) );
  OAI211_X1 U20719 ( .C1(n17578), .C2(n17873), .A(n17561), .B(n17877), .ZN(
        P3_U2828) );
  OAI21_X1 U20720 ( .B1(n17563), .B2(n17571), .A(n17562), .ZN(n17891) );
  NAND2_X1 U20721 ( .A1(n18546), .A2(n17572), .ZN(n17564) );
  XNOR2_X1 U20722 ( .A(n17564), .B(n17563), .ZN(n17884) );
  AOI22_X1 U20723 ( .A1(n17565), .A2(n17884), .B1(n17896), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17570) );
  AOI22_X1 U20724 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17568), .B1(
        n17567), .B2(n17566), .ZN(n17569) );
  OAI211_X1 U20725 ( .C1(n17577), .C2(n17891), .A(n17570), .B(n17569), .ZN(
        P3_U2829) );
  AOI21_X1 U20726 ( .B1(n17572), .B2(n18546), .A(n17571), .ZN(n17901) );
  INV_X1 U20727 ( .A(n17901), .ZN(n17899) );
  NAND3_X1 U20728 ( .A1(n18426), .A2(n17574), .A3(n17573), .ZN(n17575) );
  AOI22_X1 U20729 ( .A1(n17896), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17575), .ZN(n17576) );
  OAI221_X1 U20730 ( .B1(n17901), .B2(n17578), .C1(n17899), .C2(n17577), .A(
        n17576), .ZN(P3_U2830) );
  AOI22_X1 U20731 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17888), .B1(
        n17896), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n17590) );
  INV_X1 U20732 ( .A(n18380), .ZN(n18354) );
  NOR2_X1 U20733 ( .A1(n18354), .A2(n18378), .ZN(n17865) );
  NOR2_X1 U20734 ( .A1(n17579), .A2(n17865), .ZN(n17580) );
  AOI211_X1 U20735 ( .C1(n18563), .C2(n17582), .A(n17581), .B(n17580), .ZN(
        n17583) );
  NAND2_X1 U20736 ( .A1(n18378), .A2(n18546), .ZN(n17866) );
  OR4_X1 U20737 ( .A1(n17678), .A2(n17643), .A3(n17641), .A4(n17849), .ZN(
        n17645) );
  NAND2_X1 U20738 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17598) );
  INV_X1 U20739 ( .A(n17865), .ZN(n17803) );
  OAI21_X1 U20740 ( .B1(n17645), .B2(n17598), .A(n17803), .ZN(n17604) );
  OAI211_X1 U20741 ( .C1(n17584), .C2(n17770), .A(n17583), .B(n17604), .ZN(
        n17594) );
  OAI22_X1 U20742 ( .A1(n17586), .A2(n17585), .B1(n17588), .B2(n17886), .ZN(
        n17587) );
  OAI21_X1 U20743 ( .B1(n17588), .B2(n17594), .A(n17587), .ZN(n17589) );
  OAI211_X1 U20744 ( .C1(n17591), .C2(n17788), .A(n17590), .B(n17589), .ZN(
        P3_U2835) );
  AOI22_X1 U20745 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17888), .B1(
        n17896), .B2(P3_REIP_REG_26__SCAN_IN), .ZN(n17597) );
  AOI22_X1 U20746 ( .A1(n17814), .A2(n17593), .B1(n17613), .B2(n17592), .ZN(
        n17596) );
  NAND3_X1 U20747 ( .A1(n17892), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n17594), .ZN(n17595) );
  NAND3_X1 U20748 ( .A1(n17597), .A2(n17596), .A3(n17595), .ZN(P3_U2836) );
  NAND2_X1 U20749 ( .A1(n17627), .A2(n17679), .ZN(n17618) );
  AOI221_X1 U20750 ( .B1(n17598), .B2(n18404), .C1(n17618), .C2(n18404), .A(
        n17599), .ZN(n17605) );
  OAI21_X1 U20751 ( .B1(n17601), .B2(n17600), .A(n17599), .ZN(n17602) );
  INV_X1 U20752 ( .A(n17602), .ZN(n17603) );
  AOI211_X1 U20753 ( .C1(n17605), .C2(n17604), .A(n17603), .B(n17886), .ZN(
        n17606) );
  AOI211_X1 U20754 ( .C1(n17888), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17607), .B(n17606), .ZN(n17611) );
  AOI22_X1 U20755 ( .A1(n17816), .A2(n17609), .B1(n17814), .B2(n17608), .ZN(
        n17610) );
  OAI211_X1 U20756 ( .C1(n17900), .C2(n17612), .A(n17611), .B(n17610), .ZN(
        P3_U2837) );
  INV_X1 U20757 ( .A(n17613), .ZN(n17634) );
  NOR2_X1 U20758 ( .A1(n17614), .A2(n17636), .ZN(n17616) );
  NOR2_X1 U20759 ( .A1(n17638), .A2(n17614), .ZN(n17615) );
  OAI22_X1 U20760 ( .A1(n17616), .A2(n17770), .B1(n17615), .B2(n17769), .ZN(
        n17617) );
  AOI211_X1 U20761 ( .C1(n17803), .C2(n17645), .A(n17888), .B(n17617), .ZN(
        n17621) );
  AOI21_X1 U20762 ( .B1(n18404), .B2(n17618), .A(n20685), .ZN(n17619) );
  AOI21_X1 U20763 ( .B1(n17621), .B2(n17619), .A(n17896), .ZN(n17629) );
  AOI21_X1 U20764 ( .B1(n17703), .B2(n17621), .A(n17620), .ZN(n17622) );
  AOI22_X1 U20765 ( .A1(n17814), .A2(n17623), .B1(n17629), .B2(n17622), .ZN(
        n17625) );
  NAND2_X1 U20766 ( .A1(n17896), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17624) );
  OAI211_X1 U20767 ( .C1(n17626), .C2(n17634), .A(n17625), .B(n17624), .ZN(
        P3_U2838) );
  NAND2_X1 U20768 ( .A1(n17896), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17632) );
  AND3_X1 U20769 ( .A1(n17880), .A2(n17628), .A3(n17627), .ZN(n17630) );
  OAI21_X1 U20770 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17630), .A(
        n17629), .ZN(n17631) );
  OAI211_X1 U20771 ( .C1(n17633), .C2(n17788), .A(n17632), .B(n17631), .ZN(
        P3_U2839) );
  AOI22_X1 U20772 ( .A1(n17642), .A2(n17672), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17892), .ZN(n17650) );
  INV_X1 U20773 ( .A(n17780), .ZN(n17748) );
  AOI22_X1 U20774 ( .A1(n18563), .A2(n17638), .B1(n17637), .B2(n17636), .ZN(
        n17653) );
  NAND2_X1 U20775 ( .A1(n17769), .A2(n17770), .ZN(n17764) );
  AOI21_X1 U20776 ( .B1(n17652), .B2(n17679), .A(n18374), .ZN(n17639) );
  AOI221_X1 U20777 ( .B1(n17678), .B2(n18354), .C1(n17666), .C2(n18354), .A(
        n17639), .ZN(n17668) );
  OAI21_X1 U20778 ( .B1(n18380), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17668), .ZN(n17640) );
  AOI21_X1 U20779 ( .B1(n17641), .B2(n17764), .A(n17640), .ZN(n17655) );
  OAI211_X1 U20780 ( .C1(n17748), .C2(n17642), .A(n17653), .B(n17655), .ZN(
        n17644) );
  AOI211_X1 U20781 ( .C1(n17645), .C2(n18378), .A(n17644), .B(n17643), .ZN(
        n17649) );
  AOI22_X1 U20782 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17888), .B1(
        n17814), .B2(n17646), .ZN(n17648) );
  OAI211_X1 U20783 ( .C1(n17650), .C2(n17649), .A(n17648), .B(n17647), .ZN(
        P3_U2840) );
  INV_X1 U20784 ( .A(n17651), .ZN(n17656) );
  NOR2_X1 U20785 ( .A1(n18404), .A2(n18378), .ZN(n17887) );
  AOI21_X1 U20786 ( .B1(n17652), .B2(n17700), .A(n17773), .ZN(n17654) );
  NAND2_X1 U20787 ( .A1(n17892), .A2(n17653), .ZN(n17699) );
  NOR2_X1 U20788 ( .A1(n17654), .A2(n17699), .ZN(n17664) );
  OAI211_X1 U20789 ( .C1(n17656), .C2(n17887), .A(n17655), .B(n17664), .ZN(
        n17657) );
  NAND2_X1 U20790 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17657), .ZN(
        n17661) );
  AOI22_X1 U20791 ( .A1(n17814), .A2(n17659), .B1(n17658), .B2(n17672), .ZN(
        n17660) );
  OAI221_X1 U20792 ( .B1(n17896), .B2(n17661), .C1(n17894), .C2(n18491), .A(
        n17660), .ZN(P3_U2841) );
  AOI22_X1 U20793 ( .A1(n17814), .A2(n17663), .B1(n17662), .B2(n17672), .ZN(
        n17671) );
  INV_X1 U20794 ( .A(n17664), .ZN(n17665) );
  AOI21_X1 U20795 ( .B1(n17666), .B2(n17764), .A(n17665), .ZN(n17667) );
  AOI21_X1 U20796 ( .B1(n17668), .B2(n17667), .A(n17896), .ZN(n17674) );
  NOR3_X1 U20797 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17887), .A3(
        n18415), .ZN(n17669) );
  OAI21_X1 U20798 ( .B1(n17674), .B2(n17669), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17670) );
  OAI211_X1 U20799 ( .C1(n18488), .C2(n17894), .A(n17671), .B(n17670), .ZN(
        P3_U2842) );
  INV_X1 U20800 ( .A(n17672), .ZN(n17677) );
  AOI22_X1 U20801 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17674), .B1(
        n17814), .B2(n17673), .ZN(n17676) );
  OAI211_X1 U20802 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17677), .A(
        n17676), .B(n17675), .ZN(P3_U2843) );
  NOR2_X1 U20803 ( .A1(n17849), .A2(n17678), .ZN(n17684) );
  AOI21_X1 U20804 ( .B1(n17680), .B2(n17679), .A(n18374), .ZN(n17681) );
  AOI211_X1 U20805 ( .C1(n17682), .C2(n17764), .A(n17681), .B(n17699), .ZN(
        n17683) );
  OAI221_X1 U20806 ( .B1(n17865), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), 
        .C1(n17865), .C2(n17684), .A(n17683), .ZN(n17695) );
  OAI221_X1 U20807 ( .B1(n17695), .B2(n17685), .C1(n17695), .C2(n17803), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17693) );
  INV_X1 U20808 ( .A(n17869), .ZN(n17846) );
  AOI22_X1 U20809 ( .A1(n18404), .A2(n17846), .B1(n17847), .B2(n17864), .ZN(
        n17857) );
  NOR2_X1 U20810 ( .A1(n17857), .A2(n17686), .ZN(n17821) );
  NAND2_X1 U20811 ( .A1(n17687), .A2(n17821), .ZN(n17730) );
  NAND2_X1 U20812 ( .A1(n17688), .A2(n17730), .ZN(n17755) );
  NAND2_X1 U20813 ( .A1(n17892), .A2(n17755), .ZN(n17801) );
  NOR2_X1 U20814 ( .A1(n17689), .A2(n17801), .ZN(n17705) );
  AOI22_X1 U20815 ( .A1(n17814), .A2(n17691), .B1(n17690), .B2(n17705), .ZN(
        n17692) );
  OAI221_X1 U20816 ( .B1(n17896), .B2(n17693), .C1(n17894), .C2(n18484), .A(
        n17692), .ZN(P3_U2844) );
  AOI22_X1 U20817 ( .A1(n17896), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17705), 
        .B2(n17694), .ZN(n17697) );
  NAND3_X1 U20818 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17894), .A3(
        n17695), .ZN(n17696) );
  OAI211_X1 U20819 ( .C1(n17698), .C2(n17788), .A(n17697), .B(n17696), .ZN(
        P3_U2845) );
  INV_X1 U20820 ( .A(n17699), .ZN(n17702) );
  OAI21_X1 U20821 ( .B1(n17802), .B2(n17804), .A(n18354), .ZN(n17793) );
  OAI21_X1 U20822 ( .B1(n18380), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n17793), .ZN(n17781) );
  NAND2_X1 U20823 ( .A1(n18404), .A2(n17726), .ZN(n17794) );
  OAI211_X1 U20824 ( .C1(n17700), .C2(n17773), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17794), .ZN(n17701) );
  AOI211_X1 U20825 ( .C1(n17780), .C2(n17712), .A(n17781), .B(n17701), .ZN(
        n17711) );
  AOI221_X1 U20826 ( .B1(n17703), .B2(n17702), .C1(n17711), .C2(n17702), .A(
        n17896), .ZN(n17706) );
  AOI22_X1 U20827 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17706), .B1(
        n17705), .B2(n17704), .ZN(n17708) );
  NAND2_X1 U20828 ( .A1(n17896), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17707) );
  OAI211_X1 U20829 ( .C1(n17709), .C2(n17788), .A(n17708), .B(n17707), .ZN(
        P3_U2846) );
  NOR2_X1 U20830 ( .A1(n17710), .A2(n17770), .ZN(n17715) );
  AOI221_X1 U20831 ( .B1(n17712), .B2(n17718), .C1(n17730), .C2(n17718), .A(
        n17711), .ZN(n17713) );
  AOI21_X1 U20832 ( .B1(n17715), .B2(n17714), .A(n17713), .ZN(n17723) );
  NOR3_X1 U20833 ( .A1(n17717), .A2(n17716), .A3(n17900), .ZN(n17720) );
  OAI22_X1 U20834 ( .A1(n17718), .A2(n17880), .B1(n17894), .B2(n18478), .ZN(
        n17719) );
  AOI211_X1 U20835 ( .C1(n17721), .C2(n17814), .A(n17720), .B(n17719), .ZN(
        n17722) );
  OAI21_X1 U20836 ( .B1(n17723), .B2(n17886), .A(n17722), .ZN(P3_U2847) );
  AOI21_X1 U20837 ( .B1(n17725), .B2(n17724), .A(n18380), .ZN(n17729) );
  AOI221_X1 U20838 ( .B1(n17741), .B2(n18404), .C1(n17726), .C2(n18404), .A(
        n20690), .ZN(n17727) );
  OAI21_X1 U20839 ( .B1(n17741), .B2(n17790), .A(n18378), .ZN(n17746) );
  OAI211_X1 U20840 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n17887), .A(
        n17727), .B(n17746), .ZN(n17728) );
  OAI21_X1 U20841 ( .B1(n17729), .B2(n17728), .A(n17892), .ZN(n17733) );
  OR2_X1 U20842 ( .A1(n17731), .A2(n17730), .ZN(n17732) );
  AOI222_X1 U20843 ( .A1(n20690), .A2(n17733), .B1(n20690), .B2(n17732), .C1(
        n17733), .C2(n17880), .ZN(n17734) );
  AOI21_X1 U20844 ( .B1(n17896), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17734), 
        .ZN(n17738) );
  AOI22_X1 U20845 ( .A1(n17885), .A2(n17736), .B1(n17814), .B2(n17735), .ZN(
        n17737) );
  OAI211_X1 U20846 ( .C1(n17740), .C2(n17739), .A(n17738), .B(n17737), .ZN(
        P3_U2848) );
  NOR3_X1 U20847 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17741), .A3(
        n17801), .ZN(n17742) );
  AOI21_X1 U20848 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n17896), .A(n17742), 
        .ZN(n17751) );
  OAI22_X1 U20849 ( .A1(n17769), .A2(n17744), .B1(n17770), .B2(n17743), .ZN(
        n17745) );
  INV_X1 U20850 ( .A(n17745), .ZN(n17747) );
  OAI21_X1 U20851 ( .B1(n17753), .B2(n17781), .A(n17780), .ZN(n17772) );
  NAND4_X1 U20852 ( .A1(n17747), .A2(n17794), .A3(n17746), .A4(n17772), .ZN(
        n17754) );
  OAI21_X1 U20853 ( .B1(n17748), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17892), .ZN(n17749) );
  OAI211_X1 U20854 ( .C1(n17754), .C2(n17749), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17894), .ZN(n17750) );
  OAI211_X1 U20855 ( .C1(n17752), .C2(n17788), .A(n17751), .B(n17750), .ZN(
        P3_U2849) );
  INV_X1 U20856 ( .A(n17753), .ZN(n17756) );
  OAI222_X1 U20857 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17756), 
        .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17755), .C1(n17754), 
        .C2(n17758), .ZN(n17762) );
  OAI22_X1 U20858 ( .A1(n17758), .A2(n17880), .B1(n17788), .B2(n17757), .ZN(
        n17759) );
  INV_X1 U20859 ( .A(n17759), .ZN(n17760) );
  OAI211_X1 U20860 ( .C1(n17886), .C2(n17762), .A(n17761), .B(n17760), .ZN(
        P3_U2850) );
  AOI22_X1 U20861 ( .A1(n17896), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17814), 
        .B2(n17763), .ZN(n17776) );
  INV_X1 U20862 ( .A(n17764), .ZN(n17766) );
  OAI21_X1 U20863 ( .B1(n17800), .B2(n17790), .A(n18378), .ZN(n17765) );
  OAI211_X1 U20864 ( .C1(n17767), .C2(n17766), .A(n17765), .B(n17794), .ZN(
        n17778) );
  OAI22_X1 U20865 ( .A1(n17771), .A2(n17770), .B1(n17769), .B2(n17768), .ZN(
        n17779) );
  NOR2_X1 U20866 ( .A1(n17886), .A2(n17779), .ZN(n17795) );
  OAI211_X1 U20867 ( .C1(n17773), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17795), .B(n17772), .ZN(n17774) );
  OAI211_X1 U20868 ( .C1(n17778), .C2(n17774), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17894), .ZN(n17775) );
  OAI211_X1 U20869 ( .C1(n17777), .C2(n17801), .A(n17776), .B(n17775), .ZN(
        P3_U2851) );
  NOR3_X1 U20870 ( .A1(n17888), .A2(n17779), .A3(n17778), .ZN(n17784) );
  OAI21_X1 U20871 ( .B1(n17800), .B2(n17781), .A(n17780), .ZN(n17783) );
  AOI21_X1 U20872 ( .B1(n17784), .B2(n17783), .A(n17782), .ZN(n17786) );
  NOR3_X1 U20873 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17800), .A3(
        n17801), .ZN(n17785) );
  AOI221_X1 U20874 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17896), .C1(n17786), 
        .C2(n17894), .A(n17785), .ZN(n17787) );
  OAI21_X1 U20875 ( .B1(n17789), .B2(n17788), .A(n17787), .ZN(P3_U2852) );
  NOR2_X1 U20876 ( .A1(n18380), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17791) );
  OAI21_X1 U20877 ( .B1(n17791), .B2(n18378), .A(n17790), .ZN(n17792) );
  NAND4_X1 U20878 ( .A1(n17795), .A2(n17794), .A3(n17793), .A4(n17792), .ZN(
        n17796) );
  NAND2_X1 U20879 ( .A1(n17894), .A2(n17796), .ZN(n17799) );
  AOI22_X1 U20880 ( .A1(n17896), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17814), 
        .B2(n17797), .ZN(n17798) );
  OAI221_X1 U20881 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17801), .C1(
        n17800), .C2(n17799), .A(n17798), .ZN(P3_U2853) );
  NOR3_X1 U20882 ( .A1(n17857), .A2(n17886), .A3(n15483), .ZN(n17853) );
  NAND3_X1 U20883 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n17853), .ZN(n17837) );
  NOR2_X1 U20884 ( .A1(n17802), .A2(n17837), .ZN(n17812) );
  AOI21_X1 U20885 ( .B1(n17804), .B2(n17803), .A(n17849), .ZN(n17805) );
  OAI21_X1 U20886 ( .B1(n17806), .B2(n18374), .A(n17805), .ZN(n17829) );
  AOI211_X1 U20887 ( .C1(n17808), .C2(n17836), .A(n17807), .B(n17829), .ZN(
        n17823) );
  OAI21_X1 U20888 ( .B1(n17823), .B2(n17881), .A(n17880), .ZN(n17810) );
  AOI221_X1 U20889 ( .B1(n17812), .B2(n17811), .C1(n17810), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n17809), .ZN(n17818) );
  AOI22_X1 U20890 ( .A1(n17816), .A2(n17815), .B1(n17814), .B2(n17813), .ZN(
        n17817) );
  OAI211_X1 U20891 ( .C1(n17900), .C2(n17819), .A(n17818), .B(n17817), .ZN(
        P3_U2854) );
  AOI21_X1 U20892 ( .B1(n17888), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17820), .ZN(n17827) );
  AOI21_X1 U20893 ( .B1(n17821), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17822) );
  NOR2_X1 U20894 ( .A1(n17823), .A2(n17822), .ZN(n17825) );
  AOI22_X1 U20895 ( .A1(n17892), .A2(n17825), .B1(n17885), .B2(n17824), .ZN(
        n17826) );
  OAI211_X1 U20896 ( .C1(n17898), .C2(n17828), .A(n17827), .B(n17826), .ZN(
        P3_U2855) );
  OAI21_X1 U20897 ( .B1(n17886), .B2(n17829), .A(n17894), .ZN(n17839) );
  INV_X1 U20898 ( .A(n17830), .ZN(n17833) );
  OAI22_X1 U20899 ( .A1(n17894), .A2(n20750), .B1(n17900), .B2(n17831), .ZN(
        n17832) );
  AOI21_X1 U20900 ( .B1(n17834), .B2(n17833), .A(n17832), .ZN(n17835) );
  OAI221_X1 U20901 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17837), .C1(
        n17836), .C2(n17839), .A(n17835), .ZN(P3_U2856) );
  NOR2_X1 U20902 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20762), .ZN(
        n17842) );
  OAI22_X1 U20903 ( .A1(n17840), .A2(n17839), .B1(n17898), .B2(n17838), .ZN(
        n17841) );
  AOI21_X1 U20904 ( .B1(n17842), .B2(n17853), .A(n17841), .ZN(n17844) );
  OAI211_X1 U20905 ( .C1(n17845), .C2(n17900), .A(n17844), .B(n17843), .ZN(
        P3_U2857) );
  OAI22_X1 U20906 ( .A1(n17847), .A2(n17865), .B1(n18374), .B2(n17846), .ZN(
        n17848) );
  NOR3_X1 U20907 ( .A1(n17849), .A2(n15483), .A3(n17848), .ZN(n17856) );
  OAI21_X1 U20908 ( .B1(n17856), .B2(n17881), .A(n17880), .ZN(n17852) );
  OAI22_X1 U20909 ( .A1(n17894), .A2(n18458), .B1(n17900), .B2(n17850), .ZN(
        n17851) );
  AOI221_X1 U20910 ( .B1(n17853), .B2(n20762), .C1(n17852), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n17851), .ZN(n17854) );
  OAI21_X1 U20911 ( .B1(n17898), .B2(n17855), .A(n17854), .ZN(P3_U2858) );
  AOI211_X1 U20912 ( .C1(n17857), .C2(n15483), .A(n17856), .B(n17886), .ZN(
        n17861) );
  OAI22_X1 U20913 ( .A1(n17898), .A2(n17859), .B1(n17900), .B2(n17858), .ZN(
        n17860) );
  NOR2_X1 U20914 ( .A1(n17861), .A2(n17860), .ZN(n17863) );
  OAI211_X1 U20915 ( .C1(n17880), .C2(n15483), .A(n17863), .B(n17862), .ZN(
        P3_U2859) );
  NAND2_X1 U20916 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17864), .ZN(
        n17872) );
  NOR2_X1 U20917 ( .A1(n18546), .A2(n15467), .ZN(n17868) );
  AOI21_X1 U20918 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17866), .A(
        n17865), .ZN(n17867) );
  AOI21_X1 U20919 ( .B1(n17868), .B2(n18404), .A(n17867), .ZN(n17871) );
  NAND2_X1 U20920 ( .A1(n18404), .A2(n17869), .ZN(n17870) );
  OAI221_X1 U20921 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n17872), .C1(
        n17879), .C2(n17871), .A(n17870), .ZN(n17876) );
  OAI22_X1 U20922 ( .A1(n17898), .A2(n17874), .B1(n17900), .B2(n17873), .ZN(
        n17875) );
  AOI21_X1 U20923 ( .B1(n17892), .B2(n17876), .A(n17875), .ZN(n17878) );
  OAI211_X1 U20924 ( .C1(n17880), .C2(n17879), .A(n17878), .B(n17877), .ZN(
        P3_U2860) );
  NOR2_X1 U20925 ( .A1(n17894), .A2(n18551), .ZN(n17883) );
  AOI211_X1 U20926 ( .C1(n18380), .C2(n18546), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n17881), .ZN(n17882) );
  AOI211_X1 U20927 ( .C1(n17885), .C2(n17884), .A(n17883), .B(n17882), .ZN(
        n17890) );
  NOR3_X1 U20928 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17887), .A3(
        n17886), .ZN(n17893) );
  OAI21_X1 U20929 ( .B1(n17888), .B2(n17893), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17889) );
  OAI211_X1 U20930 ( .C1(n17891), .C2(n17898), .A(n17890), .B(n17889), .ZN(
        P3_U2861) );
  AOI21_X1 U20931 ( .B1(n18380), .B2(n17892), .A(n18546), .ZN(n17895) );
  AOI221_X1 U20932 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n17896), .C1(n17895), 
        .C2(n17894), .A(n17893), .ZN(n17897) );
  OAI221_X1 U20933 ( .B1(n17901), .B2(n17900), .C1(n17899), .C2(n17898), .A(
        n17897), .ZN(P3_U2862) );
  AOI21_X1 U20934 ( .B1(n17904), .B2(n17903), .A(n17902), .ZN(n18416) );
  OAI21_X1 U20935 ( .B1(n18416), .B2(n17905), .A(n17910), .ZN(n17906) );
  OAI221_X1 U20936 ( .B1(n18166), .B2(n18568), .C1(n18166), .C2(n17910), .A(
        n17906), .ZN(P3_U2863) );
  INV_X1 U20937 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18398) );
  NOR2_X1 U20938 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18390), .ZN(
        n18095) );
  NOR2_X1 U20939 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18398), .ZN(
        n18189) );
  NOR2_X1 U20940 ( .A1(n18095), .A2(n18189), .ZN(n17908) );
  OAI22_X1 U20941 ( .A1(n17909), .A2(n18398), .B1(n17908), .B2(n17907), .ZN(
        P3_U2866) );
  NOR2_X1 U20942 ( .A1(n18399), .A2(n17910), .ZN(P3_U2867) );
  NAND2_X1 U20943 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18385), .ZN(
        n18146) );
  INV_X1 U20944 ( .A(n18146), .ZN(n18049) );
  NOR2_X1 U20945 ( .A1(n18390), .A2(n18398), .ZN(n18238) );
  NAND2_X1 U20946 ( .A1(n18049), .A2(n18238), .ZN(n18323) );
  INV_X1 U20947 ( .A(n18323), .ZN(n18343) );
  NOR2_X1 U20948 ( .A1(n18398), .A2(n18071), .ZN(n18297) );
  NAND2_X1 U20949 ( .A1(n18297), .A2(n18166), .ZN(n18293) );
  INV_X1 U20950 ( .A(n18293), .ZN(n18277) );
  NOR2_X1 U20951 ( .A1(n18343), .A2(n18277), .ZN(n18260) );
  NOR2_X1 U20952 ( .A1(n18166), .A2(n18520), .ZN(n17911) );
  NAND2_X1 U20953 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18384) );
  INV_X1 U20954 ( .A(n18384), .ZN(n18190) );
  NAND2_X1 U20955 ( .A1(n18190), .A2(n18238), .ZN(n18352) );
  INV_X1 U20956 ( .A(n18352), .ZN(n18319) );
  NAND2_X1 U20957 ( .A1(n18385), .A2(n18166), .ZN(n18386) );
  NAND2_X1 U20958 ( .A1(n18390), .A2(n18398), .ZN(n17985) );
  OR2_X1 U20959 ( .A1(n18386), .A2(n17985), .ZN(n17992) );
  NOR2_X1 U20960 ( .A1(n18319), .A2(n18024), .ZN(n17986) );
  OAI22_X1 U20961 ( .A1(n18261), .A2(n18260), .B1(n17911), .B2(n17986), .ZN(
        n17912) );
  AND2_X1 U20962 ( .A1(n17912), .A2(n18264), .ZN(n17965) );
  NAND2_X1 U20963 ( .A1(n18299), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18303) );
  NOR2_X2 U20964 ( .A1(n18119), .A2(n17913), .ZN(n18295) );
  NOR2_X1 U20965 ( .A1(n18429), .A2(n17986), .ZN(n17956) );
  AOI22_X1 U20966 ( .A1(n18259), .A2(n18277), .B1(n18295), .B2(n17956), .ZN(
        n17919) );
  NOR2_X1 U20967 ( .A1(n17915), .A2(n17914), .ZN(n17960) );
  INV_X1 U20968 ( .A(n17960), .ZN(n17932) );
  NOR2_X1 U20969 ( .A1(n17916), .A2(n17932), .ZN(n18300) );
  NOR2_X2 U20970 ( .A1(n17917), .A2(n17958), .ZN(n18294) );
  AOI22_X1 U20971 ( .A1(n18300), .A2(n18024), .B1(n18294), .B2(n18343), .ZN(
        n17918) );
  OAI211_X1 U20972 ( .C1(n17965), .C2(n17920), .A(n17919), .B(n17918), .ZN(
        P3_U2868) );
  AND2_X1 U20973 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18299), .ZN(n18306) );
  NOR2_X2 U20974 ( .A1(n18119), .A2(n17921), .ZN(n18304) );
  AOI22_X1 U20975 ( .A1(n18306), .A2(n18343), .B1(n18304), .B2(n17956), .ZN(
        n17924) );
  NAND2_X1 U20976 ( .A1(n17960), .A2(n17922), .ZN(n18309) );
  INV_X1 U20977 ( .A(n18309), .ZN(n18268) );
  NAND2_X1 U20978 ( .A1(n18299), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18271) );
  INV_X1 U20979 ( .A(n18271), .ZN(n18305) );
  AOI22_X1 U20980 ( .A1(n18268), .A2(n18024), .B1(n18305), .B2(n18277), .ZN(
        n17923) );
  OAI211_X1 U20981 ( .C1(n17965), .C2(n17925), .A(n17924), .B(n17923), .ZN(
        P3_U2869) );
  NAND2_X1 U20982 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18299), .ZN(n18316) );
  INV_X1 U20983 ( .A(n18316), .ZN(n18272) );
  NOR2_X2 U20984 ( .A1(n18119), .A2(n17926), .ZN(n18310) );
  AOI22_X1 U20985 ( .A1(n18272), .A2(n18343), .B1(n18310), .B2(n17956), .ZN(
        n17929) );
  NAND2_X1 U20986 ( .A1(n18299), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18275) );
  INV_X1 U20987 ( .A(n18275), .ZN(n18311) );
  NOR2_X2 U20988 ( .A1(n17927), .A2(n17932), .ZN(n18312) );
  AOI22_X1 U20989 ( .A1(n18311), .A2(n18277), .B1(n18312), .B2(n18024), .ZN(
        n17928) );
  OAI211_X1 U20990 ( .C1(n17965), .C2(n17930), .A(n17929), .B(n17928), .ZN(
        P3_U2870) );
  NAND2_X1 U20991 ( .A1(n18299), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18324) );
  INV_X1 U20992 ( .A(n18324), .ZN(n18276) );
  NOR2_X2 U20993 ( .A1(n18119), .A2(n17931), .ZN(n18317) );
  AOI22_X1 U20994 ( .A1(n18276), .A2(n18277), .B1(n18317), .B2(n17956), .ZN(
        n17935) );
  NOR2_X2 U20995 ( .A1(n17933), .A2(n17932), .ZN(n18320) );
  NOR2_X1 U20996 ( .A1(n19015), .A2(n17958), .ZN(n18318) );
  AOI22_X1 U20997 ( .A1(n18320), .A2(n18024), .B1(n18318), .B2(n18343), .ZN(
        n17934) );
  OAI211_X1 U20998 ( .C1(n17965), .C2(n17936), .A(n17935), .B(n17934), .ZN(
        P3_U2871) );
  NOR2_X2 U20999 ( .A1(n18119), .A2(n17937), .ZN(n18325) );
  NOR2_X2 U21000 ( .A1(n17958), .A2(n19020), .ZN(n18327) );
  AOI22_X1 U21001 ( .A1(n18325), .A2(n17956), .B1(n18327), .B2(n18277), .ZN(
        n17940) );
  AND2_X1 U21002 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18299), .ZN(n18326) );
  NAND2_X1 U21003 ( .A1(n17960), .A2(n17938), .ZN(n18330) );
  INV_X1 U21004 ( .A(n18330), .ZN(n18132) );
  AOI22_X1 U21005 ( .A1(n18326), .A2(n18343), .B1(n18132), .B2(n18024), .ZN(
        n17939) );
  OAI211_X1 U21006 ( .C1(n17965), .C2(n17941), .A(n17940), .B(n17939), .ZN(
        P3_U2872) );
  NOR2_X2 U21007 ( .A1(n14790), .A2(n17958), .ZN(n18333) );
  NOR2_X2 U21008 ( .A1(n18119), .A2(n17942), .ZN(n18331) );
  AOI22_X1 U21009 ( .A1(n18333), .A2(n18343), .B1(n18331), .B2(n17956), .ZN(
        n17947) );
  NAND2_X1 U21010 ( .A1(n17960), .A2(n17943), .ZN(n18336) );
  INV_X1 U21011 ( .A(n18336), .ZN(n17945) );
  NOR2_X2 U21012 ( .A1(n17958), .A2(n17944), .ZN(n18332) );
  AOI22_X1 U21013 ( .A1(n17945), .A2(n18024), .B1(n18332), .B2(n18277), .ZN(
        n17946) );
  OAI211_X1 U21014 ( .C1(n17965), .C2(n17948), .A(n17947), .B(n17946), .ZN(
        P3_U2873) );
  NOR2_X2 U21015 ( .A1(n12527), .A2(n17958), .ZN(n18338) );
  NOR2_X2 U21016 ( .A1(n18119), .A2(n17949), .ZN(n18337) );
  AOI22_X1 U21017 ( .A1(n18338), .A2(n18343), .B1(n18337), .B2(n17956), .ZN(
        n17953) );
  NAND2_X1 U21018 ( .A1(n17960), .A2(n17950), .ZN(n18342) );
  INV_X1 U21019 ( .A(n18342), .ZN(n17951) );
  AND2_X1 U21020 ( .A1(n18299), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U21021 ( .A1(n17951), .A2(n18024), .B1(n18339), .B2(n18277), .ZN(
        n17952) );
  OAI211_X1 U21022 ( .C1(n17965), .C2(n17954), .A(n17953), .B(n17952), .ZN(
        P3_U2874) );
  NOR2_X2 U21023 ( .A1(n17955), .A2(n18119), .ZN(n18346) );
  NOR2_X2 U21024 ( .A1(n19038), .A2(n17958), .ZN(n18344) );
  AOI22_X1 U21025 ( .A1(n18346), .A2(n17956), .B1(n18344), .B2(n18277), .ZN(
        n17963) );
  NOR2_X2 U21026 ( .A1(n17958), .A2(n17957), .ZN(n18348) );
  NAND2_X1 U21027 ( .A1(n17960), .A2(n17959), .ZN(n18353) );
  INV_X1 U21028 ( .A(n18353), .ZN(n17961) );
  AOI22_X1 U21029 ( .A1(n18348), .A2(n18343), .B1(n17961), .B2(n18024), .ZN(
        n17962) );
  OAI211_X1 U21030 ( .C1(n17965), .C2(n17964), .A(n17963), .B(n17962), .ZN(
        P3_U2875) );
  NAND2_X1 U21031 ( .A1(n18385), .A2(n18419), .ZN(n18235) );
  NOR2_X1 U21032 ( .A1(n17985), .A2(n18235), .ZN(n17981) );
  AOI22_X1 U21033 ( .A1(n18295), .A2(n17981), .B1(n18294), .B2(n18277), .ZN(
        n17968) );
  INV_X1 U21034 ( .A(n17985), .ZN(n18007) );
  NAND2_X1 U21035 ( .A1(n18264), .A2(n17966), .ZN(n18191) );
  NOR2_X1 U21036 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18191), .ZN(
        n18237) );
  AOI22_X1 U21037 ( .A1(n18299), .A2(n18297), .B1(n18007), .B2(n18237), .ZN(
        n17982) );
  NOR2_X2 U21038 ( .A1(n17985), .A2(n18146), .ZN(n18045) );
  AOI22_X1 U21039 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n17982), .B1(
        n18045), .B2(n18300), .ZN(n17967) );
  OAI211_X1 U21040 ( .C1(n18303), .C2(n18352), .A(n17968), .B(n17967), .ZN(
        P3_U2876) );
  AOI22_X1 U21041 ( .A1(n18306), .A2(n18277), .B1(n18304), .B2(n17981), .ZN(
        n17970) );
  AOI22_X1 U21042 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17982), .B1(
        n18045), .B2(n18268), .ZN(n17969) );
  OAI211_X1 U21043 ( .C1(n18271), .C2(n18352), .A(n17970), .B(n17969), .ZN(
        P3_U2877) );
  AOI22_X1 U21044 ( .A1(n18311), .A2(n18319), .B1(n18310), .B2(n17981), .ZN(
        n17972) );
  AOI22_X1 U21045 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n17982), .B1(
        n18045), .B2(n18312), .ZN(n17971) );
  OAI211_X1 U21046 ( .C1(n18316), .C2(n18293), .A(n17972), .B(n17971), .ZN(
        P3_U2878) );
  AOI22_X1 U21047 ( .A1(n18276), .A2(n18319), .B1(n18317), .B2(n17981), .ZN(
        n17974) );
  AOI22_X1 U21048 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n17982), .B1(
        n18045), .B2(n18320), .ZN(n17973) );
  OAI211_X1 U21049 ( .C1(n18281), .C2(n18293), .A(n17974), .B(n17973), .ZN(
        P3_U2879) );
  INV_X1 U21050 ( .A(n18045), .ZN(n18016) );
  AOI22_X1 U21051 ( .A1(n18326), .A2(n18277), .B1(n18325), .B2(n17981), .ZN(
        n17976) );
  AOI22_X1 U21052 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n17982), .B1(
        n18327), .B2(n18319), .ZN(n17975) );
  OAI211_X1 U21053 ( .C1(n18016), .C2(n18330), .A(n17976), .B(n17975), .ZN(
        P3_U2880) );
  AOI22_X1 U21054 ( .A1(n18332), .A2(n18319), .B1(n18331), .B2(n17981), .ZN(
        n17978) );
  AOI22_X1 U21055 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n17982), .B1(
        n18333), .B2(n18277), .ZN(n17977) );
  OAI211_X1 U21056 ( .C1(n18016), .C2(n18336), .A(n17978), .B(n17977), .ZN(
        P3_U2881) );
  AOI22_X1 U21057 ( .A1(n18338), .A2(n18277), .B1(n18337), .B2(n17981), .ZN(
        n17980) );
  AOI22_X1 U21058 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n17982), .B1(
        n18339), .B2(n18319), .ZN(n17979) );
  OAI211_X1 U21059 ( .C1(n18016), .C2(n18342), .A(n17980), .B(n17979), .ZN(
        P3_U2882) );
  AOI22_X1 U21060 ( .A1(n18346), .A2(n17981), .B1(n18344), .B2(n18319), .ZN(
        n17984) );
  AOI22_X1 U21061 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17982), .B1(
        n18348), .B2(n18277), .ZN(n17983) );
  OAI211_X1 U21062 ( .C1(n18016), .C2(n18353), .A(n17984), .B(n17983), .ZN(
        P3_U2883) );
  NOR2_X1 U21063 ( .A1(n18385), .A2(n17985), .ZN(n18050) );
  NAND2_X1 U21064 ( .A1(n18050), .A2(n18166), .ZN(n18057) );
  NOR2_X1 U21065 ( .A1(n18067), .A2(n18045), .ZN(n18028) );
  NOR2_X1 U21066 ( .A1(n18429), .A2(n18028), .ZN(n18003) );
  AOI22_X1 U21067 ( .A1(n18295), .A2(n18003), .B1(n18294), .B2(n18319), .ZN(
        n17989) );
  OAI21_X1 U21068 ( .B1(n17986), .B2(n18261), .A(n18028), .ZN(n17987) );
  OAI211_X1 U21069 ( .C1(n18067), .C2(n18520), .A(n18264), .B(n17987), .ZN(
        n18004) );
  AOI22_X1 U21070 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18004), .B1(
        n18067), .B2(n18300), .ZN(n17988) );
  OAI211_X1 U21071 ( .C1(n18303), .C2(n17992), .A(n17989), .B(n17988), .ZN(
        P3_U2884) );
  AOI22_X1 U21072 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18004), .B1(
        n18304), .B2(n18003), .ZN(n17991) );
  AOI22_X1 U21073 ( .A1(n18067), .A2(n18268), .B1(n18306), .B2(n18319), .ZN(
        n17990) );
  OAI211_X1 U21074 ( .C1(n18271), .C2(n17992), .A(n17991), .B(n17990), .ZN(
        P3_U2885) );
  AOI22_X1 U21075 ( .A1(n18311), .A2(n18024), .B1(n18310), .B2(n18003), .ZN(
        n17994) );
  AOI22_X1 U21076 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18004), .B1(
        n18067), .B2(n18312), .ZN(n17993) );
  OAI211_X1 U21077 ( .C1(n18316), .C2(n18352), .A(n17994), .B(n17993), .ZN(
        P3_U2886) );
  AOI22_X1 U21078 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18004), .B1(
        n18317), .B2(n18003), .ZN(n17996) );
  AOI22_X1 U21079 ( .A1(n18067), .A2(n18320), .B1(n18276), .B2(n18024), .ZN(
        n17995) );
  OAI211_X1 U21080 ( .C1(n18281), .C2(n18352), .A(n17996), .B(n17995), .ZN(
        P3_U2887) );
  AOI22_X1 U21081 ( .A1(n18325), .A2(n18003), .B1(n18327), .B2(n18024), .ZN(
        n17998) );
  AOI22_X1 U21082 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18004), .B1(
        n18326), .B2(n18319), .ZN(n17997) );
  OAI211_X1 U21083 ( .C1(n18057), .C2(n18330), .A(n17998), .B(n17997), .ZN(
        P3_U2888) );
  AOI22_X1 U21084 ( .A1(n18333), .A2(n18319), .B1(n18331), .B2(n18003), .ZN(
        n18000) );
  AOI22_X1 U21085 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18004), .B1(
        n18332), .B2(n18024), .ZN(n17999) );
  OAI211_X1 U21086 ( .C1(n18057), .C2(n18336), .A(n18000), .B(n17999), .ZN(
        P3_U2889) );
  AOI22_X1 U21087 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18004), .B1(
        n18337), .B2(n18003), .ZN(n18002) );
  AOI22_X1 U21088 ( .A1(n18338), .A2(n18319), .B1(n18339), .B2(n18024), .ZN(
        n18001) );
  OAI211_X1 U21089 ( .C1(n18057), .C2(n18342), .A(n18002), .B(n18001), .ZN(
        P3_U2890) );
  AOI22_X1 U21090 ( .A1(n18348), .A2(n18319), .B1(n18346), .B2(n18003), .ZN(
        n18006) );
  AOI22_X1 U21091 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18004), .B1(
        n18344), .B2(n18024), .ZN(n18005) );
  OAI211_X1 U21092 ( .C1(n18057), .C2(n18353), .A(n18006), .B(n18005), .ZN(
        P3_U2891) );
  NAND2_X1 U21093 ( .A1(n18190), .A2(n18007), .ZN(n18082) );
  INV_X1 U21094 ( .A(n18300), .ZN(n18267) );
  AND2_X1 U21095 ( .A1(n18419), .A2(n18050), .ZN(n18023) );
  AOI22_X1 U21096 ( .A1(n18295), .A2(n18023), .B1(n18294), .B2(n18024), .ZN(
        n18009) );
  AOI21_X1 U21097 ( .B1(n18385), .B2(n18261), .A(n18191), .ZN(n18094) );
  NAND2_X1 U21098 ( .A1(n18007), .A2(n18094), .ZN(n18025) );
  AOI22_X1 U21099 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18025), .B1(
        n18259), .B2(n18045), .ZN(n18008) );
  OAI211_X1 U21100 ( .C1(n18082), .C2(n18267), .A(n18009), .B(n18008), .ZN(
        P3_U2892) );
  AOI22_X1 U21101 ( .A1(n18306), .A2(n18024), .B1(n18304), .B2(n18023), .ZN(
        n18011) );
  AOI22_X1 U21102 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18025), .B1(
        n18045), .B2(n18305), .ZN(n18010) );
  OAI211_X1 U21103 ( .C1(n18082), .C2(n18309), .A(n18011), .B(n18010), .ZN(
        P3_U2893) );
  AOI22_X1 U21104 ( .A1(n18272), .A2(n18024), .B1(n18310), .B2(n18023), .ZN(
        n18013) );
  AOI22_X1 U21105 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18025), .B1(
        n18090), .B2(n18312), .ZN(n18012) );
  OAI211_X1 U21106 ( .C1(n18016), .C2(n18275), .A(n18013), .B(n18012), .ZN(
        P3_U2894) );
  AOI22_X1 U21107 ( .A1(n18318), .A2(n18024), .B1(n18317), .B2(n18023), .ZN(
        n18015) );
  AOI22_X1 U21108 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18025), .B1(
        n18090), .B2(n18320), .ZN(n18014) );
  OAI211_X1 U21109 ( .C1(n18016), .C2(n18324), .A(n18015), .B(n18014), .ZN(
        P3_U2895) );
  AOI22_X1 U21110 ( .A1(n18045), .A2(n18327), .B1(n18325), .B2(n18023), .ZN(
        n18018) );
  AOI22_X1 U21111 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18025), .B1(
        n18326), .B2(n18024), .ZN(n18017) );
  OAI211_X1 U21112 ( .C1(n18082), .C2(n18330), .A(n18018), .B(n18017), .ZN(
        P3_U2896) );
  AOI22_X1 U21113 ( .A1(n18045), .A2(n18332), .B1(n18331), .B2(n18023), .ZN(
        n18020) );
  AOI22_X1 U21114 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18025), .B1(
        n18333), .B2(n18024), .ZN(n18019) );
  OAI211_X1 U21115 ( .C1(n18082), .C2(n18336), .A(n18020), .B(n18019), .ZN(
        P3_U2897) );
  AOI22_X1 U21116 ( .A1(n18338), .A2(n18024), .B1(n18337), .B2(n18023), .ZN(
        n18022) );
  AOI22_X1 U21117 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18025), .B1(
        n18045), .B2(n18339), .ZN(n18021) );
  OAI211_X1 U21118 ( .C1(n18082), .C2(n18342), .A(n18022), .B(n18021), .ZN(
        P3_U2898) );
  AOI22_X1 U21119 ( .A1(n18348), .A2(n18024), .B1(n18346), .B2(n18023), .ZN(
        n18027) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18025), .B1(
        n18045), .B2(n18344), .ZN(n18026) );
  OAI211_X1 U21121 ( .C1(n18082), .C2(n18353), .A(n18027), .B(n18026), .ZN(
        P3_U2899) );
  INV_X1 U21122 ( .A(n18095), .ZN(n18096) );
  NOR2_X2 U21123 ( .A1(n18386), .A2(n18096), .ZN(n18113) );
  AOI21_X1 U21124 ( .B1(n18105), .B2(n18082), .A(n18429), .ZN(n18044) );
  AOI22_X1 U21125 ( .A1(n18045), .A2(n18294), .B1(n18295), .B2(n18044), .ZN(
        n18031) );
  AOI221_X1 U21126 ( .B1(n18028), .B2(n18082), .C1(n18261), .C2(n18082), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18029) );
  OAI21_X1 U21127 ( .B1(n18113), .B2(n18029), .A(n18264), .ZN(n18046) );
  AOI22_X1 U21128 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18046), .B1(
        n18113), .B2(n18300), .ZN(n18030) );
  OAI211_X1 U21129 ( .C1(n18303), .C2(n18057), .A(n18031), .B(n18030), .ZN(
        P3_U2900) );
  AOI22_X1 U21130 ( .A1(n18067), .A2(n18305), .B1(n18044), .B2(n18304), .ZN(
        n18033) );
  AOI22_X1 U21131 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18046), .B1(
        n18045), .B2(n18306), .ZN(n18032) );
  OAI211_X1 U21132 ( .C1(n18105), .C2(n18309), .A(n18033), .B(n18032), .ZN(
        P3_U2901) );
  AOI22_X1 U21133 ( .A1(n18045), .A2(n18272), .B1(n18044), .B2(n18310), .ZN(
        n18035) );
  AOI22_X1 U21134 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18046), .B1(
        n18113), .B2(n18312), .ZN(n18034) );
  OAI211_X1 U21135 ( .C1(n18057), .C2(n18275), .A(n18035), .B(n18034), .ZN(
        P3_U2902) );
  AOI22_X1 U21136 ( .A1(n18045), .A2(n18318), .B1(n18044), .B2(n18317), .ZN(
        n18037) );
  AOI22_X1 U21137 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18046), .B1(
        n18113), .B2(n18320), .ZN(n18036) );
  OAI211_X1 U21138 ( .C1(n18057), .C2(n18324), .A(n18037), .B(n18036), .ZN(
        P3_U2903) );
  AOI22_X1 U21139 ( .A1(n18067), .A2(n18327), .B1(n18044), .B2(n18325), .ZN(
        n18039) );
  AOI22_X1 U21140 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18046), .B1(
        n18045), .B2(n18326), .ZN(n18038) );
  OAI211_X1 U21141 ( .C1(n18105), .C2(n18330), .A(n18039), .B(n18038), .ZN(
        P3_U2904) );
  AOI22_X1 U21142 ( .A1(n18067), .A2(n18332), .B1(n18044), .B2(n18331), .ZN(
        n18041) );
  AOI22_X1 U21143 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18046), .B1(
        n18045), .B2(n18333), .ZN(n18040) );
  OAI211_X1 U21144 ( .C1(n18105), .C2(n18336), .A(n18041), .B(n18040), .ZN(
        P3_U2905) );
  AOI22_X1 U21145 ( .A1(n18067), .A2(n18339), .B1(n18044), .B2(n18337), .ZN(
        n18043) );
  AOI22_X1 U21146 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18046), .B1(
        n18045), .B2(n18338), .ZN(n18042) );
  OAI211_X1 U21147 ( .C1(n18105), .C2(n18342), .A(n18043), .B(n18042), .ZN(
        P3_U2906) );
  AOI22_X1 U21148 ( .A1(n18067), .A2(n18344), .B1(n18044), .B2(n18346), .ZN(
        n18048) );
  AOI22_X1 U21149 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18046), .B1(
        n18045), .B2(n18348), .ZN(n18047) );
  OAI211_X1 U21150 ( .C1(n18105), .C2(n18353), .A(n18048), .B(n18047), .ZN(
        P3_U2907) );
  NAND2_X1 U21151 ( .A1(n18095), .A2(n18049), .ZN(n18131) );
  NOR2_X1 U21152 ( .A1(n18096), .A2(n18235), .ZN(n18066) );
  AOI22_X1 U21153 ( .A1(n18067), .A2(n18294), .B1(n18295), .B2(n18066), .ZN(
        n18052) );
  AOI22_X1 U21154 ( .A1(n18299), .A2(n18050), .B1(n18095), .B2(n18237), .ZN(
        n18068) );
  AOI22_X1 U21155 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18068), .B1(
        n18259), .B2(n18090), .ZN(n18051) );
  OAI211_X1 U21156 ( .C1(n18267), .C2(n18131), .A(n18052), .B(n18051), .ZN(
        P3_U2908) );
  AOI22_X1 U21157 ( .A1(n18067), .A2(n18306), .B1(n18304), .B2(n18066), .ZN(
        n18054) );
  AOI22_X1 U21158 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18068), .B1(
        n18090), .B2(n18305), .ZN(n18053) );
  OAI211_X1 U21159 ( .C1(n18309), .C2(n18131), .A(n18054), .B(n18053), .ZN(
        P3_U2909) );
  AOI22_X1 U21160 ( .A1(n18090), .A2(n18311), .B1(n18310), .B2(n18066), .ZN(
        n18056) );
  AOI22_X1 U21161 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18068), .B1(
        n18312), .B2(n18141), .ZN(n18055) );
  OAI211_X1 U21162 ( .C1(n18057), .C2(n18316), .A(n18056), .B(n18055), .ZN(
        P3_U2910) );
  AOI22_X1 U21163 ( .A1(n18067), .A2(n18318), .B1(n18317), .B2(n18066), .ZN(
        n18059) );
  AOI22_X1 U21164 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18068), .B1(
        n18320), .B2(n18141), .ZN(n18058) );
  OAI211_X1 U21165 ( .C1(n18082), .C2(n18324), .A(n18059), .B(n18058), .ZN(
        P3_U2911) );
  AOI22_X1 U21166 ( .A1(n18067), .A2(n18326), .B1(n18325), .B2(n18066), .ZN(
        n18061) );
  AOI22_X1 U21167 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18068), .B1(
        n18090), .B2(n18327), .ZN(n18060) );
  OAI211_X1 U21168 ( .C1(n18330), .C2(n18131), .A(n18061), .B(n18060), .ZN(
        P3_U2912) );
  AOI22_X1 U21169 ( .A1(n18067), .A2(n18333), .B1(n18331), .B2(n18066), .ZN(
        n18063) );
  AOI22_X1 U21170 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18068), .B1(
        n18090), .B2(n18332), .ZN(n18062) );
  OAI211_X1 U21171 ( .C1(n18336), .C2(n18131), .A(n18063), .B(n18062), .ZN(
        P3_U2913) );
  AOI22_X1 U21172 ( .A1(n18067), .A2(n18338), .B1(n18337), .B2(n18066), .ZN(
        n18065) );
  AOI22_X1 U21173 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18068), .B1(
        n18090), .B2(n18339), .ZN(n18064) );
  OAI211_X1 U21174 ( .C1(n18342), .C2(n18131), .A(n18065), .B(n18064), .ZN(
        P3_U2914) );
  AOI22_X1 U21175 ( .A1(n18090), .A2(n18344), .B1(n18346), .B2(n18066), .ZN(
        n18070) );
  AOI22_X1 U21176 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18068), .B1(
        n18067), .B2(n18348), .ZN(n18069) );
  OAI211_X1 U21177 ( .C1(n18353), .C2(n18131), .A(n18070), .B(n18069), .ZN(
        P3_U2915) );
  NOR2_X1 U21178 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18071), .ZN(
        n18145) );
  NAND2_X1 U21179 ( .A1(n18145), .A2(n18166), .ZN(n18128) );
  AOI21_X1 U21180 ( .B1(n18131), .B2(n18128), .A(n18429), .ZN(n18089) );
  AOI22_X1 U21181 ( .A1(n18259), .A2(n18113), .B1(n18295), .B2(n18089), .ZN(
        n18075) );
  NOR2_X1 U21182 ( .A1(n18113), .A2(n18090), .ZN(n18072) );
  AOI221_X1 U21183 ( .B1(n18072), .B2(n18131), .C1(n18261), .C2(n18131), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18073) );
  OAI21_X1 U21184 ( .B1(n18161), .B2(n18073), .A(n18264), .ZN(n18091) );
  AOI22_X1 U21185 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18091), .B1(
        n18090), .B2(n18294), .ZN(n18074) );
  OAI211_X1 U21186 ( .C1(n18267), .C2(n18128), .A(n18075), .B(n18074), .ZN(
        P3_U2916) );
  AOI22_X1 U21187 ( .A1(n18113), .A2(n18305), .B1(n18304), .B2(n18089), .ZN(
        n18077) );
  AOI22_X1 U21188 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18091), .B1(
        n18090), .B2(n18306), .ZN(n18076) );
  OAI211_X1 U21189 ( .C1(n18309), .C2(n18128), .A(n18077), .B(n18076), .ZN(
        P3_U2917) );
  AOI22_X1 U21190 ( .A1(n18090), .A2(n18272), .B1(n18310), .B2(n18089), .ZN(
        n18079) );
  AOI22_X1 U21191 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18091), .B1(
        n18312), .B2(n18161), .ZN(n18078) );
  OAI211_X1 U21192 ( .C1(n18105), .C2(n18275), .A(n18079), .B(n18078), .ZN(
        P3_U2918) );
  AOI22_X1 U21193 ( .A1(n18113), .A2(n18276), .B1(n18317), .B2(n18089), .ZN(
        n18081) );
  AOI22_X1 U21194 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18091), .B1(
        n18320), .B2(n18161), .ZN(n18080) );
  OAI211_X1 U21195 ( .C1(n18082), .C2(n18281), .A(n18081), .B(n18080), .ZN(
        P3_U2919) );
  AOI22_X1 U21196 ( .A1(n18113), .A2(n18327), .B1(n18325), .B2(n18089), .ZN(
        n18084) );
  AOI22_X1 U21197 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18091), .B1(
        n18090), .B2(n18326), .ZN(n18083) );
  OAI211_X1 U21198 ( .C1(n18330), .C2(n18128), .A(n18084), .B(n18083), .ZN(
        P3_U2920) );
  AOI22_X1 U21199 ( .A1(n18113), .A2(n18332), .B1(n18331), .B2(n18089), .ZN(
        n18086) );
  AOI22_X1 U21200 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18091), .B1(
        n18090), .B2(n18333), .ZN(n18085) );
  OAI211_X1 U21201 ( .C1(n18336), .C2(n18128), .A(n18086), .B(n18085), .ZN(
        P3_U2921) );
  AOI22_X1 U21202 ( .A1(n18090), .A2(n18338), .B1(n18337), .B2(n18089), .ZN(
        n18088) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18091), .B1(
        n18113), .B2(n18339), .ZN(n18087) );
  OAI211_X1 U21204 ( .C1(n18342), .C2(n18128), .A(n18088), .B(n18087), .ZN(
        P3_U2922) );
  AOI22_X1 U21205 ( .A1(n18113), .A2(n18344), .B1(n18346), .B2(n18089), .ZN(
        n18093) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18091), .B1(
        n18090), .B2(n18348), .ZN(n18092) );
  OAI211_X1 U21207 ( .C1(n18353), .C2(n18128), .A(n18093), .B(n18092), .ZN(
        P3_U2923) );
  AND2_X1 U21208 ( .A1(n18419), .A2(n18145), .ZN(n18112) );
  AOI22_X1 U21209 ( .A1(n18113), .A2(n18294), .B1(n18295), .B2(n18112), .ZN(
        n18098) );
  NAND2_X1 U21210 ( .A1(n18095), .A2(n18094), .ZN(n18114) );
  NOR2_X2 U21211 ( .A1(n18384), .A2(n18096), .ZN(n18185) );
  AOI22_X1 U21212 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18114), .B1(
        n18300), .B2(n18185), .ZN(n18097) );
  OAI211_X1 U21213 ( .C1(n18303), .C2(n18131), .A(n18098), .B(n18097), .ZN(
        P3_U2924) );
  AOI22_X1 U21214 ( .A1(n18305), .A2(n18141), .B1(n18304), .B2(n18112), .ZN(
        n18100) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18114), .B1(
        n18113), .B2(n18306), .ZN(n18099) );
  OAI211_X1 U21216 ( .C1(n18309), .C2(n18177), .A(n18100), .B(n18099), .ZN(
        P3_U2925) );
  AOI22_X1 U21217 ( .A1(n18113), .A2(n18272), .B1(n18310), .B2(n18112), .ZN(
        n18102) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18114), .B1(
        n18312), .B2(n18185), .ZN(n18101) );
  OAI211_X1 U21219 ( .C1(n18275), .C2(n18131), .A(n18102), .B(n18101), .ZN(
        P3_U2926) );
  AOI22_X1 U21220 ( .A1(n18276), .A2(n18141), .B1(n18317), .B2(n18112), .ZN(
        n18104) );
  AOI22_X1 U21221 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18114), .B1(
        n18320), .B2(n18185), .ZN(n18103) );
  OAI211_X1 U21222 ( .C1(n18105), .C2(n18281), .A(n18104), .B(n18103), .ZN(
        P3_U2927) );
  AOI22_X1 U21223 ( .A1(n18113), .A2(n18326), .B1(n18325), .B2(n18112), .ZN(
        n18107) );
  AOI22_X1 U21224 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18114), .B1(
        n18327), .B2(n18141), .ZN(n18106) );
  OAI211_X1 U21225 ( .C1(n18330), .C2(n18177), .A(n18107), .B(n18106), .ZN(
        P3_U2928) );
  AOI22_X1 U21226 ( .A1(n18113), .A2(n18333), .B1(n18331), .B2(n18112), .ZN(
        n18109) );
  AOI22_X1 U21227 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18114), .B1(
        n18332), .B2(n18141), .ZN(n18108) );
  OAI211_X1 U21228 ( .C1(n18336), .C2(n18177), .A(n18109), .B(n18108), .ZN(
        P3_U2929) );
  AOI22_X1 U21229 ( .A1(n18113), .A2(n18338), .B1(n18337), .B2(n18112), .ZN(
        n18111) );
  AOI22_X1 U21230 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18114), .B1(
        n18339), .B2(n18141), .ZN(n18110) );
  OAI211_X1 U21231 ( .C1(n18342), .C2(n18177), .A(n18111), .B(n18110), .ZN(
        P3_U2930) );
  AOI22_X1 U21232 ( .A1(n18113), .A2(n18348), .B1(n18346), .B2(n18112), .ZN(
        n18116) );
  AOI22_X1 U21233 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18114), .B1(
        n18344), .B2(n18141), .ZN(n18115) );
  OAI211_X1 U21234 ( .C1(n18353), .C2(n18177), .A(n18116), .B(n18115), .ZN(
        P3_U2931) );
  NOR2_X2 U21235 ( .A1(n18386), .A2(n18165), .ZN(n18210) );
  NAND2_X1 U21236 ( .A1(n18131), .A2(n18128), .ZN(n18117) );
  NAND2_X1 U21237 ( .A1(n18177), .A2(n18202), .ZN(n18121) );
  AOI21_X1 U21238 ( .B1(n18118), .B2(n18117), .A(n18121), .ZN(n18120) );
  AOI211_X1 U21239 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n18202), .A(n18120), 
        .B(n18119), .ZN(n18135) );
  INV_X1 U21240 ( .A(n18121), .ZN(n18167) );
  NOR2_X1 U21241 ( .A1(n18429), .A2(n18167), .ZN(n18140) );
  AOI22_X1 U21242 ( .A1(n18295), .A2(n18140), .B1(n18294), .B2(n18141), .ZN(
        n18123) );
  AOI22_X1 U21243 ( .A1(n18259), .A2(n18161), .B1(n18300), .B2(n18210), .ZN(
        n18122) );
  OAI211_X1 U21244 ( .C1(n18135), .C2(n20659), .A(n18123), .B(n18122), .ZN(
        P3_U2932) );
  AOI22_X1 U21245 ( .A1(n18305), .A2(n18161), .B1(n18304), .B2(n18140), .ZN(
        n18125) );
  INV_X1 U21246 ( .A(n18135), .ZN(n18142) );
  AOI22_X1 U21247 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18142), .B1(
        n18306), .B2(n18141), .ZN(n18124) );
  OAI211_X1 U21248 ( .C1(n18309), .C2(n18202), .A(n18125), .B(n18124), .ZN(
        P3_U2933) );
  AOI22_X1 U21249 ( .A1(n18272), .A2(n18141), .B1(n18310), .B2(n18140), .ZN(
        n18127) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18142), .B1(
        n18312), .B2(n18210), .ZN(n18126) );
  OAI211_X1 U21251 ( .C1(n18275), .C2(n18128), .A(n18127), .B(n18126), .ZN(
        P3_U2934) );
  AOI22_X1 U21252 ( .A1(n18276), .A2(n18161), .B1(n18317), .B2(n18140), .ZN(
        n18130) );
  AOI22_X1 U21253 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18142), .B1(
        n18320), .B2(n18210), .ZN(n18129) );
  OAI211_X1 U21254 ( .C1(n18281), .C2(n18131), .A(n18130), .B(n18129), .ZN(
        P3_U2935) );
  AOI22_X1 U21255 ( .A1(n18326), .A2(n18141), .B1(n18325), .B2(n18140), .ZN(
        n18134) );
  AOI22_X1 U21256 ( .A1(n18132), .A2(n18210), .B1(n18327), .B2(n18161), .ZN(
        n18133) );
  OAI211_X1 U21257 ( .C1(n18135), .C2(n20698), .A(n18134), .B(n18133), .ZN(
        P3_U2936) );
  AOI22_X1 U21258 ( .A1(n18332), .A2(n18161), .B1(n18331), .B2(n18140), .ZN(
        n18137) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18142), .B1(
        n18333), .B2(n18141), .ZN(n18136) );
  OAI211_X1 U21260 ( .C1(n18336), .C2(n18202), .A(n18137), .B(n18136), .ZN(
        P3_U2937) );
  AOI22_X1 U21261 ( .A1(n18337), .A2(n18140), .B1(n18339), .B2(n18161), .ZN(
        n18139) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18142), .B1(
        n18338), .B2(n18141), .ZN(n18138) );
  OAI211_X1 U21263 ( .C1(n18342), .C2(n18202), .A(n18139), .B(n18138), .ZN(
        P3_U2938) );
  AOI22_X1 U21264 ( .A1(n18348), .A2(n18141), .B1(n18346), .B2(n18140), .ZN(
        n18144) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18142), .B1(
        n18344), .B2(n18161), .ZN(n18143) );
  OAI211_X1 U21266 ( .C1(n18353), .C2(n18202), .A(n18144), .B(n18143), .ZN(
        P3_U2939) );
  NOR2_X1 U21267 ( .A1(n18165), .A2(n18235), .ZN(n18192) );
  AOI22_X1 U21268 ( .A1(n18295), .A2(n18192), .B1(n18294), .B2(n18161), .ZN(
        n18148) );
  AOI22_X1 U21269 ( .A1(n18299), .A2(n18145), .B1(n18189), .B2(n18237), .ZN(
        n18162) );
  NOR2_X2 U21270 ( .A1(n18146), .A2(n18165), .ZN(n18231) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18162), .B1(
        n18300), .B2(n18231), .ZN(n18147) );
  OAI211_X1 U21272 ( .C1(n18303), .C2(n18177), .A(n18148), .B(n18147), .ZN(
        P3_U2940) );
  INV_X1 U21273 ( .A(n18231), .ZN(n18199) );
  AOI22_X1 U21274 ( .A1(n18305), .A2(n18185), .B1(n18304), .B2(n18192), .ZN(
        n18150) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18162), .B1(
        n18306), .B2(n18161), .ZN(n18149) );
  OAI211_X1 U21276 ( .C1(n18309), .C2(n18199), .A(n18150), .B(n18149), .ZN(
        P3_U2941) );
  AOI22_X1 U21277 ( .A1(n18272), .A2(n18161), .B1(n18310), .B2(n18192), .ZN(
        n18152) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18162), .B1(
        n18312), .B2(n18231), .ZN(n18151) );
  OAI211_X1 U21279 ( .C1(n18275), .C2(n18177), .A(n18152), .B(n18151), .ZN(
        P3_U2942) );
  AOI22_X1 U21280 ( .A1(n18318), .A2(n18161), .B1(n18317), .B2(n18192), .ZN(
        n18154) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18162), .B1(
        n18320), .B2(n18231), .ZN(n18153) );
  OAI211_X1 U21282 ( .C1(n18324), .C2(n18177), .A(n18154), .B(n18153), .ZN(
        P3_U2943) );
  AOI22_X1 U21283 ( .A1(n18325), .A2(n18192), .B1(n18327), .B2(n18185), .ZN(
        n18156) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18162), .B1(
        n18326), .B2(n18161), .ZN(n18155) );
  OAI211_X1 U21285 ( .C1(n18330), .C2(n18199), .A(n18156), .B(n18155), .ZN(
        P3_U2944) );
  AOI22_X1 U21286 ( .A1(n18333), .A2(n18161), .B1(n18331), .B2(n18192), .ZN(
        n18158) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18162), .B1(
        n18332), .B2(n18185), .ZN(n18157) );
  OAI211_X1 U21288 ( .C1(n18336), .C2(n18199), .A(n18158), .B(n18157), .ZN(
        P3_U2945) );
  AOI22_X1 U21289 ( .A1(n18338), .A2(n18161), .B1(n18337), .B2(n18192), .ZN(
        n18160) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18162), .B1(
        n18339), .B2(n18185), .ZN(n18159) );
  OAI211_X1 U21291 ( .C1(n18342), .C2(n18199), .A(n18160), .B(n18159), .ZN(
        P3_U2946) );
  AOI22_X1 U21292 ( .A1(n18348), .A2(n18161), .B1(n18346), .B2(n18192), .ZN(
        n18164) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18162), .B1(
        n18344), .B2(n18185), .ZN(n18163) );
  OAI211_X1 U21294 ( .C1(n18353), .C2(n18199), .A(n18164), .B(n18163), .ZN(
        P3_U2947) );
  NOR2_X1 U21295 ( .A1(n18385), .A2(n18165), .ZN(n18239) );
  NAND2_X1 U21296 ( .A1(n18166), .A2(n18239), .ZN(n18248) );
  INV_X1 U21297 ( .A(n18248), .ZN(n18255) );
  NOR2_X1 U21298 ( .A1(n18231), .A2(n18255), .ZN(n18214) );
  NOR2_X1 U21299 ( .A1(n18429), .A2(n18214), .ZN(n18184) );
  AOI22_X1 U21300 ( .A1(n18295), .A2(n18184), .B1(n18294), .B2(n18185), .ZN(
        n18170) );
  OAI21_X1 U21301 ( .B1(n18167), .B2(n18261), .A(n18214), .ZN(n18168) );
  OAI211_X1 U21302 ( .C1(n18255), .C2(n18520), .A(n18264), .B(n18168), .ZN(
        n18186) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18186), .B1(
        n18300), .B2(n18255), .ZN(n18169) );
  OAI211_X1 U21304 ( .C1(n18303), .C2(n18202), .A(n18170), .B(n18169), .ZN(
        P3_U2948) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18186), .B1(
        n18304), .B2(n18184), .ZN(n18172) );
  AOI22_X1 U21306 ( .A1(n18306), .A2(n18185), .B1(n18268), .B2(n18255), .ZN(
        n18171) );
  OAI211_X1 U21307 ( .C1(n18271), .C2(n18202), .A(n18172), .B(n18171), .ZN(
        P3_U2949) );
  AOI22_X1 U21308 ( .A1(n18272), .A2(n18185), .B1(n18310), .B2(n18184), .ZN(
        n18174) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18186), .B1(
        n18312), .B2(n18255), .ZN(n18173) );
  OAI211_X1 U21310 ( .C1(n18275), .C2(n18202), .A(n18174), .B(n18173), .ZN(
        P3_U2950) );
  AOI22_X1 U21311 ( .A1(n18276), .A2(n18210), .B1(n18317), .B2(n18184), .ZN(
        n18176) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18186), .B1(
        n18320), .B2(n18255), .ZN(n18175) );
  OAI211_X1 U21313 ( .C1(n18281), .C2(n18177), .A(n18176), .B(n18175), .ZN(
        P3_U2951) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18186), .B1(
        n18325), .B2(n18184), .ZN(n18179) );
  AOI22_X1 U21315 ( .A1(n18326), .A2(n18185), .B1(n18327), .B2(n18210), .ZN(
        n18178) );
  OAI211_X1 U21316 ( .C1(n18330), .C2(n18248), .A(n18179), .B(n18178), .ZN(
        P3_U2952) );
  AOI22_X1 U21317 ( .A1(n18332), .A2(n18210), .B1(n18331), .B2(n18184), .ZN(
        n18181) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18186), .B1(
        n18333), .B2(n18185), .ZN(n18180) );
  OAI211_X1 U21319 ( .C1(n18336), .C2(n18248), .A(n18181), .B(n18180), .ZN(
        P3_U2953) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18186), .B1(
        n18337), .B2(n18184), .ZN(n18183) );
  AOI22_X1 U21321 ( .A1(n18338), .A2(n18185), .B1(n18339), .B2(n18210), .ZN(
        n18182) );
  OAI211_X1 U21322 ( .C1(n18342), .C2(n18248), .A(n18183), .B(n18182), .ZN(
        P3_U2954) );
  AOI22_X1 U21323 ( .A1(n18346), .A2(n18184), .B1(n18344), .B2(n18210), .ZN(
        n18188) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18186), .B1(
        n18348), .B2(n18185), .ZN(n18187) );
  OAI211_X1 U21325 ( .C1(n18353), .C2(n18248), .A(n18188), .B(n18187), .ZN(
        P3_U2955) );
  NAND2_X1 U21326 ( .A1(n18190), .A2(n18189), .ZN(n18280) );
  AND2_X1 U21327 ( .A1(n18419), .A2(n18239), .ZN(n18209) );
  AOI22_X1 U21328 ( .A1(n18259), .A2(n18231), .B1(n18295), .B2(n18209), .ZN(
        n18194) );
  INV_X1 U21329 ( .A(n18191), .ZN(n18296) );
  AOI22_X1 U21330 ( .A1(n18299), .A2(n18192), .B1(n18239), .B2(n18296), .ZN(
        n18211) );
  AOI22_X1 U21331 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18211), .B1(
        n18294), .B2(n18210), .ZN(n18193) );
  OAI211_X1 U21332 ( .C1(n18267), .C2(n18280), .A(n18194), .B(n18193), .ZN(
        P3_U2956) );
  AOI22_X1 U21333 ( .A1(n18305), .A2(n18231), .B1(n18304), .B2(n18209), .ZN(
        n18196) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18211), .B1(
        n18306), .B2(n18210), .ZN(n18195) );
  OAI211_X1 U21335 ( .C1(n18309), .C2(n18280), .A(n18196), .B(n18195), .ZN(
        P3_U2957) );
  AOI22_X1 U21336 ( .A1(n18272), .A2(n18210), .B1(n18310), .B2(n18209), .ZN(
        n18198) );
  INV_X1 U21337 ( .A(n18280), .ZN(n18289) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18211), .B1(
        n18312), .B2(n18289), .ZN(n18197) );
  OAI211_X1 U21339 ( .C1(n18275), .C2(n18199), .A(n18198), .B(n18197), .ZN(
        P3_U2958) );
  AOI22_X1 U21340 ( .A1(n18276), .A2(n18231), .B1(n18317), .B2(n18209), .ZN(
        n18201) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18211), .B1(
        n18320), .B2(n18289), .ZN(n18200) );
  OAI211_X1 U21342 ( .C1(n18281), .C2(n18202), .A(n18201), .B(n18200), .ZN(
        P3_U2959) );
  AOI22_X1 U21343 ( .A1(n18325), .A2(n18209), .B1(n18327), .B2(n18231), .ZN(
        n18204) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18211), .B1(
        n18326), .B2(n18210), .ZN(n18203) );
  OAI211_X1 U21345 ( .C1(n18330), .C2(n18280), .A(n18204), .B(n18203), .ZN(
        P3_U2960) );
  AOI22_X1 U21346 ( .A1(n18332), .A2(n18231), .B1(n18331), .B2(n18209), .ZN(
        n18206) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18211), .B1(
        n18333), .B2(n18210), .ZN(n18205) );
  OAI211_X1 U21348 ( .C1(n18336), .C2(n18280), .A(n18206), .B(n18205), .ZN(
        P3_U2961) );
  AOI22_X1 U21349 ( .A1(n18337), .A2(n18209), .B1(n18339), .B2(n18231), .ZN(
        n18208) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18211), .B1(
        n18338), .B2(n18210), .ZN(n18207) );
  OAI211_X1 U21351 ( .C1(n18342), .C2(n18280), .A(n18208), .B(n18207), .ZN(
        P3_U2962) );
  AOI22_X1 U21352 ( .A1(n18346), .A2(n18209), .B1(n18344), .B2(n18231), .ZN(
        n18213) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18211), .B1(
        n18348), .B2(n18210), .ZN(n18212) );
  OAI211_X1 U21354 ( .C1(n18353), .C2(n18280), .A(n18213), .B(n18212), .ZN(
        P3_U2963) );
  INV_X1 U21355 ( .A(n18238), .ZN(n18236) );
  NOR2_X2 U21356 ( .A1(n18386), .A2(n18236), .ZN(n18347) );
  AOI21_X1 U21357 ( .B1(n18315), .B2(n18280), .A(n18429), .ZN(n18230) );
  AOI22_X1 U21358 ( .A1(n18259), .A2(n18255), .B1(n18295), .B2(n18230), .ZN(
        n18217) );
  AOI221_X1 U21359 ( .B1(n18214), .B2(n18280), .C1(n18261), .C2(n18280), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18215) );
  OAI21_X1 U21360 ( .B1(n18347), .B2(n18215), .A(n18264), .ZN(n18232) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18232), .B1(
        n18294), .B2(n18231), .ZN(n18216) );
  OAI211_X1 U21362 ( .C1(n18267), .C2(n18315), .A(n18217), .B(n18216), .ZN(
        P3_U2964) );
  AOI22_X1 U21363 ( .A1(n18306), .A2(n18231), .B1(n18304), .B2(n18230), .ZN(
        n18219) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18232), .B1(
        n18305), .B2(n18255), .ZN(n18218) );
  OAI211_X1 U21365 ( .C1(n18309), .C2(n18315), .A(n18219), .B(n18218), .ZN(
        P3_U2965) );
  AOI22_X1 U21366 ( .A1(n18272), .A2(n18231), .B1(n18310), .B2(n18230), .ZN(
        n18221) );
  AOI22_X1 U21367 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18232), .B1(
        n18312), .B2(n18347), .ZN(n18220) );
  OAI211_X1 U21368 ( .C1(n18275), .C2(n18248), .A(n18221), .B(n18220), .ZN(
        P3_U2966) );
  AOI22_X1 U21369 ( .A1(n18318), .A2(n18231), .B1(n18317), .B2(n18230), .ZN(
        n18223) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18232), .B1(
        n18320), .B2(n18347), .ZN(n18222) );
  OAI211_X1 U21371 ( .C1(n18324), .C2(n18248), .A(n18223), .B(n18222), .ZN(
        P3_U2967) );
  AOI22_X1 U21372 ( .A1(n18325), .A2(n18230), .B1(n18327), .B2(n18255), .ZN(
        n18225) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18232), .B1(
        n18326), .B2(n18231), .ZN(n18224) );
  OAI211_X1 U21374 ( .C1(n18330), .C2(n18315), .A(n18225), .B(n18224), .ZN(
        P3_U2968) );
  AOI22_X1 U21375 ( .A1(n18332), .A2(n18255), .B1(n18331), .B2(n18230), .ZN(
        n18227) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18232), .B1(
        n18333), .B2(n18231), .ZN(n18226) );
  OAI211_X1 U21377 ( .C1(n18336), .C2(n18315), .A(n18227), .B(n18226), .ZN(
        P3_U2969) );
  AOI22_X1 U21378 ( .A1(n18337), .A2(n18230), .B1(n18339), .B2(n18255), .ZN(
        n18229) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18232), .B1(
        n18338), .B2(n18231), .ZN(n18228) );
  OAI211_X1 U21380 ( .C1(n18342), .C2(n18315), .A(n18229), .B(n18228), .ZN(
        P3_U2970) );
  AOI22_X1 U21381 ( .A1(n18348), .A2(n18231), .B1(n18346), .B2(n18230), .ZN(
        n18234) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18232), .B1(
        n18344), .B2(n18255), .ZN(n18233) );
  OAI211_X1 U21383 ( .C1(n18353), .C2(n18315), .A(n18234), .B(n18233), .ZN(
        P3_U2971) );
  NOR2_X1 U21384 ( .A1(n18236), .A2(n18235), .ZN(n18298) );
  AOI22_X1 U21385 ( .A1(n18259), .A2(n18289), .B1(n18295), .B2(n18298), .ZN(
        n18241) );
  AOI22_X1 U21386 ( .A1(n18299), .A2(n18239), .B1(n18238), .B2(n18237), .ZN(
        n18256) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18256), .B1(
        n18294), .B2(n18255), .ZN(n18240) );
  OAI211_X1 U21388 ( .C1(n18267), .C2(n18323), .A(n18241), .B(n18240), .ZN(
        P3_U2972) );
  AOI22_X1 U21389 ( .A1(n18306), .A2(n18255), .B1(n18304), .B2(n18298), .ZN(
        n18243) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18256), .B1(
        n18268), .B2(n18343), .ZN(n18242) );
  OAI211_X1 U21391 ( .C1(n18271), .C2(n18280), .A(n18243), .B(n18242), .ZN(
        P3_U2973) );
  AOI22_X1 U21392 ( .A1(n18311), .A2(n18289), .B1(n18310), .B2(n18298), .ZN(
        n18245) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18256), .B1(
        n18312), .B2(n18343), .ZN(n18244) );
  OAI211_X1 U21394 ( .C1(n18316), .C2(n18248), .A(n18245), .B(n18244), .ZN(
        P3_U2974) );
  AOI22_X1 U21395 ( .A1(n18276), .A2(n18289), .B1(n18317), .B2(n18298), .ZN(
        n18247) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18256), .B1(
        n18320), .B2(n18343), .ZN(n18246) );
  OAI211_X1 U21397 ( .C1(n18281), .C2(n18248), .A(n18247), .B(n18246), .ZN(
        P3_U2975) );
  AOI22_X1 U21398 ( .A1(n18326), .A2(n18255), .B1(n18325), .B2(n18298), .ZN(
        n18250) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18256), .B1(
        n18327), .B2(n18289), .ZN(n18249) );
  OAI211_X1 U21400 ( .C1(n18330), .C2(n18323), .A(n18250), .B(n18249), .ZN(
        P3_U2976) );
  AOI22_X1 U21401 ( .A1(n18332), .A2(n18289), .B1(n18331), .B2(n18298), .ZN(
        n18252) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18256), .B1(
        n18333), .B2(n18255), .ZN(n18251) );
  OAI211_X1 U21403 ( .C1(n18336), .C2(n18323), .A(n18252), .B(n18251), .ZN(
        P3_U2977) );
  AOI22_X1 U21404 ( .A1(n18337), .A2(n18298), .B1(n18339), .B2(n18289), .ZN(
        n18254) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18256), .B1(
        n18338), .B2(n18255), .ZN(n18253) );
  OAI211_X1 U21406 ( .C1(n18342), .C2(n18323), .A(n18254), .B(n18253), .ZN(
        P3_U2978) );
  AOI22_X1 U21407 ( .A1(n18346), .A2(n18298), .B1(n18344), .B2(n18289), .ZN(
        n18258) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18256), .B1(
        n18348), .B2(n18255), .ZN(n18257) );
  OAI211_X1 U21409 ( .C1(n18353), .C2(n18323), .A(n18258), .B(n18257), .ZN(
        P3_U2979) );
  NOR2_X1 U21410 ( .A1(n18429), .A2(n18260), .ZN(n18288) );
  AOI22_X1 U21411 ( .A1(n18259), .A2(n18347), .B1(n18295), .B2(n18288), .ZN(
        n18266) );
  NOR2_X1 U21412 ( .A1(n18347), .A2(n18289), .ZN(n18262) );
  OAI21_X1 U21413 ( .B1(n18262), .B2(n18261), .A(n18260), .ZN(n18263) );
  OAI211_X1 U21414 ( .C1(n18277), .C2(n18520), .A(n18264), .B(n18263), .ZN(
        n18290) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18290), .B1(
        n18294), .B2(n18289), .ZN(n18265) );
  OAI211_X1 U21416 ( .C1(n18267), .C2(n18293), .A(n18266), .B(n18265), .ZN(
        P3_U2980) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18290), .B1(
        n18304), .B2(n18288), .ZN(n18270) );
  AOI22_X1 U21418 ( .A1(n18306), .A2(n18289), .B1(n18268), .B2(n18277), .ZN(
        n18269) );
  OAI211_X1 U21419 ( .C1(n18271), .C2(n18315), .A(n18270), .B(n18269), .ZN(
        P3_U2981) );
  AOI22_X1 U21420 ( .A1(n18272), .A2(n18289), .B1(n18310), .B2(n18288), .ZN(
        n18274) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18290), .B1(
        n18312), .B2(n18277), .ZN(n18273) );
  OAI211_X1 U21422 ( .C1(n18275), .C2(n18315), .A(n18274), .B(n18273), .ZN(
        P3_U2982) );
  AOI22_X1 U21423 ( .A1(n18276), .A2(n18347), .B1(n18317), .B2(n18288), .ZN(
        n18279) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18290), .B1(
        n18320), .B2(n18277), .ZN(n18278) );
  OAI211_X1 U21425 ( .C1(n18281), .C2(n18280), .A(n18279), .B(n18278), .ZN(
        P3_U2983) );
  AOI22_X1 U21426 ( .A1(n18326), .A2(n18289), .B1(n18325), .B2(n18288), .ZN(
        n18283) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18290), .B1(
        n18327), .B2(n18347), .ZN(n18282) );
  OAI211_X1 U21428 ( .C1(n18330), .C2(n18293), .A(n18283), .B(n18282), .ZN(
        P3_U2984) );
  AOI22_X1 U21429 ( .A1(n18333), .A2(n18289), .B1(n18331), .B2(n18288), .ZN(
        n18285) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18290), .B1(
        n18332), .B2(n18347), .ZN(n18284) );
  OAI211_X1 U21431 ( .C1(n18336), .C2(n18293), .A(n18285), .B(n18284), .ZN(
        P3_U2985) );
  AOI22_X1 U21432 ( .A1(n18337), .A2(n18288), .B1(n18339), .B2(n18347), .ZN(
        n18287) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18290), .B1(
        n18338), .B2(n18289), .ZN(n18286) );
  OAI211_X1 U21434 ( .C1(n18342), .C2(n18293), .A(n18287), .B(n18286), .ZN(
        P3_U2986) );
  AOI22_X1 U21435 ( .A1(n18346), .A2(n18288), .B1(n18344), .B2(n18347), .ZN(
        n18292) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18290), .B1(
        n18348), .B2(n18289), .ZN(n18291) );
  OAI211_X1 U21437 ( .C1(n18353), .C2(n18293), .A(n18292), .B(n18291), .ZN(
        P3_U2987) );
  AND2_X1 U21438 ( .A1(n18419), .A2(n18297), .ZN(n18345) );
  AOI22_X1 U21439 ( .A1(n18295), .A2(n18345), .B1(n18294), .B2(n18347), .ZN(
        n18302) );
  AOI22_X1 U21440 ( .A1(n18299), .A2(n18298), .B1(n18297), .B2(n18296), .ZN(
        n18349) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18349), .B1(
        n18300), .B2(n18319), .ZN(n18301) );
  OAI211_X1 U21442 ( .C1(n18303), .C2(n18323), .A(n18302), .B(n18301), .ZN(
        P3_U2988) );
  AOI22_X1 U21443 ( .A1(n18305), .A2(n18343), .B1(n18304), .B2(n18345), .ZN(
        n18308) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18349), .B1(
        n18306), .B2(n18347), .ZN(n18307) );
  OAI211_X1 U21445 ( .C1(n18309), .C2(n18352), .A(n18308), .B(n18307), .ZN(
        P3_U2989) );
  AOI22_X1 U21446 ( .A1(n18311), .A2(n18343), .B1(n18310), .B2(n18345), .ZN(
        n18314) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18349), .B1(
        n18312), .B2(n18319), .ZN(n18313) );
  OAI211_X1 U21448 ( .C1(n18316), .C2(n18315), .A(n18314), .B(n18313), .ZN(
        P3_U2990) );
  AOI22_X1 U21449 ( .A1(n18318), .A2(n18347), .B1(n18317), .B2(n18345), .ZN(
        n18322) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18349), .B1(
        n18320), .B2(n18319), .ZN(n18321) );
  OAI211_X1 U21451 ( .C1(n18324), .C2(n18323), .A(n18322), .B(n18321), .ZN(
        P3_U2991) );
  AOI22_X1 U21452 ( .A1(n18326), .A2(n18347), .B1(n18325), .B2(n18345), .ZN(
        n18329) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18349), .B1(
        n18327), .B2(n18343), .ZN(n18328) );
  OAI211_X1 U21454 ( .C1(n18330), .C2(n18352), .A(n18329), .B(n18328), .ZN(
        P3_U2992) );
  AOI22_X1 U21455 ( .A1(n18332), .A2(n18343), .B1(n18331), .B2(n18345), .ZN(
        n18335) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18349), .B1(
        n18333), .B2(n18347), .ZN(n18334) );
  OAI211_X1 U21457 ( .C1(n18336), .C2(n18352), .A(n18335), .B(n18334), .ZN(
        P3_U2993) );
  AOI22_X1 U21458 ( .A1(n18338), .A2(n18347), .B1(n18337), .B2(n18345), .ZN(
        n18341) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18349), .B1(
        n18339), .B2(n18343), .ZN(n18340) );
  OAI211_X1 U21460 ( .C1(n18342), .C2(n18352), .A(n18341), .B(n18340), .ZN(
        P3_U2994) );
  AOI22_X1 U21461 ( .A1(n18346), .A2(n18345), .B1(n18344), .B2(n18343), .ZN(
        n18351) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18349), .B1(
        n18348), .B2(n18347), .ZN(n18350) );
  OAI211_X1 U21463 ( .C1(n18353), .C2(n18352), .A(n18351), .B(n18350), .ZN(
        P3_U2995) );
  NAND2_X1 U21464 ( .A1(n18535), .A2(n18371), .ZN(n18360) );
  NOR2_X1 U21465 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18354), .ZN(
        n18381) );
  INV_X1 U21466 ( .A(n18381), .ZN(n18355) );
  AOI22_X1 U21467 ( .A1(n18404), .A2(n18360), .B1(n18366), .B2(n18355), .ZN(
        n18523) );
  NOR2_X1 U21468 ( .A1(n18388), .A2(n18523), .ZN(n18365) );
  OAI21_X1 U21469 ( .B1(n18358), .B2(n18357), .A(n18356), .ZN(n18369) );
  AOI21_X1 U21470 ( .B1(n18368), .B2(n18359), .A(n18366), .ZN(n18362) );
  INV_X1 U21471 ( .A(n18360), .ZN(n18361) );
  AOI211_X1 U21472 ( .C1(n18363), .C2(n18369), .A(n18362), .B(n18361), .ZN(
        n18521) );
  NAND2_X1 U21473 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18521), .ZN(
        n18364) );
  OAI22_X1 U21474 ( .A1(n18365), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18388), .B2(n18364), .ZN(n18406) );
  AOI211_X1 U21475 ( .C1(n18535), .C2(n18542), .A(n18366), .B(n18400), .ZN(
        n18377) );
  NAND2_X1 U21476 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18378), .ZN(
        n18367) );
  AOI211_X1 U21477 ( .C1(n18368), .C2(n18367), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18542), .ZN(n18376) );
  AOI21_X1 U21478 ( .B1(n18542), .B2(n18370), .A(n18369), .ZN(n18373) );
  NAND2_X1 U21479 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18371), .ZN(
        n18372) );
  OAI22_X1 U21480 ( .A1(n18533), .A2(n18374), .B1(n18373), .B2(n18372), .ZN(
        n18375) );
  NOR3_X1 U21481 ( .A1(n18377), .A2(n18376), .A3(n18375), .ZN(n18531) );
  INV_X1 U21482 ( .A(n18388), .ZN(n18396) );
  AOI22_X1 U21483 ( .A1(n18388), .A2(n18535), .B1(n18531), .B2(n18396), .ZN(
        n18397) );
  NOR2_X1 U21484 ( .A1(n18379), .A2(n18378), .ZN(n18383) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18380), .B1(
        n18383), .B2(n18549), .ZN(n18544) );
  OAI22_X1 U21486 ( .A1(n18383), .A2(n18382), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18381), .ZN(n18540) );
  AOI222_X1 U21487 ( .A1(n18544), .A2(n18540), .B1(n18544), .B2(n18385), .C1(
        n18540), .C2(n18384), .ZN(n18387) );
  OAI21_X1 U21488 ( .B1(n18388), .B2(n18387), .A(n18386), .ZN(n18389) );
  AOI222_X1 U21489 ( .A1(n18390), .A2(n18397), .B1(n18390), .B2(n18389), .C1(
        n18397), .C2(n18389), .ZN(n18391) );
  AOI211_X1 U21490 ( .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n18406), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n18391), .ZN(n18410) );
  OAI21_X1 U21491 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18392), .ZN(n18394) );
  OAI211_X1 U21492 ( .C1(n18396), .C2(n18395), .A(n18394), .B(n18393), .ZN(
        n18409) );
  AOI21_X1 U21493 ( .B1(n18399), .B2(n18398), .A(n18397), .ZN(n18407) );
  NAND2_X1 U21494 ( .A1(n18401), .A2(n18400), .ZN(n18402) );
  AOI22_X1 U21495 ( .A1(n18404), .A2(n18562), .B1(n18403), .B2(n18402), .ZN(
        n18565) );
  OAI211_X1 U21496 ( .C1(n18407), .C2(n18406), .A(n18565), .B(n18405), .ZN(
        n18408) );
  NOR4_X1 U21497 ( .A1(n18563), .A2(n18410), .A3(n18409), .A4(n18408), .ZN(
        n18423) );
  INV_X1 U21498 ( .A(n18411), .ZN(n18579) );
  AOI22_X1 U21499 ( .A1(n18543), .A2(n18579), .B1(n18571), .B2(n17160), .ZN(
        n18412) );
  INV_X1 U21500 ( .A(n18412), .ZN(n18418) );
  OAI211_X1 U21501 ( .C1(n18414), .C2(n18413), .A(n18569), .B(n18423), .ZN(
        n18519) );
  NAND2_X1 U21502 ( .A1(n18571), .A2(n18415), .ZN(n18424) );
  NAND2_X1 U21503 ( .A1(n18519), .A2(n18424), .ZN(n18427) );
  NOR2_X1 U21504 ( .A1(n18416), .A2(n18427), .ZN(n18417) );
  MUX2_X1 U21505 ( .A(n18418), .B(n18417), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18421) );
  OR2_X1 U21506 ( .A1(n18428), .A2(n18419), .ZN(n18420) );
  OAI211_X1 U21507 ( .C1(n18423), .C2(n18422), .A(n18421), .B(n18420), .ZN(
        P3_U2996) );
  NOR2_X1 U21508 ( .A1(n18577), .A2(n18570), .ZN(n18431) );
  NOR3_X1 U21509 ( .A1(n18426), .A2(n18425), .A3(n18424), .ZN(n18434) );
  NOR3_X1 U21510 ( .A1(n18429), .A2(n18428), .A3(n18427), .ZN(n18430) );
  OR4_X1 U21511 ( .A1(n18432), .A2(n18431), .A3(n18434), .A4(n18430), .ZN(
        P3_U2997) );
  NOR4_X1 U21512 ( .A1(n18579), .A2(n18435), .A3(n18434), .A4(n18433), .ZN(
        P3_U2998) );
  AND2_X1 U21513 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18436), .ZN(
        P3_U2999) );
  AND2_X1 U21514 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18436), .ZN(
        P3_U3000) );
  AND2_X1 U21515 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18436), .ZN(
        P3_U3001) );
  AND2_X1 U21516 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18436), .ZN(
        P3_U3002) );
  AND2_X1 U21517 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18436), .ZN(
        P3_U3003) );
  INV_X1 U21518 ( .A(P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20658) );
  NOR2_X1 U21519 ( .A1(n20658), .A2(n18517), .ZN(P3_U3004) );
  AND2_X1 U21520 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18436), .ZN(
        P3_U3005) );
  AND2_X1 U21521 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18436), .ZN(
        P3_U3006) );
  INV_X1 U21522 ( .A(P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20672) );
  NOR2_X1 U21523 ( .A1(n20672), .A2(n18517), .ZN(P3_U3007) );
  AND2_X1 U21524 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18436), .ZN(
        P3_U3008) );
  AND2_X1 U21525 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18436), .ZN(
        P3_U3009) );
  AND2_X1 U21526 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18436), .ZN(
        P3_U3010) );
  AND2_X1 U21527 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18436), .ZN(
        P3_U3011) );
  AND2_X1 U21528 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18436), .ZN(
        P3_U3012) );
  AND2_X1 U21529 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18436), .ZN(
        P3_U3013) );
  AND2_X1 U21530 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18436), .ZN(
        P3_U3014) );
  AND2_X1 U21531 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18436), .ZN(
        P3_U3015) );
  AND2_X1 U21532 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18436), .ZN(
        P3_U3016) );
  AND2_X1 U21533 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18436), .ZN(
        P3_U3017) );
  INV_X1 U21534 ( .A(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20653) );
  NOR2_X1 U21535 ( .A1(n20653), .A2(n18517), .ZN(P3_U3018) );
  AND2_X1 U21536 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18436), .ZN(
        P3_U3019) );
  AND2_X1 U21537 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18436), .ZN(
        P3_U3020) );
  AND2_X1 U21538 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18436), .ZN(P3_U3021) );
  AND2_X1 U21539 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18436), .ZN(P3_U3022) );
  AND2_X1 U21540 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18436), .ZN(P3_U3023) );
  AND2_X1 U21541 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18436), .ZN(P3_U3024) );
  AND2_X1 U21542 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18436), .ZN(P3_U3025) );
  AND2_X1 U21543 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18436), .ZN(P3_U3026) );
  AND2_X1 U21544 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18436), .ZN(P3_U3027) );
  AND2_X1 U21545 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18436), .ZN(P3_U3028) );
  NOR2_X1 U21546 ( .A1(n18452), .A2(n19627), .ZN(n18447) );
  INV_X1 U21547 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18440) );
  AOI211_X1 U21548 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n18447), .B(
        n18440), .ZN(n18439) );
  NAND2_X1 U21549 ( .A1(n18571), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18445) );
  AND2_X1 U21550 ( .A1(n18445), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18451) );
  INV_X1 U21551 ( .A(NA), .ZN(n20540) );
  OAI21_X1 U21552 ( .B1(n20540), .B2(n18437), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18450) );
  INV_X1 U21553 ( .A(n18450), .ZN(n18438) );
  OAI22_X1 U21554 ( .A1(n18584), .A2(n18439), .B1(n18451), .B2(n18438), .ZN(
        P3_U3029) );
  NOR2_X1 U21555 ( .A1(n18447), .A2(n18440), .ZN(n18443) );
  NOR2_X1 U21556 ( .A1(n18441), .A2(n19627), .ZN(n18442) );
  AOI22_X1 U21557 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18443), .B1(n18442), 
        .B2(n18452), .ZN(n18444) );
  NAND3_X1 U21558 ( .A1(n18444), .A2(n18574), .A3(n18445), .ZN(P3_U3030) );
  OAI22_X1 U21559 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18445), .ZN(n18446) );
  OAI22_X1 U21560 ( .A1(n18447), .A2(n18446), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18448) );
  OAI22_X1 U21561 ( .A1(n18451), .A2(n18450), .B1(n18449), .B2(n18448), .ZN(
        P3_U3031) );
  INV_X1 U21562 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18454) );
  NAND2_X1 U21563 ( .A1(n18584), .A2(n18452), .ZN(n18498) );
  CLKBUF_X1 U21564 ( .A(n18498), .Z(n18509) );
  OAI222_X1 U21565 ( .A1(n18551), .A2(n18513), .B1(n18453), .B2(n18584), .C1(
        n18454), .C2(n18509), .ZN(P3_U3032) );
  OAI222_X1 U21566 ( .A1(n18509), .A2(n18456), .B1(n18455), .B2(n18584), .C1(
        n18454), .C2(n18513), .ZN(P3_U3033) );
  OAI222_X1 U21567 ( .A1(n18498), .A2(n18458), .B1(n18457), .B2(n18584), .C1(
        n18456), .C2(n18513), .ZN(P3_U3034) );
  OAI222_X1 U21568 ( .A1(n18498), .A2(n18460), .B1(n18459), .B2(n18584), .C1(
        n18458), .C2(n18513), .ZN(P3_U3035) );
  OAI222_X1 U21569 ( .A1(n18498), .A2(n20750), .B1(n18461), .B2(n18584), .C1(
        n18460), .C2(n18513), .ZN(P3_U3036) );
  OAI222_X1 U21570 ( .A1(n18498), .A2(n18463), .B1(n18462), .B2(n18584), .C1(
        n20750), .C2(n18513), .ZN(P3_U3037) );
  OAI222_X1 U21571 ( .A1(n18498), .A2(n18465), .B1(n18464), .B2(n18584), .C1(
        n18463), .C2(n18513), .ZN(P3_U3038) );
  OAI222_X1 U21572 ( .A1(n18509), .A2(n18467), .B1(n18466), .B2(n18584), .C1(
        n18465), .C2(n18513), .ZN(P3_U3039) );
  OAI222_X1 U21573 ( .A1(n18509), .A2(n18469), .B1(n18468), .B2(n18584), .C1(
        n18467), .C2(n18513), .ZN(P3_U3040) );
  INV_X1 U21574 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18471) );
  OAI222_X1 U21575 ( .A1(n18509), .A2(n18471), .B1(n18470), .B2(n18584), .C1(
        n18469), .C2(n18513), .ZN(P3_U3041) );
  OAI222_X1 U21576 ( .A1(n18509), .A2(n18472), .B1(n20733), .B2(n18584), .C1(
        n18471), .C2(n18513), .ZN(P3_U3042) );
  OAI222_X1 U21577 ( .A1(n18509), .A2(n18474), .B1(n18473), .B2(n18584), .C1(
        n18472), .C2(n18513), .ZN(P3_U3043) );
  OAI222_X1 U21578 ( .A1(n18509), .A2(n18477), .B1(n18475), .B2(n18584), .C1(
        n18474), .C2(n18513), .ZN(P3_U3044) );
  OAI222_X1 U21579 ( .A1(n18477), .A2(n18513), .B1(n18476), .B2(n18584), .C1(
        n18478), .C2(n18509), .ZN(P3_U3045) );
  OAI222_X1 U21580 ( .A1(n18498), .A2(n18480), .B1(n18479), .B2(n18584), .C1(
        n18478), .C2(n18513), .ZN(P3_U3046) );
  INV_X1 U21581 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18482) );
  OAI222_X1 U21582 ( .A1(n18498), .A2(n18482), .B1(n18481), .B2(n18584), .C1(
        n18480), .C2(n18513), .ZN(P3_U3047) );
  OAI222_X1 U21583 ( .A1(n18498), .A2(n18484), .B1(n18483), .B2(n18584), .C1(
        n18482), .C2(n18513), .ZN(P3_U3048) );
  INV_X1 U21584 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18486) );
  OAI222_X1 U21585 ( .A1(n18498), .A2(n18486), .B1(n18485), .B2(n18584), .C1(
        n18484), .C2(n18513), .ZN(P3_U3049) );
  OAI222_X1 U21586 ( .A1(n18498), .A2(n18488), .B1(n18487), .B2(n18584), .C1(
        n18486), .C2(n18513), .ZN(P3_U3050) );
  OAI222_X1 U21587 ( .A1(n18498), .A2(n18491), .B1(n18489), .B2(n18584), .C1(
        n18488), .C2(n18513), .ZN(P3_U3051) );
  INV_X1 U21588 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18492) );
  OAI222_X1 U21589 ( .A1(n18491), .A2(n18513), .B1(n18490), .B2(n18584), .C1(
        n18492), .C2(n18509), .ZN(P3_U3052) );
  OAI222_X1 U21590 ( .A1(n18509), .A2(n18495), .B1(n18493), .B2(n18584), .C1(
        n18492), .C2(n18513), .ZN(P3_U3053) );
  OAI222_X1 U21591 ( .A1(n18495), .A2(n18513), .B1(n18494), .B2(n18584), .C1(
        n18496), .C2(n18509), .ZN(P3_U3054) );
  OAI222_X1 U21592 ( .A1(n18498), .A2(n18499), .B1(n18497), .B2(n18584), .C1(
        n18496), .C2(n18513), .ZN(P3_U3055) );
  OAI222_X1 U21593 ( .A1(n18509), .A2(n18501), .B1(n18500), .B2(n18584), .C1(
        n18499), .C2(n18513), .ZN(P3_U3056) );
  OAI222_X1 U21594 ( .A1(n18509), .A2(n18503), .B1(n18502), .B2(n18584), .C1(
        n18501), .C2(n18513), .ZN(P3_U3057) );
  OAI222_X1 U21595 ( .A1(n18509), .A2(n18506), .B1(n18504), .B2(n18584), .C1(
        n18503), .C2(n18513), .ZN(P3_U3058) );
  OAI222_X1 U21596 ( .A1(n18506), .A2(n18513), .B1(n18505), .B2(n18584), .C1(
        n18507), .C2(n18509), .ZN(P3_U3059) );
  OAI222_X1 U21597 ( .A1(n18509), .A2(n18512), .B1(n18508), .B2(n18584), .C1(
        n18507), .C2(n18513), .ZN(P3_U3060) );
  OAI222_X1 U21598 ( .A1(n18513), .A2(n18512), .B1(n18511), .B2(n18584), .C1(
        n18510), .C2(n18509), .ZN(P3_U3061) );
  MUX2_X1 U21599 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n18584), .Z(P3_U3274) );
  MUX2_X1 U21600 ( .A(P3_BE_N_REG_2__SCAN_IN), .B(P3_BYTEENABLE_REG_2__SCAN_IN), .S(n18584), .Z(P3_U3275) );
  MUX2_X1 U21601 ( .A(P3_BE_N_REG_1__SCAN_IN), .B(P3_BYTEENABLE_REG_1__SCAN_IN), .S(n18584), .Z(P3_U3276) );
  INV_X1 U21602 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18558) );
  INV_X1 U21603 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18514) );
  AOI22_X1 U21604 ( .A1(n18584), .A2(n18558), .B1(n18514), .B2(n18585), .ZN(
        P3_U3277) );
  OAI21_X1 U21605 ( .B1(n18517), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18516), 
        .ZN(n18515) );
  INV_X1 U21606 ( .A(n18515), .ZN(P3_U3280) );
  INV_X1 U21607 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20699) );
  OAI21_X1 U21608 ( .B1(n18517), .B2(n20699), .A(n18516), .ZN(P3_U3281) );
  OAI221_X1 U21609 ( .B1(n18520), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18520), 
        .C2(n18519), .A(n18518), .ZN(P3_U3282) );
  NOR2_X1 U21610 ( .A1(n18521), .A2(n18530), .ZN(n18522) );
  NOR2_X1 U21611 ( .A1(n18522), .A2(n18550), .ZN(n18527) );
  NOR3_X1 U21612 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18523), .A3(
        n18530), .ZN(n18524) );
  AOI21_X1 U21613 ( .B1(n18543), .B2(n18525), .A(n18524), .ZN(n18526) );
  OAI22_X1 U21614 ( .A1(n18528), .A2(n18527), .B1(n18550), .B2(n18526), .ZN(
        P3_U3285) );
  AOI22_X1 U21615 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15467), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18529), .ZN(n18538) );
  NAND2_X1 U21616 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18536) );
  OAI22_X1 U21617 ( .A1(n18531), .A2(n18530), .B1(n18538), .B2(n18536), .ZN(
        n18532) );
  AOI21_X1 U21618 ( .B1(n18543), .B2(n18533), .A(n18532), .ZN(n18534) );
  AOI22_X1 U21619 ( .A1(n18550), .A2(n18535), .B1(n18534), .B2(n18547), .ZN(
        P3_U3288) );
  INV_X1 U21620 ( .A(n18536), .ZN(n18537) );
  AOI222_X1 U21621 ( .A1(n18540), .A2(n18545), .B1(n18543), .B2(n18539), .C1(
        n18538), .C2(n18537), .ZN(n18541) );
  AOI22_X1 U21622 ( .A1(n18550), .A2(n18542), .B1(n18541), .B2(n18547), .ZN(
        P3_U3289) );
  AOI222_X1 U21623 ( .A1(n18546), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18545), 
        .B2(n18544), .C1(n18549), .C2(n18543), .ZN(n18548) );
  AOI22_X1 U21624 ( .A1(n18550), .A2(n18549), .B1(n18548), .B2(n18547), .ZN(
        P3_U3290) );
  AOI22_X1 U21625 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18552), .B2(n18551), .ZN(n18556) );
  NOR2_X1 U21626 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n18553), .ZN(n18557) );
  NAND2_X1 U21627 ( .A1(P3_DATAWIDTH_REG_0__SCAN_IN), .A2(n18557), .ZN(n18555)
         );
  NAND2_X1 U21628 ( .A1(n18559), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18554) );
  OAI211_X1 U21629 ( .C1(n18559), .C2(n18556), .A(n18555), .B(n18554), .ZN(
        P3_U3292) );
  AOI21_X1 U21630 ( .B1(n18559), .B2(n18558), .A(n18557), .ZN(P3_U3293) );
  INV_X1 U21631 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n20732) );
  AOI22_X1 U21632 ( .A1(n18584), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n20732), 
        .B2(n18585), .ZN(P3_U3294) );
  AOI22_X1 U21633 ( .A1(n18563), .A2(n18562), .B1(n18561), .B2(n18560), .ZN(
        n18564) );
  NAND2_X1 U21634 ( .A1(n18565), .A2(n18564), .ZN(n18567) );
  MUX2_X1 U21635 ( .A(P3_MORE_REG_SCAN_IN), .B(n18567), .S(n18566), .Z(
        P3_U3295) );
  OAI22_X1 U21636 ( .A1(n18571), .A2(n18570), .B1(n18569), .B2(n18568), .ZN(
        n18572) );
  NOR2_X1 U21637 ( .A1(n18573), .A2(n18572), .ZN(n18583) );
  AOI21_X1 U21638 ( .B1(n18576), .B2(n18575), .A(n18574), .ZN(n18578) );
  OAI211_X1 U21639 ( .C1(n18588), .C2(n18578), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18577), .ZN(n18580) );
  AOI21_X1 U21640 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18580), .A(n18579), 
        .ZN(n18582) );
  NAND2_X1 U21641 ( .A1(n18583), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18581) );
  OAI21_X1 U21642 ( .B1(n18583), .B2(n18582), .A(n18581), .ZN(P3_U3296) );
  OAI22_X1 U21643 ( .A1(n18585), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18584), .ZN(n18586) );
  INV_X1 U21644 ( .A(n18586), .ZN(P3_U3297) );
  NAND2_X1 U21645 ( .A1(n18587), .A2(n18589), .ZN(n18592) );
  OAI22_X1 U21646 ( .A1(n18592), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18589), 
        .B2(n18588), .ZN(n18590) );
  INV_X1 U21647 ( .A(n18590), .ZN(P3_U3298) );
  OAI21_X1 U21648 ( .B1(n18592), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18591), 
        .ZN(n18593) );
  INV_X1 U21649 ( .A(n18593), .ZN(P3_U3299) );
  INV_X1 U21650 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18594) );
  NAND2_X1 U21651 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19639), .ZN(n19626) );
  AOI22_X1 U21652 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19626), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19621), .ZN(n19687) );
  OAI21_X1 U21653 ( .B1(n19621), .B2(n18594), .A(n19616), .ZN(P2_U2815) );
  INV_X1 U21654 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18597) );
  OAI22_X1 U21655 ( .A1(n18598), .A2(n18597), .B1(n18596), .B2(n18595), .ZN(
        P2_U2816) );
  AOI21_X1 U21656 ( .B1(n19621), .B2(n19639), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18599) );
  AOI22_X1 U21657 ( .A1(n19672), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18599), 
        .B2(n19735), .ZN(P2_U2817) );
  OAI21_X1 U21658 ( .B1(n19630), .B2(BS16), .A(n19687), .ZN(n19685) );
  OAI21_X1 U21659 ( .B1(n19687), .B2(n18993), .A(n19685), .ZN(P2_U2818) );
  NOR4_X1 U21660 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18603) );
  NOR4_X1 U21661 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18602) );
  NOR4_X1 U21662 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18601) );
  NOR4_X1 U21663 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18600) );
  NAND4_X1 U21664 ( .A1(n18603), .A2(n18602), .A3(n18601), .A4(n18600), .ZN(
        n18609) );
  NOR4_X1 U21665 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18607) );
  AOI211_X1 U21666 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18606) );
  NOR4_X1 U21667 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18605) );
  NOR4_X1 U21668 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18604) );
  NAND4_X1 U21669 ( .A1(n18607), .A2(n18606), .A3(n18605), .A4(n18604), .ZN(
        n18608) );
  NOR2_X1 U21670 ( .A1(n18609), .A2(n18608), .ZN(n18617) );
  INV_X1 U21671 ( .A(n18617), .ZN(n18610) );
  NOR2_X1 U21672 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18610), .ZN(n18612) );
  INV_X1 U21673 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19683) );
  AOI22_X1 U21674 ( .A1(n18612), .A2(n18826), .B1(n18610), .B2(n19683), .ZN(
        P2_U2820) );
  NOR2_X1 U21675 ( .A1(n18617), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18611)
         );
  OR4_X1 U21676 ( .A1(n18610), .A2(P2_REIP_REG_0__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A4(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18615) );
  OAI21_X1 U21677 ( .B1(n18612), .B2(n18611), .A(n18615), .ZN(P2_U2821) );
  INV_X1 U21678 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19686) );
  NAND2_X1 U21679 ( .A1(n18612), .A2(n19686), .ZN(n18616) );
  OAI21_X1 U21680 ( .B1(n18826), .B2(n19640), .A(n18617), .ZN(n18613) );
  OAI21_X1 U21681 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18617), .A(n18613), 
        .ZN(n18614) );
  OAI221_X1 U21682 ( .B1(n18616), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18616), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18614), .ZN(P2_U2822) );
  INV_X1 U21683 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20718) );
  OAI211_X1 U21684 ( .C1(n18617), .C2(n20718), .A(n18616), .B(n18615), .ZN(
        P2_U2823) );
  AOI22_X1 U21685 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18802), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18807), .ZN(n18629) );
  AOI22_X1 U21686 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n18803), .B1(n18618), 
        .B2(n18775), .ZN(n18628) );
  INV_X1 U21687 ( .A(n18619), .ZN(n18620) );
  AOI22_X1 U21688 ( .A1(n18621), .A2(n18831), .B1(n18620), .B2(n18759), .ZN(
        n18627) );
  AOI21_X1 U21689 ( .B1(n18624), .B2(n18623), .A(n18622), .ZN(n18625) );
  NAND2_X1 U21690 ( .A1(n18819), .A2(n18625), .ZN(n18626) );
  NAND4_X1 U21691 ( .A1(n18629), .A2(n18628), .A3(n18627), .A4(n18626), .ZN(
        P2_U2835) );
  AOI211_X1 U21692 ( .C1(n18632), .C2(n18631), .A(n18630), .B(n18811), .ZN(
        n18637) );
  AOI21_X1 U21693 ( .B1(P2_REIP_REG_19__SCAN_IN), .B2(n18807), .A(n18791), 
        .ZN(n18634) );
  AOI22_X1 U21694 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n18803), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18802), .ZN(n18633) );
  OAI211_X1 U21695 ( .C1(n18635), .C2(n18822), .A(n18634), .B(n18633), .ZN(
        n18636) );
  AOI211_X1 U21696 ( .C1(n18759), .C2(n18638), .A(n18637), .B(n18636), .ZN(
        n18639) );
  OAI21_X1 U21697 ( .B1(n18640), .B2(n18796), .A(n18639), .ZN(P2_U2836) );
  AOI211_X1 U21698 ( .C1(n18642), .C2(n18650), .A(n18641), .B(n18811), .ZN(
        n18647) );
  AOI21_X1 U21699 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n18807), .A(n18791), 
        .ZN(n18644) );
  AOI22_X1 U21700 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n18803), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18802), .ZN(n18643) );
  OAI211_X1 U21701 ( .C1(n18645), .C2(n18822), .A(n18644), .B(n18643), .ZN(
        n18646) );
  AOI211_X1 U21702 ( .C1(n18831), .C2(n10111), .A(n18647), .B(n18646), .ZN(
        n18648) );
  OAI21_X1 U21703 ( .B1(n18649), .B2(n18823), .A(n18648), .ZN(P2_U2837) );
  AOI22_X1 U21704 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n18803), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18802), .ZN(n18653) );
  OAI211_X1 U21705 ( .C1(n18651), .C2(n18661), .A(n18819), .B(n18650), .ZN(
        n18652) );
  OAI211_X1 U21706 ( .C1(n18822), .C2(n18654), .A(n18653), .B(n18652), .ZN(
        n18655) );
  AOI211_X1 U21707 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n18807), .A(n18791), 
        .B(n18655), .ZN(n18659) );
  AOI22_X1 U21708 ( .A1(n18657), .A2(n18759), .B1(n18656), .B2(n18831), .ZN(
        n18658) );
  OAI211_X1 U21709 ( .C1(n18661), .C2(n18660), .A(n18659), .B(n18658), .ZN(
        P2_U2838) );
  NAND2_X1 U21710 ( .A1(n9969), .A2(n18662), .ZN(n18663) );
  XOR2_X1 U21711 ( .A(n18664), .B(n18663), .Z(n18671) );
  AOI22_X1 U21712 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n18803), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18802), .ZN(n18665) );
  OAI21_X1 U21713 ( .B1(n18666), .B2(n18822), .A(n18665), .ZN(n18667) );
  AOI211_X1 U21714 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18807), .A(n18791), 
        .B(n18667), .ZN(n18670) );
  INV_X1 U21715 ( .A(n18863), .ZN(n18668) );
  AOI22_X1 U21716 ( .A1(n18668), .A2(n18759), .B1(n18841), .B2(n18831), .ZN(
        n18669) );
  OAI211_X1 U21717 ( .C1(n18811), .C2(n18671), .A(n18670), .B(n18669), .ZN(
        P2_U2839) );
  OAI22_X1 U21718 ( .A1(n18828), .A2(n18673), .B1(n18672), .B2(n18822), .ZN(
        n18674) );
  AOI211_X1 U21719 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18807), .A(n18791), 
        .B(n18674), .ZN(n18684) );
  NOR2_X1 U21720 ( .A1(n18676), .A2(n18675), .ZN(n18677) );
  XNOR2_X1 U21721 ( .A(n18678), .B(n18677), .ZN(n18682) );
  OAI22_X1 U21722 ( .A1(n18680), .A2(n18796), .B1(n18679), .B2(n18823), .ZN(
        n18681) );
  AOI21_X1 U21723 ( .B1(n18682), .B2(n18819), .A(n18681), .ZN(n18683) );
  OAI211_X1 U21724 ( .C1(n18685), .C2(n18833), .A(n18684), .B(n18683), .ZN(
        P2_U2840) );
  NAND2_X1 U21725 ( .A1(n9969), .A2(n18686), .ZN(n18687) );
  XNOR2_X1 U21726 ( .A(n18688), .B(n18687), .ZN(n18695) );
  AOI22_X1 U21727 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18802), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n18803), .ZN(n18689) );
  OAI21_X1 U21728 ( .B1(n18690), .B2(n18822), .A(n18689), .ZN(n18691) );
  AOI211_X1 U21729 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18807), .A(n18791), 
        .B(n18691), .ZN(n18694) );
  AOI22_X1 U21730 ( .A1(n18692), .A2(n18831), .B1(n18868), .B2(n18759), .ZN(
        n18693) );
  OAI211_X1 U21731 ( .C1(n18811), .C2(n18695), .A(n18694), .B(n18693), .ZN(
        P2_U2841) );
  OAI22_X1 U21732 ( .A1(n18697), .A2(n18833), .B1(n18696), .B2(n18822), .ZN(
        n18698) );
  AOI211_X1 U21733 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18807), .A(n18791), 
        .B(n18698), .ZN(n18707) );
  NOR2_X1 U21734 ( .A1(n18676), .A2(n18699), .ZN(n18700) );
  XNOR2_X1 U21735 ( .A(n18701), .B(n18700), .ZN(n18705) );
  OAI22_X1 U21736 ( .A1(n18703), .A2(n18796), .B1(n18702), .B2(n18823), .ZN(
        n18704) );
  AOI21_X1 U21737 ( .B1(n18705), .B2(n18819), .A(n18704), .ZN(n18706) );
  OAI211_X1 U21738 ( .C1(n18828), .C2(n10792), .A(n18707), .B(n18706), .ZN(
        P2_U2842) );
  NAND2_X1 U21739 ( .A1(n9969), .A2(n18708), .ZN(n18709) );
  XNOR2_X1 U21740 ( .A(n18710), .B(n18709), .ZN(n18718) );
  AOI22_X1 U21741 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(n18803), .B1(n18711), 
        .B2(n18775), .ZN(n18712) );
  OAI21_X1 U21742 ( .B1(n20739), .B2(n18833), .A(n18712), .ZN(n18713) );
  AOI211_X1 U21743 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n18807), .A(n18791), 
        .B(n18713), .ZN(n18717) );
  AOI22_X1 U21744 ( .A1(n18715), .A2(n18831), .B1(n18714), .B2(n18759), .ZN(
        n18716) );
  OAI211_X1 U21745 ( .C1(n18811), .C2(n18718), .A(n18717), .B(n18716), .ZN(
        P2_U2843) );
  NOR2_X1 U21746 ( .A1(n18676), .A2(n18719), .ZN(n18721) );
  XNOR2_X1 U21747 ( .A(n18721), .B(n18720), .ZN(n18728) );
  AOI22_X1 U21748 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18802), .B1(
        n18722), .B2(n18775), .ZN(n18723) );
  OAI211_X1 U21749 ( .C1(n10635), .C2(n18825), .A(n18723), .B(n15891), .ZN(
        n18726) );
  OAI22_X1 U21750 ( .A1(n18724), .A2(n18796), .B1(n18873), .B2(n18823), .ZN(
        n18725) );
  AOI211_X1 U21751 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n18803), .A(n18726), .B(
        n18725), .ZN(n18727) );
  OAI21_X1 U21752 ( .B1(n18811), .B2(n18728), .A(n18727), .ZN(P2_U2844) );
  AOI22_X1 U21753 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18802), .B1(
        P2_EBX_REG_10__SCAN_IN), .B2(n18803), .ZN(n18729) );
  OAI21_X1 U21754 ( .B1(n18730), .B2(n18822), .A(n18729), .ZN(n18731) );
  AOI211_X1 U21755 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n18807), .A(n18791), 
        .B(n18731), .ZN(n18738) );
  NAND2_X1 U21756 ( .A1(n9969), .A2(n18732), .ZN(n18733) );
  XNOR2_X1 U21757 ( .A(n18734), .B(n18733), .ZN(n18735) );
  AOI22_X1 U21758 ( .A1(n18736), .A2(n18831), .B1(n18819), .B2(n18735), .ZN(
        n18737) );
  OAI211_X1 U21759 ( .C1(n18876), .C2(n18823), .A(n18738), .B(n18737), .ZN(
        P2_U2845) );
  AOI22_X1 U21760 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(n18803), .B1(n18775), .B2(
        n18739), .ZN(n18740) );
  OAI21_X1 U21761 ( .B1(n18741), .B2(n18833), .A(n18740), .ZN(n18742) );
  AOI211_X1 U21762 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18807), .A(n18791), .B(
        n18742), .ZN(n18749) );
  NOR2_X1 U21763 ( .A1(n18676), .A2(n18743), .ZN(n18745) );
  XNOR2_X1 U21764 ( .A(n18745), .B(n18744), .ZN(n18746) );
  AOI22_X1 U21765 ( .A1(n18747), .A2(n18831), .B1(n18819), .B2(n18746), .ZN(
        n18748) );
  OAI211_X1 U21766 ( .C1(n18750), .C2(n18823), .A(n18749), .B(n18748), .ZN(
        P2_U2846) );
  NAND2_X1 U21767 ( .A1(n9969), .A2(n18751), .ZN(n18752) );
  XOR2_X1 U21768 ( .A(n18753), .B(n18752), .Z(n18762) );
  AOI22_X1 U21769 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(n18803), .B1(n18754), .B2(
        n18775), .ZN(n18755) );
  OAI21_X1 U21770 ( .B1(n18756), .B2(n18833), .A(n18755), .ZN(n18757) );
  AOI211_X1 U21771 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n18807), .A(n18791), .B(
        n18757), .ZN(n18761) );
  AOI22_X1 U21772 ( .A1(n18759), .A2(n18877), .B1(n18831), .B2(n18758), .ZN(
        n18760) );
  OAI211_X1 U21773 ( .C1(n18811), .C2(n18762), .A(n18761), .B(n18760), .ZN(
        P2_U2847) );
  NOR2_X1 U21774 ( .A1(n18764), .A2(n18763), .ZN(n18765) );
  XOR2_X1 U21775 ( .A(n18766), .B(n18765), .Z(n18774) );
  AOI22_X1 U21776 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18802), .B1(
        n18767), .B2(n18775), .ZN(n18768) );
  OAI211_X1 U21777 ( .C1(n10622), .C2(n18825), .A(n18768), .B(n15891), .ZN(
        n18772) );
  OAI22_X1 U21778 ( .A1(n18823), .A2(n18770), .B1(n18796), .B2(n18769), .ZN(
        n18771) );
  AOI211_X1 U21779 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n18803), .A(n18772), .B(
        n18771), .ZN(n18773) );
  OAI21_X1 U21780 ( .B1(n18811), .B2(n18774), .A(n18773), .ZN(P2_U2848) );
  OAI21_X1 U21781 ( .B1(n10618), .B2(n18825), .A(n15891), .ZN(n18779) );
  AOI22_X1 U21782 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18802), .B1(
        n18776), .B2(n18775), .ZN(n18777) );
  INV_X1 U21783 ( .A(n18777), .ZN(n18778) );
  AOI211_X1 U21784 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n18803), .A(n18779), .B(
        n18778), .ZN(n18786) );
  NAND2_X1 U21785 ( .A1(n9969), .A2(n18780), .ZN(n18781) );
  XNOR2_X1 U21786 ( .A(n18782), .B(n18781), .ZN(n18784) );
  AOI22_X1 U21787 ( .A1(n18819), .A2(n18784), .B1(n18831), .B2(n18783), .ZN(
        n18785) );
  OAI211_X1 U21788 ( .C1(n18823), .C2(n18787), .A(n18786), .B(n18785), .ZN(
        P2_U2849) );
  INV_X1 U21789 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18801) );
  OAI22_X1 U21790 ( .A1(n18789), .A2(n18833), .B1(n18788), .B2(n18822), .ZN(
        n18790) );
  AOI211_X1 U21791 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18807), .A(n18791), .B(
        n18790), .ZN(n18800) );
  NOR2_X1 U21792 ( .A1(n18676), .A2(n18792), .ZN(n18793) );
  XNOR2_X1 U21793 ( .A(n18794), .B(n18793), .ZN(n18798) );
  OAI22_X1 U21794 ( .A1(n18823), .A2(n18889), .B1(n18796), .B2(n18795), .ZN(
        n18797) );
  AOI21_X1 U21795 ( .B1(n18798), .B2(n18819), .A(n18797), .ZN(n18799) );
  OAI211_X1 U21796 ( .C1(n18828), .C2(n18801), .A(n18800), .B(n18799), .ZN(
        P2_U2850) );
  AOI22_X1 U21797 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n18803), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18802), .ZN(n18818) );
  OAI22_X1 U21798 ( .A1(n18805), .A2(n18822), .B1(n18823), .B2(n18804), .ZN(
        n18806) );
  AOI211_X1 U21799 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n18807), .A(n18791), .B(
        n18806), .ZN(n18817) );
  INV_X1 U21800 ( .A(n18808), .ZN(n18885) );
  INV_X1 U21801 ( .A(n18809), .ZN(n18847) );
  AOI22_X1 U21802 ( .A1(n18885), .A2(n18834), .B1(n18847), .B2(n18831), .ZN(
        n18816) );
  AND2_X1 U21803 ( .A1(n9969), .A2(n18810), .ZN(n18813) );
  AOI21_X1 U21804 ( .B1(n18814), .B2(n18813), .A(n18811), .ZN(n18812) );
  OAI21_X1 U21805 ( .B1(n18814), .B2(n18813), .A(n18812), .ZN(n18815) );
  NAND4_X1 U21806 ( .A1(n18818), .A2(n18817), .A3(n18816), .A4(n18815), .ZN(
        P2_U2851) );
  INV_X1 U21807 ( .A(n18820), .ZN(n18821) );
  OAI22_X1 U21808 ( .A1(n18824), .A2(n18823), .B1(n18822), .B2(n18821), .ZN(
        n18830) );
  OAI22_X1 U21809 ( .A1(n18828), .A2(n18827), .B1(n18826), .B2(n18825), .ZN(
        n18829) );
  AOI211_X1 U21810 ( .C1(n18832), .C2(n18831), .A(n18830), .B(n18829), .ZN(
        n18836) );
  AOI22_X1 U21811 ( .A1(n18802), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19276), .B2(n18834), .ZN(n18835) );
  OAI211_X1 U21812 ( .C1(n18837), .C2(n18811), .A(n18836), .B(n18835), .ZN(
        P2_U2855) );
  OR2_X1 U21813 ( .A1(n18839), .A2(n18838), .ZN(n18840) );
  NAND2_X1 U21814 ( .A1(n13603), .A2(n18840), .ZN(n18860) );
  INV_X1 U21815 ( .A(n18841), .ZN(n18842) );
  OAI22_X1 U21816 ( .A1(n18860), .A2(n18844), .B1(n18843), .B2(n18842), .ZN(
        n18845) );
  INV_X1 U21817 ( .A(n18845), .ZN(n18846) );
  OAI21_X1 U21818 ( .B1(n18851), .B2(n10807), .A(n18846), .ZN(P2_U2871) );
  INV_X1 U21819 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18850) );
  AOI22_X1 U21820 ( .A1(n18885), .A2(n18848), .B1(n18851), .B2(n18847), .ZN(
        n18849) );
  OAI21_X1 U21821 ( .B1(n18851), .B2(n18850), .A(n18849), .ZN(P2_U2883) );
  AOI22_X1 U21822 ( .A1(n18853), .A2(n18852), .B1(n18858), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18855) );
  AOI22_X1 U21823 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n18881), .B1(n18859), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n18854) );
  NAND2_X1 U21824 ( .A1(n18855), .A2(n18854), .ZN(P2_U2888) );
  AOI22_X1 U21825 ( .A1(n18857), .A2(n18856), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n18881), .ZN(n18867) );
  AOI22_X1 U21826 ( .A1(n18859), .A2(BUF1_REG_16__SCAN_IN), .B1(n18858), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18866) );
  OAI22_X1 U21827 ( .A1(n18863), .A2(n18862), .B1(n18861), .B2(n18860), .ZN(
        n18864) );
  INV_X1 U21828 ( .A(n18864), .ZN(n18865) );
  NAND3_X1 U21829 ( .A1(n18867), .A2(n18866), .A3(n18865), .ZN(P2_U2903) );
  INV_X1 U21830 ( .A(n18868), .ZN(n18870) );
  AOI22_X1 U21831 ( .A1(n18883), .A2(n18954), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n18881), .ZN(n18869) );
  OAI21_X1 U21832 ( .B1(n18890), .B2(n18870), .A(n18869), .ZN(P2_U2905) );
  AOI22_X1 U21833 ( .A1(n18883), .A2(n18871), .B1(P2_EAX_REG_11__SCAN_IN), 
        .B2(n18881), .ZN(n18872) );
  OAI21_X1 U21834 ( .B1(n18890), .B2(n18873), .A(n18872), .ZN(P2_U2908) );
  AOI22_X1 U21835 ( .A1(n18883), .A2(n18874), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n18881), .ZN(n18875) );
  OAI21_X1 U21836 ( .B1(n18890), .B2(n18876), .A(n18875), .ZN(P2_U2909) );
  INV_X1 U21837 ( .A(n18877), .ZN(n18880) );
  AOI22_X1 U21838 ( .A1(n18883), .A2(n18878), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n18881), .ZN(n18879) );
  OAI21_X1 U21839 ( .B1(n18890), .B2(n18880), .A(n18879), .ZN(P2_U2911) );
  AOI22_X1 U21840 ( .A1(n18883), .A2(n18882), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n18881), .ZN(n18888) );
  NAND3_X1 U21841 ( .A1(n18886), .A2(n18885), .A3(n18884), .ZN(n18887) );
  OAI211_X1 U21842 ( .C1(n18890), .C2(n18889), .A(n18888), .B(n18887), .ZN(
        P2_U2914) );
  NOR2_X1 U21843 ( .A1(n18911), .A2(n18891), .ZN(P2_U2920) );
  AOI22_X1 U21844 ( .A1(n18924), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18892) );
  OAI21_X1 U21845 ( .B1(n18893), .B2(n18926), .A(n18892), .ZN(P2_U2936) );
  AOI22_X1 U21846 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n18894), .B1(n18924), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n18895) );
  OAI21_X1 U21847 ( .B1(n20771), .B2(n18911), .A(n18895), .ZN(P2_U2937) );
  AOI22_X1 U21848 ( .A1(n18924), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18896) );
  OAI21_X1 U21849 ( .B1(n18897), .B2(n18926), .A(n18896), .ZN(P2_U2938) );
  AOI22_X1 U21850 ( .A1(n18924), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18898) );
  OAI21_X1 U21851 ( .B1(n18899), .B2(n18926), .A(n18898), .ZN(P2_U2939) );
  AOI22_X1 U21852 ( .A1(n18924), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18900) );
  OAI21_X1 U21853 ( .B1(n18901), .B2(n18926), .A(n18900), .ZN(P2_U2940) );
  AOI22_X1 U21854 ( .A1(n18924), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18902) );
  OAI21_X1 U21855 ( .B1(n18903), .B2(n18926), .A(n18902), .ZN(P2_U2941) );
  AOI22_X1 U21856 ( .A1(n18924), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18904) );
  OAI21_X1 U21857 ( .B1(n18905), .B2(n18926), .A(n18904), .ZN(P2_U2942) );
  AOI22_X1 U21858 ( .A1(n18924), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18906) );
  OAI21_X1 U21859 ( .B1(n18907), .B2(n18926), .A(n18906), .ZN(P2_U2943) );
  INV_X1 U21860 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n18908) );
  OAI222_X1 U21861 ( .A1(n18911), .A2(n20671), .B1(n18926), .B2(n18910), .C1(
        n18909), .C2(n18908), .ZN(P2_U2944) );
  AOI22_X1 U21862 ( .A1(n18924), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18912) );
  OAI21_X1 U21863 ( .B1(n18913), .B2(n18926), .A(n18912), .ZN(P2_U2945) );
  INV_X1 U21864 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n20763) );
  AOI22_X1 U21865 ( .A1(n18924), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18914) );
  OAI21_X1 U21866 ( .B1(n20763), .B2(n18926), .A(n18914), .ZN(P2_U2946) );
  INV_X1 U21867 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n18916) );
  AOI22_X1 U21868 ( .A1(n18924), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18915) );
  OAI21_X1 U21869 ( .B1(n18916), .B2(n18926), .A(n18915), .ZN(P2_U2947) );
  INV_X1 U21870 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18918) );
  AOI22_X1 U21871 ( .A1(n18924), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18917) );
  OAI21_X1 U21872 ( .B1(n18918), .B2(n18926), .A(n18917), .ZN(P2_U2948) );
  INV_X1 U21873 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18920) );
  AOI22_X1 U21874 ( .A1(n18924), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18919) );
  OAI21_X1 U21875 ( .B1(n18920), .B2(n18926), .A(n18919), .ZN(P2_U2949) );
  INV_X1 U21876 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18922) );
  AOI22_X1 U21877 ( .A1(n18924), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18921) );
  OAI21_X1 U21878 ( .B1(n18922), .B2(n18926), .A(n18921), .ZN(P2_U2950) );
  AOI22_X1 U21879 ( .A1(n18924), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18923), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18925) );
  OAI21_X1 U21880 ( .B1(n11028), .B2(n18926), .A(n18925), .ZN(P2_U2951) );
  AOI22_X1 U21881 ( .A1(n18959), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n18958), .ZN(n18927) );
  OAI21_X1 U21882 ( .B1(n18940), .B2(n18961), .A(n18927), .ZN(P2_U2952) );
  AOI22_X1 U21883 ( .A1(n18959), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n18928) );
  OAI21_X1 U21884 ( .B1(n19007), .B2(n18961), .A(n18928), .ZN(P2_U2953) );
  AOI22_X1 U21885 ( .A1(n18959), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n18958), .ZN(n18929) );
  OAI21_X1 U21886 ( .B1(n19011), .B2(n18961), .A(n18929), .ZN(P2_U2954) );
  AOI22_X1 U21887 ( .A1(n18959), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_19__SCAN_IN), .B2(n18958), .ZN(n18930) );
  OAI21_X1 U21888 ( .B1(n19017), .B2(n18961), .A(n18930), .ZN(P2_U2955) );
  INV_X1 U21889 ( .A(n18931), .ZN(n19024) );
  AOI22_X1 U21890 ( .A1(n18959), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n18958), .ZN(n18932) );
  OAI21_X1 U21891 ( .B1(n19024), .B2(n18961), .A(n18932), .ZN(P2_U2956) );
  AOI22_X1 U21892 ( .A1(n18959), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_21__SCAN_IN), .B2(n18958), .ZN(n18933) );
  OAI21_X1 U21893 ( .B1(n19029), .B2(n18961), .A(n18933), .ZN(P2_U2957) );
  AOI22_X1 U21894 ( .A1(n18959), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n18958), .ZN(n18934) );
  OAI21_X1 U21895 ( .B1(n19034), .B2(n18961), .A(n18934), .ZN(P2_U2958) );
  AOI22_X1 U21896 ( .A1(n18959), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n18935) );
  OAI21_X1 U21897 ( .B1(n19047), .B2(n18961), .A(n18935), .ZN(P2_U2959) );
  AOI22_X1 U21898 ( .A1(n18959), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n18958), .ZN(n18936) );
  OAI21_X1 U21899 ( .B1(n18949), .B2(n18961), .A(n18936), .ZN(P2_U2961) );
  AOI22_X1 U21900 ( .A1(n18959), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n18958), .ZN(n18937) );
  OAI21_X1 U21901 ( .B1(n18951), .B2(n18961), .A(n18937), .ZN(P2_U2964) );
  AOI22_X1 U21902 ( .A1(n18959), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n18958), .ZN(n18938) );
  OAI21_X1 U21903 ( .B1(n18953), .B2(n18961), .A(n18938), .ZN(P2_U2965) );
  AOI22_X1 U21904 ( .A1(n18959), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n18958), .ZN(n18939) );
  OAI21_X1 U21905 ( .B1(n18940), .B2(n18961), .A(n18939), .ZN(P2_U2967) );
  AOI22_X1 U21906 ( .A1(n18959), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n18941) );
  OAI21_X1 U21907 ( .B1(n19007), .B2(n18961), .A(n18941), .ZN(P2_U2968) );
  AOI22_X1 U21908 ( .A1(n18959), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n18942) );
  OAI21_X1 U21909 ( .B1(n19011), .B2(n18961), .A(n18942), .ZN(P2_U2969) );
  AOI22_X1 U21910 ( .A1(n18959), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n18958), .ZN(n18943) );
  OAI21_X1 U21911 ( .B1(n19017), .B2(n18961), .A(n18943), .ZN(P2_U2970) );
  AOI22_X1 U21912 ( .A1(n18959), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n18958), .ZN(n18944) );
  OAI21_X1 U21913 ( .B1(n19024), .B2(n18961), .A(n18944), .ZN(P2_U2971) );
  AOI22_X1 U21914 ( .A1(n18959), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n18958), .ZN(n18945) );
  OAI21_X1 U21915 ( .B1(n19029), .B2(n18961), .A(n18945), .ZN(P2_U2972) );
  AOI22_X1 U21916 ( .A1(n18959), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n18946) );
  OAI21_X1 U21917 ( .B1(n19034), .B2(n18961), .A(n18946), .ZN(P2_U2973) );
  AOI22_X1 U21918 ( .A1(n18959), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n18947) );
  OAI21_X1 U21919 ( .B1(n19047), .B2(n18961), .A(n18947), .ZN(P2_U2974) );
  AOI22_X1 U21920 ( .A1(n18959), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n18948) );
  OAI21_X1 U21921 ( .B1(n18949), .B2(n18961), .A(n18948), .ZN(P2_U2976) );
  AOI22_X1 U21922 ( .A1(n18959), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n18950) );
  OAI21_X1 U21923 ( .B1(n18951), .B2(n18961), .A(n18950), .ZN(P2_U2979) );
  AOI22_X1 U21924 ( .A1(n18959), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n18952) );
  OAI21_X1 U21925 ( .B1(n18953), .B2(n18961), .A(n18952), .ZN(P2_U2980) );
  AOI22_X1 U21926 ( .A1(n18959), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n18957) );
  NAND2_X1 U21927 ( .A1(n18955), .A2(n18954), .ZN(n18956) );
  NAND2_X1 U21928 ( .A1(n18957), .A2(n18956), .ZN(P2_U2981) );
  AOI22_X1 U21929 ( .A1(n18959), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18958), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n18960) );
  OAI21_X1 U21930 ( .B1(n18962), .B2(n18961), .A(n18960), .ZN(P2_U2982) );
  AOI21_X1 U21931 ( .B1(n18964), .B2(n18965), .A(n18963), .ZN(n18991) );
  INV_X1 U21932 ( .A(n18965), .ZN(n18966) );
  NAND2_X1 U21933 ( .A1(n18967), .A2(n18966), .ZN(n18981) );
  INV_X1 U21934 ( .A(n18968), .ZN(n18969) );
  OAI21_X1 U21935 ( .B1(n18970), .B2(n10276), .A(n18969), .ZN(n18971) );
  AOI21_X1 U21936 ( .B1(n18973), .B2(n18972), .A(n18971), .ZN(n18980) );
  NAND3_X1 U21937 ( .A1(n11303), .A2(n18975), .A3(n18974), .ZN(n18979) );
  NAND2_X1 U21938 ( .A1(n18977), .A2(n18976), .ZN(n18978) );
  AND4_X1 U21939 ( .A1(n18981), .A2(n18980), .A3(n18979), .A4(n18978), .ZN(
        n18985) );
  NAND2_X1 U21940 ( .A1(n18983), .A2(n18982), .ZN(n18984) );
  OAI211_X1 U21941 ( .C1(n18987), .C2(n18986), .A(n18985), .B(n18984), .ZN(
        n18988) );
  INV_X1 U21942 ( .A(n18988), .ZN(n18989) );
  OAI21_X1 U21943 ( .B1(n18991), .B2(n18990), .A(n18989), .ZN(P2_U3044) );
  NOR2_X1 U21944 ( .A1(n19278), .A2(n19083), .ZN(n19045) );
  AOI22_X1 U21945 ( .A1(n19555), .A2(n19599), .B1(n19546), .B2(n19045), .ZN(
        n19005) );
  NOR3_X1 U21946 ( .A1(n19599), .A2(n19692), .A3(n19078), .ZN(n18995) );
  NAND2_X1 U21947 ( .A1(n19688), .A2(n18993), .ZN(n19690) );
  INV_X1 U21948 ( .A(n19690), .ZN(n18994) );
  NOR2_X1 U21949 ( .A1(n18995), .A2(n18994), .ZN(n19003) );
  NOR2_X1 U21950 ( .A1(n18996), .A2(n13264), .ZN(n19580) );
  NOR2_X1 U21951 ( .A1(n19580), .A2(n19045), .ZN(n19002) );
  INV_X1 U21952 ( .A(n19002), .ZN(n19000) );
  INV_X1 U21953 ( .A(n19045), .ZN(n18997) );
  OAI211_X1 U21954 ( .C1(n18998), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19692), 
        .B(n18997), .ZN(n18999) );
  OAI211_X1 U21955 ( .C1(n19003), .C2(n19000), .A(n19553), .B(n18999), .ZN(
        n19049) );
  OAI21_X1 U21956 ( .B1(n10496), .B2(n19045), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19001) );
  AOI22_X1 U21957 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19049), .B1(
        n19547), .B2(n19048), .ZN(n19004) );
  OAI211_X1 U21958 ( .C1(n19558), .C2(n19074), .A(n19005), .B(n19004), .ZN(
        P2_U3048) );
  AOI22_X1 U21959 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19041), .ZN(n19426) );
  AOI22_X1 U21960 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19041), .ZN(n19565) );
  AOI22_X1 U21961 ( .A1(n19599), .A2(n19503), .B1(n19502), .B2(n19045), .ZN(
        n19009) );
  AOI22_X1 U21962 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19049), .B1(
        n19504), .B2(n19048), .ZN(n19008) );
  OAI211_X1 U21963 ( .C1(n19426), .C2(n19074), .A(n19009), .B(n19008), .ZN(
        P2_U3049) );
  AOI22_X1 U21964 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19041), .ZN(n19463) );
  AOI22_X1 U21965 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19041), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19042), .ZN(n19572) );
  AOI22_X1 U21966 ( .A1(n19599), .A2(n19508), .B1(n19507), .B2(n19045), .ZN(
        n19013) );
  AOI22_X1 U21967 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19049), .B1(
        n19509), .B2(n19048), .ZN(n19012) );
  OAI211_X1 U21968 ( .C1(n19463), .C2(n19074), .A(n19013), .B(n19012), .ZN(
        P2_U3050) );
  AOI22_X2 U21969 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19041), .ZN(n19579) );
  OAI22_X2 U21970 ( .A1(n19015), .A2(n19037), .B1(n19014), .B2(n19039), .ZN(
        n19576) );
  AOI22_X1 U21971 ( .A1(n19576), .A2(n19599), .B1(n19513), .B2(n19045), .ZN(
        n19019) );
  AOI22_X1 U21972 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19049), .B1(
        n19515), .B2(n19048), .ZN(n19018) );
  OAI211_X1 U21973 ( .C1(n19579), .C2(n19074), .A(n19019), .B(n19018), .ZN(
        P2_U3051) );
  AOI22_X1 U21974 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19041), .ZN(n19396) );
  NOR2_X2 U21975 ( .A1(n19023), .A2(n19022), .ZN(n19581) );
  AOI22_X1 U21976 ( .A1(n19599), .A2(n19584), .B1(n19581), .B2(n19045), .ZN(
        n19026) );
  NOR2_X2 U21977 ( .A1(n19024), .A2(n19046), .ZN(n19582) );
  AOI22_X1 U21978 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19049), .B1(
        n19582), .B2(n19048), .ZN(n19025) );
  OAI211_X1 U21979 ( .C1(n19587), .C2(n19074), .A(n19026), .B(n19025), .ZN(
        P2_U3052) );
  AOI22_X2 U21980 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19041), .ZN(n19594) );
  OAI22_X2 U21981 ( .A1(n19027), .A2(n19039), .B1(n14790), .B2(n19037), .ZN(
        n19591) );
  AOI22_X1 U21982 ( .A1(n19591), .A2(n19599), .B1(n19522), .B2(n19045), .ZN(
        n19031) );
  AOI22_X1 U21983 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19049), .B1(
        n19525), .B2(n19048), .ZN(n19030) );
  OAI211_X1 U21984 ( .C1(n19594), .C2(n19074), .A(n19031), .B(n19030), .ZN(
        P2_U3053) );
  AOI22_X2 U21985 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19041), .ZN(n19438) );
  OAI22_X2 U21986 ( .A1(n19032), .A2(n19039), .B1(n12527), .B2(n19037), .ZN(
        n19435) );
  AOI22_X1 U21987 ( .A1(n19435), .A2(n19599), .B1(n19528), .B2(n19045), .ZN(
        n19036) );
  AOI22_X1 U21988 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19049), .B1(
        n19529), .B2(n19048), .ZN(n19035) );
  OAI211_X1 U21989 ( .C1(n19438), .C2(n19074), .A(n19036), .B(n19035), .ZN(
        P2_U3054) );
  AOI22_X1 U21990 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19042), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19041), .ZN(n19541) );
  AOI22_X1 U21991 ( .A1(n19599), .A2(n19609), .B1(n19533), .B2(n19045), .ZN(
        n19051) );
  AOI22_X1 U21992 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19049), .B1(
        n19536), .B2(n19048), .ZN(n19050) );
  OAI211_X1 U21993 ( .C1(n19615), .C2(n19074), .A(n19051), .B(n19050), .ZN(
        P2_U3055) );
  INV_X1 U21994 ( .A(n19504), .ZN(n19560) );
  INV_X1 U21995 ( .A(n19502), .ZN(n19559) );
  OAI22_X1 U21996 ( .A1(n19076), .A2(n19560), .B1(n19075), .B2(n19559), .ZN(
        n19052) );
  INV_X1 U21997 ( .A(n19052), .ZN(n19054) );
  INV_X1 U21998 ( .A(n19426), .ZN(n19562) );
  AOI22_X1 U21999 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19071), .B1(
        n19108), .B2(n19562), .ZN(n19053) );
  OAI211_X1 U22000 ( .C1(n19565), .C2(n19074), .A(n19054), .B(n19053), .ZN(
        P2_U3057) );
  INV_X1 U22001 ( .A(n19509), .ZN(n19567) );
  INV_X1 U22002 ( .A(n19507), .ZN(n19566) );
  OAI22_X1 U22003 ( .A1(n19076), .A2(n19567), .B1(n19075), .B2(n19566), .ZN(
        n19055) );
  INV_X1 U22004 ( .A(n19055), .ZN(n19057) );
  INV_X1 U22005 ( .A(n19463), .ZN(n19569) );
  AOI22_X1 U22006 ( .A1(n19078), .A2(n19508), .B1(n19108), .B2(n19569), .ZN(
        n19056) );
  OAI211_X1 U22007 ( .C1(n19082), .C2(n19058), .A(n19057), .B(n19056), .ZN(
        P2_U3058) );
  INV_X1 U22008 ( .A(n19515), .ZN(n19574) );
  INV_X1 U22009 ( .A(n19513), .ZN(n19573) );
  OAI22_X1 U22010 ( .A1(n19076), .A2(n19574), .B1(n19075), .B2(n19573), .ZN(
        n19059) );
  INV_X1 U22011 ( .A(n19059), .ZN(n19061) );
  AOI22_X1 U22012 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19071), .B1(
        n19078), .B2(n19576), .ZN(n19060) );
  OAI211_X1 U22013 ( .C1(n19579), .C2(n19069), .A(n19061), .B(n19060), .ZN(
        P2_U3059) );
  INV_X1 U22014 ( .A(n19075), .ZN(n19062) );
  AOI22_X1 U22015 ( .A1(n19063), .A2(n19582), .B1(n19062), .B2(n19581), .ZN(
        n19065) );
  AOI22_X1 U22016 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19071), .B1(
        n19078), .B2(n19584), .ZN(n19064) );
  OAI211_X1 U22017 ( .C1(n19587), .C2(n19069), .A(n19065), .B(n19064), .ZN(
        P2_U3060) );
  INV_X1 U22018 ( .A(n19525), .ZN(n19589) );
  INV_X1 U22019 ( .A(n19522), .ZN(n19588) );
  OAI22_X1 U22020 ( .A1(n19076), .A2(n19589), .B1(n19075), .B2(n19588), .ZN(
        n19066) );
  INV_X1 U22021 ( .A(n19066), .ZN(n19068) );
  AOI22_X1 U22022 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19071), .B1(
        n19078), .B2(n19591), .ZN(n19067) );
  OAI211_X1 U22023 ( .C1(n19594), .C2(n19069), .A(n19068), .B(n19067), .ZN(
        P2_U3061) );
  INV_X1 U22024 ( .A(n19435), .ZN(n19603) );
  INV_X1 U22025 ( .A(n19529), .ZN(n19596) );
  INV_X1 U22026 ( .A(n19528), .ZN(n19595) );
  OAI22_X1 U22027 ( .A1(n19076), .A2(n19596), .B1(n19075), .B2(n19595), .ZN(
        n19070) );
  INV_X1 U22028 ( .A(n19070), .ZN(n19073) );
  INV_X1 U22029 ( .A(n19438), .ZN(n19598) );
  AOI22_X1 U22030 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19071), .B1(
        n19108), .B2(n19598), .ZN(n19072) );
  OAI211_X1 U22031 ( .C1(n19603), .C2(n19074), .A(n19073), .B(n19072), .ZN(
        P2_U3062) );
  INV_X1 U22032 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n19081) );
  INV_X1 U22033 ( .A(n19536), .ZN(n19606) );
  INV_X1 U22034 ( .A(n19533), .ZN(n19605) );
  OAI22_X1 U22035 ( .A1(n19076), .A2(n19606), .B1(n19075), .B2(n19605), .ZN(
        n19077) );
  INV_X1 U22036 ( .A(n19077), .ZN(n19080) );
  AOI22_X1 U22037 ( .A1(n19108), .A2(n19534), .B1(n19078), .B2(n19609), .ZN(
        n19079) );
  OAI211_X1 U22038 ( .C1(n19082), .C2(n19081), .A(n19080), .B(n19079), .ZN(
        P2_U3063) );
  NOR3_X2 U22039 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10562), .A3(
        n19083), .ZN(n19106) );
  OAI21_X1 U22040 ( .B1(n19084), .B2(n19106), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19086) );
  NAND2_X1 U22041 ( .A1(n19208), .A2(n19085), .ZN(n19088) );
  NAND2_X1 U22042 ( .A1(n19086), .A2(n19088), .ZN(n19107) );
  AOI22_X1 U22043 ( .A1(n19107), .A2(n19547), .B1(n19546), .B2(n19106), .ZN(
        n19093) );
  AOI21_X1 U22044 ( .B1(n19087), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19091) );
  OAI21_X1 U22045 ( .B1(n19131), .B2(n19108), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19089) );
  NAND3_X1 U22046 ( .A1(n19089), .A2(n19688), .A3(n19088), .ZN(n19090) );
  OAI211_X1 U22047 ( .C1(n19106), .C2(n19091), .A(n19090), .B(n19553), .ZN(
        n19109) );
  AOI22_X1 U22048 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19109), .B1(
        n19108), .B2(n19555), .ZN(n19092) );
  OAI211_X1 U22049 ( .C1(n19558), .C2(n19112), .A(n19093), .B(n19092), .ZN(
        P2_U3064) );
  AOI22_X1 U22050 ( .A1(n19107), .A2(n19504), .B1(n19502), .B2(n19106), .ZN(
        n19095) );
  AOI22_X1 U22051 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19109), .B1(
        n19108), .B2(n19503), .ZN(n19094) );
  OAI211_X1 U22052 ( .C1(n19426), .C2(n19112), .A(n19095), .B(n19094), .ZN(
        P2_U3065) );
  AOI22_X1 U22053 ( .A1(n19107), .A2(n19509), .B1(n19507), .B2(n19106), .ZN(
        n19097) );
  AOI22_X1 U22054 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19109), .B1(
        n19108), .B2(n19508), .ZN(n19096) );
  OAI211_X1 U22055 ( .C1(n19463), .C2(n19112), .A(n19097), .B(n19096), .ZN(
        P2_U3066) );
  AOI22_X1 U22056 ( .A1(n19107), .A2(n19515), .B1(n19513), .B2(n19106), .ZN(
        n19099) );
  AOI22_X1 U22057 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19109), .B1(
        n19108), .B2(n19576), .ZN(n19098) );
  OAI211_X1 U22058 ( .C1(n19579), .C2(n19112), .A(n19099), .B(n19098), .ZN(
        P2_U3067) );
  AOI22_X1 U22059 ( .A1(n19107), .A2(n19582), .B1(n19581), .B2(n19106), .ZN(
        n19101) );
  AOI22_X1 U22060 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19109), .B1(
        n19108), .B2(n19584), .ZN(n19100) );
  OAI211_X1 U22061 ( .C1(n19587), .C2(n19112), .A(n19101), .B(n19100), .ZN(
        P2_U3068) );
  AOI22_X1 U22062 ( .A1(n19107), .A2(n19525), .B1(n19522), .B2(n19106), .ZN(
        n19103) );
  AOI22_X1 U22063 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19109), .B1(
        n19108), .B2(n19591), .ZN(n19102) );
  OAI211_X1 U22064 ( .C1(n19594), .C2(n19112), .A(n19103), .B(n19102), .ZN(
        P2_U3069) );
  AOI22_X1 U22065 ( .A1(n19107), .A2(n19529), .B1(n19528), .B2(n19106), .ZN(
        n19105) );
  AOI22_X1 U22066 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19109), .B1(
        n19108), .B2(n19435), .ZN(n19104) );
  OAI211_X1 U22067 ( .C1(n19438), .C2(n19112), .A(n19105), .B(n19104), .ZN(
        P2_U3070) );
  AOI22_X1 U22068 ( .A1(n19107), .A2(n19536), .B1(n19533), .B2(n19106), .ZN(
        n19111) );
  AOI22_X1 U22069 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19109), .B1(
        n19108), .B2(n19609), .ZN(n19110) );
  OAI211_X1 U22070 ( .C1(n19615), .C2(n19112), .A(n19111), .B(n19110), .ZN(
        P2_U3071) );
  INV_X1 U22071 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n19115) );
  AOI22_X1 U22072 ( .A1(n19131), .A2(n19503), .B1(n19130), .B2(n19502), .ZN(
        n19114) );
  AOI22_X1 U22073 ( .A1(n19504), .A2(n19132), .B1(n19166), .B2(n19562), .ZN(
        n19113) );
  OAI211_X1 U22074 ( .C1(n19125), .C2(n19115), .A(n19114), .B(n19113), .ZN(
        P2_U3073) );
  INV_X1 U22075 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n19118) );
  AOI22_X1 U22076 ( .A1(n19569), .A2(n19166), .B1(n19130), .B2(n19507), .ZN(
        n19117) );
  AOI22_X1 U22077 ( .A1(n19509), .A2(n19132), .B1(n19131), .B2(n19508), .ZN(
        n19116) );
  OAI211_X1 U22078 ( .C1(n19125), .C2(n19118), .A(n19117), .B(n19116), .ZN(
        P2_U3074) );
  INV_X1 U22079 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n19121) );
  AOI22_X1 U22080 ( .A1(n19576), .A2(n19131), .B1(n19130), .B2(n19513), .ZN(
        n19120) );
  INV_X1 U22081 ( .A(n19579), .ZN(n19514) );
  AOI22_X1 U22082 ( .A1(n19515), .A2(n19132), .B1(n19166), .B2(n19514), .ZN(
        n19119) );
  OAI211_X1 U22083 ( .C1(n19125), .C2(n19121), .A(n19120), .B(n19119), .ZN(
        P2_U3075) );
  INV_X1 U22084 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n19124) );
  AOI22_X1 U22085 ( .A1(n19131), .A2(n19584), .B1(n19130), .B2(n19581), .ZN(
        n19123) );
  AOI22_X1 U22086 ( .A1(n19582), .A2(n19132), .B1(n19166), .B2(n19518), .ZN(
        n19122) );
  OAI211_X1 U22087 ( .C1(n19125), .C2(n19124), .A(n19123), .B(n19122), .ZN(
        P2_U3076) );
  INV_X1 U22088 ( .A(n19166), .ZN(n19153) );
  AOI22_X1 U22089 ( .A1(n19591), .A2(n19131), .B1(n19130), .B2(n19522), .ZN(
        n19127) );
  AOI22_X1 U22090 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19133), .B1(
        n19525), .B2(n19132), .ZN(n19126) );
  OAI211_X1 U22091 ( .C1(n19594), .C2(n19153), .A(n19127), .B(n19126), .ZN(
        P2_U3077) );
  AOI22_X1 U22092 ( .A1(n19435), .A2(n19131), .B1(n19130), .B2(n19528), .ZN(
        n19129) );
  AOI22_X1 U22093 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19133), .B1(
        n19529), .B2(n19132), .ZN(n19128) );
  OAI211_X1 U22094 ( .C1(n19438), .C2(n19153), .A(n19129), .B(n19128), .ZN(
        P2_U3078) );
  AOI22_X1 U22095 ( .A1(n19131), .A2(n19609), .B1(n19130), .B2(n19533), .ZN(
        n19135) );
  AOI22_X1 U22096 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19133), .B1(
        n19536), .B2(n19132), .ZN(n19134) );
  OAI211_X1 U22097 ( .C1(n19615), .C2(n19153), .A(n19135), .B(n19134), .ZN(
        P2_U3079) );
  NOR2_X1 U22098 ( .A1(n19170), .A2(n19278), .ZN(n19164) );
  NOR2_X1 U22099 ( .A1(n19688), .A2(n19164), .ZN(n19136) );
  OAI21_X1 U22100 ( .B1(n19137), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19136), 
        .ZN(n19144) );
  NOR2_X1 U22101 ( .A1(n19138), .A2(n19213), .ZN(n19413) );
  NAND2_X1 U22102 ( .A1(n19413), .A2(n13264), .ZN(n19147) );
  INV_X1 U22103 ( .A(n19207), .ZN(n19140) );
  OAI21_X1 U22104 ( .B1(n19166), .B2(n19202), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19141) );
  NAND2_X1 U22105 ( .A1(n19147), .A2(n19141), .ZN(n19142) );
  AND2_X1 U22106 ( .A1(n19553), .A2(n19142), .ZN(n19143) );
  INV_X1 U22107 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n20725) );
  OAI21_X1 U22108 ( .B1(n19145), .B2(n19164), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19146) );
  OAI21_X1 U22109 ( .B1(n19147), .B2(n19692), .A(n19146), .ZN(n19165) );
  AOI22_X1 U22110 ( .A1(n19165), .A2(n19547), .B1(n19546), .B2(n19164), .ZN(
        n19149) );
  AOI22_X1 U22111 ( .A1(n19166), .A2(n19555), .B1(n19202), .B2(n19493), .ZN(
        n19148) );
  OAI211_X1 U22112 ( .C1(n19150), .C2(n20725), .A(n19149), .B(n19148), .ZN(
        P2_U3080) );
  AOI22_X1 U22113 ( .A1(n19165), .A2(n19504), .B1(n19502), .B2(n19164), .ZN(
        n19152) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19167), .B1(
        n19202), .B2(n19562), .ZN(n19151) );
  OAI211_X1 U22115 ( .C1(n19565), .C2(n19153), .A(n19152), .B(n19151), .ZN(
        P2_U3081) );
  AOI22_X1 U22116 ( .A1(n19165), .A2(n19509), .B1(n19507), .B2(n19164), .ZN(
        n19155) );
  AOI22_X1 U22117 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19508), .ZN(n19154) );
  OAI211_X1 U22118 ( .C1(n19463), .C2(n19196), .A(n19155), .B(n19154), .ZN(
        P2_U3082) );
  AOI22_X1 U22119 ( .A1(n19165), .A2(n19515), .B1(n19513), .B2(n19164), .ZN(
        n19157) );
  AOI22_X1 U22120 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19576), .ZN(n19156) );
  OAI211_X1 U22121 ( .C1(n19579), .C2(n19196), .A(n19157), .B(n19156), .ZN(
        P2_U3083) );
  AOI22_X1 U22122 ( .A1(n19165), .A2(n19582), .B1(n19581), .B2(n19164), .ZN(
        n19159) );
  AOI22_X1 U22123 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19584), .ZN(n19158) );
  OAI211_X1 U22124 ( .C1(n19587), .C2(n19196), .A(n19159), .B(n19158), .ZN(
        P2_U3084) );
  AOI22_X1 U22125 ( .A1(n19165), .A2(n19525), .B1(n19522), .B2(n19164), .ZN(
        n19161) );
  AOI22_X1 U22126 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19591), .ZN(n19160) );
  OAI211_X1 U22127 ( .C1(n19594), .C2(n19196), .A(n19161), .B(n19160), .ZN(
        P2_U3085) );
  AOI22_X1 U22128 ( .A1(n19165), .A2(n19529), .B1(n19528), .B2(n19164), .ZN(
        n19163) );
  AOI22_X1 U22129 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19435), .ZN(n19162) );
  OAI211_X1 U22130 ( .C1(n19438), .C2(n19196), .A(n19163), .B(n19162), .ZN(
        P2_U3086) );
  AOI22_X1 U22131 ( .A1(n19165), .A2(n19536), .B1(n19533), .B2(n19164), .ZN(
        n19169) );
  AOI22_X1 U22132 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19167), .B1(
        n19166), .B2(n19609), .ZN(n19168) );
  OAI211_X1 U22133 ( .C1(n19615), .C2(n19196), .A(n19169), .B(n19168), .ZN(
        P2_U3087) );
  NAND2_X1 U22134 ( .A1(n19179), .A2(n19544), .ZN(n19172) );
  NOR3_X2 U22135 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19720), .A3(
        n19170), .ZN(n19201) );
  INV_X1 U22136 ( .A(n19201), .ZN(n19171) );
  NAND2_X1 U22137 ( .A1(n19172), .A2(n19171), .ZN(n19175) );
  NAND2_X1 U22138 ( .A1(n19245), .A2(n19450), .ZN(n19173) );
  NAND2_X1 U22139 ( .A1(n19212), .A2(n10562), .ZN(n19177) );
  NAND2_X1 U22140 ( .A1(n19173), .A2(n19177), .ZN(n19174) );
  MUX2_X1 U22141 ( .A(n19175), .B(n19174), .S(n19688), .Z(n19176) );
  AND2_X1 U22142 ( .A1(n19176), .A2(n19553), .ZN(n19193) );
  INV_X1 U22143 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19184) );
  AOI22_X1 U22144 ( .A1(n19202), .A2(n19555), .B1(n19546), .B2(n19201), .ZN(
        n19183) );
  INV_X1 U22145 ( .A(n19177), .ZN(n19178) );
  NAND2_X1 U22146 ( .A1(n19178), .A2(n19688), .ZN(n19181) );
  OAI21_X1 U22147 ( .B1(n19179), .B2(n19201), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19180) );
  NAND2_X1 U22148 ( .A1(n19181), .A2(n19180), .ZN(n19203) );
  AOI22_X1 U22149 ( .A1(n19547), .A2(n19203), .B1(n19234), .B2(n19493), .ZN(
        n19182) );
  OAI211_X1 U22150 ( .C1(n19193), .C2(n19184), .A(n19183), .B(n19182), .ZN(
        P2_U3088) );
  INV_X1 U22151 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19187) );
  AOI22_X1 U22152 ( .A1(n19202), .A2(n19503), .B1(n19201), .B2(n19502), .ZN(
        n19186) );
  AOI22_X1 U22153 ( .A1(n19504), .A2(n19203), .B1(n19234), .B2(n19562), .ZN(
        n19185) );
  OAI211_X1 U22154 ( .C1(n19193), .C2(n19187), .A(n19186), .B(n19185), .ZN(
        P2_U3089) );
  AOI22_X1 U22155 ( .A1(n19569), .A2(n19234), .B1(n19201), .B2(n19507), .ZN(
        n19189) );
  AOI22_X1 U22156 ( .A1(n19509), .A2(n19203), .B1(n19202), .B2(n19508), .ZN(
        n19188) );
  OAI211_X1 U22157 ( .C1(n19193), .C2(n20737), .A(n19189), .B(n19188), .ZN(
        P2_U3090) );
  INV_X1 U22158 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n19192) );
  AOI22_X1 U22159 ( .A1(n19202), .A2(n19576), .B1(n19201), .B2(n19513), .ZN(
        n19191) );
  AOI22_X1 U22160 ( .A1(n19515), .A2(n19203), .B1(n19234), .B2(n19514), .ZN(
        n19190) );
  OAI211_X1 U22161 ( .C1(n19193), .C2(n19192), .A(n19191), .B(n19190), .ZN(
        P2_U3091) );
  AOI22_X1 U22162 ( .A1(n19518), .A2(n19234), .B1(n19201), .B2(n19581), .ZN(
        n19195) );
  INV_X1 U22163 ( .A(n19193), .ZN(n19204) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19204), .B1(
        n19582), .B2(n19203), .ZN(n19194) );
  OAI211_X1 U22165 ( .C1(n19396), .C2(n19196), .A(n19195), .B(n19194), .ZN(
        P2_U3092) );
  AOI22_X1 U22166 ( .A1(n19202), .A2(n19591), .B1(n19201), .B2(n19522), .ZN(
        n19198) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19204), .B1(
        n19525), .B2(n19203), .ZN(n19197) );
  OAI211_X1 U22168 ( .C1(n19594), .C2(n19215), .A(n19198), .B(n19197), .ZN(
        P2_U3093) );
  AOI22_X1 U22169 ( .A1(n19202), .A2(n19435), .B1(n19201), .B2(n19528), .ZN(
        n19200) );
  AOI22_X1 U22170 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19204), .B1(
        n19529), .B2(n19203), .ZN(n19199) );
  OAI211_X1 U22171 ( .C1(n19438), .C2(n19215), .A(n19200), .B(n19199), .ZN(
        P2_U3094) );
  AOI22_X1 U22172 ( .A1(n19202), .A2(n19609), .B1(n19201), .B2(n19533), .ZN(
        n19206) );
  AOI22_X1 U22173 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19204), .B1(
        n19536), .B2(n19203), .ZN(n19205) );
  OAI211_X1 U22174 ( .C1(n19615), .C2(n19215), .A(n19206), .B(n19205), .ZN(
        P2_U3095) );
  INV_X1 U22175 ( .A(n19208), .ZN(n19341) );
  NAND3_X1 U22176 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n13264), .ZN(n19246) );
  NOR2_X1 U22177 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19246), .ZN(
        n19232) );
  OAI21_X1 U22178 ( .B1(n19209), .B2(n19232), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19210) );
  OAI21_X1 U22179 ( .B1(n19341), .B2(n19170), .A(n19210), .ZN(n19233) );
  AOI22_X1 U22180 ( .A1(n19233), .A2(n19547), .B1(n19546), .B2(n19232), .ZN(
        n19219) );
  AOI21_X1 U22181 ( .B1(n19211), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19217) );
  NAND2_X1 U22182 ( .A1(n19213), .A2(n19212), .ZN(n19214) );
  OAI221_X1 U22183 ( .B1(n18993), .B2(n19215), .C1(n18993), .C2(n19275), .A(
        n19214), .ZN(n19216) );
  OAI211_X1 U22184 ( .C1(n19232), .C2(n19217), .A(n19216), .B(n19553), .ZN(
        n19235) );
  AOI22_X1 U22185 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19235), .B1(
        n19234), .B2(n19555), .ZN(n19218) );
  OAI211_X1 U22186 ( .C1(n19558), .C2(n19275), .A(n19219), .B(n19218), .ZN(
        P2_U3096) );
  AOI22_X1 U22187 ( .A1(n19233), .A2(n19504), .B1(n19502), .B2(n19232), .ZN(
        n19221) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19235), .B1(
        n19234), .B2(n19503), .ZN(n19220) );
  OAI211_X1 U22189 ( .C1(n19426), .C2(n19275), .A(n19221), .B(n19220), .ZN(
        P2_U3097) );
  AOI22_X1 U22190 ( .A1(n19233), .A2(n19509), .B1(n19507), .B2(n19232), .ZN(
        n19223) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19235), .B1(
        n19234), .B2(n19508), .ZN(n19222) );
  OAI211_X1 U22192 ( .C1(n19463), .C2(n19275), .A(n19223), .B(n19222), .ZN(
        P2_U3098) );
  AOI22_X1 U22193 ( .A1(n19233), .A2(n19515), .B1(n19513), .B2(n19232), .ZN(
        n19225) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19235), .B1(
        n19234), .B2(n19576), .ZN(n19224) );
  OAI211_X1 U22195 ( .C1(n19579), .C2(n19275), .A(n19225), .B(n19224), .ZN(
        P2_U3099) );
  AOI22_X1 U22196 ( .A1(n19233), .A2(n19582), .B1(n19581), .B2(n19232), .ZN(
        n19227) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19235), .B1(
        n19234), .B2(n19584), .ZN(n19226) );
  OAI211_X1 U22198 ( .C1(n19587), .C2(n19275), .A(n19227), .B(n19226), .ZN(
        P2_U3100) );
  AOI22_X1 U22199 ( .A1(n19233), .A2(n19525), .B1(n19522), .B2(n19232), .ZN(
        n19229) );
  AOI22_X1 U22200 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19235), .B1(
        n19234), .B2(n19591), .ZN(n19228) );
  OAI211_X1 U22201 ( .C1(n19594), .C2(n19275), .A(n19229), .B(n19228), .ZN(
        P2_U3101) );
  AOI22_X1 U22202 ( .A1(n19233), .A2(n19529), .B1(n19528), .B2(n19232), .ZN(
        n19231) );
  AOI22_X1 U22203 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19235), .B1(
        n19234), .B2(n19435), .ZN(n19230) );
  OAI211_X1 U22204 ( .C1(n19438), .C2(n19275), .A(n19231), .B(n19230), .ZN(
        P2_U3102) );
  AOI22_X1 U22205 ( .A1(n19233), .A2(n19536), .B1(n19533), .B2(n19232), .ZN(
        n19237) );
  AOI22_X1 U22206 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19235), .B1(
        n19234), .B2(n19609), .ZN(n19236) );
  OAI211_X1 U22207 ( .C1(n19615), .C2(n19275), .A(n19237), .B(n19236), .ZN(
        P2_U3103) );
  NAND2_X1 U22208 ( .A1(n19281), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19239) );
  INV_X1 U22209 ( .A(n19246), .ZN(n19241) );
  NOR2_X1 U22210 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19241), .ZN(n19242) );
  NOR2_X1 U22211 ( .A1(n19243), .A2(n19242), .ZN(n19244) );
  NAND2_X1 U22212 ( .A1(n19248), .A2(n19244), .ZN(n19270) );
  INV_X1 U22213 ( .A(n19270), .ZN(n19260) );
  INV_X1 U22214 ( .A(n19281), .ZN(n19284) );
  AOI22_X1 U22215 ( .A1(n19260), .A2(n19547), .B1(n19284), .B2(n19546), .ZN(
        n19250) );
  NAND2_X1 U22216 ( .A1(n19548), .A2(n19245), .ZN(n19693) );
  AOI22_X1 U22217 ( .A1(n19281), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19246), 
        .B2(n19693), .ZN(n19247) );
  NAND3_X1 U22218 ( .A1(n19248), .A2(n19247), .A3(n19553), .ZN(n19272) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19272), .B1(
        n19267), .B2(n19555), .ZN(n19249) );
  OAI211_X1 U22220 ( .C1(n19558), .C2(n19307), .A(n19250), .B(n19249), .ZN(
        P2_U3104) );
  OAI22_X1 U22221 ( .A1(n19270), .A2(n19560), .B1(n19281), .B2(n19559), .ZN(
        n19251) );
  INV_X1 U22222 ( .A(n19251), .ZN(n19253) );
  AOI22_X1 U22223 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19272), .B1(
        n19267), .B2(n19503), .ZN(n19252) );
  OAI211_X1 U22224 ( .C1(n19426), .C2(n19307), .A(n19253), .B(n19252), .ZN(
        P2_U3105) );
  OAI22_X1 U22225 ( .A1(n19270), .A2(n19567), .B1(n19281), .B2(n19566), .ZN(
        n19254) );
  INV_X1 U22226 ( .A(n19254), .ZN(n19256) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19272), .B1(
        n19299), .B2(n19569), .ZN(n19255) );
  OAI211_X1 U22228 ( .C1(n19572), .C2(n19275), .A(n19256), .B(n19255), .ZN(
        P2_U3106) );
  OAI22_X1 U22229 ( .A1(n19270), .A2(n19574), .B1(n19281), .B2(n19573), .ZN(
        n19257) );
  INV_X1 U22230 ( .A(n19257), .ZN(n19259) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19272), .B1(
        n19267), .B2(n19576), .ZN(n19258) );
  OAI211_X1 U22232 ( .C1(n19579), .C2(n19307), .A(n19259), .B(n19258), .ZN(
        P2_U3107) );
  AOI22_X1 U22233 ( .A1(n19260), .A2(n19582), .B1(n19284), .B2(n19581), .ZN(
        n19262) );
  AOI22_X1 U22234 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19272), .B1(
        n19267), .B2(n19584), .ZN(n19261) );
  OAI211_X1 U22235 ( .C1(n19587), .C2(n19307), .A(n19262), .B(n19261), .ZN(
        P2_U3108) );
  OAI22_X1 U22236 ( .A1(n19270), .A2(n19589), .B1(n19281), .B2(n19588), .ZN(
        n19263) );
  INV_X1 U22237 ( .A(n19263), .ZN(n19265) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19272), .B1(
        n19267), .B2(n19591), .ZN(n19264) );
  OAI211_X1 U22239 ( .C1(n19594), .C2(n19307), .A(n19265), .B(n19264), .ZN(
        P2_U3109) );
  OAI22_X1 U22240 ( .A1(n19270), .A2(n19596), .B1(n19281), .B2(n19595), .ZN(
        n19266) );
  INV_X1 U22241 ( .A(n19266), .ZN(n19269) );
  AOI22_X1 U22242 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19272), .B1(
        n19267), .B2(n19435), .ZN(n19268) );
  OAI211_X1 U22243 ( .C1(n19438), .C2(n19307), .A(n19269), .B(n19268), .ZN(
        P2_U3110) );
  OAI22_X1 U22244 ( .A1(n19270), .A2(n19606), .B1(n19281), .B2(n19605), .ZN(
        n19271) );
  INV_X1 U22245 ( .A(n19271), .ZN(n19274) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19272), .B1(
        n19299), .B2(n19534), .ZN(n19273) );
  OAI211_X1 U22247 ( .C1(n19541), .C2(n19275), .A(n19274), .B(n19273), .ZN(
        P2_U3111) );
  NAND2_X1 U22248 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12211), .ZN(
        n19371) );
  NOR2_X1 U22249 ( .A1(n19278), .A2(n19371), .ZN(n19302) );
  AOI22_X1 U22250 ( .A1(n19555), .A2(n19299), .B1(n19546), .B2(n19302), .ZN(
        n19288) );
  NAND3_X1 U22251 ( .A1(n19324), .A2(n19688), .A3(n19307), .ZN(n19279) );
  NAND2_X1 U22252 ( .A1(n19279), .A2(n19690), .ZN(n19283) );
  OAI21_X1 U22253 ( .B1(n10473), .B2(n13409), .A(n19544), .ZN(n19280) );
  AOI21_X1 U22254 ( .B1(n19283), .B2(n19281), .A(n19280), .ZN(n19282) );
  OAI21_X1 U22255 ( .B1(n19302), .B2(n19282), .A(n19553), .ZN(n19304) );
  OAI21_X1 U22256 ( .B1(n19284), .B2(n19302), .A(n19283), .ZN(n19286) );
  OAI21_X1 U22257 ( .B1(n10473), .B2(n19302), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19285) );
  NAND2_X1 U22258 ( .A1(n19286), .A2(n19285), .ZN(n19303) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19304), .B1(
        n19547), .B2(n19303), .ZN(n19287) );
  OAI211_X1 U22260 ( .C1(n19558), .C2(n19324), .A(n19288), .B(n19287), .ZN(
        P2_U3112) );
  AOI22_X1 U22261 ( .A1(n19333), .A2(n19562), .B1(n19502), .B2(n19302), .ZN(
        n19290) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19504), .ZN(n19289) );
  OAI211_X1 U22263 ( .C1(n19565), .C2(n19307), .A(n19290), .B(n19289), .ZN(
        P2_U3113) );
  AOI22_X1 U22264 ( .A1(n19299), .A2(n19508), .B1(n19302), .B2(n19507), .ZN(
        n19292) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19509), .ZN(n19291) );
  OAI211_X1 U22266 ( .C1(n19463), .C2(n19324), .A(n19292), .B(n19291), .ZN(
        P2_U3114) );
  AOI22_X1 U22267 ( .A1(n19576), .A2(n19299), .B1(n19513), .B2(n19302), .ZN(
        n19294) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19515), .ZN(n19293) );
  OAI211_X1 U22269 ( .C1(n19579), .C2(n19324), .A(n19294), .B(n19293), .ZN(
        P2_U3115) );
  AOI22_X1 U22270 ( .A1(n19333), .A2(n19518), .B1(n19581), .B2(n19302), .ZN(
        n19296) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19582), .ZN(n19295) );
  OAI211_X1 U22272 ( .C1(n19396), .C2(n19307), .A(n19296), .B(n19295), .ZN(
        P2_U3116) );
  AOI22_X1 U22273 ( .A1(n19591), .A2(n19299), .B1(n19522), .B2(n19302), .ZN(
        n19298) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19525), .ZN(n19297) );
  OAI211_X1 U22275 ( .C1(n19594), .C2(n19324), .A(n19298), .B(n19297), .ZN(
        P2_U3117) );
  AOI22_X1 U22276 ( .A1(n19435), .A2(n19299), .B1(n19528), .B2(n19302), .ZN(
        n19301) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19529), .ZN(n19300) );
  OAI211_X1 U22278 ( .C1(n19438), .C2(n19324), .A(n19301), .B(n19300), .ZN(
        P2_U3118) );
  AOI22_X1 U22279 ( .A1(n19333), .A2(n19534), .B1(n19533), .B2(n19302), .ZN(
        n19306) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19536), .ZN(n19305) );
  OAI211_X1 U22281 ( .C1(n19541), .C2(n19307), .A(n19306), .B(n19305), .ZN(
        P2_U3119) );
  NOR3_X2 U22282 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19720), .A3(
        n19371), .ZN(n19342) );
  AOI22_X1 U22283 ( .A1(n19333), .A2(n19555), .B1(n19546), .B2(n19342), .ZN(
        n19319) );
  NAND2_X1 U22284 ( .A1(n19696), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19374) );
  OAI21_X1 U22285 ( .B1(n19374), .B2(n19309), .A(n19688), .ZN(n19317) );
  NOR2_X1 U22286 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19371), .ZN(
        n19313) );
  INV_X1 U22287 ( .A(n19342), .ZN(n19310) );
  OAI211_X1 U22288 ( .C1(n19311), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19692), 
        .B(n19310), .ZN(n19312) );
  OAI211_X1 U22289 ( .C1(n19317), .C2(n19313), .A(n19553), .B(n19312), .ZN(
        n19335) );
  INV_X1 U22290 ( .A(n19313), .ZN(n19316) );
  OAI21_X1 U22291 ( .B1(n19314), .B2(n19342), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19315) );
  OAI21_X1 U22292 ( .B1(n19317), .B2(n19316), .A(n19315), .ZN(n19334) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19335), .B1(
        n19547), .B2(n19334), .ZN(n19318) );
  OAI211_X1 U22294 ( .C1(n19558), .C2(n19338), .A(n19319), .B(n19318), .ZN(
        P2_U3120) );
  AOI22_X1 U22295 ( .A1(n19333), .A2(n19503), .B1(n19502), .B2(n19342), .ZN(
        n19321) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19335), .B1(
        n19504), .B2(n19334), .ZN(n19320) );
  OAI211_X1 U22297 ( .C1(n19426), .C2(n19338), .A(n19321), .B(n19320), .ZN(
        P2_U3121) );
  AOI22_X1 U22298 ( .A1(n19363), .A2(n19569), .B1(n19507), .B2(n19342), .ZN(
        n19323) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19335), .B1(
        n19509), .B2(n19334), .ZN(n19322) );
  OAI211_X1 U22300 ( .C1(n19572), .C2(n19324), .A(n19323), .B(n19322), .ZN(
        P2_U3122) );
  AOI22_X1 U22301 ( .A1(n19333), .A2(n19576), .B1(n19513), .B2(n19342), .ZN(
        n19326) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19335), .B1(
        n19515), .B2(n19334), .ZN(n19325) );
  OAI211_X1 U22303 ( .C1(n19579), .C2(n19338), .A(n19326), .B(n19325), .ZN(
        P2_U3123) );
  AOI22_X1 U22304 ( .A1(n19333), .A2(n19584), .B1(n19581), .B2(n19342), .ZN(
        n19328) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19335), .B1(
        n19582), .B2(n19334), .ZN(n19327) );
  OAI211_X1 U22306 ( .C1(n19587), .C2(n19338), .A(n19328), .B(n19327), .ZN(
        P2_U3124) );
  AOI22_X1 U22307 ( .A1(n19333), .A2(n19591), .B1(n19522), .B2(n19342), .ZN(
        n19330) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19335), .B1(
        n19525), .B2(n19334), .ZN(n19329) );
  OAI211_X1 U22309 ( .C1(n19594), .C2(n19338), .A(n19330), .B(n19329), .ZN(
        P2_U3125) );
  AOI22_X1 U22310 ( .A1(n19333), .A2(n19435), .B1(n19528), .B2(n19342), .ZN(
        n19332) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19335), .B1(
        n19529), .B2(n19334), .ZN(n19331) );
  OAI211_X1 U22312 ( .C1(n19438), .C2(n19338), .A(n19332), .B(n19331), .ZN(
        P2_U3126) );
  AOI22_X1 U22313 ( .A1(n19333), .A2(n19609), .B1(n19533), .B2(n19342), .ZN(
        n19337) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19335), .B1(
        n19536), .B2(n19334), .ZN(n19336) );
  OAI211_X1 U22315 ( .C1(n19615), .C2(n19338), .A(n19337), .B(n19336), .ZN(
        P2_U3127) );
  NOR3_X2 U22316 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10562), .A3(
        n19371), .ZN(n19361) );
  OAI21_X1 U22317 ( .B1(n19339), .B2(n19361), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19340) );
  OAI21_X1 U22318 ( .B1(n19371), .B2(n19341), .A(n19340), .ZN(n19362) );
  AOI22_X1 U22319 ( .A1(n19362), .A2(n19547), .B1(n19546), .B2(n19361), .ZN(
        n19348) );
  AOI221_X1 U22320 ( .B1(n19363), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19406), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19342), .ZN(n19344) );
  MUX2_X1 U22321 ( .A(n19344), .B(n19343), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19345) );
  NOR2_X1 U22322 ( .A1(n19345), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19346) );
  OAI21_X1 U22323 ( .B1(n19346), .B2(n19361), .A(n19553), .ZN(n19364) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19555), .ZN(n19347) );
  OAI211_X1 U22325 ( .C1(n19558), .C2(n19395), .A(n19348), .B(n19347), .ZN(
        P2_U3128) );
  AOI22_X1 U22326 ( .A1(n19362), .A2(n19504), .B1(n19502), .B2(n19361), .ZN(
        n19350) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19503), .ZN(n19349) );
  OAI211_X1 U22328 ( .C1(n19426), .C2(n19395), .A(n19350), .B(n19349), .ZN(
        P2_U3129) );
  AOI22_X1 U22329 ( .A1(n19362), .A2(n19509), .B1(n19507), .B2(n19361), .ZN(
        n19352) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19508), .ZN(n19351) );
  OAI211_X1 U22331 ( .C1(n19463), .C2(n19395), .A(n19352), .B(n19351), .ZN(
        P2_U3130) );
  AOI22_X1 U22332 ( .A1(n19362), .A2(n19515), .B1(n19513), .B2(n19361), .ZN(
        n19354) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19576), .ZN(n19353) );
  OAI211_X1 U22334 ( .C1(n19579), .C2(n19395), .A(n19354), .B(n19353), .ZN(
        P2_U3131) );
  AOI22_X1 U22335 ( .A1(n19362), .A2(n19582), .B1(n19581), .B2(n19361), .ZN(
        n19356) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19584), .ZN(n19355) );
  OAI211_X1 U22337 ( .C1(n19587), .C2(n19395), .A(n19356), .B(n19355), .ZN(
        P2_U3132) );
  AOI22_X1 U22338 ( .A1(n19362), .A2(n19525), .B1(n19522), .B2(n19361), .ZN(
        n19358) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19591), .ZN(n19357) );
  OAI211_X1 U22340 ( .C1(n19594), .C2(n19395), .A(n19358), .B(n19357), .ZN(
        P2_U3133) );
  AOI22_X1 U22341 ( .A1(n19362), .A2(n19529), .B1(n19528), .B2(n19361), .ZN(
        n19360) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19435), .ZN(n19359) );
  OAI211_X1 U22343 ( .C1(n19438), .C2(n19395), .A(n19360), .B(n19359), .ZN(
        P2_U3134) );
  AOI22_X1 U22344 ( .A1(n19362), .A2(n19536), .B1(n19533), .B2(n19361), .ZN(
        n19366) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19364), .B1(
        n19363), .B2(n19609), .ZN(n19365) );
  OAI211_X1 U22346 ( .C1(n19615), .C2(n19395), .A(n19366), .B(n19365), .ZN(
        P2_U3135) );
  INV_X1 U22347 ( .A(n19375), .ZN(n19689) );
  NOR2_X2 U22348 ( .A1(n19446), .A2(n19689), .ZN(n19441) );
  INV_X1 U22349 ( .A(n19441), .ZN(n19410) );
  INV_X1 U22350 ( .A(n19371), .ZN(n19367) );
  AND2_X1 U22351 ( .A1(n19368), .A2(n19367), .ZN(n19391) );
  INV_X1 U22352 ( .A(n19391), .ZN(n19403) );
  NAND2_X1 U22353 ( .A1(n19403), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19369) );
  NOR2_X1 U22354 ( .A1(n19370), .A2(n19369), .ZN(n19376) );
  OR2_X1 U22355 ( .A1(n10562), .A2(n19371), .ZN(n19377) );
  INV_X1 U22356 ( .A(n19377), .ZN(n19372) );
  AOI21_X1 U22357 ( .B1(n19544), .B2(n19372), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19373) );
  INV_X1 U22358 ( .A(n19404), .ZN(n19392) );
  AOI22_X1 U22359 ( .A1(n19392), .A2(n19547), .B1(n19546), .B2(n19391), .ZN(
        n19381) );
  INV_X1 U22360 ( .A(n19374), .ZN(n19549) );
  NAND2_X1 U22361 ( .A1(n19549), .A2(n19375), .ZN(n19378) );
  AOI21_X1 U22362 ( .B1(n19378), .B2(n19377), .A(n19376), .ZN(n19379) );
  OAI211_X1 U22363 ( .C1(n19391), .C2(n19544), .A(n19379), .B(n19553), .ZN(
        n19407) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19407), .B1(
        n19406), .B2(n19555), .ZN(n19380) );
  OAI211_X1 U22365 ( .C1(n19558), .C2(n19410), .A(n19381), .B(n19380), .ZN(
        P2_U3136) );
  OAI22_X1 U22366 ( .A1(n19404), .A2(n19560), .B1(n19559), .B2(n19403), .ZN(
        n19382) );
  INV_X1 U22367 ( .A(n19382), .ZN(n19384) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19407), .B1(
        n19441), .B2(n19562), .ZN(n19383) );
  OAI211_X1 U22369 ( .C1(n19565), .C2(n19395), .A(n19384), .B(n19383), .ZN(
        P2_U3137) );
  OAI22_X1 U22370 ( .A1(n19404), .A2(n19567), .B1(n19566), .B2(n19403), .ZN(
        n19385) );
  INV_X1 U22371 ( .A(n19385), .ZN(n19387) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19407), .B1(
        n19441), .B2(n19569), .ZN(n19386) );
  OAI211_X1 U22373 ( .C1(n19572), .C2(n19395), .A(n19387), .B(n19386), .ZN(
        P2_U3138) );
  OAI22_X1 U22374 ( .A1(n19404), .A2(n19574), .B1(n19573), .B2(n19403), .ZN(
        n19388) );
  INV_X1 U22375 ( .A(n19388), .ZN(n19390) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19407), .B1(
        n19406), .B2(n19576), .ZN(n19389) );
  OAI211_X1 U22377 ( .C1(n19579), .C2(n19410), .A(n19390), .B(n19389), .ZN(
        P2_U3139) );
  AOI22_X1 U22378 ( .A1(n19392), .A2(n19582), .B1(n19581), .B2(n19391), .ZN(
        n19394) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19407), .B1(
        n19441), .B2(n19518), .ZN(n19393) );
  OAI211_X1 U22380 ( .C1(n19396), .C2(n19395), .A(n19394), .B(n19393), .ZN(
        P2_U3140) );
  OAI22_X1 U22381 ( .A1(n19404), .A2(n19589), .B1(n19588), .B2(n19403), .ZN(
        n19397) );
  INV_X1 U22382 ( .A(n19397), .ZN(n19399) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19407), .B1(
        n19406), .B2(n19591), .ZN(n19398) );
  OAI211_X1 U22384 ( .C1(n19594), .C2(n19410), .A(n19399), .B(n19398), .ZN(
        P2_U3141) );
  OAI22_X1 U22385 ( .A1(n19404), .A2(n19596), .B1(n19595), .B2(n19403), .ZN(
        n19400) );
  INV_X1 U22386 ( .A(n19400), .ZN(n19402) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19407), .B1(
        n19406), .B2(n19435), .ZN(n19401) );
  OAI211_X1 U22388 ( .C1(n19438), .C2(n19410), .A(n19402), .B(n19401), .ZN(
        P2_U3142) );
  OAI22_X1 U22389 ( .A1(n19404), .A2(n19606), .B1(n19605), .B2(n19403), .ZN(
        n19405) );
  INV_X1 U22390 ( .A(n19405), .ZN(n19409) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19407), .B1(
        n19406), .B2(n19609), .ZN(n19408) );
  OAI211_X1 U22392 ( .C1(n19615), .C2(n19410), .A(n19409), .B(n19408), .ZN(
        P2_U3143) );
  INV_X1 U22393 ( .A(n19412), .ZN(n19416) );
  INV_X1 U22394 ( .A(n19413), .ZN(n19419) );
  NAND3_X1 U22395 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n10562), .ZN(n19452) );
  NOR2_X1 U22396 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19452), .ZN(
        n19439) );
  OAI21_X1 U22397 ( .B1(n19414), .B2(n19439), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19415) );
  OAI21_X1 U22398 ( .B1(n19416), .B2(n19419), .A(n19415), .ZN(n19440) );
  AOI22_X1 U22399 ( .A1(n19440), .A2(n19547), .B1(n19546), .B2(n19439), .ZN(
        n19423) );
  AOI21_X1 U22400 ( .B1(n19417), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19421) );
  OAI21_X1 U22401 ( .B1(n19471), .B2(n19441), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19418) );
  OAI21_X1 U22402 ( .B1(n19419), .B2(n13264), .A(n19418), .ZN(n19420) );
  OAI211_X1 U22403 ( .C1(n19439), .C2(n19421), .A(n19420), .B(n19553), .ZN(
        n19442) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19555), .ZN(n19422) );
  OAI211_X1 U22405 ( .C1(n19558), .C2(n19483), .A(n19423), .B(n19422), .ZN(
        P2_U3144) );
  AOI22_X1 U22406 ( .A1(n19440), .A2(n19504), .B1(n19502), .B2(n19439), .ZN(
        n19425) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19503), .ZN(n19424) );
  OAI211_X1 U22408 ( .C1(n19426), .C2(n19483), .A(n19425), .B(n19424), .ZN(
        P2_U3145) );
  AOI22_X1 U22409 ( .A1(n19440), .A2(n19509), .B1(n19507), .B2(n19439), .ZN(
        n19428) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19508), .ZN(n19427) );
  OAI211_X1 U22411 ( .C1(n19463), .C2(n19483), .A(n19428), .B(n19427), .ZN(
        P2_U3146) );
  AOI22_X1 U22412 ( .A1(n19440), .A2(n19515), .B1(n19513), .B2(n19439), .ZN(
        n19430) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19576), .ZN(n19429) );
  OAI211_X1 U22414 ( .C1(n19579), .C2(n19483), .A(n19430), .B(n19429), .ZN(
        P2_U3147) );
  AOI22_X1 U22415 ( .A1(n19440), .A2(n19582), .B1(n19581), .B2(n19439), .ZN(
        n19432) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19584), .ZN(n19431) );
  OAI211_X1 U22417 ( .C1(n19587), .C2(n19483), .A(n19432), .B(n19431), .ZN(
        P2_U3148) );
  AOI22_X1 U22418 ( .A1(n19440), .A2(n19525), .B1(n19522), .B2(n19439), .ZN(
        n19434) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19591), .ZN(n19433) );
  OAI211_X1 U22420 ( .C1(n19594), .C2(n19483), .A(n19434), .B(n19433), .ZN(
        P2_U3149) );
  AOI22_X1 U22421 ( .A1(n19440), .A2(n19529), .B1(n19528), .B2(n19439), .ZN(
        n19437) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19435), .ZN(n19436) );
  OAI211_X1 U22423 ( .C1(n19438), .C2(n19483), .A(n19437), .B(n19436), .ZN(
        P2_U3150) );
  AOI22_X1 U22424 ( .A1(n19440), .A2(n19536), .B1(n19533), .B2(n19439), .ZN(
        n19444) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19442), .B1(
        n19441), .B2(n19609), .ZN(n19443) );
  OAI211_X1 U22426 ( .C1(n19615), .C2(n19483), .A(n19444), .B(n19443), .ZN(
        P2_U3151) );
  INV_X1 U22427 ( .A(n19523), .ZN(n19540) );
  NOR2_X1 U22428 ( .A1(n19720), .A2(n19452), .ZN(n19487) );
  INV_X1 U22429 ( .A(n19487), .ZN(n19477) );
  NAND2_X1 U22430 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19477), .ZN(n19447) );
  NOR2_X1 U22431 ( .A1(n10354), .A2(n19447), .ZN(n19451) );
  INV_X1 U22432 ( .A(n19452), .ZN(n19448) );
  AOI21_X1 U22433 ( .B1(n19544), .B2(n19448), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19449) );
  OR2_X1 U22434 ( .A1(n19451), .A2(n19449), .ZN(n19478) );
  INV_X1 U22435 ( .A(n19478), .ZN(n19467) );
  AOI22_X1 U22436 ( .A1(n19467), .A2(n19547), .B1(n19546), .B2(n19487), .ZN(
        n19456) );
  NAND2_X1 U22437 ( .A1(n19549), .A2(n19450), .ZN(n19453) );
  AOI21_X1 U22438 ( .B1(n19453), .B2(n19452), .A(n19451), .ZN(n19454) );
  OAI211_X1 U22439 ( .C1(n19487), .C2(n19544), .A(n19454), .B(n19553), .ZN(
        n19480) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19480), .B1(
        n19471), .B2(n19555), .ZN(n19455) );
  OAI211_X1 U22441 ( .C1(n19558), .C2(n19540), .A(n19456), .B(n19455), .ZN(
        P2_U3152) );
  OAI22_X1 U22442 ( .A1(n19478), .A2(n19560), .B1(n19559), .B2(n19477), .ZN(
        n19457) );
  INV_X1 U22443 ( .A(n19457), .ZN(n19459) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19480), .B1(
        n19523), .B2(n19562), .ZN(n19458) );
  OAI211_X1 U22445 ( .C1(n19565), .C2(n19483), .A(n19459), .B(n19458), .ZN(
        P2_U3153) );
  OAI22_X1 U22446 ( .A1(n19478), .A2(n19567), .B1(n19566), .B2(n19477), .ZN(
        n19460) );
  INV_X1 U22447 ( .A(n19460), .ZN(n19462) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19480), .B1(
        n19471), .B2(n19508), .ZN(n19461) );
  OAI211_X1 U22449 ( .C1(n19463), .C2(n19540), .A(n19462), .B(n19461), .ZN(
        P2_U3154) );
  OAI22_X1 U22450 ( .A1(n19478), .A2(n19574), .B1(n19573), .B2(n19477), .ZN(
        n19464) );
  INV_X1 U22451 ( .A(n19464), .ZN(n19466) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19480), .B1(
        n19471), .B2(n19576), .ZN(n19465) );
  OAI211_X1 U22453 ( .C1(n19579), .C2(n19540), .A(n19466), .B(n19465), .ZN(
        P2_U3155) );
  AOI22_X1 U22454 ( .A1(n19467), .A2(n19582), .B1(n19581), .B2(n19487), .ZN(
        n19469) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19480), .B1(
        n19471), .B2(n19584), .ZN(n19468) );
  OAI211_X1 U22456 ( .C1(n19587), .C2(n19540), .A(n19469), .B(n19468), .ZN(
        P2_U3156) );
  OAI22_X1 U22457 ( .A1(n19478), .A2(n19589), .B1(n19588), .B2(n19477), .ZN(
        n19470) );
  INV_X1 U22458 ( .A(n19470), .ZN(n19473) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19480), .B1(
        n19471), .B2(n19591), .ZN(n19472) );
  OAI211_X1 U22460 ( .C1(n19594), .C2(n19540), .A(n19473), .B(n19472), .ZN(
        P2_U3157) );
  OAI22_X1 U22461 ( .A1(n19478), .A2(n19596), .B1(n19595), .B2(n19477), .ZN(
        n19474) );
  INV_X1 U22462 ( .A(n19474), .ZN(n19476) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19480), .B1(
        n19523), .B2(n19598), .ZN(n19475) );
  OAI211_X1 U22464 ( .C1(n19603), .C2(n19483), .A(n19476), .B(n19475), .ZN(
        P2_U3158) );
  OAI22_X1 U22465 ( .A1(n19478), .A2(n19606), .B1(n19605), .B2(n19477), .ZN(
        n19479) );
  INV_X1 U22466 ( .A(n19479), .ZN(n19482) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19480), .B1(
        n19523), .B2(n19534), .ZN(n19481) );
  OAI211_X1 U22468 ( .C1(n19541), .C2(n19483), .A(n19482), .B(n19481), .ZN(
        P2_U3159) );
  OR2_X1 U22469 ( .A1(n19523), .A2(n19692), .ZN(n19486) );
  OAI21_X1 U22470 ( .B1(n19486), .B2(n19610), .A(n19690), .ZN(n19494) );
  NAND3_X1 U22471 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19551) );
  NOR2_X1 U22472 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19551), .ZN(
        n19532) );
  NOR2_X1 U22473 ( .A1(n19532), .A2(n19487), .ZN(n19497) );
  NAND2_X1 U22474 ( .A1(n19494), .A2(n19497), .ZN(n19492) );
  INV_X1 U22475 ( .A(n19532), .ZN(n19488) );
  OAI211_X1 U22476 ( .C1(n19489), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19692), 
        .B(n19488), .ZN(n19490) );
  AND2_X1 U22477 ( .A1(n19490), .A2(n19553), .ZN(n19491) );
  AOI22_X1 U22478 ( .A1(n19493), .A2(n19610), .B1(n19546), .B2(n19532), .ZN(
        n19500) );
  INV_X1 U22479 ( .A(n19494), .ZN(n19498) );
  OAI21_X1 U22480 ( .B1(n19495), .B2(n19532), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19496) );
  AOI22_X1 U22481 ( .A1(n19547), .A2(n19535), .B1(n19523), .B2(n19555), .ZN(
        n19499) );
  OAI211_X1 U22482 ( .C1(n19524), .C2(n19501), .A(n19500), .B(n19499), .ZN(
        P2_U3160) );
  AOI22_X1 U22483 ( .A1(n19610), .A2(n19562), .B1(n19502), .B2(n19532), .ZN(
        n19506) );
  AOI22_X1 U22484 ( .A1(n19504), .A2(n19535), .B1(n19523), .B2(n19503), .ZN(
        n19505) );
  OAI211_X1 U22485 ( .C1(n19524), .C2(n10363), .A(n19506), .B(n19505), .ZN(
        P2_U3161) );
  INV_X1 U22486 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19512) );
  AOI22_X1 U22487 ( .A1(n19610), .A2(n19569), .B1(n19507), .B2(n19532), .ZN(
        n19511) );
  AOI22_X1 U22488 ( .A1(n19509), .A2(n19535), .B1(n19523), .B2(n19508), .ZN(
        n19510) );
  OAI211_X1 U22489 ( .C1(n19524), .C2(n19512), .A(n19511), .B(n19510), .ZN(
        P2_U3162) );
  AOI22_X1 U22490 ( .A1(n19514), .A2(n19610), .B1(n19513), .B2(n19532), .ZN(
        n19517) );
  AOI22_X1 U22491 ( .A1(n19515), .A2(n19535), .B1(n19523), .B2(n19576), .ZN(
        n19516) );
  OAI211_X1 U22492 ( .C1(n19524), .C2(n10316), .A(n19517), .B(n19516), .ZN(
        P2_U3163) );
  INV_X1 U22493 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19521) );
  AOI22_X1 U22494 ( .A1(n19523), .A2(n19584), .B1(n19581), .B2(n19532), .ZN(
        n19520) );
  AOI22_X1 U22495 ( .A1(n19582), .A2(n19535), .B1(n19610), .B2(n19518), .ZN(
        n19519) );
  OAI211_X1 U22496 ( .C1(n19524), .C2(n19521), .A(n19520), .B(n19519), .ZN(
        P2_U3164) );
  INV_X1 U22497 ( .A(n19610), .ZN(n19602) );
  AOI22_X1 U22498 ( .A1(n19591), .A2(n19523), .B1(n19522), .B2(n19532), .ZN(
        n19527) );
  INV_X1 U22499 ( .A(n19524), .ZN(n19537) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19537), .B1(
        n19525), .B2(n19535), .ZN(n19526) );
  OAI211_X1 U22501 ( .C1(n19594), .C2(n19602), .A(n19527), .B(n19526), .ZN(
        P2_U3165) );
  AOI22_X1 U22502 ( .A1(n19598), .A2(n19610), .B1(n19528), .B2(n19532), .ZN(
        n19531) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19537), .B1(
        n19529), .B2(n19535), .ZN(n19530) );
  OAI211_X1 U22504 ( .C1(n19603), .C2(n19540), .A(n19531), .B(n19530), .ZN(
        P2_U3166) );
  AOI22_X1 U22505 ( .A1(n19534), .A2(n19610), .B1(n19533), .B2(n19532), .ZN(
        n19539) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19535), .ZN(n19538) );
  OAI211_X1 U22507 ( .C1(n19541), .C2(n19540), .A(n19539), .B(n19538), .ZN(
        P2_U3167) );
  INV_X1 U22508 ( .A(n19599), .ZN(n19614) );
  OR2_X1 U22509 ( .A1(n19580), .A2(n13409), .ZN(n19542) );
  NOR2_X1 U22510 ( .A1(n10353), .A2(n19542), .ZN(n19550) );
  INV_X1 U22511 ( .A(n19551), .ZN(n19543) );
  AOI21_X1 U22512 ( .B1(n19544), .B2(n19543), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19545) );
  INV_X1 U22513 ( .A(n19607), .ZN(n19583) );
  AOI22_X1 U22514 ( .A1(n19583), .A2(n19547), .B1(n19546), .B2(n19580), .ZN(
        n19557) );
  NAND2_X1 U22515 ( .A1(n19549), .A2(n19548), .ZN(n19552) );
  AOI21_X1 U22516 ( .B1(n19552), .B2(n19551), .A(n19550), .ZN(n19554) );
  OAI211_X1 U22517 ( .C1(n19580), .C2(n19544), .A(n19554), .B(n19553), .ZN(
        n19611) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19555), .ZN(n19556) );
  OAI211_X1 U22519 ( .C1(n19558), .C2(n19614), .A(n19557), .B(n19556), .ZN(
        P2_U3168) );
  INV_X1 U22520 ( .A(n19580), .ZN(n19604) );
  OAI22_X1 U22521 ( .A1(n19607), .A2(n19560), .B1(n19559), .B2(n19604), .ZN(
        n19561) );
  INV_X1 U22522 ( .A(n19561), .ZN(n19564) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19611), .B1(
        n19599), .B2(n19562), .ZN(n19563) );
  OAI211_X1 U22524 ( .C1(n19565), .C2(n19602), .A(n19564), .B(n19563), .ZN(
        P2_U3169) );
  OAI22_X1 U22525 ( .A1(n19607), .A2(n19567), .B1(n19566), .B2(n19604), .ZN(
        n19568) );
  INV_X1 U22526 ( .A(n19568), .ZN(n19571) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19611), .B1(
        n19599), .B2(n19569), .ZN(n19570) );
  OAI211_X1 U22528 ( .C1(n19572), .C2(n19602), .A(n19571), .B(n19570), .ZN(
        P2_U3170) );
  OAI22_X1 U22529 ( .A1(n19607), .A2(n19574), .B1(n19573), .B2(n19604), .ZN(
        n19575) );
  INV_X1 U22530 ( .A(n19575), .ZN(n19578) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19576), .ZN(n19577) );
  OAI211_X1 U22532 ( .C1(n19579), .C2(n19614), .A(n19578), .B(n19577), .ZN(
        P2_U3171) );
  AOI22_X1 U22533 ( .A1(n19583), .A2(n19582), .B1(n19581), .B2(n19580), .ZN(
        n19586) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19584), .ZN(n19585) );
  OAI211_X1 U22535 ( .C1(n19587), .C2(n19614), .A(n19586), .B(n19585), .ZN(
        P2_U3172) );
  OAI22_X1 U22536 ( .A1(n19607), .A2(n19589), .B1(n19588), .B2(n19604), .ZN(
        n19590) );
  INV_X1 U22537 ( .A(n19590), .ZN(n19593) );
  AOI22_X1 U22538 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19591), .ZN(n19592) );
  OAI211_X1 U22539 ( .C1(n19594), .C2(n19614), .A(n19593), .B(n19592), .ZN(
        P2_U3173) );
  OAI22_X1 U22540 ( .A1(n19607), .A2(n19596), .B1(n19595), .B2(n19604), .ZN(
        n19597) );
  INV_X1 U22541 ( .A(n19597), .ZN(n19601) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19611), .B1(
        n19599), .B2(n19598), .ZN(n19600) );
  OAI211_X1 U22543 ( .C1(n19603), .C2(n19602), .A(n19601), .B(n19600), .ZN(
        P2_U3174) );
  OAI22_X1 U22544 ( .A1(n19607), .A2(n19606), .B1(n19605), .B2(n19604), .ZN(
        n19608) );
  INV_X1 U22545 ( .A(n19608), .ZN(n19613) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19611), .B1(
        n19610), .B2(n19609), .ZN(n19612) );
  OAI211_X1 U22547 ( .C1(n19615), .C2(n19614), .A(n19613), .B(n19612), .ZN(
        P2_U3175) );
  AND2_X1 U22548 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19616), .ZN(
        P2_U3179) );
  AND2_X1 U22549 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19616), .ZN(
        P2_U3180) );
  AND2_X1 U22550 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19616), .ZN(
        P2_U3181) );
  AND2_X1 U22551 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19616), .ZN(
        P2_U3182) );
  AND2_X1 U22552 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19616), .ZN(
        P2_U3183) );
  AND2_X1 U22553 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19616), .ZN(
        P2_U3184) );
  AND2_X1 U22554 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19616), .ZN(
        P2_U3185) );
  AND2_X1 U22555 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19616), .ZN(
        P2_U3186) );
  AND2_X1 U22556 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19616), .ZN(
        P2_U3187) );
  AND2_X1 U22557 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19616), .ZN(
        P2_U3188) );
  AND2_X1 U22558 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19616), .ZN(
        P2_U3189) );
  AND2_X1 U22559 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19616), .ZN(
        P2_U3190) );
  AND2_X1 U22560 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19616), .ZN(
        P2_U3191) );
  AND2_X1 U22561 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19616), .ZN(
        P2_U3192) );
  AND2_X1 U22562 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19616), .ZN(
        P2_U3193) );
  AND2_X1 U22563 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19616), .ZN(
        P2_U3194) );
  AND2_X1 U22564 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19616), .ZN(
        P2_U3195) );
  AND2_X1 U22565 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19616), .ZN(
        P2_U3196) );
  AND2_X1 U22566 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19616), .ZN(
        P2_U3197) );
  AND2_X1 U22567 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19616), .ZN(
        P2_U3198) );
  AND2_X1 U22568 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19616), .ZN(
        P2_U3199) );
  AND2_X1 U22569 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19616), .ZN(
        P2_U3200) );
  AND2_X1 U22570 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19616), .ZN(P2_U3201) );
  AND2_X1 U22571 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19616), .ZN(P2_U3202) );
  AND2_X1 U22572 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19616), .ZN(P2_U3203) );
  AND2_X1 U22573 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19616), .ZN(P2_U3204) );
  AND2_X1 U22574 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19616), .ZN(P2_U3205) );
  AND2_X1 U22575 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19616), .ZN(P2_U3206) );
  AND2_X1 U22576 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19616), .ZN(P2_U3207) );
  AND2_X1 U22577 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19616), .ZN(P2_U3208) );
  INV_X1 U22578 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19631) );
  NOR2_X1 U22579 ( .A1(n19617), .A2(n19631), .ZN(n19628) );
  OR3_X1 U22580 ( .A1(n19628), .A2(n19629), .A3(n19621), .ZN(n19619) );
  AOI211_X1 U22581 ( .C1(n19627), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19630), .B(n19672), .ZN(n19618) );
  NOR3_X1 U22582 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20540), .ZN(n19636) );
  AOI211_X1 U22583 ( .C1(n19639), .C2(n19619), .A(n19618), .B(n19636), .ZN(
        n19620) );
  INV_X1 U22584 ( .A(n19620), .ZN(P2_U3209) );
  AOI21_X1 U22585 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19627), .A(n19639), 
        .ZN(n19632) );
  INV_X1 U22586 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19621) );
  NOR3_X1 U22587 ( .A1(n19632), .A2(n19629), .A3(n19621), .ZN(n19622) );
  NOR2_X1 U22588 ( .A1(n19622), .A2(n19628), .ZN(n19625) );
  INV_X1 U22589 ( .A(n19623), .ZN(n19624) );
  OAI211_X1 U22590 ( .C1(n19627), .C2(n19626), .A(n19625), .B(n19624), .ZN(
        P2_U3210) );
  AOI22_X1 U22591 ( .A1(n19630), .A2(n19629), .B1(n19628), .B2(n20540), .ZN(
        n19638) );
  OAI21_X1 U22592 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19637) );
  NOR2_X1 U22593 ( .A1(n19631), .A2(n19639), .ZN(n19634) );
  AOI21_X1 U22594 ( .B1(n19634), .B2(n19633), .A(n19632), .ZN(n19635) );
  OAI22_X1 U22595 ( .A1(n19638), .A2(n19637), .B1(n19636), .B2(n19635), .ZN(
        P2_U3211) );
  NAND2_X1 U22596 ( .A1(n19672), .A2(n19639), .ZN(n19681) );
  CLKBUF_X1 U22597 ( .A(n19681), .Z(n19678) );
  NAND2_X2 U22598 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19672), .ZN(n19679) );
  OAI222_X1 U22599 ( .A1(n19678), .A2(n10276), .B1(n19641), .B2(n19672), .C1(
        n19640), .C2(n19679), .ZN(P2_U3212) );
  OAI222_X1 U22600 ( .A1(n19679), .A2(n10276), .B1(n19642), .B2(n19672), .C1(
        n10292), .C2(n19678), .ZN(P2_U3213) );
  OAI222_X1 U22601 ( .A1(n19679), .A2(n10292), .B1(n19643), .B2(n19672), .C1(
        n10613), .C2(n19678), .ZN(P2_U3214) );
  OAI222_X1 U22602 ( .A1(n19681), .A2(n13626), .B1(n19644), .B2(n19672), .C1(
        n10613), .C2(n19679), .ZN(P2_U3215) );
  OAI222_X1 U22603 ( .A1(n19681), .A2(n10618), .B1(n19645), .B2(n19672), .C1(
        n13626), .C2(n19679), .ZN(P2_U3216) );
  OAI222_X1 U22604 ( .A1(n19681), .A2(n10622), .B1(n19646), .B2(n19672), .C1(
        n10618), .C2(n19679), .ZN(P2_U3217) );
  OAI222_X1 U22605 ( .A1(n19681), .A2(n11092), .B1(n19647), .B2(n19672), .C1(
        n10622), .C2(n19679), .ZN(P2_U3218) );
  OAI222_X1 U22606 ( .A1(n19681), .A2(n15320), .B1(n19648), .B2(n19672), .C1(
        n11092), .C2(n19679), .ZN(P2_U3219) );
  OAI222_X1 U22607 ( .A1(n19678), .A2(n10631), .B1(n19649), .B2(n19672), .C1(
        n15320), .C2(n19679), .ZN(P2_U3220) );
  OAI222_X1 U22608 ( .A1(n19678), .A2(n10635), .B1(n19650), .B2(n19672), .C1(
        n10631), .C2(n19679), .ZN(P2_U3221) );
  OAI222_X1 U22609 ( .A1(n19678), .A2(n11151), .B1(n19651), .B2(n19672), .C1(
        n10635), .C2(n19679), .ZN(P2_U3222) );
  OAI222_X1 U22610 ( .A1(n19678), .A2(n10602), .B1(n20705), .B2(n19672), .C1(
        n11151), .C2(n19679), .ZN(P2_U3223) );
  OAI222_X1 U22611 ( .A1(n19678), .A2(n11025), .B1(n19652), .B2(n19672), .C1(
        n10602), .C2(n19679), .ZN(P2_U3224) );
  OAI222_X1 U22612 ( .A1(n19678), .A2(n15042), .B1(n19653), .B2(n19672), .C1(
        n11025), .C2(n19679), .ZN(P2_U3225) );
  INV_X1 U22613 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20674) );
  OAI222_X1 U22614 ( .A1(n19681), .A2(n20674), .B1(n19654), .B2(n19672), .C1(
        n15042), .C2(n19679), .ZN(P2_U3226) );
  OAI222_X1 U22615 ( .A1(n19681), .A2(n19656), .B1(n19655), .B2(n19672), .C1(
        n20674), .C2(n19679), .ZN(P2_U3227) );
  OAI222_X1 U22616 ( .A1(n19681), .A2(n19658), .B1(n19657), .B2(n19672), .C1(
        n19656), .C2(n19679), .ZN(P2_U3228) );
  OAI222_X1 U22617 ( .A1(n19681), .A2(n19660), .B1(n19659), .B2(n19672), .C1(
        n19658), .C2(n19679), .ZN(P2_U3229) );
  OAI222_X1 U22618 ( .A1(n19681), .A2(n19661), .B1(n20704), .B2(n19672), .C1(
        n19660), .C2(n19679), .ZN(P2_U3230) );
  OAI222_X1 U22619 ( .A1(n19681), .A2(n20723), .B1(n19662), .B2(n19672), .C1(
        n19661), .C2(n19679), .ZN(P2_U3231) );
  OAI222_X1 U22620 ( .A1(n19678), .A2(n14942), .B1(n19663), .B2(n19672), .C1(
        n20723), .C2(n19679), .ZN(P2_U3232) );
  OAI222_X1 U22621 ( .A1(n19678), .A2(n19665), .B1(n19664), .B2(n19672), .C1(
        n14942), .C2(n19679), .ZN(P2_U3233) );
  OAI222_X1 U22622 ( .A1(n19678), .A2(n19667), .B1(n19666), .B2(n19672), .C1(
        n19665), .C2(n19679), .ZN(P2_U3234) );
  OAI222_X1 U22623 ( .A1(n19678), .A2(n19669), .B1(n19668), .B2(n19672), .C1(
        n19667), .C2(n19679), .ZN(P2_U3235) );
  OAI222_X1 U22624 ( .A1(n19678), .A2(n14898), .B1(n19670), .B2(n19672), .C1(
        n19669), .C2(n19679), .ZN(P2_U3236) );
  OAI222_X1 U22625 ( .A1(n19678), .A2(n19674), .B1(n19671), .B2(n19672), .C1(
        n14898), .C2(n19679), .ZN(P2_U3237) );
  INV_X1 U22626 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19675) );
  OAI222_X1 U22627 ( .A1(n19679), .A2(n19674), .B1(n19673), .B2(n19672), .C1(
        n19675), .C2(n19678), .ZN(P2_U3238) );
  OAI222_X1 U22628 ( .A1(n19678), .A2(n20752), .B1(n19676), .B2(n19672), .C1(
        n19675), .C2(n19679), .ZN(P2_U3239) );
  OAI222_X1 U22629 ( .A1(n19678), .A2(n11209), .B1(n19677), .B2(n19672), .C1(
        n20752), .C2(n19679), .ZN(P2_U3240) );
  OAI222_X1 U22630 ( .A1(n19681), .A2(n10714), .B1(n19680), .B2(n19672), .C1(
        n11209), .C2(n19679), .ZN(P2_U3241) );
  INV_X1 U22631 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19682) );
  AOI22_X1 U22632 ( .A1(n19672), .A2(n20718), .B1(n19682), .B2(n19735), .ZN(
        P2_U3585) );
  MUX2_X1 U22633 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19672), .Z(P2_U3586) );
  MUX2_X1 U22634 ( .A(P2_BE_N_REG_1__SCAN_IN), .B(P2_BYTEENABLE_REG_1__SCAN_IN), .S(n19672), .Z(P2_U3587) );
  INV_X1 U22635 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20662) );
  AOI22_X1 U22636 ( .A1(n19672), .A2(n19683), .B1(n20662), .B2(n19735), .ZN(
        P2_U3588) );
  OAI21_X1 U22637 ( .B1(n19687), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19685), 
        .ZN(n19684) );
  INV_X1 U22638 ( .A(n19684), .ZN(P2_U3591) );
  OAI21_X1 U22639 ( .B1(n19687), .B2(n19686), .A(n19685), .ZN(P2_U3592) );
  NAND2_X1 U22640 ( .A1(n19688), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19708) );
  NOR2_X1 U22641 ( .A1(n19689), .A2(n19708), .ZN(n19702) );
  OAI211_X1 U22642 ( .C1(n19709), .C2(n19692), .A(n19691), .B(n19690), .ZN(
        n19700) );
  OR2_X1 U22643 ( .A1(n19702), .A2(n19700), .ZN(n19697) );
  OAI22_X1 U22644 ( .A1(n19694), .A2(n19544), .B1(n19693), .B2(n19692), .ZN(
        n19695) );
  AOI21_X1 U22645 ( .B1(n19697), .B2(n19696), .A(n19695), .ZN(n19698) );
  AOI22_X1 U22646 ( .A1(n19721), .A2(n13264), .B1(n19698), .B2(n19718), .ZN(
        P2_U3602) );
  AOI22_X1 U22647 ( .A1(n19701), .A2(n19700), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19699), .ZN(n19704) );
  NOR2_X1 U22648 ( .A1(n19721), .A2(n19702), .ZN(n19703) );
  AOI22_X1 U22649 ( .A1(n12211), .A2(n19721), .B1(n19704), .B2(n19703), .ZN(
        P2_U3603) );
  INV_X1 U22650 ( .A(n19705), .ZN(n19706) );
  NAND3_X1 U22651 ( .A1(n19709), .A2(n19713), .A3(n19706), .ZN(n19707) );
  OAI21_X1 U22652 ( .B1(n19709), .B2(n19708), .A(n19707), .ZN(n19710) );
  AOI21_X1 U22653 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19711), .A(n19710), 
        .ZN(n19712) );
  AOI22_X1 U22654 ( .A1(n19721), .A2(n10562), .B1(n19712), .B2(n19718), .ZN(
        P2_U3604) );
  INV_X1 U22655 ( .A(n19713), .ZN(n19714) );
  OAI22_X1 U22656 ( .A1(n19715), .A2(n19714), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19544), .ZN(n19716) );
  AOI21_X1 U22657 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19717), .A(n19716), 
        .ZN(n19719) );
  AOI22_X1 U22658 ( .A1(n19721), .A2(n19720), .B1(n19719), .B2(n19718), .ZN(
        P2_U3605) );
  INV_X1 U22659 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19722) );
  AOI22_X1 U22660 ( .A1(n19672), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19722), 
        .B2(n19735), .ZN(P2_U3608) );
  INV_X1 U22661 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19734) );
  INV_X1 U22662 ( .A(n19723), .ZN(n19733) );
  AOI21_X1 U22663 ( .B1(n19726), .B2(n19725), .A(n19724), .ZN(n19727) );
  AOI21_X1 U22664 ( .B1(n19729), .B2(n19728), .A(n19727), .ZN(n19732) );
  NOR2_X1 U22665 ( .A1(n19733), .A2(n19730), .ZN(n19731) );
  AOI22_X1 U22666 ( .A1(n19734), .A2(n19733), .B1(n19732), .B2(n19731), .ZN(
        P2_U3609) );
  INV_X1 U22667 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19736) );
  AOI22_X1 U22668 ( .A1(n19672), .A2(n19737), .B1(n19736), .B2(n19735), .ZN(
        P2_U3611) );
  NOR2_X1 U22669 ( .A1(n20532), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20543) );
  NOR2_X1 U22670 ( .A1(n20543), .A2(n12697), .ZN(n19746) );
  INV_X1 U22671 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19738) );
  OR2_X1 U22672 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20532), .ZN(n20634) );
  INV_X2 U22673 ( .A(n20634), .ZN(n20637) );
  AOI21_X1 U22674 ( .B1(n19746), .B2(n19738), .A(n20637), .ZN(P1_U2802) );
  INV_X1 U22675 ( .A(n19739), .ZN(n19742) );
  OAI211_X1 U22676 ( .C1(n19742), .C2(n19741), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .B(n19740), .ZN(n19743) );
  OAI21_X1 U22677 ( .B1(n19744), .B2(n20611), .A(n19743), .ZN(P1_U2803) );
  NOR2_X1 U22678 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19747) );
  OAI21_X1 U22679 ( .B1(n19747), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20634), .ZN(
        n19745) );
  OAI21_X1 U22680 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20634), .A(n19745), 
        .ZN(P1_U2804) );
  NOR2_X1 U22681 ( .A1(n20637), .A2(n19746), .ZN(n20606) );
  OAI21_X1 U22682 ( .B1(BS16), .B2(n19747), .A(n20606), .ZN(n20604) );
  OAI21_X1 U22683 ( .B1(n20606), .B2(n20429), .A(n20604), .ZN(P1_U2805) );
  OAI21_X1 U22684 ( .B1(n19750), .B2(n19749), .A(n19748), .ZN(P1_U2806) );
  NOR4_X1 U22685 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19754) );
  NOR4_X1 U22686 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19753) );
  NOR4_X1 U22687 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19752) );
  NOR4_X1 U22688 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19751) );
  NAND4_X1 U22689 ( .A1(n19754), .A2(n19753), .A3(n19752), .A4(n19751), .ZN(
        n19760) );
  NOR4_X1 U22690 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19758) );
  AOI211_X1 U22691 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_4__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19757) );
  NOR4_X1 U22692 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19756) );
  NOR4_X1 U22693 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19755) );
  NAND4_X1 U22694 ( .A1(n19758), .A2(n19757), .A3(n19756), .A4(n19755), .ZN(
        n19759) );
  NOR2_X1 U22695 ( .A1(n19760), .A2(n19759), .ZN(n20621) );
  INV_X1 U22696 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20601) );
  NOR3_X1 U22697 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19762) );
  OAI21_X1 U22698 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19762), .A(n20621), .ZN(
        n19761) );
  OAI21_X1 U22699 ( .B1(n20621), .B2(n20601), .A(n19761), .ZN(P1_U2807) );
  NAND2_X1 U22700 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n20621), .ZN(n20617) );
  NOR2_X1 U22701 ( .A1(n19762), .A2(n20617), .ZN(n19764) );
  NOR2_X1 U22702 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(n20621), .ZN(n19763)
         );
  AOI211_X1 U22703 ( .C1(n20621), .C2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n19764), 
        .B(n19763), .ZN(P1_U2808) );
  AOI22_X1 U22704 ( .A1(n19832), .A2(n19765), .B1(n19834), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19766) );
  OAI211_X1 U22705 ( .C1(n19782), .C2(n19767), .A(n19766), .B(n19921), .ZN(
        n19768) );
  AOI21_X1 U22706 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n19769), .A(n19768), .ZN(
        n19775) );
  OAI22_X1 U22707 ( .A1(n19772), .A2(n19771), .B1(n19770), .B2(n19843), .ZN(
        n19773) );
  INV_X1 U22708 ( .A(n19773), .ZN(n19774) );
  OAI211_X1 U22709 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n19776), .A(n19775), .B(
        n19774), .ZN(P1_U2831) );
  INV_X1 U22710 ( .A(n19802), .ZN(n19779) );
  AOI21_X1 U22711 ( .B1(n19779), .B2(n19778), .A(n19777), .ZN(n19788) );
  AOI22_X1 U22712 ( .A1(n19832), .A2(n19844), .B1(n19834), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n19780) );
  OAI211_X1 U22713 ( .C1(n19782), .C2(n19781), .A(n19780), .B(n19921), .ZN(
        n19783) );
  AOI21_X1 U22714 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n19788), .A(n19783), .ZN(
        n19786) );
  NOR4_X1 U22715 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19817), .A3(n20554), .A4(
        n19807), .ZN(n19784) );
  AOI22_X1 U22716 ( .A1(n19847), .A2(n19796), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n19784), .ZN(n19785) );
  OAI211_X1 U22717 ( .C1(n19787), .C2(n19843), .A(n19786), .B(n19785), .ZN(
        P1_U2833) );
  INV_X1 U22718 ( .A(n19788), .ZN(n19793) );
  OAI222_X1 U22719 ( .A1(n19793), .A2(n20556), .B1(n19792), .B2(n19791), .C1(
        n19790), .C2(n19789), .ZN(n19794) );
  AOI211_X1 U22720 ( .C1(n19830), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19819), .B(n19794), .ZN(n19799) );
  NOR3_X1 U22721 ( .A1(n19817), .A2(n20554), .A3(n19807), .ZN(n19795) );
  AOI22_X1 U22722 ( .A1(n19797), .A2(n19796), .B1(n19795), .B2(n20556), .ZN(
        n19798) );
  OAI211_X1 U22723 ( .C1(n19800), .C2(n19843), .A(n19799), .B(n19798), .ZN(
        P1_U2834) );
  OAI21_X1 U22724 ( .B1(n19802), .B2(n19807), .A(n19801), .ZN(n19813) );
  OR2_X1 U22725 ( .A1(n19813), .A2(n20554), .ZN(n19806) );
  AOI22_X1 U22726 ( .A1(n19834), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n19830), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19805) );
  NAND2_X1 U22727 ( .A1(n19832), .A2(n19803), .ZN(n19804) );
  AND4_X1 U22728 ( .A1(n19806), .A2(n19805), .A3(n19921), .A4(n19804), .ZN(
        n19811) );
  NOR2_X1 U22729 ( .A1(n19817), .A2(n19807), .ZN(n19808) );
  AOI22_X1 U22730 ( .A1(n19809), .A2(n19840), .B1(n20554), .B2(n19808), .ZN(
        n19810) );
  OAI211_X1 U22731 ( .C1(n19812), .C2(n19843), .A(n19811), .B(n19810), .ZN(
        P1_U2835) );
  INV_X1 U22732 ( .A(n19813), .ZN(n19816) );
  INV_X1 U22733 ( .A(n19814), .ZN(n19833) );
  AOI22_X1 U22734 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19816), .B1(n19815), 
        .B2(n19833), .ZN(n19828) );
  NOR3_X1 U22735 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19817), .A3(n20550), .ZN(
        n19818) );
  AOI211_X1 U22736 ( .C1(n19830), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19819), .B(n19818), .ZN(n19827) );
  INV_X1 U22737 ( .A(n19820), .ZN(n19821) );
  AOI22_X1 U22738 ( .A1(n19832), .A2(n19821), .B1(n19834), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U22739 ( .A1(n19824), .A2(n19840), .B1(n19823), .B2(n19822), .ZN(
        n19825) );
  NAND4_X1 U22740 ( .A1(n19828), .A2(n19827), .A3(n19826), .A4(n19825), .ZN(
        P1_U2836) );
  NOR2_X1 U22741 ( .A1(n19829), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19838) );
  AOI22_X1 U22742 ( .A1(n19832), .A2(n19831), .B1(n19830), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19836) );
  INV_X1 U22743 ( .A(n13879), .ZN(n20431) );
  AOI22_X1 U22744 ( .A1(n19834), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n20431), .B2(
        n19833), .ZN(n19835) );
  OAI211_X1 U22745 ( .C1(n19838), .C2(n19837), .A(n19836), .B(n19835), .ZN(
        n19839) );
  AOI21_X1 U22746 ( .B1(n19841), .B2(n19840), .A(n19839), .ZN(n19842) );
  OAI21_X1 U22747 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19843), .A(
        n19842), .ZN(P1_U2839) );
  AOI22_X1 U22748 ( .A1(n19847), .A2(n19846), .B1(n19845), .B2(n19844), .ZN(
        n19848) );
  OAI21_X1 U22749 ( .B1(n19850), .B2(n19849), .A(n19848), .ZN(P1_U2865) );
  INV_X1 U22750 ( .A(n19851), .ZN(n19852) );
  AOI22_X1 U22751 ( .A1(n19882), .A2(P1_DATAO_REG_26__SCAN_IN), .B1(n19852), 
        .B2(P1_EAX_REG_26__SCAN_IN), .ZN(n19853) );
  OAI21_X1 U22752 ( .B1(n20677), .B2(n20630), .A(n19853), .ZN(P1_U2910) );
  OAI222_X1 U22753 ( .A1(n20630), .A2(n19855), .B1(n19885), .B2(n19854), .C1(
        n20688), .C2(n19862), .ZN(P1_U2921) );
  INV_X1 U22754 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19857) );
  AOI22_X1 U22755 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19856) );
  OAI21_X1 U22756 ( .B1(n19857), .B2(n19885), .A(n19856), .ZN(P1_U2922) );
  INV_X1 U22757 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U22758 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19858) );
  OAI21_X1 U22759 ( .B1(n19859), .B2(n19885), .A(n19858), .ZN(P1_U2923) );
  AOI22_X1 U22760 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n19860), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19883), .ZN(n19861) );
  OAI21_X1 U22761 ( .B1(n20753), .B2(n19862), .A(n19861), .ZN(P1_U2924) );
  AOI22_X1 U22762 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19863) );
  OAI21_X1 U22763 ( .B1(n19864), .B2(n19885), .A(n19863), .ZN(P1_U2925) );
  INV_X1 U22764 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U22765 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19865) );
  OAI21_X1 U22766 ( .B1(n19866), .B2(n19885), .A(n19865), .ZN(P1_U2926) );
  AOI22_X1 U22767 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19867) );
  OAI21_X1 U22768 ( .B1(n13600), .B2(n19885), .A(n19867), .ZN(P1_U2927) );
  INV_X1 U22769 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19869) );
  AOI22_X1 U22770 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19868) );
  OAI21_X1 U22771 ( .B1(n19869), .B2(n19885), .A(n19868), .ZN(P1_U2928) );
  INV_X1 U22772 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19871) );
  AOI22_X1 U22773 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U22774 ( .B1(n19871), .B2(n19885), .A(n19870), .ZN(P1_U2929) );
  AOI22_X1 U22775 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19872) );
  OAI21_X1 U22776 ( .B1(n11679), .B2(n19885), .A(n19872), .ZN(P1_U2930) );
  AOI22_X1 U22777 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19873) );
  OAI21_X1 U22778 ( .B1(n11611), .B2(n19885), .A(n19873), .ZN(P1_U2931) );
  AOI22_X1 U22779 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U22780 ( .B1(n19875), .B2(n19885), .A(n19874), .ZN(P1_U2932) );
  AOI22_X1 U22781 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19876) );
  OAI21_X1 U22782 ( .B1(n19877), .B2(n19885), .A(n19876), .ZN(P1_U2933) );
  AOI22_X1 U22783 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U22784 ( .B1(n19879), .B2(n19885), .A(n19878), .ZN(P1_U2934) );
  AOI22_X1 U22785 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U22786 ( .B1(n19881), .B2(n19885), .A(n19880), .ZN(P1_U2935) );
  AOI22_X1 U22787 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19883), .B1(n19882), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19884) );
  OAI21_X1 U22788 ( .B1(n19886), .B2(n19885), .A(n19884), .ZN(P1_U2936) );
  AOI22_X1 U22789 ( .A1(n19905), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19904), .ZN(n19888) );
  NAND2_X1 U22790 ( .A1(n19892), .A2(n19887), .ZN(n19894) );
  NAND2_X1 U22791 ( .A1(n19888), .A2(n19894), .ZN(P1_U2945) );
  AOI22_X1 U22792 ( .A1(n19905), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n19890) );
  NAND2_X1 U22793 ( .A1(n19892), .A2(n19889), .ZN(n19900) );
  NAND2_X1 U22794 ( .A1(n19890), .A2(n19900), .ZN(P1_U2949) );
  AOI22_X1 U22795 ( .A1(n19905), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n19904), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n19893) );
  NAND2_X1 U22796 ( .A1(n19892), .A2(n19891), .ZN(n19906) );
  NAND2_X1 U22797 ( .A1(n19893), .A2(n19906), .ZN(P1_U2951) );
  AOI22_X1 U22798 ( .A1(n19905), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n19895) );
  NAND2_X1 U22799 ( .A1(n19895), .A2(n19894), .ZN(P1_U2960) );
  AOI22_X1 U22800 ( .A1(n19905), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n19904), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n19897) );
  NAND2_X1 U22801 ( .A1(n19897), .A2(n19896), .ZN(P1_U2961) );
  AOI22_X1 U22802 ( .A1(n19905), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n19899) );
  NAND2_X1 U22803 ( .A1(n19899), .A2(n19898), .ZN(P1_U2962) );
  AOI22_X1 U22804 ( .A1(n19905), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n19901) );
  NAND2_X1 U22805 ( .A1(n19901), .A2(n19900), .ZN(P1_U2964) );
  AOI22_X1 U22806 ( .A1(n19905), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n19903) );
  NAND2_X1 U22807 ( .A1(n19903), .A2(n19902), .ZN(P1_U2965) );
  AOI22_X1 U22808 ( .A1(n19905), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n19904), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n19907) );
  NAND2_X1 U22809 ( .A1(n19907), .A2(n19906), .ZN(P1_U2966) );
  INV_X1 U22810 ( .A(n19908), .ZN(n19912) );
  INV_X1 U22811 ( .A(n19909), .ZN(n19910) );
  AOI22_X1 U22812 ( .A1(n19913), .A2(n19912), .B1(n19911), .B2(n19910), .ZN(
        n19920) );
  NAND2_X1 U22813 ( .A1(n19915), .A2(n19914), .ZN(n19916) );
  OAI22_X1 U22814 ( .A1(n19918), .A2(n19917), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19916), .ZN(n19919) );
  OAI211_X1 U22815 ( .C1(n12944), .C2(n19921), .A(n19920), .B(n19919), .ZN(
        P1_U3031) );
  AND2_X1 U22816 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19922), .ZN(
        P1_U3032) );
  NOR2_X2 U22817 ( .A1(n19924), .A2(n19923), .ZN(n19973) );
  AOI22_X1 U22818 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19973), .B1(DATAI_16_), 
        .B2(n19926), .ZN(n20482) );
  INV_X1 U22819 ( .A(n20049), .ZN(n19928) );
  NAND2_X1 U22820 ( .A1(n19974), .A2(n19932), .ZN(n20271) );
  NAND2_X1 U22821 ( .A1(n20276), .A2(n20220), .ZN(n20053) );
  OR2_X1 U22822 ( .A1(n20351), .A2(n20053), .ZN(n19975) );
  OAI22_X1 U22823 ( .A1(n20515), .A2(n20364), .B1(n20271), .B2(n19975), .ZN(
        n19933) );
  INV_X1 U22824 ( .A(n19933), .ZN(n19944) );
  INV_X1 U22825 ( .A(n20008), .ZN(n19934) );
  OAI21_X1 U22826 ( .B1(n19934), .B2(n20522), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n19935) );
  NAND2_X1 U22827 ( .A1(n19935), .A2(n20398), .ZN(n19942) );
  INV_X1 U22828 ( .A(n13102), .ZN(n19936) );
  OR2_X1 U22829 ( .A1(n20221), .A2(n19936), .ZN(n20051) );
  NOR2_X1 U22830 ( .A1(n20051), .A2(n20431), .ZN(n19939) );
  NAND2_X1 U22831 ( .A1(n19940), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20428) );
  INV_X1 U22832 ( .A(n20275), .ZN(n20280) );
  OR2_X1 U22833 ( .A1(n20222), .A2(n20280), .ZN(n20088) );
  AOI22_X1 U22834 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20088), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n19975), .ZN(n19937) );
  OAI211_X1 U22835 ( .C1(n19942), .C2(n19939), .A(n20278), .B(n19937), .ZN(
        n19980) );
  NOR2_X2 U22836 ( .A1(n19938), .A2(n19986), .ZN(n20473) );
  INV_X1 U22837 ( .A(n19939), .ZN(n19941) );
  OR2_X1 U22838 ( .A1(n19940), .A2(n11609), .ZN(n20281) );
  AOI22_X1 U22839 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19980), .B1(
        n20473), .B2(n19979), .ZN(n19943) );
  OAI211_X1 U22840 ( .C1(n20482), .C2(n20008), .A(n19944), .B(n19943), .ZN(
        P1_U3033) );
  AOI22_X1 U22841 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19973), .B1(DATAI_25_), 
        .B2(n19926), .ZN(n20488) );
  NAND2_X1 U22842 ( .A1(n19974), .A2(n11424), .ZN(n20286) );
  OAI22_X1 U22843 ( .A1(n20515), .A2(n20488), .B1(n19975), .B2(n20286), .ZN(
        n19945) );
  INV_X1 U22844 ( .A(n19945), .ZN(n19948) );
  NOR2_X2 U22845 ( .A1(n19986), .A2(n19946), .ZN(n20483) );
  AOI22_X1 U22846 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19980), .B1(
        n20483), .B2(n19979), .ZN(n19947) );
  OAI211_X1 U22847 ( .C1(n20443), .C2(n20008), .A(n19948), .B(n19947), .ZN(
        P1_U3034) );
  AOI22_X1 U22848 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19973), .B1(DATAI_26_), 
        .B2(n19926), .ZN(n20372) );
  NAND2_X1 U22849 ( .A1(n19974), .A2(n19949), .ZN(n20367) );
  OAI22_X1 U22850 ( .A1(n20515), .A2(n20372), .B1(n19975), .B2(n20367), .ZN(
        n19950) );
  INV_X1 U22851 ( .A(n19950), .ZN(n19953) );
  NOR2_X2 U22852 ( .A1(n19951), .A2(n19986), .ZN(n20489) );
  AOI22_X1 U22853 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19980), .B1(
        n20489), .B2(n19979), .ZN(n19952) );
  OAI211_X1 U22854 ( .C1(n20494), .C2(n20008), .A(n19953), .B(n19952), .ZN(
        P1_U3035) );
  AOI22_X1 U22855 ( .A1(DATAI_19_), .A2(n19926), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n19973), .ZN(n20500) );
  NAND2_X1 U22856 ( .A1(n19974), .A2(n19954), .ZN(n20293) );
  OAI22_X1 U22857 ( .A1(n20515), .A2(n20376), .B1(n19975), .B2(n20293), .ZN(
        n19955) );
  INV_X1 U22858 ( .A(n19955), .ZN(n19958) );
  NOR2_X2 U22859 ( .A1(n19986), .A2(n19956), .ZN(n20495) );
  AOI22_X1 U22860 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19980), .B1(
        n20495), .B2(n19979), .ZN(n19957) );
  OAI211_X1 U22861 ( .C1(n20500), .C2(n20008), .A(n19958), .B(n19957), .ZN(
        P1_U3036) );
  AOI22_X1 U22862 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19973), .B1(DATAI_20_), 
        .B2(n19926), .ZN(n20451) );
  AOI22_X1 U22863 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19973), .B1(DATAI_28_), 
        .B2(n19926), .ZN(n20645) );
  INV_X1 U22864 ( .A(n20645), .ZN(n20448) );
  NAND2_X1 U22865 ( .A1(n19974), .A2(n11437), .ZN(n20297) );
  INV_X1 U22866 ( .A(n19975), .ZN(n19959) );
  AOI22_X1 U22867 ( .A1(n20522), .A2(n20448), .B1(n20641), .B2(n19959), .ZN(
        n19962) );
  NOR2_X2 U22868 ( .A1(n19986), .A2(n19960), .ZN(n20640) );
  AOI22_X1 U22869 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19980), .B1(
        n20640), .B2(n19979), .ZN(n19961) );
  OAI211_X1 U22870 ( .C1(n20451), .C2(n20008), .A(n19962), .B(n19961), .ZN(
        P1_U3037) );
  AOI22_X1 U22871 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19973), .B1(DATAI_29_), 
        .B2(n19926), .ZN(n20385) );
  NAND2_X1 U22872 ( .A1(n19974), .A2(n11421), .ZN(n20380) );
  OAI22_X1 U22873 ( .A1(n20515), .A2(n20385), .B1(n19975), .B2(n20380), .ZN(
        n19964) );
  INV_X1 U22874 ( .A(n19964), .ZN(n19967) );
  NOR2_X2 U22875 ( .A1(n19986), .A2(n19965), .ZN(n20503) );
  AOI22_X1 U22876 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19980), .B1(
        n20503), .B2(n19979), .ZN(n19966) );
  OAI211_X1 U22877 ( .C1(n20508), .C2(n20008), .A(n19967), .B(n19966), .ZN(
        P1_U3038) );
  AOI22_X1 U22878 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19973), .B1(DATAI_22_), 
        .B2(n19926), .ZN(n20516) );
  NAND2_X1 U22879 ( .A1(n19974), .A2(n19968), .ZN(n20304) );
  OAI22_X1 U22880 ( .A1(n20515), .A2(n20389), .B1(n19975), .B2(n20304), .ZN(
        n19969) );
  INV_X1 U22881 ( .A(n19969), .ZN(n19972) );
  NOR2_X2 U22882 ( .A1(n19986), .A2(n19970), .ZN(n20509) );
  AOI22_X1 U22883 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19980), .B1(
        n20509), .B2(n19979), .ZN(n19971) );
  OAI211_X1 U22884 ( .C1(n20516), .C2(n20008), .A(n19972), .B(n19971), .ZN(
        P1_U3039) );
  AOI22_X1 U22885 ( .A1(DATAI_23_), .A2(n19926), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n19973), .ZN(n20463) );
  NAND2_X1 U22886 ( .A1(n19974), .A2(n9938), .ZN(n20309) );
  OAI22_X1 U22887 ( .A1(n20515), .A2(n20527), .B1(n19975), .B2(n20309), .ZN(
        n19976) );
  INV_X1 U22888 ( .A(n19976), .ZN(n19982) );
  INV_X1 U22889 ( .A(n19977), .ZN(n19978) );
  NOR2_X2 U22890 ( .A1(n19986), .A2(n19978), .ZN(n20518) );
  AOI22_X1 U22891 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19980), .B1(
        n20518), .B2(n19979), .ZN(n19981) );
  OAI211_X1 U22892 ( .C1(n20463), .C2(n20008), .A(n19982), .B(n19981), .ZN(
        P1_U3040) );
  INV_X1 U22893 ( .A(n20053), .ZN(n20056) );
  NAND2_X1 U22894 ( .A1(n20056), .A2(n20467), .ZN(n19984) );
  NOR2_X1 U22895 ( .A1(n20397), .A2(n19984), .ZN(n20004) );
  INV_X1 U22896 ( .A(n20051), .ZN(n19983) );
  INV_X1 U22897 ( .A(n20399), .ZN(n20245) );
  AOI21_X1 U22898 ( .B1(n19983), .B2(n20245), .A(n20004), .ZN(n19985) );
  OAI22_X1 U22899 ( .A1(n19985), .A2(n20469), .B1(n19984), .B2(n11609), .ZN(
        n20003) );
  AOI22_X1 U22900 ( .A1(n20474), .A2(n20004), .B1(n20003), .B2(n20473), .ZN(
        n19990) );
  INV_X1 U22901 ( .A(n19984), .ZN(n19988) );
  OAI21_X1 U22902 ( .B1(n20049), .B2(n20429), .A(n19985), .ZN(n19987) );
  OAI221_X1 U22903 ( .B1(n20398), .B2(n19988), .C1(n20469), .C2(n19987), .A(
        n20476), .ZN(n20005) );
  INV_X1 U22904 ( .A(n20482), .ZN(n20352) );
  AOI22_X1 U22905 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20005), .B1(
        n20012), .B2(n20352), .ZN(n19989) );
  OAI211_X1 U22906 ( .C1(n20364), .C2(n20008), .A(n19990), .B(n19989), .ZN(
        P1_U3041) );
  AOI22_X1 U22907 ( .A1(n20484), .A2(n20004), .B1(n20483), .B2(n20003), .ZN(
        n19992) );
  INV_X1 U22908 ( .A(n20443), .ZN(n20485) );
  AOI22_X1 U22909 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20005), .B1(
        n20012), .B2(n20485), .ZN(n19991) );
  OAI211_X1 U22910 ( .C1(n20488), .C2(n20008), .A(n19992), .B(n19991), .ZN(
        P1_U3042) );
  INV_X1 U22911 ( .A(n20367), .ZN(n20490) );
  AOI22_X1 U22912 ( .A1(n20490), .A2(n20004), .B1(n20003), .B2(n20489), .ZN(
        n19994) );
  INV_X1 U22913 ( .A(n20494), .ZN(n20369) );
  AOI22_X1 U22914 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20005), .B1(
        n20012), .B2(n20369), .ZN(n19993) );
  OAI211_X1 U22915 ( .C1(n20372), .C2(n20008), .A(n19994), .B(n19993), .ZN(
        P1_U3043) );
  AOI22_X1 U22916 ( .A1(n20496), .A2(n20004), .B1(n20495), .B2(n20003), .ZN(
        n19996) );
  INV_X1 U22917 ( .A(n20500), .ZN(n20373) );
  AOI22_X1 U22918 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20005), .B1(
        n20012), .B2(n20373), .ZN(n19995) );
  OAI211_X1 U22919 ( .C1(n20376), .C2(n20008), .A(n19996), .B(n19995), .ZN(
        P1_U3044) );
  AOI22_X1 U22920 ( .A1(n20641), .A2(n20004), .B1(n20640), .B2(n20003), .ZN(
        n19998) );
  INV_X1 U22921 ( .A(n20451), .ZN(n20643) );
  AOI22_X1 U22922 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20005), .B1(
        n20012), .B2(n20643), .ZN(n19997) );
  OAI211_X1 U22923 ( .C1(n20645), .C2(n20008), .A(n19998), .B(n19997), .ZN(
        P1_U3045) );
  AOI22_X1 U22924 ( .A1(n20504), .A2(n20004), .B1(n20503), .B2(n20003), .ZN(
        n20000) );
  INV_X1 U22925 ( .A(n20508), .ZN(n20382) );
  AOI22_X1 U22926 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20005), .B1(
        n20012), .B2(n20382), .ZN(n19999) );
  OAI211_X1 U22927 ( .C1(n20385), .C2(n20008), .A(n20000), .B(n19999), .ZN(
        P1_U3046) );
  AOI22_X1 U22928 ( .A1(n20510), .A2(n20004), .B1(n20509), .B2(n20003), .ZN(
        n20002) );
  INV_X1 U22929 ( .A(n20516), .ZN(n20386) );
  AOI22_X1 U22930 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20005), .B1(
        n20012), .B2(n20386), .ZN(n20001) );
  OAI211_X1 U22931 ( .C1(n20389), .C2(n20008), .A(n20002), .B(n20001), .ZN(
        P1_U3047) );
  AOI22_X1 U22932 ( .A1(n20520), .A2(n20004), .B1(n20518), .B2(n20003), .ZN(
        n20007) );
  INV_X1 U22933 ( .A(n20463), .ZN(n20521) );
  AOI22_X1 U22934 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20005), .B1(
        n20012), .B2(n20521), .ZN(n20006) );
  OAI211_X1 U22935 ( .C1(n20527), .C2(n20008), .A(n20007), .B(n20006), .ZN(
        P1_U3048) );
  NAND2_X1 U22936 ( .A1(n20010), .A2(n20009), .ZN(n20149) );
  OR3_X1 U22937 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20467), .A3(
        n20053), .ZN(n20040) );
  OAI22_X1 U22938 ( .A1(n20041), .A2(n20364), .B1(n20271), .B2(n20040), .ZN(
        n20011) );
  INV_X1 U22939 ( .A(n20011), .ZN(n20021) );
  INV_X1 U22940 ( .A(n20081), .ZN(n20013) );
  OAI21_X1 U22941 ( .B1(n20013), .B2(n20012), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20014) );
  NAND2_X1 U22942 ( .A1(n20014), .A2(n20398), .ZN(n20019) );
  NOR2_X1 U22943 ( .A1(n20051), .A2(n13879), .ZN(n20016) );
  NOR2_X1 U22944 ( .A1(n20275), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20017) );
  NOR2_X1 U22945 ( .A1(n20017), .A2(n11609), .ZN(n20154) );
  AOI21_X1 U22946 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20040), .A(n20154), 
        .ZN(n20015) );
  OAI211_X1 U22947 ( .C1(n20019), .C2(n20016), .A(n20278), .B(n20015), .ZN(
        n20044) );
  INV_X1 U22948 ( .A(n20016), .ZN(n20018) );
  INV_X1 U22949 ( .A(n20017), .ZN(n20158) );
  AOI22_X1 U22950 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20044), .B1(
        n20473), .B2(n20043), .ZN(n20020) );
  OAI211_X1 U22951 ( .C1(n20482), .C2(n20081), .A(n20021), .B(n20020), .ZN(
        P1_U3049) );
  OAI22_X1 U22952 ( .A1(n20081), .A2(n20443), .B1(n20286), .B2(n20040), .ZN(
        n20022) );
  INV_X1 U22953 ( .A(n20022), .ZN(n20024) );
  AOI22_X1 U22954 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20044), .B1(
        n20483), .B2(n20043), .ZN(n20023) );
  OAI211_X1 U22955 ( .C1(n20488), .C2(n20041), .A(n20024), .B(n20023), .ZN(
        P1_U3050) );
  OAI22_X1 U22956 ( .A1(n20081), .A2(n20494), .B1(n20367), .B2(n20040), .ZN(
        n20025) );
  INV_X1 U22957 ( .A(n20025), .ZN(n20027) );
  AOI22_X1 U22958 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20044), .B1(
        n20489), .B2(n20043), .ZN(n20026) );
  OAI211_X1 U22959 ( .C1(n20372), .C2(n20041), .A(n20027), .B(n20026), .ZN(
        P1_U3051) );
  OAI22_X1 U22960 ( .A1(n20041), .A2(n20376), .B1(n20293), .B2(n20040), .ZN(
        n20028) );
  INV_X1 U22961 ( .A(n20028), .ZN(n20030) );
  AOI22_X1 U22962 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20044), .B1(
        n20495), .B2(n20043), .ZN(n20029) );
  OAI211_X1 U22963 ( .C1(n20500), .C2(n20081), .A(n20030), .B(n20029), .ZN(
        P1_U3052) );
  OAI22_X1 U22964 ( .A1(n20041), .A2(n20645), .B1(n20297), .B2(n20040), .ZN(
        n20031) );
  INV_X1 U22965 ( .A(n20031), .ZN(n20033) );
  AOI22_X1 U22966 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20044), .B1(
        n20640), .B2(n20043), .ZN(n20032) );
  OAI211_X1 U22967 ( .C1(n20451), .C2(n20081), .A(n20033), .B(n20032), .ZN(
        P1_U3053) );
  OAI22_X1 U22968 ( .A1(n20081), .A2(n20508), .B1(n20380), .B2(n20040), .ZN(
        n20034) );
  INV_X1 U22969 ( .A(n20034), .ZN(n20036) );
  AOI22_X1 U22970 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20044), .B1(
        n20503), .B2(n20043), .ZN(n20035) );
  OAI211_X1 U22971 ( .C1(n20385), .C2(n20041), .A(n20036), .B(n20035), .ZN(
        P1_U3054) );
  OAI22_X1 U22972 ( .A1(n20041), .A2(n20389), .B1(n20304), .B2(n20040), .ZN(
        n20037) );
  INV_X1 U22973 ( .A(n20037), .ZN(n20039) );
  AOI22_X1 U22974 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20044), .B1(
        n20509), .B2(n20043), .ZN(n20038) );
  OAI211_X1 U22975 ( .C1(n20516), .C2(n20081), .A(n20039), .B(n20038), .ZN(
        P1_U3055) );
  OAI22_X1 U22976 ( .A1(n20041), .A2(n20527), .B1(n20309), .B2(n20040), .ZN(
        n20042) );
  INV_X1 U22977 ( .A(n20042), .ZN(n20046) );
  AOI22_X1 U22978 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20044), .B1(
        n20518), .B2(n20043), .ZN(n20045) );
  OAI211_X1 U22979 ( .C1(n20463), .C2(n20081), .A(n20046), .B(n20045), .ZN(
        P1_U3056) );
  INV_X1 U22980 ( .A(n20326), .ZN(n20047) );
  NAND2_X1 U22981 ( .A1(n20465), .A2(n20056), .ZN(n20080) );
  OAI22_X1 U22982 ( .A1(n20094), .A2(n20482), .B1(n20080), .B2(n20271), .ZN(
        n20048) );
  INV_X1 U22983 ( .A(n20048), .ZN(n20061) );
  OAI21_X1 U22984 ( .B1(n20049), .B2(n20322), .A(n20398), .ZN(n20058) );
  NAND2_X1 U22985 ( .A1(n11631), .A2(n20050), .ZN(n20471) );
  OR2_X1 U22986 ( .A1(n20051), .A2(n20471), .ZN(n20052) );
  INV_X1 U22987 ( .A(n20059), .ZN(n20055) );
  OAI21_X1 U22988 ( .B1(n20467), .B2(n20053), .A(n20469), .ZN(n20054) );
  OAI211_X1 U22989 ( .C1(n20058), .C2(n20055), .A(n20476), .B(n20054), .ZN(
        n20084) );
  NAND2_X1 U22990 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20056), .ZN(
        n20057) );
  OAI22_X1 U22991 ( .A1(n20059), .A2(n20058), .B1(n11609), .B2(n20057), .ZN(
        n20083) );
  AOI22_X1 U22992 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20084), .B1(
        n20473), .B2(n20083), .ZN(n20060) );
  OAI211_X1 U22993 ( .C1(n20364), .C2(n20081), .A(n20061), .B(n20060), .ZN(
        P1_U3057) );
  OAI22_X1 U22994 ( .A1(n20094), .A2(n20443), .B1(n20080), .B2(n20286), .ZN(
        n20062) );
  INV_X1 U22995 ( .A(n20062), .ZN(n20064) );
  AOI22_X1 U22996 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20084), .B1(
        n20483), .B2(n20083), .ZN(n20063) );
  OAI211_X1 U22997 ( .C1(n20488), .C2(n20081), .A(n20064), .B(n20063), .ZN(
        P1_U3058) );
  OAI22_X1 U22998 ( .A1(n20081), .A2(n20372), .B1(n20367), .B2(n20080), .ZN(
        n20065) );
  INV_X1 U22999 ( .A(n20065), .ZN(n20067) );
  AOI22_X1 U23000 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20084), .B1(
        n20489), .B2(n20083), .ZN(n20066) );
  OAI211_X1 U23001 ( .C1(n20494), .C2(n20094), .A(n20067), .B(n20066), .ZN(
        P1_U3059) );
  OAI22_X1 U23002 ( .A1(n20081), .A2(n20376), .B1(n20293), .B2(n20080), .ZN(
        n20068) );
  INV_X1 U23003 ( .A(n20068), .ZN(n20070) );
  AOI22_X1 U23004 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20084), .B1(
        n20495), .B2(n20083), .ZN(n20069) );
  OAI211_X1 U23005 ( .C1(n20500), .C2(n20094), .A(n20070), .B(n20069), .ZN(
        P1_U3060) );
  OAI22_X1 U23006 ( .A1(n20081), .A2(n20645), .B1(n20297), .B2(n20080), .ZN(
        n20071) );
  INV_X1 U23007 ( .A(n20071), .ZN(n20073) );
  AOI22_X1 U23008 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20084), .B1(
        n20640), .B2(n20083), .ZN(n20072) );
  OAI211_X1 U23009 ( .C1(n20451), .C2(n20094), .A(n20073), .B(n20072), .ZN(
        P1_U3061) );
  OAI22_X1 U23010 ( .A1(n20094), .A2(n20508), .B1(n20380), .B2(n20080), .ZN(
        n20074) );
  INV_X1 U23011 ( .A(n20074), .ZN(n20076) );
  AOI22_X1 U23012 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20084), .B1(
        n20503), .B2(n20083), .ZN(n20075) );
  OAI211_X1 U23013 ( .C1(n20385), .C2(n20081), .A(n20076), .B(n20075), .ZN(
        P1_U3062) );
  OAI22_X1 U23014 ( .A1(n20081), .A2(n20389), .B1(n20304), .B2(n20080), .ZN(
        n20077) );
  INV_X1 U23015 ( .A(n20077), .ZN(n20079) );
  AOI22_X1 U23016 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20084), .B1(
        n20509), .B2(n20083), .ZN(n20078) );
  OAI211_X1 U23017 ( .C1(n20516), .C2(n20094), .A(n20079), .B(n20078), .ZN(
        P1_U3063) );
  OAI22_X1 U23018 ( .A1(n20081), .A2(n20527), .B1(n20309), .B2(n20080), .ZN(
        n20082) );
  INV_X1 U23019 ( .A(n20082), .ZN(n20086) );
  AOI22_X1 U23020 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20084), .B1(
        n20518), .B2(n20083), .ZN(n20085) );
  OAI211_X1 U23021 ( .C1(n20463), .C2(n20094), .A(n20086), .B(n20085), .ZN(
        P1_U3064) );
  OR2_X1 U23022 ( .A1(n20351), .A2(n20150), .ZN(n20104) );
  OR2_X1 U23023 ( .A1(n13102), .A2(n20087), .ZN(n20188) );
  NAND2_X1 U23024 ( .A1(n13879), .A2(n20398), .ZN(n20092) );
  INV_X1 U23025 ( .A(n20088), .ZN(n20090) );
  INV_X1 U23026 ( .A(n20428), .ZN(n20089) );
  NAND2_X1 U23027 ( .A1(n20090), .A2(n20089), .ZN(n20091) );
  OAI21_X1 U23028 ( .B1(n20188), .B2(n20092), .A(n20091), .ZN(n20116) );
  INV_X1 U23029 ( .A(n20116), .ZN(n20103) );
  INV_X1 U23030 ( .A(n20473), .ZN(n20192) );
  OAI22_X1 U23031 ( .A1(n20271), .A2(n20104), .B1(n20103), .B2(n20192), .ZN(
        n20093) );
  INV_X1 U23032 ( .A(n20093), .ZN(n20100) );
  INV_X1 U23033 ( .A(n20104), .ZN(n20117) );
  INV_X1 U23034 ( .A(n20148), .ZN(n20095) );
  OAI21_X1 U23035 ( .B1(n20118), .B2(n20095), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20096) );
  OAI21_X1 U23036 ( .B1(n20431), .B2(n20188), .A(n20096), .ZN(n20098) );
  INV_X1 U23037 ( .A(n20364), .ZN(n20479) );
  AOI22_X1 U23038 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20119), .B1(
        n20118), .B2(n20479), .ZN(n20099) );
  OAI211_X1 U23039 ( .C1(n20482), .C2(n20148), .A(n20100), .B(n20099), .ZN(
        P1_U3065) );
  AOI22_X1 U23040 ( .A1(n20484), .A2(n20117), .B1(n20483), .B2(n20116), .ZN(
        n20102) );
  INV_X1 U23041 ( .A(n20488), .ZN(n20440) );
  AOI22_X1 U23042 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20119), .B1(
        n20118), .B2(n20440), .ZN(n20101) );
  OAI211_X1 U23043 ( .C1(n20443), .C2(n20148), .A(n20102), .B(n20101), .ZN(
        P1_U3066) );
  INV_X1 U23044 ( .A(n20489), .ZN(n20204) );
  OAI22_X1 U23045 ( .A1(n20367), .A2(n20104), .B1(n20103), .B2(n20204), .ZN(
        n20105) );
  INV_X1 U23046 ( .A(n20105), .ZN(n20107) );
  INV_X1 U23047 ( .A(n20372), .ZN(n20491) );
  AOI22_X1 U23048 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20119), .B1(
        n20118), .B2(n20491), .ZN(n20106) );
  OAI211_X1 U23049 ( .C1(n20494), .C2(n20148), .A(n20107), .B(n20106), .ZN(
        P1_U3067) );
  AOI22_X1 U23050 ( .A1(n20496), .A2(n20117), .B1(n20495), .B2(n20116), .ZN(
        n20109) );
  INV_X1 U23051 ( .A(n20376), .ZN(n20497) );
  AOI22_X1 U23052 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20119), .B1(
        n20118), .B2(n20497), .ZN(n20108) );
  OAI211_X1 U23053 ( .C1(n20500), .C2(n20148), .A(n20109), .B(n20108), .ZN(
        P1_U3068) );
  AOI22_X1 U23054 ( .A1(n20641), .A2(n20117), .B1(n20640), .B2(n20116), .ZN(
        n20111) );
  AOI22_X1 U23055 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20119), .B1(
        n20118), .B2(n20448), .ZN(n20110) );
  OAI211_X1 U23056 ( .C1(n20451), .C2(n20148), .A(n20111), .B(n20110), .ZN(
        P1_U3069) );
  AOI22_X1 U23057 ( .A1(n20504), .A2(n20117), .B1(n20503), .B2(n20116), .ZN(
        n20113) );
  INV_X1 U23058 ( .A(n20385), .ZN(n20505) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20119), .B1(
        n20118), .B2(n20505), .ZN(n20112) );
  OAI211_X1 U23060 ( .C1(n20508), .C2(n20148), .A(n20113), .B(n20112), .ZN(
        P1_U3070) );
  AOI22_X1 U23061 ( .A1(n20510), .A2(n20117), .B1(n20509), .B2(n20116), .ZN(
        n20115) );
  INV_X1 U23062 ( .A(n20389), .ZN(n20511) );
  AOI22_X1 U23063 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20119), .B1(
        n20118), .B2(n20511), .ZN(n20114) );
  OAI211_X1 U23064 ( .C1(n20516), .C2(n20148), .A(n20115), .B(n20114), .ZN(
        P1_U3071) );
  AOI22_X1 U23065 ( .A1(n20520), .A2(n20117), .B1(n20518), .B2(n20116), .ZN(
        n20121) );
  INV_X1 U23066 ( .A(n20527), .ZN(n20458) );
  AOI22_X1 U23067 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20119), .B1(
        n20118), .B2(n20458), .ZN(n20120) );
  OAI211_X1 U23068 ( .C1(n20463), .C2(n20148), .A(n20121), .B(n20120), .ZN(
        P1_U3072) );
  NOR2_X1 U23069 ( .A1(n20150), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20126) );
  INV_X1 U23070 ( .A(n20126), .ZN(n20122) );
  NOR2_X1 U23071 ( .A1(n20397), .A2(n20122), .ZN(n20143) );
  INV_X1 U23072 ( .A(n20188), .ZN(n20153) );
  AOI21_X1 U23073 ( .B1(n20153), .B2(n20245), .A(n20143), .ZN(n20123) );
  OAI22_X1 U23074 ( .A1(n20123), .A2(n20469), .B1(n20122), .B2(n11609), .ZN(
        n20142) );
  AOI22_X1 U23075 ( .A1(n20474), .A2(n20143), .B1(n20473), .B2(n20142), .ZN(
        n20129) );
  INV_X1 U23076 ( .A(n20199), .ZN(n20124) );
  OAI21_X1 U23077 ( .B1(n20124), .B2(n20429), .A(n20123), .ZN(n20125) );
  OAI221_X1 U23078 ( .B1(n20398), .B2(n20126), .C1(n20469), .C2(n20125), .A(
        n20476), .ZN(n20145) );
  AOI22_X1 U23079 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20145), .B1(
        n20144), .B2(n20352), .ZN(n20128) );
  OAI211_X1 U23080 ( .C1(n20364), .C2(n20148), .A(n20129), .B(n20128), .ZN(
        P1_U3073) );
  AOI22_X1 U23081 ( .A1(n20484), .A2(n20143), .B1(n20483), .B2(n20142), .ZN(
        n20131) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20145), .B1(
        n20144), .B2(n20485), .ZN(n20130) );
  OAI211_X1 U23083 ( .C1(n20488), .C2(n20148), .A(n20131), .B(n20130), .ZN(
        P1_U3074) );
  AOI22_X1 U23084 ( .A1(n20490), .A2(n20143), .B1(n20489), .B2(n20142), .ZN(
        n20133) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20145), .B1(
        n20144), .B2(n20369), .ZN(n20132) );
  OAI211_X1 U23086 ( .C1(n20372), .C2(n20148), .A(n20133), .B(n20132), .ZN(
        P1_U3075) );
  AOI22_X1 U23087 ( .A1(n20496), .A2(n20143), .B1(n20495), .B2(n20142), .ZN(
        n20135) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20145), .B1(
        n20144), .B2(n20373), .ZN(n20134) );
  OAI211_X1 U23089 ( .C1(n20376), .C2(n20148), .A(n20135), .B(n20134), .ZN(
        P1_U3076) );
  AOI22_X1 U23090 ( .A1(n20641), .A2(n20143), .B1(n20640), .B2(n20142), .ZN(
        n20137) );
  AOI22_X1 U23091 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20145), .B1(
        n20144), .B2(n20643), .ZN(n20136) );
  OAI211_X1 U23092 ( .C1(n20645), .C2(n20148), .A(n20137), .B(n20136), .ZN(
        P1_U3077) );
  AOI22_X1 U23093 ( .A1(n20504), .A2(n20143), .B1(n20503), .B2(n20142), .ZN(
        n20139) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20145), .B1(
        n20144), .B2(n20382), .ZN(n20138) );
  OAI211_X1 U23095 ( .C1(n20385), .C2(n20148), .A(n20139), .B(n20138), .ZN(
        P1_U3078) );
  AOI22_X1 U23096 ( .A1(n20510), .A2(n20143), .B1(n20509), .B2(n20142), .ZN(
        n20141) );
  AOI22_X1 U23097 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20145), .B1(
        n20144), .B2(n20386), .ZN(n20140) );
  OAI211_X1 U23098 ( .C1(n20389), .C2(n20148), .A(n20141), .B(n20140), .ZN(
        P1_U3079) );
  AOI22_X1 U23099 ( .A1(n20520), .A2(n20143), .B1(n20518), .B2(n20142), .ZN(
        n20147) );
  AOI22_X1 U23100 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20145), .B1(
        n20144), .B2(n20521), .ZN(n20146) );
  OAI211_X1 U23101 ( .C1(n20527), .C2(n20148), .A(n20147), .B(n20146), .ZN(
        P1_U3080) );
  NOR2_X1 U23102 ( .A1(n20467), .A2(n20150), .ZN(n20195) );
  AND2_X1 U23103 ( .A1(n20397), .A2(n20195), .ZN(n20156) );
  INV_X1 U23104 ( .A(n20156), .ZN(n20181) );
  OAI22_X1 U23105 ( .A1(n20187), .A2(n20364), .B1(n20271), .B2(n20181), .ZN(
        n20151) );
  INV_X1 U23106 ( .A(n20151), .ZN(n20162) );
  NAND3_X1 U23107 ( .A1(n20646), .A2(n20187), .A3(n20398), .ZN(n20152) );
  NAND2_X1 U23108 ( .A1(n20398), .A2(n20429), .ZN(n20353) );
  NAND2_X1 U23109 ( .A1(n20152), .A2(n20353), .ZN(n20157) );
  NAND2_X1 U23110 ( .A1(n20153), .A2(n20431), .ZN(n20159) );
  AOI21_X1 U23111 ( .B1(n20157), .B2(n20159), .A(n20154), .ZN(n20155) );
  OAI211_X1 U23112 ( .C1(n20156), .C2(n20357), .A(n20435), .B(n20155), .ZN(
        n20184) );
  INV_X1 U23113 ( .A(n20157), .ZN(n20160) );
  OAI22_X1 U23114 ( .A1(n20160), .A2(n20159), .B1(n20158), .B2(n20428), .ZN(
        n20183) );
  AOI22_X1 U23115 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20184), .B1(
        n20473), .B2(n20183), .ZN(n20161) );
  OAI211_X1 U23116 ( .C1(n20482), .C2(n20646), .A(n20162), .B(n20161), .ZN(
        P1_U3081) );
  OAI22_X1 U23117 ( .A1(n20646), .A2(n20443), .B1(n20286), .B2(n20181), .ZN(
        n20163) );
  INV_X1 U23118 ( .A(n20163), .ZN(n20165) );
  AOI22_X1 U23119 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20184), .B1(
        n20483), .B2(n20183), .ZN(n20164) );
  OAI211_X1 U23120 ( .C1(n20488), .C2(n20187), .A(n20165), .B(n20164), .ZN(
        P1_U3082) );
  OAI22_X1 U23121 ( .A1(n20187), .A2(n20372), .B1(n20367), .B2(n20181), .ZN(
        n20166) );
  INV_X1 U23122 ( .A(n20166), .ZN(n20168) );
  AOI22_X1 U23123 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20184), .B1(
        n20489), .B2(n20183), .ZN(n20167) );
  OAI211_X1 U23124 ( .C1(n20494), .C2(n20646), .A(n20168), .B(n20167), .ZN(
        P1_U3083) );
  OAI22_X1 U23125 ( .A1(n20187), .A2(n20376), .B1(n20293), .B2(n20181), .ZN(
        n20169) );
  INV_X1 U23126 ( .A(n20169), .ZN(n20171) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20184), .B1(
        n20495), .B2(n20183), .ZN(n20170) );
  OAI211_X1 U23128 ( .C1(n20500), .C2(n20646), .A(n20171), .B(n20170), .ZN(
        P1_U3084) );
  OAI22_X1 U23129 ( .A1(n20187), .A2(n20645), .B1(n20297), .B2(n20181), .ZN(
        n20172) );
  INV_X1 U23130 ( .A(n20172), .ZN(n20174) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20184), .B1(
        n20640), .B2(n20183), .ZN(n20173) );
  OAI211_X1 U23132 ( .C1(n20451), .C2(n20646), .A(n20174), .B(n20173), .ZN(
        P1_U3085) );
  OAI22_X1 U23133 ( .A1(n20646), .A2(n20508), .B1(n20380), .B2(n20181), .ZN(
        n20175) );
  INV_X1 U23134 ( .A(n20175), .ZN(n20177) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20184), .B1(
        n20503), .B2(n20183), .ZN(n20176) );
  OAI211_X1 U23136 ( .C1(n20385), .C2(n20187), .A(n20177), .B(n20176), .ZN(
        P1_U3086) );
  OAI22_X1 U23137 ( .A1(n20187), .A2(n20389), .B1(n20304), .B2(n20181), .ZN(
        n20178) );
  INV_X1 U23138 ( .A(n20178), .ZN(n20180) );
  AOI22_X1 U23139 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20184), .B1(
        n20509), .B2(n20183), .ZN(n20179) );
  OAI211_X1 U23140 ( .C1(n20516), .C2(n20646), .A(n20180), .B(n20179), .ZN(
        P1_U3087) );
  OAI22_X1 U23141 ( .A1(n20646), .A2(n20463), .B1(n20309), .B2(n20181), .ZN(
        n20182) );
  INV_X1 U23142 ( .A(n20182), .ZN(n20186) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20184), .B1(
        n20518), .B2(n20183), .ZN(n20185) );
  OAI211_X1 U23144 ( .C1(n20527), .C2(n20187), .A(n20186), .B(n20185), .ZN(
        P1_U3088) );
  OAI21_X1 U23145 ( .B1(n20188), .B2(n20471), .A(n20206), .ZN(n20189) );
  NAND2_X1 U23146 ( .A1(n20189), .A2(n20398), .ZN(n20191) );
  NAND2_X1 U23147 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20195), .ZN(n20190) );
  NAND2_X1 U23148 ( .A1(n20191), .A2(n20190), .ZN(n20639) );
  INV_X1 U23149 ( .A(n20639), .ZN(n20205) );
  OAI22_X1 U23150 ( .A1(n20271), .A2(n20206), .B1(n20205), .B2(n20192), .ZN(
        n20193) );
  INV_X1 U23151 ( .A(n20193), .ZN(n20201) );
  INV_X1 U23152 ( .A(n20195), .ZN(n20196) );
  OAI21_X1 U23153 ( .B1(n20475), .B2(n20197), .A(n20196), .ZN(n20198) );
  NAND2_X1 U23154 ( .A1(n20198), .A2(n20476), .ZN(n20638) );
  AOI22_X1 U23155 ( .A1(n20638), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n20644), .B2(n20352), .ZN(n20200) );
  OAI211_X1 U23156 ( .C1(n20364), .C2(n20646), .A(n20201), .B(n20200), .ZN(
        P1_U3089) );
  INV_X1 U23157 ( .A(n20644), .ZN(n20215) );
  INV_X1 U23158 ( .A(n20206), .ZN(n20642) );
  AOI22_X1 U23159 ( .A1(n20642), .A2(n20484), .B1(n20483), .B2(n20639), .ZN(
        n20203) );
  INV_X1 U23160 ( .A(n20646), .ZN(n20212) );
  AOI22_X1 U23161 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20638), .B1(
        n20212), .B2(n20440), .ZN(n20202) );
  OAI211_X1 U23162 ( .C1(n20443), .C2(n20215), .A(n20203), .B(n20202), .ZN(
        P1_U3090) );
  OAI22_X1 U23163 ( .A1(n20367), .A2(n20206), .B1(n20205), .B2(n20204), .ZN(
        n20207) );
  INV_X1 U23164 ( .A(n20207), .ZN(n20209) );
  AOI22_X1 U23165 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20638), .B1(
        n20212), .B2(n20491), .ZN(n20208) );
  OAI211_X1 U23166 ( .C1(n20494), .C2(n20215), .A(n20209), .B(n20208), .ZN(
        P1_U3091) );
  AOI22_X1 U23167 ( .A1(n20642), .A2(n20496), .B1(n20495), .B2(n20639), .ZN(
        n20211) );
  AOI22_X1 U23168 ( .A1(n20638), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n20644), .B2(n20373), .ZN(n20210) );
  OAI211_X1 U23169 ( .C1(n20376), .C2(n20646), .A(n20211), .B(n20210), .ZN(
        P1_U3092) );
  AOI22_X1 U23170 ( .A1(n20642), .A2(n20504), .B1(n20503), .B2(n20639), .ZN(
        n20214) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20638), .B1(
        n20212), .B2(n20505), .ZN(n20213) );
  OAI211_X1 U23172 ( .C1(n20508), .C2(n20215), .A(n20214), .B(n20213), .ZN(
        P1_U3094) );
  AOI22_X1 U23173 ( .A1(n20642), .A2(n20510), .B1(n20509), .B2(n20639), .ZN(
        n20217) );
  AOI22_X1 U23174 ( .A1(n20638), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n20644), .B2(n20386), .ZN(n20216) );
  OAI211_X1 U23175 ( .C1(n20389), .C2(n20646), .A(n20217), .B(n20216), .ZN(
        P1_U3095) );
  AOI22_X1 U23176 ( .A1(n20642), .A2(n20520), .B1(n20518), .B2(n20639), .ZN(
        n20219) );
  AOI22_X1 U23177 ( .A1(n20638), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n20644), .B2(n20521), .ZN(n20218) );
  OAI211_X1 U23178 ( .C1(n20527), .C2(n20646), .A(n20219), .B(n20218), .ZN(
        P1_U3096) );
  NAND2_X1 U23179 ( .A1(n20220), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20316) );
  NAND2_X1 U23180 ( .A1(n20221), .A2(n13102), .ZN(n20274) );
  AOI21_X1 U23181 ( .B1(n20319), .B2(n13879), .A(n10124), .ZN(n20224) );
  NAND2_X1 U23182 ( .A1(n20222), .A2(n20275), .ZN(n20359) );
  OAI22_X1 U23183 ( .A1(n20224), .A2(n20469), .B1(n20359), .B2(n20281), .ZN(
        n20241) );
  AOI22_X1 U23184 ( .A1(n20474), .A2(n10124), .B1(n20241), .B2(n20473), .ZN(
        n20228) );
  INV_X1 U23185 ( .A(n20270), .ZN(n20223) );
  OAI21_X1 U23186 ( .B1(n20223), .B2(n20644), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20225) );
  NAND2_X1 U23187 ( .A1(n20225), .A2(n20224), .ZN(n20226) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20242), .B1(
        n20644), .B2(n20479), .ZN(n20227) );
  OAI211_X1 U23189 ( .C1(n20482), .C2(n20270), .A(n20228), .B(n20227), .ZN(
        P1_U3097) );
  AOI22_X1 U23190 ( .A1(n10124), .A2(n20484), .B1(n20483), .B2(n20241), .ZN(
        n20230) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20242), .B1(
        n20644), .B2(n20440), .ZN(n20229) );
  OAI211_X1 U23192 ( .C1(n20443), .C2(n20270), .A(n20230), .B(n20229), .ZN(
        P1_U3098) );
  AOI22_X1 U23193 ( .A1(n20490), .A2(n10124), .B1(n20241), .B2(n20489), .ZN(
        n20232) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20242), .B1(
        n20644), .B2(n20491), .ZN(n20231) );
  OAI211_X1 U23195 ( .C1(n20494), .C2(n20270), .A(n20232), .B(n20231), .ZN(
        P1_U3099) );
  AOI22_X1 U23196 ( .A1(n10124), .A2(n20496), .B1(n20495), .B2(n20241), .ZN(
        n20234) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20242), .B1(
        n20644), .B2(n20497), .ZN(n20233) );
  OAI211_X1 U23198 ( .C1(n20500), .C2(n20270), .A(n20234), .B(n20233), .ZN(
        P1_U3100) );
  AOI22_X1 U23199 ( .A1(n20641), .A2(n10124), .B1(n20640), .B2(n20241), .ZN(
        n20236) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20242), .B1(
        n20644), .B2(n20448), .ZN(n20235) );
  OAI211_X1 U23201 ( .C1(n20451), .C2(n20270), .A(n20236), .B(n20235), .ZN(
        P1_U3101) );
  AOI22_X1 U23202 ( .A1(n10124), .A2(n20504), .B1(n20503), .B2(n20241), .ZN(
        n20238) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20242), .B1(
        n20644), .B2(n20505), .ZN(n20237) );
  OAI211_X1 U23204 ( .C1(n20508), .C2(n20270), .A(n20238), .B(n20237), .ZN(
        P1_U3102) );
  AOI22_X1 U23205 ( .A1(n10124), .A2(n20510), .B1(n20509), .B2(n20241), .ZN(
        n20240) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20242), .B1(
        n20644), .B2(n20511), .ZN(n20239) );
  OAI211_X1 U23207 ( .C1(n20516), .C2(n20270), .A(n20240), .B(n20239), .ZN(
        P1_U3103) );
  AOI22_X1 U23208 ( .A1(n10124), .A2(n20520), .B1(n20518), .B2(n20241), .ZN(
        n20244) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20242), .B1(
        n20644), .B2(n20458), .ZN(n20243) );
  OAI211_X1 U23210 ( .C1(n20463), .C2(n20270), .A(n20244), .B(n20243), .ZN(
        P1_U3104) );
  NOR2_X1 U23211 ( .A1(n20316), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20249) );
  INV_X1 U23212 ( .A(n20249), .ZN(n20246) );
  NOR2_X1 U23213 ( .A1(n20397), .A2(n20246), .ZN(n20265) );
  AOI21_X1 U23214 ( .B1(n20319), .B2(n20245), .A(n20265), .ZN(n20247) );
  OAI22_X1 U23215 ( .A1(n20247), .A2(n20469), .B1(n20246), .B2(n11609), .ZN(
        n20264) );
  AOI22_X1 U23216 ( .A1(n20474), .A2(n20265), .B1(n20264), .B2(n20473), .ZN(
        n20251) );
  OAI21_X1 U23217 ( .B1(n20323), .B2(n20429), .A(n20247), .ZN(n20248) );
  OAI221_X1 U23218 ( .B1(n20398), .B2(n20249), .C1(n20469), .C2(n20248), .A(
        n20476), .ZN(n20267) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20267), .B1(
        n20266), .B2(n20352), .ZN(n20250) );
  OAI211_X1 U23220 ( .C1(n20364), .C2(n20270), .A(n20251), .B(n20250), .ZN(
        P1_U3105) );
  AOI22_X1 U23221 ( .A1(n20484), .A2(n20265), .B1(n20483), .B2(n20264), .ZN(
        n20253) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20267), .B1(
        n20266), .B2(n20485), .ZN(n20252) );
  OAI211_X1 U23223 ( .C1(n20488), .C2(n20270), .A(n20253), .B(n20252), .ZN(
        P1_U3106) );
  AOI22_X1 U23224 ( .A1(n20490), .A2(n20265), .B1(n20264), .B2(n20489), .ZN(
        n20255) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20267), .B1(
        n20266), .B2(n20369), .ZN(n20254) );
  OAI211_X1 U23226 ( .C1(n20372), .C2(n20270), .A(n20255), .B(n20254), .ZN(
        P1_U3107) );
  AOI22_X1 U23227 ( .A1(n20496), .A2(n20265), .B1(n20495), .B2(n20264), .ZN(
        n20257) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20267), .B1(
        n20266), .B2(n20373), .ZN(n20256) );
  OAI211_X1 U23229 ( .C1(n20376), .C2(n20270), .A(n20257), .B(n20256), .ZN(
        P1_U3108) );
  AOI22_X1 U23230 ( .A1(n20641), .A2(n20265), .B1(n20640), .B2(n20264), .ZN(
        n20259) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20267), .B1(
        n20266), .B2(n20643), .ZN(n20258) );
  OAI211_X1 U23232 ( .C1(n20645), .C2(n20270), .A(n20259), .B(n20258), .ZN(
        P1_U3109) );
  AOI22_X1 U23233 ( .A1(n20504), .A2(n20265), .B1(n20503), .B2(n20264), .ZN(
        n20261) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20267), .B1(
        n20266), .B2(n20382), .ZN(n20260) );
  OAI211_X1 U23235 ( .C1(n20385), .C2(n20270), .A(n20261), .B(n20260), .ZN(
        P1_U3110) );
  AOI22_X1 U23236 ( .A1(n20510), .A2(n20265), .B1(n20509), .B2(n20264), .ZN(
        n20263) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20267), .B1(
        n20266), .B2(n20386), .ZN(n20262) );
  OAI211_X1 U23238 ( .C1(n20389), .C2(n20270), .A(n20263), .B(n20262), .ZN(
        P1_U3111) );
  AOI22_X1 U23239 ( .A1(n20520), .A2(n20265), .B1(n20518), .B2(n20264), .ZN(
        n20269) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20267), .B1(
        n20266), .B2(n20521), .ZN(n20268) );
  OAI211_X1 U23241 ( .C1(n20527), .C2(n20270), .A(n20269), .B(n20268), .ZN(
        P1_U3112) );
  NOR2_X1 U23242 ( .A1(n20467), .A2(n20316), .ZN(n20325) );
  INV_X1 U23243 ( .A(n20325), .ZN(n20320) );
  OR2_X1 U23244 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20320), .ZN(
        n20308) );
  OAI22_X1 U23245 ( .A1(n20310), .A2(n20364), .B1(n20271), .B2(n20308), .ZN(
        n20272) );
  INV_X1 U23246 ( .A(n20272), .ZN(n20285) );
  NAND3_X1 U23247 ( .A1(n20343), .A2(n20310), .A3(n20398), .ZN(n20273) );
  NAND2_X1 U23248 ( .A1(n20273), .A2(n20353), .ZN(n20279) );
  OR2_X1 U23249 ( .A1(n20274), .A2(n13879), .ZN(n20282) );
  AOI22_X1 U23250 ( .A1(n20279), .A2(n20282), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20308), .ZN(n20277) );
  OAI21_X1 U23251 ( .B1(n20276), .B2(n20275), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20434) );
  NAND3_X1 U23252 ( .A1(n20278), .A2(n20277), .A3(n20434), .ZN(n20313) );
  INV_X1 U23253 ( .A(n20279), .ZN(n20283) );
  NAND2_X1 U23254 ( .A1(n20280), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20427) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20313), .B1(
        n20473), .B2(n20312), .ZN(n20284) );
  OAI211_X1 U23256 ( .C1(n20482), .C2(n20343), .A(n20285), .B(n20284), .ZN(
        P1_U3113) );
  OAI22_X1 U23257 ( .A1(n20343), .A2(n20443), .B1(n20286), .B2(n20308), .ZN(
        n20287) );
  INV_X1 U23258 ( .A(n20287), .ZN(n20289) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20313), .B1(
        n20483), .B2(n20312), .ZN(n20288) );
  OAI211_X1 U23260 ( .C1(n20488), .C2(n20310), .A(n20289), .B(n20288), .ZN(
        P1_U3114) );
  OAI22_X1 U23261 ( .A1(n20343), .A2(n20494), .B1(n20367), .B2(n20308), .ZN(
        n20290) );
  INV_X1 U23262 ( .A(n20290), .ZN(n20292) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20313), .B1(
        n20489), .B2(n20312), .ZN(n20291) );
  OAI211_X1 U23264 ( .C1(n20372), .C2(n20310), .A(n20292), .B(n20291), .ZN(
        P1_U3115) );
  OAI22_X1 U23265 ( .A1(n20343), .A2(n20500), .B1(n20293), .B2(n20308), .ZN(
        n20294) );
  INV_X1 U23266 ( .A(n20294), .ZN(n20296) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20313), .B1(
        n20495), .B2(n20312), .ZN(n20295) );
  OAI211_X1 U23268 ( .C1(n20376), .C2(n20310), .A(n20296), .B(n20295), .ZN(
        P1_U3116) );
  OAI22_X1 U23269 ( .A1(n20310), .A2(n20645), .B1(n20297), .B2(n20308), .ZN(
        n20298) );
  INV_X1 U23270 ( .A(n20298), .ZN(n20300) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20313), .B1(
        n20640), .B2(n20312), .ZN(n20299) );
  OAI211_X1 U23272 ( .C1(n20451), .C2(n20343), .A(n20300), .B(n20299), .ZN(
        P1_U3117) );
  OAI22_X1 U23273 ( .A1(n20310), .A2(n20385), .B1(n20380), .B2(n20308), .ZN(
        n20301) );
  INV_X1 U23274 ( .A(n20301), .ZN(n20303) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20313), .B1(
        n20503), .B2(n20312), .ZN(n20302) );
  OAI211_X1 U23276 ( .C1(n20508), .C2(n20343), .A(n20303), .B(n20302), .ZN(
        P1_U3118) );
  OAI22_X1 U23277 ( .A1(n20343), .A2(n20516), .B1(n20304), .B2(n20308), .ZN(
        n20305) );
  INV_X1 U23278 ( .A(n20305), .ZN(n20307) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20313), .B1(
        n20509), .B2(n20312), .ZN(n20306) );
  OAI211_X1 U23280 ( .C1(n20389), .C2(n20310), .A(n20307), .B(n20306), .ZN(
        P1_U3119) );
  OAI22_X1 U23281 ( .A1(n20310), .A2(n20527), .B1(n20309), .B2(n20308), .ZN(
        n20311) );
  INV_X1 U23282 ( .A(n20311), .ZN(n20315) );
  AOI22_X1 U23283 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20313), .B1(
        n20518), .B2(n20312), .ZN(n20314) );
  OAI211_X1 U23284 ( .C1(n20463), .C2(n20343), .A(n20315), .B(n20314), .ZN(
        P1_U3120) );
  NOR2_X1 U23285 ( .A1(n20317), .A2(n20316), .ZN(n20345) );
  INV_X1 U23286 ( .A(n20471), .ZN(n20318) );
  AOI21_X1 U23287 ( .B1(n20319), .B2(n20318), .A(n20345), .ZN(n20321) );
  OAI22_X1 U23288 ( .A1(n20321), .A2(n20469), .B1(n20320), .B2(n11609), .ZN(
        n20344) );
  AOI22_X1 U23289 ( .A1(n20474), .A2(n20345), .B1(n20344), .B2(n20473), .ZN(
        n20329) );
  OAI21_X1 U23290 ( .B1(n20323), .B2(n20322), .A(n20321), .ZN(n20324) );
  OAI221_X1 U23291 ( .B1(n20398), .B2(n20325), .C1(n20469), .C2(n20324), .A(
        n20476), .ZN(n20347) );
  INV_X1 U23292 ( .A(n20395), .ZN(n20340) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20347), .B1(
        n20340), .B2(n20352), .ZN(n20328) );
  OAI211_X1 U23294 ( .C1(n20364), .C2(n20343), .A(n20329), .B(n20328), .ZN(
        P1_U3121) );
  AOI22_X1 U23295 ( .A1(n20484), .A2(n20345), .B1(n20483), .B2(n20344), .ZN(
        n20331) );
  INV_X1 U23296 ( .A(n20343), .ZN(n20346) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20440), .ZN(n20330) );
  OAI211_X1 U23298 ( .C1(n20443), .C2(n20395), .A(n20331), .B(n20330), .ZN(
        P1_U3122) );
  AOI22_X1 U23299 ( .A1(n20490), .A2(n20345), .B1(n20344), .B2(n20489), .ZN(
        n20333) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20347), .B1(
        n20340), .B2(n20369), .ZN(n20332) );
  OAI211_X1 U23301 ( .C1(n20372), .C2(n20343), .A(n20333), .B(n20332), .ZN(
        P1_U3123) );
  AOI22_X1 U23302 ( .A1(n20496), .A2(n20345), .B1(n20495), .B2(n20344), .ZN(
        n20335) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20347), .B1(
        n20340), .B2(n20373), .ZN(n20334) );
  OAI211_X1 U23304 ( .C1(n20376), .C2(n20343), .A(n20335), .B(n20334), .ZN(
        P1_U3124) );
  AOI22_X1 U23305 ( .A1(n20641), .A2(n20345), .B1(n20640), .B2(n20344), .ZN(
        n20337) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20448), .ZN(n20336) );
  OAI211_X1 U23307 ( .C1(n20451), .C2(n20395), .A(n20337), .B(n20336), .ZN(
        P1_U3125) );
  AOI22_X1 U23308 ( .A1(n20504), .A2(n20345), .B1(n20503), .B2(n20344), .ZN(
        n20339) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20347), .B1(
        n20340), .B2(n20382), .ZN(n20338) );
  OAI211_X1 U23310 ( .C1(n20385), .C2(n20343), .A(n20339), .B(n20338), .ZN(
        P1_U3126) );
  AOI22_X1 U23311 ( .A1(n20510), .A2(n20345), .B1(n20509), .B2(n20344), .ZN(
        n20342) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20347), .B1(
        n20340), .B2(n20386), .ZN(n20341) );
  OAI211_X1 U23313 ( .C1(n20389), .C2(n20343), .A(n20342), .B(n20341), .ZN(
        P1_U3127) );
  AOI22_X1 U23314 ( .A1(n20520), .A2(n20345), .B1(n20518), .B2(n20344), .ZN(
        n20349) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20347), .B1(
        n20346), .B2(n20458), .ZN(n20348) );
  OAI211_X1 U23316 ( .C1(n20463), .C2(n20395), .A(n20349), .B(n20348), .ZN(
        P1_U3128) );
  NAND2_X1 U23317 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20466) );
  OR2_X1 U23318 ( .A1(n20351), .A2(n20466), .ZN(n20379) );
  INV_X1 U23319 ( .A(n20379), .ZN(n20390) );
  AOI22_X1 U23320 ( .A1(n20421), .A2(n20352), .B1(n20474), .B2(n20390), .ZN(
        n20363) );
  NAND2_X1 U23321 ( .A1(n20395), .A2(n20398), .ZN(n20354) );
  OAI21_X1 U23322 ( .B1(n20354), .B2(n20421), .A(n20353), .ZN(n20358) );
  NOR2_X1 U23323 ( .A1(n13102), .A2(n20355), .ZN(n20432) );
  NAND2_X1 U23324 ( .A1(n20432), .A2(n13879), .ZN(n20360) );
  AOI22_X1 U23325 ( .A1(n20358), .A2(n20360), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20359), .ZN(n20356) );
  INV_X1 U23326 ( .A(n20358), .ZN(n20361) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20392), .B1(
        n20473), .B2(n20391), .ZN(n20362) );
  OAI211_X1 U23328 ( .C1(n20364), .C2(n20395), .A(n20363), .B(n20362), .ZN(
        P1_U3129) );
  AOI22_X1 U23329 ( .A1(n20421), .A2(n20485), .B1(n20484), .B2(n20390), .ZN(
        n20366) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20392), .B1(
        n20483), .B2(n20391), .ZN(n20365) );
  OAI211_X1 U23331 ( .C1(n20488), .C2(n20395), .A(n20366), .B(n20365), .ZN(
        P1_U3130) );
  NOR2_X1 U23332 ( .A1(n20367), .A2(n20379), .ZN(n20368) );
  AOI21_X1 U23333 ( .B1(n20421), .B2(n20369), .A(n20368), .ZN(n20371) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20392), .B1(
        n20489), .B2(n20391), .ZN(n20370) );
  OAI211_X1 U23335 ( .C1(n20372), .C2(n20395), .A(n20371), .B(n20370), .ZN(
        P1_U3131) );
  AOI22_X1 U23336 ( .A1(n20421), .A2(n20373), .B1(n20496), .B2(n20390), .ZN(
        n20375) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20392), .B1(
        n20495), .B2(n20391), .ZN(n20374) );
  OAI211_X1 U23338 ( .C1(n20376), .C2(n20395), .A(n20375), .B(n20374), .ZN(
        P1_U3132) );
  AOI22_X1 U23339 ( .A1(n20421), .A2(n20643), .B1(n20641), .B2(n20390), .ZN(
        n20378) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20392), .B1(
        n20640), .B2(n20391), .ZN(n20377) );
  OAI211_X1 U23341 ( .C1(n20645), .C2(n20395), .A(n20378), .B(n20377), .ZN(
        P1_U3133) );
  NOR2_X1 U23342 ( .A1(n20380), .A2(n20379), .ZN(n20381) );
  AOI21_X1 U23343 ( .B1(n20421), .B2(n20382), .A(n20381), .ZN(n20384) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20392), .B1(
        n20503), .B2(n20391), .ZN(n20383) );
  OAI211_X1 U23345 ( .C1(n20385), .C2(n20395), .A(n20384), .B(n20383), .ZN(
        P1_U3134) );
  AOI22_X1 U23346 ( .A1(n20421), .A2(n20386), .B1(n20510), .B2(n20390), .ZN(
        n20388) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20392), .B1(
        n20509), .B2(n20391), .ZN(n20387) );
  OAI211_X1 U23348 ( .C1(n20389), .C2(n20395), .A(n20388), .B(n20387), .ZN(
        P1_U3135) );
  AOI22_X1 U23349 ( .A1(n20421), .A2(n20521), .B1(n20520), .B2(n20390), .ZN(
        n20394) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20392), .B1(
        n20518), .B2(n20391), .ZN(n20393) );
  OAI211_X1 U23351 ( .C1(n20527), .C2(n20395), .A(n20394), .B(n20393), .ZN(
        P1_U3136) );
  NOR3_X2 U23352 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20397), .A3(
        n20466), .ZN(n20420) );
  INV_X1 U23353 ( .A(n20420), .ZN(n20401) );
  NOR2_X1 U23354 ( .A1(n20466), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20403) );
  INV_X1 U23355 ( .A(n20403), .ZN(n20400) );
  NAND2_X1 U23356 ( .A1(n20432), .A2(n20398), .ZN(n20472) );
  OAI222_X1 U23357 ( .A1(n20401), .A2(n20469), .B1(n11609), .B2(n20400), .C1(
        n20399), .C2(n20472), .ZN(n20419) );
  AOI22_X1 U23358 ( .A1(n20474), .A2(n20420), .B1(n20473), .B2(n20419), .ZN(
        n20406) );
  NOR3_X1 U23359 ( .A1(n20402), .A2(n20429), .A3(n20469), .ZN(n20404) );
  OAI21_X1 U23360 ( .B1(n20404), .B2(n20403), .A(n20476), .ZN(n20422) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20479), .ZN(n20405) );
  OAI211_X1 U23362 ( .C1(n20482), .C2(n20437), .A(n20406), .B(n20405), .ZN(
        P1_U3137) );
  AOI22_X1 U23363 ( .A1(n20484), .A2(n20420), .B1(n20483), .B2(n20419), .ZN(
        n20408) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20440), .ZN(n20407) );
  OAI211_X1 U23365 ( .C1(n20443), .C2(n20437), .A(n20408), .B(n20407), .ZN(
        P1_U3138) );
  AOI22_X1 U23366 ( .A1(n20490), .A2(n20420), .B1(n20489), .B2(n20419), .ZN(
        n20410) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20491), .ZN(n20409) );
  OAI211_X1 U23368 ( .C1(n20494), .C2(n20437), .A(n20410), .B(n20409), .ZN(
        P1_U3139) );
  AOI22_X1 U23369 ( .A1(n20496), .A2(n20420), .B1(n20495), .B2(n20419), .ZN(
        n20412) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20497), .ZN(n20411) );
  OAI211_X1 U23371 ( .C1(n20500), .C2(n20437), .A(n20412), .B(n20411), .ZN(
        P1_U3140) );
  AOI22_X1 U23372 ( .A1(n20641), .A2(n20420), .B1(n20640), .B2(n20419), .ZN(
        n20414) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20448), .ZN(n20413) );
  OAI211_X1 U23374 ( .C1(n20451), .C2(n20437), .A(n20414), .B(n20413), .ZN(
        P1_U3141) );
  AOI22_X1 U23375 ( .A1(n20504), .A2(n20420), .B1(n20503), .B2(n20419), .ZN(
        n20416) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20505), .ZN(n20415) );
  OAI211_X1 U23377 ( .C1(n20508), .C2(n20437), .A(n20416), .B(n20415), .ZN(
        P1_U3142) );
  AOI22_X1 U23378 ( .A1(n20510), .A2(n20420), .B1(n20509), .B2(n20419), .ZN(
        n20418) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20511), .ZN(n20417) );
  OAI211_X1 U23380 ( .C1(n20516), .C2(n20437), .A(n20418), .B(n20417), .ZN(
        P1_U3143) );
  AOI22_X1 U23381 ( .A1(n20520), .A2(n20420), .B1(n20518), .B2(n20419), .ZN(
        n20424) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20422), .B1(
        n20421), .B2(n20458), .ZN(n20423) );
  OAI211_X1 U23383 ( .C1(n20463), .C2(n20437), .A(n20424), .B(n20423), .ZN(
        P1_U3144) );
  NOR3_X2 U23384 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20467), .A3(
        n20466), .ZN(n20457) );
  OAI22_X1 U23385 ( .A1(n20472), .A2(n13879), .B1(n20428), .B2(n20427), .ZN(
        n20456) );
  AOI22_X1 U23386 ( .A1(n20474), .A2(n20457), .B1(n20473), .B2(n20456), .ZN(
        n20439) );
  AOI21_X1 U23387 ( .B1(n20526), .B2(n20437), .A(n20429), .ZN(n20430) );
  AOI21_X1 U23388 ( .B1(n20432), .B2(n20431), .A(n20430), .ZN(n20433) );
  NOR2_X1 U23389 ( .A1(n20433), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20436) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20460), .B1(
        n20459), .B2(n20479), .ZN(n20438) );
  OAI211_X1 U23391 ( .C1(n20482), .C2(n20526), .A(n20439), .B(n20438), .ZN(
        P1_U3145) );
  AOI22_X1 U23392 ( .A1(n20484), .A2(n20457), .B1(n20483), .B2(n20456), .ZN(
        n20442) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20460), .B1(
        n20459), .B2(n20440), .ZN(n20441) );
  OAI211_X1 U23394 ( .C1(n20443), .C2(n20526), .A(n20442), .B(n20441), .ZN(
        P1_U3146) );
  AOI22_X1 U23395 ( .A1(n20490), .A2(n20457), .B1(n20489), .B2(n20456), .ZN(
        n20445) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20460), .B1(
        n20459), .B2(n20491), .ZN(n20444) );
  OAI211_X1 U23397 ( .C1(n20494), .C2(n20526), .A(n20445), .B(n20444), .ZN(
        P1_U3147) );
  AOI22_X1 U23398 ( .A1(n20496), .A2(n20457), .B1(n20495), .B2(n20456), .ZN(
        n20447) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20460), .B1(
        n20459), .B2(n20497), .ZN(n20446) );
  OAI211_X1 U23400 ( .C1(n20500), .C2(n20526), .A(n20447), .B(n20446), .ZN(
        P1_U3148) );
  AOI22_X1 U23401 ( .A1(n20641), .A2(n20457), .B1(n20640), .B2(n20456), .ZN(
        n20450) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20460), .B1(
        n20459), .B2(n20448), .ZN(n20449) );
  OAI211_X1 U23403 ( .C1(n20451), .C2(n20526), .A(n20450), .B(n20449), .ZN(
        P1_U3149) );
  AOI22_X1 U23404 ( .A1(n20504), .A2(n20457), .B1(n20503), .B2(n20456), .ZN(
        n20453) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20460), .B1(
        n20459), .B2(n20505), .ZN(n20452) );
  OAI211_X1 U23406 ( .C1(n20508), .C2(n20526), .A(n20453), .B(n20452), .ZN(
        P1_U3150) );
  AOI22_X1 U23407 ( .A1(n20510), .A2(n20457), .B1(n20509), .B2(n20456), .ZN(
        n20455) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20460), .B1(
        n20459), .B2(n20511), .ZN(n20454) );
  OAI211_X1 U23409 ( .C1(n20516), .C2(n20526), .A(n20455), .B(n20454), .ZN(
        P1_U3151) );
  AOI22_X1 U23410 ( .A1(n20520), .A2(n20457), .B1(n20518), .B2(n20456), .ZN(
        n20462) );
  AOI22_X1 U23411 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20460), .B1(
        n20459), .B2(n20458), .ZN(n20461) );
  OAI211_X1 U23412 ( .C1(n20463), .C2(n20526), .A(n20462), .B(n20461), .ZN(
        P1_U3152) );
  INV_X1 U23413 ( .A(n20466), .ZN(n20464) );
  NAND2_X1 U23414 ( .A1(n20465), .A2(n20464), .ZN(n20468) );
  INV_X1 U23415 ( .A(n20468), .ZN(n20519) );
  NOR2_X1 U23416 ( .A1(n20467), .A2(n20466), .ZN(n20477) );
  INV_X1 U23417 ( .A(n20477), .ZN(n20470) );
  OAI222_X1 U23418 ( .A1(n20472), .A2(n20471), .B1(n11609), .B2(n20470), .C1(
        n20469), .C2(n20468), .ZN(n20517) );
  AOI22_X1 U23419 ( .A1(n20474), .A2(n20519), .B1(n20473), .B2(n20517), .ZN(
        n20481) );
  NOR2_X1 U23420 ( .A1(n20475), .A2(n13137), .ZN(n20478) );
  OAI21_X1 U23421 ( .B1(n20478), .B2(n20477), .A(n20476), .ZN(n20523) );
  INV_X1 U23422 ( .A(n20526), .ZN(n20512) );
  AOI22_X1 U23423 ( .A1(n20523), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n20512), .B2(n20479), .ZN(n20480) );
  OAI211_X1 U23424 ( .C1(n20482), .C2(n20515), .A(n20481), .B(n20480), .ZN(
        P1_U3153) );
  AOI22_X1 U23425 ( .A1(n20484), .A2(n20519), .B1(n20483), .B2(n20517), .ZN(
        n20487) );
  AOI22_X1 U23426 ( .A1(n20523), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n20522), .B2(n20485), .ZN(n20486) );
  OAI211_X1 U23427 ( .C1(n20488), .C2(n20526), .A(n20487), .B(n20486), .ZN(
        P1_U3154) );
  AOI22_X1 U23428 ( .A1(n20490), .A2(n20519), .B1(n20489), .B2(n20517), .ZN(
        n20493) );
  AOI22_X1 U23429 ( .A1(n20523), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n20512), .B2(n20491), .ZN(n20492) );
  OAI211_X1 U23430 ( .C1(n20494), .C2(n20515), .A(n20493), .B(n20492), .ZN(
        P1_U3155) );
  AOI22_X1 U23431 ( .A1(n20496), .A2(n20519), .B1(n20495), .B2(n20517), .ZN(
        n20499) );
  AOI22_X1 U23432 ( .A1(n20523), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n20512), .B2(n20497), .ZN(n20498) );
  OAI211_X1 U23433 ( .C1(n20500), .C2(n20515), .A(n20499), .B(n20498), .ZN(
        P1_U3156) );
  AOI22_X1 U23434 ( .A1(n20641), .A2(n20519), .B1(n20640), .B2(n20517), .ZN(
        n20502) );
  AOI22_X1 U23435 ( .A1(n20523), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n20522), .B2(n20643), .ZN(n20501) );
  OAI211_X1 U23436 ( .C1(n20645), .C2(n20526), .A(n20502), .B(n20501), .ZN(
        P1_U3157) );
  AOI22_X1 U23437 ( .A1(n20504), .A2(n20519), .B1(n20503), .B2(n20517), .ZN(
        n20507) );
  AOI22_X1 U23438 ( .A1(n20523), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n20512), .B2(n20505), .ZN(n20506) );
  OAI211_X1 U23439 ( .C1(n20508), .C2(n20515), .A(n20507), .B(n20506), .ZN(
        P1_U3158) );
  AOI22_X1 U23440 ( .A1(n20510), .A2(n20519), .B1(n20509), .B2(n20517), .ZN(
        n20514) );
  AOI22_X1 U23441 ( .A1(n20523), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n20512), .B2(n20511), .ZN(n20513) );
  OAI211_X1 U23442 ( .C1(n20516), .C2(n20515), .A(n20514), .B(n20513), .ZN(
        P1_U3159) );
  AOI22_X1 U23443 ( .A1(n20520), .A2(n20519), .B1(n20518), .B2(n20517), .ZN(
        n20525) );
  AOI22_X1 U23444 ( .A1(n20523), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n20522), .B2(n20521), .ZN(n20524) );
  OAI211_X1 U23445 ( .C1(n20527), .C2(n20526), .A(n20525), .B(n20524), .ZN(
        P1_U3160) );
  OR2_X1 U23446 ( .A1(n20529), .A2(n20528), .ZN(P1_U3163) );
  AND2_X1 U23447 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20530), .ZN(
        P1_U3164) );
  AND2_X1 U23448 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20530), .ZN(
        P1_U3165) );
  AND2_X1 U23449 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20530), .ZN(
        P1_U3166) );
  AND2_X1 U23450 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20530), .ZN(
        P1_U3167) );
  AND2_X1 U23451 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20530), .ZN(
        P1_U3168) );
  AND2_X1 U23452 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20530), .ZN(
        P1_U3169) );
  AND2_X1 U23453 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20530), .ZN(
        P1_U3170) );
  AND2_X1 U23454 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20530), .ZN(
        P1_U3171) );
  AND2_X1 U23455 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20530), .ZN(
        P1_U3172) );
  AND2_X1 U23456 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20530), .ZN(
        P1_U3173) );
  AND2_X1 U23457 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20530), .ZN(
        P1_U3174) );
  AND2_X1 U23458 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20530), .ZN(
        P1_U3175) );
  AND2_X1 U23459 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20530), .ZN(
        P1_U3176) );
  AND2_X1 U23460 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20530), .ZN(
        P1_U3177) );
  AND2_X1 U23461 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20530), .ZN(
        P1_U3178) );
  AND2_X1 U23462 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20530), .ZN(
        P1_U3179) );
  AND2_X1 U23463 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20530), .ZN(
        P1_U3180) );
  AND2_X1 U23464 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20530), .ZN(
        P1_U3181) );
  AND2_X1 U23465 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20530), .ZN(
        P1_U3182) );
  AND2_X1 U23466 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20530), .ZN(
        P1_U3183) );
  AND2_X1 U23467 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20530), .ZN(
        P1_U3184) );
  AND2_X1 U23468 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20530), .ZN(
        P1_U3185) );
  AND2_X1 U23469 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20530), .ZN(P1_U3186) );
  AND2_X1 U23470 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20530), .ZN(P1_U3187) );
  AND2_X1 U23471 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20530), .ZN(P1_U3188) );
  AND2_X1 U23472 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20530), .ZN(P1_U3189) );
  AND2_X1 U23473 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20530), .ZN(P1_U3190) );
  INV_X1 U23474 ( .A(P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20720) );
  NOR2_X1 U23475 ( .A1(n20606), .A2(n20720), .ZN(P1_U3191) );
  AND2_X1 U23476 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20530), .ZN(P1_U3192) );
  AND2_X1 U23477 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20530), .ZN(P1_U3193) );
  INV_X1 U23478 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20536) );
  AOI211_X1 U23479 ( .C1(NA), .C2(n12697), .A(n20531), .B(n20536), .ZN(n20535)
         );
  INV_X1 U23480 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20545) );
  OAI21_X1 U23481 ( .B1(n20532), .B2(n20623), .A(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20539) );
  NAND2_X1 U23482 ( .A1(n20545), .A2(n20539), .ZN(n20533) );
  OAI221_X1 U23483 ( .B1(n20637), .B2(n20535), .C1(n20637), .C2(n20534), .A(
        n20533), .ZN(P1_U3194) );
  OAI211_X1 U23484 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20536), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20544) );
  NAND2_X1 U23485 ( .A1(n20631), .A2(n20540), .ZN(n20542) );
  OAI21_X1 U23486 ( .B1(n20542), .B2(n20537), .A(n20545), .ZN(n20538) );
  OAI211_X1 U23487 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20540), .A(n20539), 
        .B(n20538), .ZN(n20541) );
  OAI221_X1 U23488 ( .B1(n20544), .B2(n20543), .C1(n20544), .C2(n20542), .A(
        n20541), .ZN(P1_U3196) );
  OAI222_X1 U23489 ( .A1(n20594), .A2(n20547), .B1(n20546), .B2(n20637), .C1(
        n20548), .C2(n20598), .ZN(P1_U3197) );
  INV_X1 U23490 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20549) );
  OAI222_X1 U23491 ( .A1(n20598), .A2(n20550), .B1(n20549), .B2(n20637), .C1(
        n20548), .C2(n20594), .ZN(P1_U3198) );
  INV_X1 U23492 ( .A(n20594), .ZN(n20596) );
  AOI222_X1 U23493 ( .A1(n20596), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20634), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20592), .ZN(n20551) );
  INV_X1 U23494 ( .A(n20551), .ZN(P1_U3199) );
  AOI222_X1 U23495 ( .A1(n20596), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20634), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20592), .ZN(n20552) );
  INV_X1 U23496 ( .A(n20552), .ZN(P1_U3200) );
  INV_X1 U23497 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20553) );
  OAI222_X1 U23498 ( .A1(n20594), .A2(n20554), .B1(n20553), .B2(n20637), .C1(
        n20556), .C2(n20598), .ZN(P1_U3201) );
  AOI22_X1 U23499 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20592), .ZN(n20555) );
  OAI21_X1 U23500 ( .B1(n20556), .B2(n20594), .A(n20555), .ZN(P1_U3202) );
  AOI22_X1 U23501 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20596), .ZN(n20557) );
  OAI21_X1 U23502 ( .B1(n20559), .B2(n20598), .A(n20557), .ZN(P1_U3203) );
  AOI22_X1 U23503 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20592), .ZN(n20558) );
  OAI21_X1 U23504 ( .B1(n20559), .B2(n20594), .A(n20558), .ZN(P1_U3204) );
  AOI22_X1 U23505 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20596), .ZN(n20560) );
  OAI21_X1 U23506 ( .B1(n20561), .B2(n20598), .A(n20560), .ZN(P1_U3205) );
  INV_X1 U23507 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20562) );
  OAI222_X1 U23508 ( .A1(n20598), .A2(n20563), .B1(n20562), .B2(n20637), .C1(
        n20561), .C2(n20594), .ZN(P1_U3206) );
  AOI222_X1 U23509 ( .A1(n20596), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20634), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20592), .ZN(n20564) );
  INV_X1 U23510 ( .A(n20564), .ZN(P1_U3207) );
  AOI222_X1 U23511 ( .A1(n20596), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20634), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20592), .ZN(n20565) );
  INV_X1 U23512 ( .A(n20565), .ZN(P1_U3208) );
  INV_X1 U23513 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20566) );
  OAI222_X1 U23514 ( .A1(n20594), .A2(n20567), .B1(n20566), .B2(n20637), .C1(
        n20568), .C2(n20598), .ZN(P1_U3209) );
  INV_X1 U23515 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20569) );
  OAI222_X1 U23516 ( .A1(n20598), .A2(n20571), .B1(n20569), .B2(n20637), .C1(
        n20568), .C2(n20594), .ZN(P1_U3210) );
  INV_X1 U23517 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20570) );
  OAI222_X1 U23518 ( .A1(n20594), .A2(n20571), .B1(n20570), .B2(n20637), .C1(
        n20573), .C2(n20598), .ZN(P1_U3211) );
  AOI22_X1 U23519 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20592), .ZN(n20572) );
  OAI21_X1 U23520 ( .B1(n20573), .B2(n20594), .A(n20572), .ZN(P1_U3212) );
  AOI22_X1 U23521 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20596), .ZN(n20574) );
  OAI21_X1 U23522 ( .B1(n14420), .B2(n20598), .A(n20574), .ZN(P1_U3213) );
  AOI22_X1 U23523 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20592), .ZN(n20575) );
  OAI21_X1 U23524 ( .B1(n14420), .B2(n20594), .A(n20575), .ZN(P1_U3214) );
  AOI22_X1 U23525 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20596), .ZN(n20576) );
  OAI21_X1 U23526 ( .B1(n20577), .B2(n20598), .A(n20576), .ZN(P1_U3215) );
  INV_X1 U23527 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20580) );
  INV_X1 U23528 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20578) );
  OAI222_X1 U23529 ( .A1(n20598), .A2(n20580), .B1(n20578), .B2(n20637), .C1(
        n20577), .C2(n20594), .ZN(P1_U3216) );
  INV_X1 U23530 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20579) );
  INV_X1 U23531 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20582) );
  OAI222_X1 U23532 ( .A1(n20594), .A2(n20580), .B1(n20579), .B2(n20637), .C1(
        n20582), .C2(n20598), .ZN(P1_U3217) );
  INV_X1 U23533 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20581) );
  OAI222_X1 U23534 ( .A1(n20594), .A2(n20582), .B1(n20581), .B2(n20637), .C1(
        n20583), .C2(n20598), .ZN(P1_U3218) );
  INV_X1 U23535 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20584) );
  OAI222_X1 U23536 ( .A1(n20598), .A2(n20586), .B1(n20584), .B2(n20637), .C1(
        n20583), .C2(n20594), .ZN(P1_U3219) );
  AOI22_X1 U23537 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n20592), .ZN(n20585) );
  OAI21_X1 U23538 ( .B1(n20586), .B2(n20594), .A(n20585), .ZN(P1_U3220) );
  INV_X1 U23539 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20587) );
  INV_X1 U23540 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20717) );
  OAI222_X1 U23541 ( .A1(n20594), .A2(n20587), .B1(n20717), .B2(n20637), .C1(
        n20588), .C2(n20598), .ZN(P1_U3221) );
  INV_X1 U23542 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20589) );
  OAI222_X1 U23543 ( .A1(n20598), .A2(n14024), .B1(n20589), .B2(n20637), .C1(
        n20588), .C2(n20594), .ZN(P1_U3222) );
  AOI22_X1 U23544 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(n20592), .ZN(n20590) );
  OAI21_X1 U23545 ( .B1(n14024), .B2(n20594), .A(n20590), .ZN(P1_U3223) );
  AOI22_X1 U23546 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(n20596), .ZN(n20591) );
  OAI21_X1 U23547 ( .B1(n20595), .B2(n20598), .A(n20591), .ZN(P1_U3224) );
  AOI22_X1 U23548 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n20592), .ZN(n20593) );
  OAI21_X1 U23549 ( .B1(n20595), .B2(n20594), .A(n20593), .ZN(P1_U3225) );
  AOI22_X1 U23550 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n20634), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n20596), .ZN(n20597) );
  OAI21_X1 U23551 ( .B1(n20599), .B2(n20598), .A(n20597), .ZN(P1_U3226) );
  MUX2_X1 U23552 ( .A(P1_BE_N_REG_3__SCAN_IN), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .S(n20637), .Z(P1_U3458) );
  MUX2_X1 U23553 ( .A(P1_BE_N_REG_2__SCAN_IN), .B(P1_BYTEENABLE_REG_2__SCAN_IN), .S(n20637), .Z(P1_U3459) );
  INV_X1 U23554 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20600) );
  AOI22_X1 U23555 ( .A1(n20637), .A2(n20601), .B1(n20600), .B2(n20634), .ZN(
        P1_U3460) );
  INV_X1 U23556 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20619) );
  INV_X1 U23557 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20602) );
  AOI22_X1 U23558 ( .A1(n20637), .A2(n20619), .B1(n20602), .B2(n20634), .ZN(
        P1_U3461) );
  OAI21_X1 U23559 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20606), .A(n20604), 
        .ZN(n20603) );
  INV_X1 U23560 ( .A(n20603), .ZN(P1_U3464) );
  INV_X1 U23561 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20605) );
  OAI21_X1 U23562 ( .B1(n20606), .B2(n20605), .A(n20604), .ZN(P1_U3465) );
  INV_X1 U23563 ( .A(n20607), .ZN(n20612) );
  INV_X1 U23564 ( .A(n20608), .ZN(n20610) );
  OAI22_X1 U23565 ( .A1(n20612), .A2(n20611), .B1(n20610), .B2(n20609), .ZN(
        n20614) );
  MUX2_X1 U23566 ( .A(n20614), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20613), .Z(P1_U3469) );
  AOI211_X1 U23567 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20615) );
  INV_X1 U23568 ( .A(n20621), .ZN(n20618) );
  AOI22_X1 U23569 ( .A1(n20621), .A2(n20615), .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n20618), .ZN(n20616) );
  OAI21_X1 U23570 ( .B1(n12944), .B2(n20617), .A(n20616), .ZN(P1_U3481) );
  NOR2_X1 U23571 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20620) );
  AOI22_X1 U23572 ( .A1(n20621), .A2(n20620), .B1(n20619), .B2(n20618), .ZN(
        P1_U3482) );
  AOI22_X1 U23573 ( .A1(n20637), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20622), 
        .B2(n20634), .ZN(P1_U3483) );
  OAI211_X1 U23574 ( .C1(n12756), .C2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .B(n20623), .ZN(n20624) );
  OAI21_X1 U23575 ( .B1(n20625), .B2(n20624), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n20627) );
  NAND2_X1 U23576 ( .A1(n20627), .A2(n20626), .ZN(n20633) );
  OAI211_X1 U23577 ( .C1(n20631), .C2(n20630), .A(n20629), .B(n20628), .ZN(
        n20632) );
  MUX2_X1 U23578 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(n20633), .S(n20632), 
        .Z(P1_U3485) );
  INV_X1 U23579 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20635) );
  AOI22_X1 U23580 ( .A1(n20637), .A2(n20636), .B1(n20635), .B2(n20634), .ZN(
        P1_U3486) );
  NAND2_X1 U23581 ( .A1(n20638), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n20650) );
  AOI22_X1 U23582 ( .A1(n20642), .A2(n20641), .B1(n20640), .B2(n20639), .ZN(
        n20649) );
  NAND2_X1 U23583 ( .A1(n20644), .A2(n20643), .ZN(n20648) );
  OR2_X1 U23584 ( .A1(n20646), .A2(n20645), .ZN(n20647) );
  AND4_X1 U23585 ( .A1(n20650), .A2(n20649), .A3(n20648), .A4(n20647), .ZN(
        n20808) );
  AOI22_X1 U23586 ( .A1(n20653), .A2(keyinput1), .B1(n20652), .B2(keyinput15), 
        .ZN(n20651) );
  OAI221_X1 U23587 ( .B1(n20653), .B2(keyinput1), .C1(n20652), .C2(keyinput15), 
        .A(n20651), .ZN(n20666) );
  INV_X1 U23588 ( .A(P3_LWORD_REG_1__SCAN_IN), .ZN(n20655) );
  AOI22_X1 U23589 ( .A1(n20656), .A2(keyinput18), .B1(keyinput13), .B2(n20655), 
        .ZN(n20654) );
  OAI221_X1 U23590 ( .B1(n20656), .B2(keyinput18), .C1(n20655), .C2(keyinput13), .A(n20654), .ZN(n20665) );
  AOI22_X1 U23591 ( .A1(n20659), .A2(keyinput14), .B1(keyinput40), .B2(n20658), 
        .ZN(n20657) );
  OAI221_X1 U23592 ( .B1(n20659), .B2(keyinput14), .C1(n20658), .C2(keyinput40), .A(n20657), .ZN(n20664) );
  INV_X1 U23593 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20661) );
  AOI22_X1 U23594 ( .A1(n20662), .A2(keyinput35), .B1(n20661), .B2(keyinput28), 
        .ZN(n20660) );
  OAI221_X1 U23595 ( .B1(n20662), .B2(keyinput35), .C1(n20661), .C2(keyinput28), .A(n20660), .ZN(n20663) );
  NOR4_X1 U23596 ( .A1(n20666), .A2(n20665), .A3(n20664), .A4(n20663), .ZN(
        n20715) );
  INV_X1 U23597 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20669) );
  AOI22_X1 U23598 ( .A1(n20669), .A2(keyinput34), .B1(n20668), .B2(keyinput50), 
        .ZN(n20667) );
  OAI221_X1 U23599 ( .B1(n20669), .B2(keyinput34), .C1(n20668), .C2(keyinput50), .A(n20667), .ZN(n20682) );
  AOI22_X1 U23600 ( .A1(n20672), .A2(keyinput11), .B1(n20671), .B2(keyinput21), 
        .ZN(n20670) );
  OAI221_X1 U23601 ( .B1(n20672), .B2(keyinput11), .C1(n20671), .C2(keyinput21), .A(n20670), .ZN(n20681) );
  INV_X1 U23602 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n20675) );
  AOI22_X1 U23603 ( .A1(n20675), .A2(keyinput58), .B1(keyinput48), .B2(n20674), 
        .ZN(n20673) );
  OAI221_X1 U23604 ( .B1(n20675), .B2(keyinput58), .C1(n20674), .C2(keyinput48), .A(n20673), .ZN(n20680) );
  AOI22_X1 U23605 ( .A1(n20678), .A2(keyinput25), .B1(keyinput47), .B2(n20677), 
        .ZN(n20676) );
  OAI221_X1 U23606 ( .B1(n20678), .B2(keyinput25), .C1(n20677), .C2(keyinput47), .A(n20676), .ZN(n20679) );
  NOR4_X1 U23607 ( .A1(n20682), .A2(n20681), .A3(n20680), .A4(n20679), .ZN(
        n20714) );
  AOI22_X1 U23608 ( .A1(n20685), .A2(keyinput22), .B1(n20684), .B2(keyinput23), 
        .ZN(n20683) );
  OAI221_X1 U23609 ( .B1(n20685), .B2(keyinput22), .C1(n20684), .C2(keyinput23), .A(n20683), .ZN(n20695) );
  AOI22_X1 U23610 ( .A1(n10726), .A2(keyinput43), .B1(keyinput57), .B2(n10276), 
        .ZN(n20686) );
  OAI221_X1 U23611 ( .B1(n10726), .B2(keyinput43), .C1(n10276), .C2(keyinput57), .A(n20686), .ZN(n20694) );
  AOI22_X1 U23612 ( .A1(n10635), .A2(keyinput49), .B1(keyinput42), .B2(n20688), 
        .ZN(n20687) );
  OAI221_X1 U23613 ( .B1(n10635), .B2(keyinput49), .C1(n20688), .C2(keyinput42), .A(n20687), .ZN(n20693) );
  INV_X1 U23614 ( .A(READY2), .ZN(n20691) );
  AOI22_X1 U23615 ( .A1(n20691), .A2(keyinput36), .B1(n20690), .B2(keyinput60), 
        .ZN(n20689) );
  OAI221_X1 U23616 ( .B1(n20691), .B2(keyinput36), .C1(n20690), .C2(keyinput60), .A(n20689), .ZN(n20692) );
  NOR4_X1 U23617 ( .A1(n20695), .A2(n20694), .A3(n20693), .A4(n20692), .ZN(
        n20713) );
  AOI22_X1 U23618 ( .A1(n20698), .A2(keyinput12), .B1(n20697), .B2(keyinput51), 
        .ZN(n20696) );
  OAI221_X1 U23619 ( .B1(n20698), .B2(keyinput12), .C1(n20697), .C2(keyinput51), .A(n20696), .ZN(n20702) );
  XNOR2_X1 U23620 ( .A(n20699), .B(keyinput33), .ZN(n20701) );
  XOR2_X1 U23621 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B(keyinput17), .Z(
        n20700) );
  OR3_X1 U23622 ( .A1(n20702), .A2(n20701), .A3(n20700), .ZN(n20711) );
  AOI22_X1 U23623 ( .A1(n20705), .A2(keyinput63), .B1(n20704), .B2(keyinput27), 
        .ZN(n20703) );
  OAI221_X1 U23624 ( .B1(n20705), .B2(keyinput63), .C1(n20704), .C2(keyinput27), .A(n20703), .ZN(n20710) );
  INV_X1 U23625 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n20707) );
  AOI22_X1 U23626 ( .A1(n20708), .A2(keyinput3), .B1(keyinput20), .B2(n20707), 
        .ZN(n20706) );
  OAI221_X1 U23627 ( .B1(n20708), .B2(keyinput3), .C1(n20707), .C2(keyinput20), 
        .A(n20706), .ZN(n20709) );
  NOR3_X1 U23628 ( .A1(n20711), .A2(n20710), .A3(n20709), .ZN(n20712) );
  NAND4_X1 U23629 ( .A1(n20715), .A2(n20714), .A3(n20713), .A4(n20712), .ZN(
        n20782) );
  AOI22_X1 U23630 ( .A1(n20718), .A2(keyinput16), .B1(n20717), .B2(keyinput0), 
        .ZN(n20716) );
  OAI221_X1 U23631 ( .B1(n20718), .B2(keyinput16), .C1(n20717), .C2(keyinput0), 
        .A(n20716), .ZN(n20730) );
  AOI22_X1 U23632 ( .A1(n20790), .A2(keyinput59), .B1(keyinput53), .B2(n20720), 
        .ZN(n20719) );
  OAI221_X1 U23633 ( .B1(n20790), .B2(keyinput59), .C1(n20720), .C2(keyinput53), .A(n20719), .ZN(n20729) );
  AOI22_X1 U23634 ( .A1(n20723), .A2(keyinput55), .B1(keyinput30), .B2(n20722), 
        .ZN(n20721) );
  OAI221_X1 U23635 ( .B1(n20723), .B2(keyinput55), .C1(n20722), .C2(keyinput30), .A(n20721), .ZN(n20728) );
  AOI22_X1 U23636 ( .A1(n20726), .A2(keyinput5), .B1(n20725), .B2(keyinput54), 
        .ZN(n20724) );
  OAI221_X1 U23637 ( .B1(n20726), .B2(keyinput5), .C1(n20725), .C2(keyinput54), 
        .A(n20724), .ZN(n20727) );
  NOR4_X1 U23638 ( .A1(n20730), .A2(n20729), .A3(n20728), .A4(n20727), .ZN(
        n20780) );
  AOI22_X1 U23639 ( .A1(n20733), .A2(keyinput19), .B1(keyinput61), .B2(n20732), 
        .ZN(n20731) );
  OAI221_X1 U23640 ( .B1(n20733), .B2(keyinput19), .C1(n20732), .C2(keyinput61), .A(n20731), .ZN(n20745) );
  AOI22_X1 U23641 ( .A1(n10562), .A2(keyinput37), .B1(keyinput29), .B2(n20735), 
        .ZN(n20734) );
  OAI221_X1 U23642 ( .B1(n10562), .B2(keyinput37), .C1(n20735), .C2(keyinput29), .A(n20734), .ZN(n20744) );
  INV_X1 U23643 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20738) );
  AOI22_X1 U23644 ( .A1(n20738), .A2(keyinput8), .B1(n20737), .B2(keyinput7), 
        .ZN(n20736) );
  OAI221_X1 U23645 ( .B1(n20738), .B2(keyinput8), .C1(n20737), .C2(keyinput7), 
        .A(n20736), .ZN(n20743) );
  XOR2_X1 U23646 ( .A(n20739), .B(keyinput9), .Z(n20741) );
  XNOR2_X1 U23647 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput46), 
        .ZN(n20740) );
  NAND2_X1 U23648 ( .A1(n20741), .A2(n20740), .ZN(n20742) );
  NOR4_X1 U23649 ( .A1(n20745), .A2(n20744), .A3(n20743), .A4(n20742), .ZN(
        n20779) );
  AOI22_X1 U23650 ( .A1(n20747), .A2(keyinput31), .B1(n9834), .B2(keyinput24), 
        .ZN(n20746) );
  OAI221_X1 U23651 ( .B1(n20747), .B2(keyinput31), .C1(n9834), .C2(keyinput24), 
        .A(n20746), .ZN(n20760) );
  INV_X1 U23652 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n20749) );
  AOI22_X1 U23653 ( .A1(n20750), .A2(keyinput41), .B1(keyinput10), .B2(n20749), 
        .ZN(n20748) );
  OAI221_X1 U23654 ( .B1(n20750), .B2(keyinput41), .C1(n20749), .C2(keyinput10), .A(n20748), .ZN(n20759) );
  AOI22_X1 U23655 ( .A1(n20753), .A2(keyinput56), .B1(n20752), .B2(keyinput26), 
        .ZN(n20751) );
  OAI221_X1 U23656 ( .B1(n20753), .B2(keyinput56), .C1(n20752), .C2(keyinput26), .A(n20751), .ZN(n20758) );
  AOI22_X1 U23657 ( .A1(n20756), .A2(keyinput62), .B1(keyinput39), .B2(n20755), 
        .ZN(n20754) );
  OAI221_X1 U23658 ( .B1(n20756), .B2(keyinput62), .C1(n20755), .C2(keyinput39), .A(n20754), .ZN(n20757) );
  NOR4_X1 U23659 ( .A1(n20760), .A2(n20759), .A3(n20758), .A4(n20757), .ZN(
        n20778) );
  AOI22_X1 U23660 ( .A1(n20763), .A2(keyinput32), .B1(keyinput45), .B2(n20762), 
        .ZN(n20761) );
  OAI221_X1 U23661 ( .B1(n20763), .B2(keyinput32), .C1(n20762), .C2(keyinput45), .A(n20761), .ZN(n20776) );
  AOI22_X1 U23662 ( .A1(n20766), .A2(keyinput2), .B1(keyinput44), .B2(n20765), 
        .ZN(n20764) );
  OAI221_X1 U23663 ( .B1(n20766), .B2(keyinput2), .C1(n20765), .C2(keyinput44), 
        .A(n20764), .ZN(n20775) );
  AOI22_X1 U23664 ( .A1(n20769), .A2(keyinput38), .B1(keyinput4), .B2(n20768), 
        .ZN(n20767) );
  OAI221_X1 U23665 ( .B1(n20769), .B2(keyinput38), .C1(n20768), .C2(keyinput4), 
        .A(n20767), .ZN(n20774) );
  INV_X1 U23666 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n20772) );
  AOI22_X1 U23667 ( .A1(n20772), .A2(keyinput6), .B1(keyinput52), .B2(n20771), 
        .ZN(n20770) );
  OAI221_X1 U23668 ( .B1(n20772), .B2(keyinput6), .C1(n20771), .C2(keyinput52), 
        .A(n20770), .ZN(n20773) );
  NOR4_X1 U23669 ( .A1(n20776), .A2(n20775), .A3(n20774), .A4(n20773), .ZN(
        n20777) );
  NAND4_X1 U23670 ( .A1(n20780), .A2(n20779), .A3(n20778), .A4(n20777), .ZN(
        n20781) );
  NOR2_X1 U23671 ( .A1(n20782), .A2(n20781), .ZN(n20806) );
  NOR4_X1 U23672 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(P1_EAX_REG_29__SCAN_IN), .A4(
        P1_EBX_REG_22__SCAN_IN), .ZN(n20804) );
  NAND4_X1 U23673 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_DATAO_REG_12__SCAN_IN), .A3(P3_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_BE_N_REG_0__SCAN_IN), .ZN(n20785) );
  NAND4_X1 U23674 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P2_DATAO_REG_14__SCAN_IN), .A4(P1_UWORD_REG_10__SCAN_IN), .ZN(
        n20784) );
  NAND4_X1 U23675 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_EBX_REG_9__SCAN_IN), .A3(P2_REIP_REG_16__SCAN_IN), .A4(
        P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20783) );
  NOR3_X1 U23676 ( .A1(n20785), .A2(n20784), .A3(n20783), .ZN(n20803) );
  NAND4_X1 U23677 ( .A1(P2_REIP_REG_21__SCAN_IN), .A2(READY2), .A3(
        P3_EAX_REG_5__SCAN_IN), .A4(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20789)
         );
  NAND4_X1 U23678 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_1__2__SCAN_IN), .A3(P3_REIP_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20788) );
  NAND4_X1 U23679 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A4(P2_DATAO_REG_17__SCAN_IN), .ZN(n20787) );
  NAND4_X1 U23680 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .A3(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A4(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20786) );
  NOR4_X1 U23681 ( .A1(n20789), .A2(n20788), .A3(n20787), .A4(n20786), .ZN(
        n20802) );
  NAND4_X1 U23682 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_2__4__SCAN_IN), .A3(P1_INSTQUEUE_REG_6__0__SCAN_IN), 
        .A4(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20800) );
  NOR4_X1 U23683 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P2_DATAO_REG_7__SCAN_IN), .A4(n20790), 
        .ZN(n20793) );
  NOR4_X1 U23684 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(BUF1_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20792) );
  NOR4_X1 U23685 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(P2_UWORD_REG_7__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(
        n20791) );
  NAND3_X1 U23686 ( .A1(n20793), .A2(n20792), .A3(n20791), .ZN(n20799) );
  NOR4_X1 U23687 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(P3_DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n20797) );
  NOR4_X1 U23688 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(
        P3_LWORD_REG_1__SCAN_IN), .A3(P3_UWORD_REG_2__SCAN_IN), .A4(
        P3_DATAO_REG_20__SCAN_IN), .ZN(n20796) );
  NOR4_X1 U23689 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(
        P2_REIP_REG_11__SCAN_IN), .A3(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n20795) );
  NOR4_X1 U23690 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A4(P2_REIP_REG_29__SCAN_IN), 
        .ZN(n20794) );
  NAND4_X1 U23691 ( .A1(n20797), .A2(n20796), .A3(n20795), .A4(n20794), .ZN(
        n20798) );
  NOR3_X1 U23692 ( .A1(n20800), .A2(n20799), .A3(n20798), .ZN(n20801) );
  NAND4_X1 U23693 ( .A1(n20804), .A2(n20803), .A3(n20802), .A4(n20801), .ZN(
        n20805) );
  XNOR2_X1 U23694 ( .A(n20806), .B(n20805), .ZN(n20807) );
  XNOR2_X1 U23695 ( .A(n20808), .B(n20807), .ZN(P1_U3093) );
  INV_X1 U11119 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10329) );
  NAND2_X1 U11296 ( .A1(n9754), .A2(n9717), .ZN(n13827) );
  CLKBUF_X2 U12736 ( .A(n15435), .Z(n16869) );
  AND2_X1 U13264 ( .A1(n12461), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10431) );
  CLKBUF_X1 U11053 ( .A(n11584), .Z(n11469) );
  CLKBUF_X2 U11094 ( .A(n11351), .Z(n11968) );
  CLKBUF_X1 U11097 ( .A(n15435), .Z(n16772) );
  CLKBUF_X1 U11110 ( .A(n15423), .Z(n9607) );
  CLKBUF_X2 U11121 ( .A(n11448), .Z(n13977) );
  CLKBUF_X1 U11134 ( .A(n11424), .Z(n13289) );
  CLKBUF_X1 U11323 ( .A(n18676), .Z(n18764) );
  CLKBUF_X1 U11326 ( .A(n11023), .Z(n12418) );
  CLKBUF_X2 U12256 ( .A(n12195), .Z(n12845) );
  NOR2_X1 U12357 ( .A1(n14096), .A2(n13970), .ZN(n14069) );
  NOR2_X1 U12777 ( .A1(n20547), .A2(n13958), .ZN(n13316) );
  XNOR2_X1 U13231 ( .A(n14311), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14544) );
  CLKBUF_X1 U14303 ( .A(n11023), .Z(n9600) );
  CLKBUF_X2 U14575 ( .A(n15048), .Z(n15313) );
  CLKBUF_X1 U16443 ( .A(n12197), .Z(n9592) );
  CLKBUF_X1 U17181 ( .A(n16156), .Z(n16163) );
endmodule

