

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653;

  INV_X2 U3684 ( .A(n4212), .ZN(n3650) );
  INV_X2 U3685 ( .A(n4221), .ZN(n4212) );
  CLKBUF_X1 U3686 ( .A(n4289), .Z(n5111) );
  CLKBUF_X2 U3687 ( .A(n3900), .Z(n4756) );
  NAND2_X1 U3688 ( .A1(n5158), .A2(n4018), .ZN(n5146) );
  OR2_X1 U3689 ( .A1(n3897), .A2(n3896), .ZN(n4044) );
  INV_X1 U3690 ( .A(n3923), .ZN(n4018) );
  AND2_X1 U3691 ( .A1(n6676), .A2(n6252), .ZN(n3661) );
  AND2_X1 U3692 ( .A1(n5072), .A2(n6671), .ZN(n3668) );
  AND2_X1 U3693 ( .A1(n5072), .A2(n6670), .ZN(n3901) );
  AND2_X1 U3694 ( .A1(n6676), .A2(n5071), .ZN(n4009) );
  AND2_X1 U3695 ( .A1(n5071), .A2(n6670), .ZN(n3900) );
  AND3_X1 U3696 ( .A1(n3949), .A2(n4962), .A3(n3924), .ZN(n3932) );
  INV_X1 U3697 ( .A(n4252), .ZN(n4269) );
  NAND2_X1 U3699 ( .A1(n4290), .A2(n4643), .ZN(n5087) );
  NAND2_X1 U3700 ( .A1(n3935), .A2(n3934), .ZN(n4055) );
  AND2_X2 U3701 ( .A1(n6266), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n6677)
         );
  NAND2_X1 U3702 ( .A1(n5019), .A2(n6328), .ZN(n5142) );
  NAND2_X1 U3703 ( .A1(n5158), .A2(n6233), .ZN(n3939) );
  AND2_X1 U3704 ( .A1(n4044), .A2(n3988), .ZN(n4914) );
  NOR2_X1 U3705 ( .A1(n6495), .A2(n4212), .ZN(n6223) );
  INV_X1 U3706 ( .A(n3988), .ZN(n3942) );
  INV_X1 U3707 ( .A(n3926), .ZN(n5158) );
  INV_X1 U3708 ( .A(n5099), .ZN(n3989) );
  INV_X1 U3710 ( .A(n3925), .ZN(n5246) );
  OR3_X1 U3711 ( .A1(n6421), .A2(n5582), .A3(n7296), .ZN(n7239) );
  AND2_X2 U3712 ( .A1(n5071), .A2(n6677), .ZN(n3908) );
  OAI21_X1 U3713 ( .B1(n5114), .B2(n4425), .A(n4300), .ZN(n5097) );
  OAI21_X1 U3714 ( .B1(n5114), .B2(n3942), .A(n4021), .ZN(n5271) );
  AND2_X4 U3715 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  OAI21_X2 U3716 ( .B1(n5035), .B2(n3743), .A(n3741), .ZN(n6222) );
  OR2_X2 U3717 ( .A1(n4079), .A2(n4078), .ZN(n5159) );
  NOR2_X2 U3718 ( .A1(n6023), .A2(n6022), .ZN(n6040) );
  AND4_X2 U3719 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3827)
         );
  XNOR2_X2 U3720 ( .A(n6071), .B(n4440), .ZN(n6142) );
  NAND2_X2 U3721 ( .A1(n3657), .A2(n5528), .ZN(n6071) );
  XNOR2_X2 U3722 ( .A(n4050), .B(n4053), .ZN(n5073) );
  NAND2_X2 U3723 ( .A1(n4000), .A2(n4051), .ZN(n4050) );
  BUF_X1 U3725 ( .A(n5110), .Z(n3662) );
  AND2_X1 U3726 ( .A1(n3899), .A2(n3898), .ZN(n3949) );
  AND2_X1 U3727 ( .A1(n3939), .A2(n5239), .ZN(n3928) );
  AND2_X2 U3729 ( .A1(n3983), .A2(n3988), .ZN(n5099) );
  BUF_X2 U3730 ( .A(n3988), .Z(n5226) );
  INV_X1 U3731 ( .A(n5239), .ZN(n3980) );
  AND4_X1 U3732 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3791)
         );
  AND4_X1 U3733 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3790)
         );
  CLKBUF_X2 U3734 ( .A(n4003), .Z(n4754) );
  BUF_X2 U3735 ( .A(n3908), .Z(n3666) );
  CLKBUF_X2 U3736 ( .A(n3901), .Z(n4755) );
  BUF_X2 U3737 ( .A(n3903), .Z(n3653) );
  BUF_X1 U3738 ( .A(n3903), .Z(n3675) );
  CLKBUF_X2 U3739 ( .A(n3961), .Z(n4761) );
  BUF_X2 U3740 ( .A(n4063), .Z(n3663) );
  BUF_X2 U3741 ( .A(n4009), .Z(n4753) );
  AND2_X2 U3742 ( .A1(n6677), .A2(n5072), .ZN(n4064) );
  CLKBUF_X2 U3743 ( .A(n3910), .Z(n4762) );
  AND2_X2 U3744 ( .A1(n6677), .A2(n5104), .ZN(n3902) );
  BUF_X4 U3745 ( .A(n3674), .Z(n3651) );
  BUF_X4 U3746 ( .A(n3908), .Z(n3652) );
  AND2_X2 U3747 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6252) );
  AOI21_X1 U3748 ( .B1(n6313), .B2(n6937), .A(n5016), .ZN(n5017) );
  XNOR2_X1 U3749 ( .A(n4797), .B(n4796), .ZN(n6313) );
  NOR2_X1 U3750 ( .A1(n4231), .A2(n6496), .ZN(n4232) );
  AND2_X1 U3751 ( .A1(n4998), .A2(n4212), .ZN(n6496) );
  AND2_X1 U3752 ( .A1(n6351), .A2(n6367), .ZN(n7514) );
  XNOR2_X1 U3753 ( .A(n4792), .B(n4781), .ZN(n6479) );
  NAND2_X1 U3754 ( .A1(n6924), .A2(n6923), .ZN(n6922) );
  OAI21_X1 U3755 ( .B1(n6222), .B2(n4228), .A(n4227), .ZN(n4229) );
  NAND2_X1 U3756 ( .A1(n3740), .A2(n3745), .ZN(n6924) );
  CLKBUF_X1 U3757 ( .A(n6364), .Z(n6365) );
  CLKBUF_X1 U3758 ( .A(n6390), .Z(n6391) );
  CLKBUF_X1 U3759 ( .A(n6446), .Z(n6447) );
  NAND2_X1 U3760 ( .A1(n4218), .A2(n4217), .ZN(n6177) );
  CLKBUF_X1 U3761 ( .A(n5994), .Z(n3656) );
  NAND2_X1 U3762 ( .A1(n5544), .A2(n4211), .ZN(n5996) );
  AND2_X1 U3763 ( .A1(n3742), .A2(n4225), .ZN(n3741) );
  OR2_X1 U3764 ( .A1(n3678), .A2(n3722), .ZN(n3721) );
  OR2_X1 U3765 ( .A1(n3677), .A2(n3743), .ZN(n3742) );
  AND2_X1 U3766 ( .A1(n3723), .A2(n3650), .ZN(n3678) );
  OR2_X1 U3767 ( .A1(n4226), .A2(n3744), .ZN(n3743) );
  OR2_X1 U3768 ( .A1(n4213), .A2(n3695), .ZN(n3723) );
  AND2_X1 U3769 ( .A1(n3650), .A2(n4219), .ZN(n6202) );
  NAND2_X1 U3770 ( .A1(n4140), .A2(n4139), .ZN(n4141) );
  OAI21_X1 U3771 ( .B1(n4325), .B2(n4202), .A(n4159), .ZN(n4160) );
  NOR2_X1 U3772 ( .A1(n3717), .A2(n6354), .ZN(n6355) );
  XNOR2_X1 U3773 ( .A(n4191), .B(n4190), .ZN(n4339) );
  NAND2_X1 U3774 ( .A1(n4178), .A2(n4177), .ZN(n4191) );
  OR2_X1 U3775 ( .A1(n5087), .A2(n5088), .ZN(n4308) );
  OR2_X1 U3776 ( .A1(n3682), .A2(n6368), .ZN(n3717) );
  NAND2_X1 U3777 ( .A1(n4077), .A2(n3738), .ZN(n5114) );
  OR2_X1 U3778 ( .A1(n3680), .A2(n6450), .ZN(n4892) );
  OR2_X1 U3779 ( .A1(n5138), .A2(n4317), .ZN(n4295) );
  AND2_X2 U3780 ( .A1(n4043), .A2(n4042), .ZN(n5161) );
  NAND2_X1 U3781 ( .A1(n4043), .A2(n3976), .ZN(n4002) );
  OR2_X1 U3782 ( .A1(n7407), .A2(n4425), .ZN(n4294) );
  NAND2_X1 U3783 ( .A1(n3739), .A2(n7313), .ZN(n4043) );
  CLKBUF_X1 U3784 ( .A(n4292), .Z(n7407) );
  AND2_X2 U3785 ( .A1(n5367), .A2(n5205), .ZN(n5487) );
  OAI21_X1 U3786 ( .B1(n3993), .B2(n4946), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3996) );
  OAI21_X1 U3787 ( .B1(n4798), .B2(n3987), .A(n4949), .ZN(n3993) );
  NAND2_X1 U3788 ( .A1(n3920), .A2(n3919), .ZN(n3977) );
  AND2_X1 U3789 ( .A1(n3982), .A2(n5183), .ZN(n5019) );
  AND2_X1 U3790 ( .A1(n3925), .A2(n4018), .ZN(n4288) );
  OR2_X1 U3792 ( .A1(n4016), .A2(n4062), .ZN(n4001) );
  OR2_X1 U3793 ( .A1(n4237), .A2(n3925), .ZN(n4252) );
  AND2_X1 U3794 ( .A1(n3980), .A2(n4044), .ZN(n3920) );
  NAND2_X2 U3795 ( .A1(n3780), .A2(n3917), .ZN(n5239) );
  AND3_X1 U3796 ( .A1(n3685), .A2(n3882), .A3(n3751), .ZN(n3752) );
  AND4_X2 U3797 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3925)
         );
  NAND2_X2 U3798 ( .A1(n3791), .A2(n3790), .ZN(n3926) );
  AND4_X1 U3799 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3866)
         );
  AND4_X1 U3800 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3882)
         );
  AND4_X1 U3801 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3847)
         );
  AND4_X1 U3802 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3917)
         );
  AND4_X1 U3803 ( .A1(n3825), .A2(n3824), .A3(n3823), .A4(n3822), .ZN(n3826)
         );
  AND4_X1 U3804 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3868)
         );
  AND4_X1 U3805 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3814)
         );
  AND4_X1 U3806 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3845)
         );
  AND4_X1 U3807 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3881)
         );
  AND4_X1 U3808 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3815)
         );
  AND4_X1 U3809 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3883)
         );
  AND4_X1 U3810 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3867)
         );
  AND4_X1 U3811 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3846)
         );
  AND4_X1 U3812 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3865)
         );
  BUF_X4 U3813 ( .A(n3902), .Z(n3664) );
  BUF_X4 U3814 ( .A(n3902), .Z(n3665) );
  BUF_X4 U3815 ( .A(n4064), .Z(n3671) );
  BUF_X4 U3816 ( .A(n4064), .Z(n3670) );
  INV_X2 U3817 ( .A(n7350), .ZN(n6947) );
  AND2_X2 U3818 ( .A1(n6676), .A2(n5104), .ZN(n3911) );
  AND2_X2 U3819 ( .A1(n6676), .A2(n6252), .ZN(n3660) );
  AND2_X2 U3820 ( .A1(n6252), .A2(n6671), .ZN(n4065) );
  AND2_X2 U3821 ( .A1(n4310), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6676)
         );
  AND2_X2 U3822 ( .A1(n6252), .A2(n6671), .ZN(n3673) );
  AND2_X2 U3823 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n6671) );
  NOR2_X2 U3824 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6670) );
  AND2_X1 U3825 ( .A1(n3778), .A2(n3725), .ZN(n3655) );
  AOI21_X1 U3826 ( .B1(n3726), .B2(n3734), .A(n3693), .ZN(n3725) );
  NAND2_X1 U3827 ( .A1(n3655), .A2(n3724), .ZN(n5035) );
  NAND2_X1 U3828 ( .A1(n5996), .A2(n5995), .ZN(n5994) );
  AND2_X1 U3829 ( .A1(n6072), .A2(n3691), .ZN(n3657) );
  AOI21_X2 U3830 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4212), .A(n6927), 
        .ZN(n6538) );
  NAND2_X1 U3831 ( .A1(n6446), .A2(n6448), .ZN(n6390) );
  AND2_X2 U3832 ( .A1(n6676), .A2(n5104), .ZN(n3658) );
  NAND2_X1 U3833 ( .A1(n4113), .A2(n5175), .ZN(n5221) );
  NOR2_X1 U3834 ( .A1(n3921), .A2(n3977), .ZN(n4962) );
  OAI222_X1 U3835 ( .A1(n6468), .A2(n6244), .B1(n6232), .B2(n6880), .C1(n6592), 
        .C2(n6876), .ZN(U2831) );
  INV_X2 U3836 ( .A(n6390), .ZN(n4603) );
  NOR2_X1 U3837 ( .A1(n6351), .A2(n3764), .ZN(n4792) );
  NOR2_X2 U3838 ( .A1(n4229), .A2(n6612), .ZN(n4997) );
  OR2_X1 U3839 ( .A1(n4002), .A2(n3748), .ZN(n3738) );
  OAI21_X1 U3840 ( .B1(n5073), .B2(STATE2_REG_0__SCAN_IN), .A(n4001), .ZN(
        n3748) );
  XNOR2_X1 U3841 ( .A(n3736), .B(n6593), .ZN(n6601) );
  XNOR2_X1 U3842 ( .A(n6339), .B(n6341), .ZN(n6504) );
  NAND2_X2 U3843 ( .A1(n4060), .A2(n7091), .ZN(n5163) );
  INV_X2 U3844 ( .A(n4292), .ZN(n3739) );
  NOR2_X2 U3845 ( .A1(n6461), .A2(n3755), .ZN(n6446) );
  NAND2_X2 U3846 ( .A1(n4494), .A2(n4493), .ZN(n6461) );
  AOI21_X1 U3847 ( .B1(n5111), .B2(n4259), .A(n4084), .ZN(n6896) );
  NOR2_X2 U3848 ( .A1(n5254), .A2(n4351), .ZN(n5527) );
  AND2_X1 U3849 ( .A1(n6676), .A2(n6252), .ZN(n4004) );
  OAI211_X1 U3850 ( .C1(n4321), .C2(n3781), .A(n4294), .B(n4293), .ZN(n5138)
         );
  AND2_X2 U3851 ( .A1(n3781), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5072)
         );
  NOR2_X2 U3852 ( .A1(n6351), .A2(n6353), .ZN(n6352) );
  XNOR2_X1 U3853 ( .A(n7091), .B(n7089), .ZN(n5110) );
  NOR2_X2 U3854 ( .A1(n5086), .A2(n5132), .ZN(n5131) );
  OAI21_X2 U3855 ( .B1(n6142), .B2(n6143), .A(n4441), .ZN(n6186) );
  AND2_X1 U3856 ( .A1(n5072), .A2(n6671), .ZN(n4063) );
  AND2_X1 U3857 ( .A1(n5072), .A2(n6671), .ZN(n3669) );
  AND2_X2 U3858 ( .A1(n3983), .A2(n3942), .ZN(n4017) );
  AND2_X1 U3859 ( .A1(n6252), .A2(n6671), .ZN(n3672) );
  AND2_X4 U3860 ( .A1(n6670), .A2(n6252), .ZN(n3912) );
  AND2_X1 U3861 ( .A1(n6677), .A2(n6252), .ZN(n3674) );
  AND2_X1 U3862 ( .A1(n6677), .A2(n6252), .ZN(n3903) );
  INV_X1 U3863 ( .A(n4317), .ZN(n4777) );
  AND2_X1 U3864 ( .A1(n3768), .A2(n3766), .ZN(n3765) );
  INV_X1 U3865 ( .A(n6353), .ZN(n3766) );
  NOR2_X1 U3866 ( .A1(n6340), .A2(n3769), .ZN(n3768) );
  INV_X1 U3867 ( .A(n6226), .ZN(n3769) );
  INV_X1 U3868 ( .A(n3745), .ZN(n3744) );
  NAND2_X1 U3869 ( .A1(n4279), .A2(n4278), .ZN(n4805) );
  NAND2_X1 U3870 ( .A1(n5367), .A2(n6327), .ZN(n5140) );
  AND2_X1 U3871 ( .A1(n3981), .A2(n3980), .ZN(n3982) );
  INV_X1 U3872 ( .A(n4643), .ZN(n4793) );
  AOI21_X1 U3873 ( .B1(n4780), .B2(n4779), .A(n4778), .ZN(n4791) );
  INV_X1 U3874 ( .A(n6366), .ZN(n4689) );
  INV_X1 U3875 ( .A(n6364), .ZN(n4690) );
  NAND2_X1 U3876 ( .A1(n4732), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4811)
         );
  AOI21_X1 U3877 ( .B1(n4777), .B2(n6237), .A(n4731), .ZN(n6226) );
  NOR2_X1 U3878 ( .A1(n6325), .A2(n7318), .ZN(n5367) );
  INV_X1 U3879 ( .A(n6864), .ZN(n3713) );
  INV_X1 U3880 ( .A(n6865), .ZN(n3712) );
  AND2_X1 U3881 ( .A1(n4975), .A2(n4974), .ZN(n6254) );
  NOR2_X1 U3882 ( .A1(n3775), .A2(n3832), .ZN(n3848) );
  INV_X2 U3883 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7295) );
  INV_X1 U3884 ( .A(n4234), .ZN(n4247) );
  AND2_X1 U3885 ( .A1(n4115), .A2(n4128), .ZN(n3749) );
  INV_X1 U3886 ( .A(n4130), .ZN(n4128) );
  OR2_X1 U3887 ( .A1(n4125), .A2(n4124), .ZN(n4137) );
  OR2_X1 U3888 ( .A1(n3971), .A2(n3970), .ZN(n4080) );
  AOI21_X1 U3889 ( .B1(n4090), .B2(n5382), .A(n3994), .ZN(n3997) );
  NAND2_X1 U3890 ( .A1(n4268), .A2(n7250), .ZN(n4806) );
  INV_X1 U3891 ( .A(n4275), .ZN(n4268) );
  INV_X1 U3892 ( .A(n6950), .ZN(n5364) );
  AND2_X1 U3893 ( .A1(n6406), .A2(n3761), .ZN(n3760) );
  INV_X1 U3894 ( .A(n6462), .ZN(n3761) );
  NOR2_X2 U3895 ( .A1(n3926), .A2(n7295), .ZN(n4468) );
  OR2_X1 U3896 ( .A1(n6443), .A2(n3718), .ZN(n3716) );
  INV_X1 U3897 ( .A(n4955), .ZN(n3718) );
  NAND2_X1 U3898 ( .A1(n3650), .A2(n3746), .ZN(n3745) );
  INV_X1 U3899 ( .A(n6644), .ZN(n3746) );
  INV_X1 U3900 ( .A(n6567), .ZN(n3727) );
  INV_X1 U3901 ( .A(n6202), .ZN(n3735) );
  AND2_X1 U3902 ( .A1(n6039), .A2(n6074), .ZN(n3706) );
  OR2_X1 U3903 ( .A1(n5134), .A2(n3711), .ZN(n3709) );
  INV_X1 U3904 ( .A(n5153), .ZN(n3711) );
  INV_X1 U3905 ( .A(n5135), .ZN(n3707) );
  OR2_X1 U3906 ( .A1(n4075), .A2(n4074), .ZN(n4105) );
  OR2_X1 U3907 ( .A1(n4015), .A2(n4014), .ZN(n4081) );
  AND2_X1 U3908 ( .A1(n4018), .A2(n5226), .ZN(n4259) );
  NAND2_X1 U3909 ( .A1(n5183), .A2(n3983), .ZN(n4909) );
  INV_X2 U3910 ( .A(n3659), .ZN(n4916) );
  AND2_X1 U3911 ( .A1(n4088), .A2(n6273), .ZN(n5285) );
  NAND2_X1 U3912 ( .A1(n3911), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3751) );
  NOR2_X1 U3913 ( .A1(n3817), .A2(n3816), .ZN(n3923) );
  NAND2_X1 U3914 ( .A1(n3815), .A2(n3814), .ZN(n3816) );
  INV_X1 U3915 ( .A(n4017), .ZN(n4957) );
  AND2_X1 U3916 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4692), .ZN(n4693)
         );
  NAND2_X1 U3917 ( .A1(n4693), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4713)
         );
  INV_X1 U3918 ( .A(n6470), .ZN(n4493) );
  AND2_X1 U3919 ( .A1(n4939), .A2(n4288), .ZN(n4947) );
  AND2_X1 U3920 ( .A1(n6355), .A2(n6230), .ZN(n6345) );
  OR2_X1 U3921 ( .A1(n3650), .A2(n4872), .ZN(n6560) );
  NOR2_X1 U3922 ( .A1(n6190), .A2(n4871), .ZN(n6472) );
  INV_X1 U3923 ( .A(n6177), .ZN(n3730) );
  AOI21_X1 U3924 ( .B1(n3733), .B2(n3676), .A(n3688), .ZN(n3732) );
  NOR2_X1 U3925 ( .A1(n6202), .A2(n6178), .ZN(n3733) );
  NAND2_X1 U3926 ( .A1(n3712), .A2(n3690), .ZN(n6023) );
  OR2_X1 U3927 ( .A1(n5258), .A2(n5328), .ZN(n6865) );
  OR2_X1 U3928 ( .A1(n4933), .A2(n3989), .ZN(n3992) );
  AND2_X1 U3929 ( .A1(n4945), .A2(n4944), .ZN(n4983) );
  AND2_X1 U3930 ( .A1(n4916), .A2(n4909), .ZN(n5121) );
  AND2_X1 U3931 ( .A1(n4285), .A2(n4284), .ZN(n6325) );
  NAND2_X1 U3932 ( .A1(n4283), .A2(n4805), .ZN(n4284) );
  OR2_X1 U3933 ( .A1(n3662), .A2(n7445), .ZN(n5387) );
  INV_X1 U3934 ( .A(n4044), .ZN(n5183) );
  NOR2_X1 U3935 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5157), .ZN(n5280) );
  AND2_X1 U3936 ( .A1(n3662), .A2(n7457), .ZN(n6093) );
  OR2_X1 U3937 ( .A1(n4933), .A2(n4957), .ZN(n7289) );
  OAI21_X1 U3938 ( .B1(n6350), .B2(REIP_REG_29__SCAN_IN), .A(n3699), .ZN(n3698) );
  NAND2_X1 U3939 ( .A1(n6348), .A2(REIP_REG_29__SCAN_IN), .ZN(n3699) );
  OR3_X1 U3940 ( .A1(n6953), .A2(n3989), .A3(n4922), .ZN(n7195) );
  OR2_X1 U3941 ( .A1(n6574), .A2(n6876), .ZN(n5027) );
  NAND2_X1 U3942 ( .A1(n5492), .A2(n5145), .ZN(n6311) );
  OAI21_X1 U3943 ( .B1(n5144), .B2(n5143), .A(n7292), .ZN(n5145) );
  XNOR2_X1 U3944 ( .A(n4812), .B(n4824), .ZN(n5581) );
  NAND2_X1 U3945 ( .A1(n3767), .A2(n3689), .ZN(n4797) );
  INV_X1 U3946 ( .A(n6340), .ZN(n6341) );
  NAND2_X1 U3947 ( .A1(n6906), .A2(n6884), .ZN(n6940) );
  NAND2_X1 U3948 ( .A1(n5367), .A2(n4947), .ZN(n7241) );
  INV_X1 U3949 ( .A(n6906), .ZN(n6932) );
  XNOR2_X1 U3950 ( .A(n6345), .B(n3701), .ZN(n6583) );
  INV_X1 U3951 ( .A(n6346), .ZN(n3701) );
  NOR2_X1 U3952 ( .A1(n6497), .A2(n6496), .ZN(n6500) );
  NOR2_X1 U3953 ( .A1(n6223), .A2(n3737), .ZN(n3736) );
  AND2_X1 U3954 ( .A1(n4981), .A2(n4980), .ZN(n7064) );
  AND2_X1 U3955 ( .A1(n7284), .A2(n7283), .ZN(n7319) );
  INV_X1 U3956 ( .A(n4114), .ZN(n3750) );
  AND2_X1 U3957 ( .A1(n4127), .A2(n4126), .ZN(n4130) );
  AND2_X1 U3958 ( .A1(n4176), .A2(n4175), .ZN(n4177) );
  INV_X1 U3959 ( .A(n4179), .ZN(n4176) );
  INV_X1 U3960 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4276) );
  OR2_X1 U3961 ( .A1(n4277), .A2(n4276), .ZN(n4275) );
  OR2_X1 U3962 ( .A1(n3983), .A2(n7313), .ZN(n4061) );
  NAND2_X1 U3963 ( .A1(n4269), .A2(n4259), .ZN(n4271) );
  AOI22_X1 U3964 ( .A1(n4003), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3788) );
  OR2_X1 U3965 ( .A1(n4032), .A2(n4031), .ZN(n4206) );
  INV_X1 U3966 ( .A(n3990), .ZN(n4800) );
  AND2_X1 U3967 ( .A1(n3763), .A2(n6381), .ZN(n3762) );
  NOR2_X1 U3968 ( .A1(n6439), .A2(n6392), .ZN(n3763) );
  NAND2_X1 U3969 ( .A1(n3756), .A2(n4563), .ZN(n3755) );
  INV_X1 U3970 ( .A(n3758), .ZN(n3756) );
  NAND2_X1 U3971 ( .A1(n3760), .A2(n3759), .ZN(n3758) );
  INV_X1 U3972 ( .A(n6870), .ZN(n3759) );
  AND2_X1 U3973 ( .A1(n4397), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4422)
         );
  INV_X1 U3974 ( .A(n6038), .ZN(n3753) );
  AND2_X1 U3975 ( .A1(n4396), .A2(n5539), .ZN(n3754) );
  INV_X1 U3976 ( .A(n6021), .ZN(n4396) );
  NOR2_X1 U3977 ( .A1(n4367), .A2(n4362), .ZN(n4381) );
  INV_X1 U3978 ( .A(n4327), .ZN(n4326) );
  AND2_X1 U3979 ( .A1(n4213), .A2(n3696), .ZN(n3722) );
  NAND2_X1 U3980 ( .A1(n3678), .A2(n3695), .ZN(n3720) );
  INV_X1 U3981 ( .A(n4906), .ZN(n4881) );
  NAND2_X1 U3982 ( .A1(n4132), .A2(n4259), .ZN(n4140) );
  AND2_X1 U3983 ( .A1(n3661), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3775) );
  INV_X1 U3984 ( .A(n4080), .ZN(n4016) );
  NAND2_X1 U3985 ( .A1(n3925), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U3986 ( .A1(n3937), .A2(n3936), .ZN(n3959) );
  INV_X1 U3987 ( .A(n4271), .ZN(n4283) );
  NAND2_X1 U3988 ( .A1(n4092), .A2(n4091), .ZN(n7089) );
  AOI21_X1 U3989 ( .B1(n7306), .B2(n7314), .A(n6689), .ZN(n5157) );
  NAND2_X1 U3990 ( .A1(n7294), .A2(n7313), .ZN(n4784) );
  AND2_X1 U3991 ( .A1(n4807), .A2(n4806), .ZN(n6317) );
  INV_X1 U3992 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6009) );
  AND2_X1 U3993 ( .A1(n4670), .A2(n4669), .ZN(n6433) );
  OR2_X1 U3994 ( .A1(n7240), .A2(n4317), .ZN(n4670) );
  INV_X1 U3995 ( .A(n3709), .ZN(n3710) );
  AND2_X1 U3996 ( .A1(n4777), .A2(n6556), .ZN(n4525) );
  NAND2_X1 U3997 ( .A1(n5369), .A2(n5368), .ZN(n6755) );
  INV_X1 U3998 ( .A(n5492), .ZN(n5475) );
  INV_X1 U3999 ( .A(n6351), .ZN(n3767) );
  AND2_X1 U4000 ( .A1(n4649), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4650)
         );
  NAND2_X1 U4001 ( .A1(n4604), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4605)
         );
  NOR2_X1 U4002 ( .A1(n4565), .A2(n4564), .ZN(n4566) );
  AND2_X1 U4003 ( .A1(n4566), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4604)
         );
  OR2_X1 U4004 ( .A1(n7213), .A2(n4317), .ZN(n4584) );
  NOR2_X1 U4005 ( .A1(n4529), .A2(n4528), .ZN(n4530) );
  NAND2_X1 U4006 ( .A1(n4530), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4565)
         );
  INV_X1 U4007 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U4008 ( .A1(n4497), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4529)
         );
  AND2_X1 U4009 ( .A1(n4459), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4478)
         );
  INV_X1 U4010 ( .A(n6211), .ZN(n4476) );
  NOR2_X1 U4011 ( .A1(n4455), .A2(n6179), .ZN(n4459) );
  CLKBUF_X1 U4012 ( .A(n6187), .Z(n6188) );
  AND2_X1 U4013 ( .A1(n4422), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4438)
         );
  AND2_X1 U4014 ( .A1(n4381), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4397)
         );
  AND2_X1 U4015 ( .A1(n4335), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4340)
         );
  AOI21_X1 U4016 ( .B1(n4332), .B2(n4468), .A(n4331), .ZN(n5256) );
  CLKBUF_X1 U4017 ( .A(n5254), .Z(n5255) );
  CLKBUF_X1 U4018 ( .A(n5149), .Z(n5150) );
  NOR2_X1 U4019 ( .A1(n4311), .A2(n6009), .ZN(n4318) );
  NAND2_X1 U4020 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4311) );
  INV_X1 U4021 ( .A(n4299), .ZN(n4300) );
  OAI21_X1 U4022 ( .B1(n4321), .B2(n4297), .A(n4298), .ZN(n4299) );
  INV_X1 U4023 ( .A(n5138), .ZN(n4296) );
  OR2_X1 U4024 ( .A1(n3650), .A2(n4224), .ZN(n4225) );
  NAND2_X1 U4025 ( .A1(n3715), .A2(n6434), .ZN(n3714) );
  INV_X1 U4026 ( .A(n3716), .ZN(n3715) );
  OR2_X1 U4027 ( .A1(n4892), .A2(n6394), .ZN(n6442) );
  NOR2_X1 U4028 ( .A1(n6442), .A2(n6443), .ZN(n6441) );
  OR3_X1 U4029 ( .A1(n6872), .A2(n5034), .A3(n3703), .ZN(n3702) );
  INV_X1 U4030 ( .A(n6455), .ZN(n3703) );
  NOR3_X1 U4031 ( .A1(n6466), .A2(n6872), .A3(n5034), .ZN(n6875) );
  NAND2_X1 U4032 ( .A1(n5035), .A2(n3677), .ZN(n3740) );
  AND2_X1 U4033 ( .A1(n4878), .A2(n4877), .ZN(n6464) );
  NAND2_X1 U4034 ( .A1(n6474), .A2(n6464), .ZN(n6466) );
  AND2_X1 U4035 ( .A1(n6472), .A2(n6471), .ZN(n6474) );
  NAND2_X1 U4036 ( .A1(n3724), .A2(n3725), .ZN(n6559) );
  NAND2_X1 U4037 ( .A1(n6040), .A2(n3679), .ZN(n6190) );
  INV_X1 U4038 ( .A(n6145), .ZN(n3705) );
  AND2_X1 U4039 ( .A1(n6040), .A2(n6039), .ZN(n6075) );
  NAND2_X1 U4040 ( .A1(n6040), .A2(n3706), .ZN(n6144) );
  NOR2_X1 U4041 ( .A1(n6865), .A2(n6864), .ZN(n6867) );
  NOR2_X1 U4042 ( .A1(n5259), .A2(n3709), .ZN(n3708) );
  XNOR2_X1 U4043 ( .A(n4141), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5222)
         );
  OR2_X1 U4044 ( .A1(n5093), .A2(n5092), .ZN(n5135) );
  NOR2_X1 U4045 ( .A1(n5135), .A2(n5134), .ZN(n5154) );
  OR2_X1 U4046 ( .A1(n4948), .A2(n5571), .ZN(n6319) );
  INV_X1 U4047 ( .A(n5316), .ZN(n6995) );
  NAND2_X1 U4048 ( .A1(n4002), .A2(n3748), .ZN(n4077) );
  INV_X1 U4049 ( .A(n5079), .ZN(n6245) );
  OR2_X1 U4050 ( .A1(n4479), .A2(n5239), .ZN(n5079) );
  NOR2_X1 U4051 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n7457) );
  OR2_X1 U4052 ( .A1(n5157), .A2(n7304), .ZN(n5213) );
  INV_X1 U4053 ( .A(n5280), .ZN(n5419) );
  AND2_X1 U4054 ( .A1(n3654), .A2(n5188), .ZN(n5421) );
  INV_X1 U4055 ( .A(n7457), .ZN(n7445) );
  AOI21_X1 U4056 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7394), .A(n5419), .ZN(
        n7459) );
  INV_X1 U4057 ( .A(n5213), .ZN(n5405) );
  OR3_X1 U4058 ( .A1(n6953), .A2(n4931), .A3(n4814), .ZN(n7192) );
  INV_X1 U4059 ( .A(n7215), .ZN(n7228) );
  AND2_X1 U4060 ( .A1(n6953), .A2(n4809), .ZN(n6421) );
  INV_X1 U4061 ( .A(n7203), .ZN(n7227) );
  INV_X1 U4062 ( .A(n7195), .ZN(n7235) );
  INV_X1 U4063 ( .A(n7112), .ZN(n7097) );
  AOI21_X1 U4064 ( .B1(n6345), .B2(n4917), .A(n5023), .ZN(n4920) );
  AND2_X1 U4065 ( .A1(n5022), .A2(n7292), .ZN(n6880) );
  INV_X1 U4066 ( .A(n6504), .ZN(n6485) );
  INV_X1 U4067 ( .A(n6311), .ZN(n7515) );
  AND2_X1 U4068 ( .A1(n6311), .A2(n6234), .ZN(n7516) );
  NAND2_X1 U4069 ( .A1(n6311), .A2(n5148), .ZN(n6219) );
  INV_X1 U4070 ( .A(n4791), .ZN(n4781) );
  INV_X1 U4071 ( .A(n3765), .ZN(n3764) );
  AND2_X1 U4072 ( .A1(n4734), .A2(n4714), .ZN(n6237) );
  INV_X1 U4073 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6179) );
  INV_X1 U4074 ( .A(n7241), .ZN(n6936) );
  AOI21_X1 U4075 ( .B1(n6345), .B2(n5024), .A(n5023), .ZN(n5026) );
  XNOR2_X1 U4076 ( .A(n5038), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6552)
         );
  NAND2_X1 U4077 ( .A1(n3728), .A2(n3732), .ZN(n6569) );
  NAND2_X1 U4078 ( .A1(n3730), .A2(n3729), .ZN(n3728) );
  NAND2_X1 U4079 ( .A1(n6177), .A2(n6178), .ZN(n3731) );
  NAND2_X1 U4080 ( .A1(n3712), .A2(n3686), .ZN(n5542) );
  AND2_X1 U4081 ( .A1(n4970), .A2(n5041), .ZN(n6992) );
  INV_X1 U4082 ( .A(n7023), .ZN(n7066) );
  INV_X1 U4083 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7394) );
  INV_X1 U4084 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7448) );
  INV_X1 U4085 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6251) );
  INV_X1 U4086 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7268) );
  INV_X1 U4087 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7296) );
  INV_X1 U4088 ( .A(n6682), .ZN(n7257) );
  NOR2_X1 U4089 ( .A1(n6325), .A2(n7305), .ZN(n6689) );
  INV_X1 U4090 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7250) );
  NOR2_X1 U4091 ( .A1(n5070), .A2(n7248), .ZN(n7244) );
  AND2_X1 U4092 ( .A1(n5342), .A2(n5341), .ZN(n6303) );
  INV_X1 U4093 ( .A(n5340), .ZN(n7647) );
  AND2_X1 U4094 ( .A1(n5170), .A2(n5169), .ZN(n6296) );
  OAI21_X1 U4095 ( .B1(n5166), .B2(n5165), .A(n5164), .ZN(n6295) );
  INV_X1 U4096 ( .A(n6290), .ZN(n7630) );
  INV_X1 U4097 ( .A(n7625), .ZN(n6283) );
  AND2_X1 U4098 ( .A1(n5289), .A2(n5288), .ZN(n6282) );
  INV_X1 U4099 ( .A(n7388), .ZN(n7612) );
  INV_X1 U4100 ( .A(n6701), .ZN(n7483) );
  INV_X1 U4101 ( .A(n6707), .ZN(n7506) );
  INV_X1 U4102 ( .A(n6719), .ZN(n7573) );
  NOR2_X1 U4103 ( .A1(n5213), .A2(n5158), .ZN(n7591) );
  INV_X1 U4104 ( .A(n6732), .ZN(n7644) );
  INV_X1 U4105 ( .A(n6706), .ZN(n7511) );
  INV_X1 U4106 ( .A(n6066), .ZN(n7538) );
  INV_X1 U4107 ( .A(n6712), .ZN(n7558) );
  INV_X1 U4108 ( .A(n6718), .ZN(n7578) );
  INV_X1 U4109 ( .A(n5430), .ZN(n6276) );
  INV_X1 U4110 ( .A(n7292), .ZN(n7318) );
  AND2_X1 U4111 ( .A1(n7291), .A2(n7290), .ZN(n7302) );
  AND2_X1 U4112 ( .A1(n4286), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7292) );
  INV_X1 U4113 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7305) );
  INV_X1 U4114 ( .A(n7333), .ZN(n6751) );
  INV_X1 U4115 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7345) );
  NAND2_X1 U4116 ( .A1(STATE_REG_1__SCAN_IN), .A2(n7345), .ZN(n7350) );
  NOR2_X1 U4117 ( .A1(n6347), .A2(n3698), .ZN(n3697) );
  OR2_X1 U4118 ( .A1(n6583), .A2(n7195), .ZN(n3700) );
  OAI21_X1 U4119 ( .B1(n6940), .B2(n5581), .A(n5015), .ZN(n5016) );
  AOI21_X1 U4120 ( .B1(n6504), .B2(n6937), .A(n6503), .ZN(n6505) );
  OAI21_X1 U4121 ( .B1(n6601), .B2(n7023), .A(n6600), .ZN(U2990) );
  INV_X1 U4122 ( .A(n3983), .ZN(n4963) );
  NAND2_X1 U4123 ( .A1(n3650), .A2(n4864), .ZN(n3676) );
  NOR2_X1 U4124 ( .A1(n6461), .A2(n6462), .ZN(n6404) );
  NAND2_X1 U4125 ( .A1(n5528), .A2(n5539), .ZN(n5538) );
  INV_X1 U4126 ( .A(n5114), .ZN(n5281) );
  AND2_X1 U4127 ( .A1(n6560), .A2(n3687), .ZN(n3677) );
  INV_X1 U4128 ( .A(n3734), .ZN(n3729) );
  NAND2_X1 U4129 ( .A1(n3735), .A2(n3676), .ZN(n3734) );
  AND2_X1 U4130 ( .A1(n3706), .A2(n3705), .ZN(n3679) );
  NAND2_X1 U4131 ( .A1(n4191), .A2(n4204), .ZN(n4221) );
  INV_X1 U4132 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4310) );
  AND2_X1 U4133 ( .A1(n5104), .A2(n6670), .ZN(n3910) );
  NAND2_X1 U4134 ( .A1(n3757), .A2(n3760), .ZN(n6405) );
  AND2_X1 U4135 ( .A1(n6676), .A2(n5072), .ZN(n4003) );
  OR2_X1 U4136 ( .A1(n6466), .A2(n3702), .ZN(n3680) );
  OR2_X1 U4137 ( .A1(n6352), .A2(n6226), .ZN(n3681) );
  OR2_X1 U4138 ( .A1(n6442), .A2(n3714), .ZN(n3682) );
  AND2_X1 U4139 ( .A1(n4603), .A2(n3762), .ZN(n6379) );
  NAND2_X1 U4140 ( .A1(n4603), .A2(n4602), .ZN(n6389) );
  NAND2_X1 U4141 ( .A1(n5035), .A2(n6560), .ZN(n5036) );
  NAND2_X1 U4142 ( .A1(n6352), .A2(n6226), .ZN(n6339) );
  AND2_X1 U4143 ( .A1(n3883), .A2(n3881), .ZN(n3683) );
  NOR2_X1 U4144 ( .A1(n3918), .A2(n5246), .ZN(n3938) );
  INV_X1 U4145 ( .A(n6461), .ZN(n3757) );
  OR2_X1 U4146 ( .A1(n6461), .A2(n3758), .ZN(n3684) );
  AND2_X1 U4147 ( .A1(n4603), .A2(n3763), .ZN(n6380) );
  AND3_X1 U4148 ( .A1(n3886), .A2(n3885), .A3(n3884), .ZN(n3685) );
  NAND2_X1 U4149 ( .A1(n3749), .A2(n3750), .ZN(n4156) );
  AND2_X1 U4150 ( .A1(n3732), .A2(n3727), .ZN(n3726) );
  INV_X1 U4151 ( .A(n4794), .ZN(n4751) );
  NAND2_X1 U4152 ( .A1(n5528), .A2(n3754), .ZN(n6019) );
  NAND2_X1 U4153 ( .A1(n3656), .A2(n4213), .ZN(n6084) );
  AND2_X1 U4154 ( .A1(n3713), .A2(n5531), .ZN(n3686) );
  OR2_X1 U4155 ( .A1(n3650), .A2(n4220), .ZN(n3687) );
  NOR2_X1 U4156 ( .A1(n3650), .A2(n4219), .ZN(n3688) );
  AND2_X1 U4157 ( .A1(n4791), .A2(n3765), .ZN(n3689) );
  AND2_X1 U4158 ( .A1(n3686), .A2(n4857), .ZN(n3690) );
  NAND2_X1 U4159 ( .A1(n3731), .A2(n3676), .ZN(n6201) );
  NOR2_X1 U4160 ( .A1(n6442), .A2(n3716), .ZN(n4954) );
  AND2_X1 U4161 ( .A1(n3754), .A2(n3753), .ZN(n3691) );
  AND2_X1 U4162 ( .A1(n6433), .A2(n3762), .ZN(n3692) );
  INV_X1 U4163 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3781) );
  INV_X1 U4164 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4297) );
  NAND2_X1 U4165 ( .A1(n3708), .A2(n3707), .ZN(n5258) );
  INV_X1 U4166 ( .A(n6878), .ZN(n6468) );
  INV_X1 U4167 ( .A(n6478), .ZN(n6878) );
  AND2_X1 U4168 ( .A1(n3650), .A2(n6662), .ZN(n3693) );
  NOR2_X1 U4169 ( .A1(n6466), .A2(n5034), .ZN(n3704) );
  OR2_X1 U4170 ( .A1(n6880), .A2(n6333), .ZN(n3694) );
  NAND2_X1 U4171 ( .A1(n3707), .A2(n3710), .ZN(n5152) );
  NAND2_X1 U4172 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3695) );
  AND2_X1 U4173 ( .A1(n4297), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5071)
         );
  NAND2_X1 U4174 ( .A1(n3992), .A2(n5074), .ZN(n4946) );
  AND2_X1 U4175 ( .A1(n4215), .A2(n4214), .ZN(n3696) );
  NOR2_X2 U4176 ( .A1(n7404), .A2(n5161), .ZN(n7622) );
  NOR2_X2 U4177 ( .A1(n7369), .A2(n5161), .ZN(n7597) );
  NOR2_X2 U4178 ( .A1(n7392), .A2(n5161), .ZN(n3771) );
  NAND2_X1 U4179 ( .A1(n4288), .A2(n4914), .ZN(n3898) );
  NAND3_X1 U4180 ( .A1(n6349), .A2(n3700), .A3(n3697), .ZN(U2798) );
  INV_X1 U4181 ( .A(n3704), .ZN(n6873) );
  NAND2_X1 U4182 ( .A1(n3719), .A2(n3720), .ZN(n4216) );
  NAND2_X1 U4183 ( .A1(n5994), .A2(n3721), .ZN(n3719) );
  NAND2_X1 U4184 ( .A1(n6177), .A2(n3726), .ZN(n3724) );
  AND2_X1 U4185 ( .A1(n6506), .A2(n6224), .ZN(n3737) );
  NAND2_X2 U4186 ( .A1(n3959), .A2(n3958), .ZN(n4053) );
  NAND2_X1 U4187 ( .A1(n3747), .A2(n6895), .ZN(n4112) );
  NAND2_X1 U4188 ( .A1(n4087), .A2(n4086), .ZN(n6895) );
  NAND2_X1 U4189 ( .A1(n6894), .A2(n6896), .ZN(n3747) );
  NAND3_X1 U4190 ( .A1(n3747), .A2(n6895), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n5174) );
  NAND2_X1 U4191 ( .A1(n3750), .A2(n4115), .ZN(n4129) );
  NAND2_X2 U4192 ( .A1(n4104), .A2(n4103), .ZN(n4115) );
  NAND2_X2 U4193 ( .A1(n3752), .A2(n3683), .ZN(n3988) );
  AND2_X1 U4194 ( .A1(n5528), .A2(n3691), .ZN(n6037) );
  NAND2_X1 U4195 ( .A1(n4603), .A2(n3692), .ZN(n6364) );
  OAI22_X2 U4196 ( .A1(n6922), .A2(n4926), .B1(n4212), .B2(n6647), .ZN(n6928)
         );
  NAND2_X1 U4197 ( .A1(n4059), .A2(n4058), .ZN(n7091) );
  AND2_X2 U4198 ( .A1(n5098), .A2(n5097), .ZN(n5088) );
  AOI22_X1 U4199 ( .A1(n3661), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3913) );
  NOR2_X1 U4200 ( .A1(n5146), .A2(n5246), .ZN(n3921) );
  OR2_X1 U4201 ( .A1(n5161), .A2(n3939), .ZN(n4291) );
  NAND2_X1 U4202 ( .A1(n5421), .A2(n5161), .ZN(n6305) );
  OR2_X1 U4203 ( .A1(n7444), .A2(n5161), .ZN(n5340) );
  INV_X1 U4204 ( .A(n5161), .ZN(n7324) );
  NAND2_X1 U4205 ( .A1(n5100), .A2(n5099), .ZN(n5102) );
  OAI21_X2 U4206 ( .B1(n5137), .B2(n4296), .A(n4295), .ZN(n5098) );
  AND2_X1 U4207 ( .A1(n4996), .A2(n3772), .ZN(n3770) );
  NAND2_X1 U4208 ( .A1(n6311), .A2(n5147), .ZN(n7352) );
  INV_X1 U4209 ( .A(n6876), .ZN(n6868) );
  INV_X1 U4210 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7313) );
  OR2_X1 U4211 ( .A1(n4995), .A2(n4994), .ZN(n3772) );
  OR2_X1 U4212 ( .A1(n7105), .A2(n6812), .ZN(n3773) );
  OR2_X1 U4213 ( .A1(n3998), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3774)
         );
  INV_X1 U4214 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4528) );
  AND3_X1 U4215 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n3776) );
  AND2_X1 U4216 ( .A1(n6498), .A2(n6578), .ZN(n3777) );
  NAND2_X1 U4217 ( .A1(n3650), .A2(n4872), .ZN(n3778) );
  INV_X1 U4218 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4086) );
  NOR2_X1 U4219 ( .A1(n5382), .A2(n5285), .ZN(n3779) );
  AND4_X1 U4220 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3780)
         );
  INV_X1 U4221 ( .A(n3984), .ZN(n3985) );
  NAND2_X1 U4222 ( .A1(n3926), .A2(n6233), .ZN(n3984) );
  NAND2_X1 U4223 ( .A1(n4258), .A2(n4257), .ZN(n4265) );
  NAND2_X1 U4224 ( .A1(n3983), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4237) );
  OR2_X1 U4225 ( .A1(n4172), .A2(n4171), .ZN(n4194) );
  OR2_X1 U4226 ( .A1(n4152), .A2(n4151), .ZN(n4182) );
  AOI22_X1 U4227 ( .A1(n4004), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3786) );
  NAND2_X1 U4228 ( .A1(n3979), .A2(n3978), .ZN(n4933) );
  INV_X1 U4229 ( .A(n3958), .ZN(n3956) );
  INV_X1 U4230 ( .A(n6454), .ZN(n4563) );
  AND2_X1 U4231 ( .A1(n4174), .A2(n4173), .ZN(n4179) );
  OR2_X1 U4232 ( .A1(n4102), .A2(n4101), .ZN(n4133) );
  NAND2_X1 U4233 ( .A1(n4062), .A2(n4061), .ZN(n4280) );
  INV_X1 U4234 ( .A(n4077), .ZN(n4078) );
  OR2_X1 U4235 ( .A1(n4933), .A2(n4963), .ZN(n4798) );
  INV_X1 U4236 ( .A(n6392), .ZN(n4602) );
  INV_X1 U4237 ( .A(n4734), .ZN(n4732) );
  OR2_X1 U4238 ( .A1(n6071), .A2(n4440), .ZN(n4441) );
  INV_X1 U4239 ( .A(n4325), .ZN(n4332) );
  NAND2_X1 U4240 ( .A1(n4916), .A2(n5099), .ZN(n4906) );
  INV_X1 U4241 ( .A(n4085), .ZN(n4087) );
  OR2_X1 U4242 ( .A1(n3954), .A2(n3953), .ZN(n4975) );
  OR2_X1 U4243 ( .A1(n4041), .A2(n4040), .ZN(n4042) );
  NAND2_X1 U4244 ( .A1(n4963), .A2(n5183), .ZN(n4799) );
  NAND2_X1 U4245 ( .A1(n6245), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4727) );
  INV_X1 U4246 ( .A(n5541), .ZN(n4857) );
  INV_X1 U4247 ( .A(n4713), .ZN(n4712) );
  AND2_X1 U4248 ( .A1(n4584), .A2(n4583), .ZN(n6448) );
  AOI21_X1 U4249 ( .B1(n4348), .B2(n4468), .A(n4347), .ZN(n5533) );
  OR2_X1 U4250 ( .A1(n3650), .A2(n6163), .ZN(n6155) );
  INV_X1 U4251 ( .A(n5387), .ZN(n6103) );
  AND2_X1 U4252 ( .A1(n7265), .A2(n7264), .ZN(n7270) );
  INV_X1 U4253 ( .A(n4798), .ZN(n6327) );
  AND2_X1 U4254 ( .A1(n4817), .A2(n7189), .ZN(n7225) );
  NAND2_X1 U4255 ( .A1(n4478), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4496)
         );
  OR2_X1 U4256 ( .A1(n4811), .A2(n4810), .ZN(n4812) );
  NAND2_X1 U4257 ( .A1(n4318), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4327)
         );
  INV_X1 U4258 ( .A(n7289), .ZN(n5205) );
  NAND2_X1 U4259 ( .A1(n4712), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4734)
         );
  NOR2_X1 U4260 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  NAND2_X1 U4261 ( .A1(n4438), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4455)
         );
  AND2_X1 U4262 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n4326), .ZN(n4335)
         );
  INV_X1 U4263 ( .A(n7059), .ZN(n7105) );
  NAND2_X1 U4264 ( .A1(n4976), .A2(n6254), .ZN(n5316) );
  OR2_X1 U4265 ( .A1(n6323), .A2(n3942), .ZN(n6682) );
  AND3_X1 U4266 ( .A1(n5069), .A2(n5068), .A3(n5067), .ZN(n7271) );
  OR2_X1 U4267 ( .A1(n7444), .A2(n7324), .ZN(n5495) );
  NOR2_X1 U4268 ( .A1(n5162), .A2(n5281), .ZN(n7420) );
  NAND2_X1 U4269 ( .A1(n5115), .A2(n5281), .ZN(n7404) );
  OR2_X1 U4270 ( .A1(n7392), .A2(n7324), .ZN(n7389) );
  AND2_X1 U4271 ( .A1(n7296), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4286) );
  NAND2_X1 U4272 ( .A1(n4800), .A2(n4967), .ZN(n6323) );
  NOR2_X1 U4273 ( .A1(n4605), .A2(n7216), .ZN(n4649) );
  AND2_X1 U4274 ( .A1(n5140), .A2(n5048), .ZN(n6953) );
  INV_X1 U4275 ( .A(n7239), .ZN(n7199) );
  INV_X1 U4276 ( .A(n7196), .ZN(n7236) );
  INV_X1 U4277 ( .A(n7192), .ZN(n7178) );
  INV_X1 U4278 ( .A(n6880), .ZN(n6475) );
  INV_X1 U4279 ( .A(n7352), .ZN(n7513) );
  NOR2_X1 U4280 ( .A1(n5206), .A2(n5487), .ZN(n5448) );
  NOR2_X1 U4281 ( .A1(n5140), .A2(READY_N), .ZN(n5206) );
  NAND2_X1 U4282 ( .A1(n4650), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4691)
         );
  AND2_X1 U4283 ( .A1(n3684), .A2(n6871), .ZN(n7356) );
  NAND2_X1 U4284 ( .A1(n4340), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4367)
         );
  INV_X1 U4285 ( .A(n6940), .ZN(n6901) );
  OR2_X1 U4286 ( .A1(n6992), .A2(n4984), .ZN(n4981) );
  INV_X1 U4287 ( .A(n7105), .ZN(n7183) );
  AND2_X1 U4288 ( .A1(n5049), .A2(n7313), .ZN(n7059) );
  INV_X1 U4289 ( .A(n4983), .ZN(n4976) );
  NOR2_X1 U4290 ( .A1(n4983), .A2(n6682), .ZN(n6974) );
  OAI21_X1 U4291 ( .B1(n5339), .B2(n5338), .A(n5337), .ZN(n6302) );
  INV_X1 U4292 ( .A(n5495), .ZN(n7646) );
  INV_X1 U4293 ( .A(n5493), .ZN(n7638) );
  INV_X1 U4294 ( .A(n5167), .ZN(n7637) );
  INV_X1 U4295 ( .A(n7422), .ZN(n7631) );
  OAI211_X1 U4296 ( .C1(n6100), .C2(n7305), .A(n6099), .B(n6098), .ZN(n6288)
         );
  NOR2_X1 U4297 ( .A1(n7404), .A2(n7324), .ZN(n7625) );
  INV_X1 U4298 ( .A(n7389), .ZN(n7617) );
  INV_X1 U4299 ( .A(n7385), .ZN(n7610) );
  AND3_X1 U4300 ( .A1(n5112), .A2(n6058), .A3(n5161), .ZN(n7604) );
  INV_X1 U4301 ( .A(n6107), .ZN(n7453) );
  INV_X1 U4302 ( .A(n6713), .ZN(n7553) );
  NOR2_X1 U4303 ( .A1(n5213), .A2(n5183), .ZN(n7533) );
  INV_X1 U4304 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7334) );
  INV_X1 U4305 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7343) );
  INV_X1 U4306 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7330) );
  OR2_X1 U4307 ( .A1(n6427), .A2(n7195), .ZN(n4923) );
  OR2_X1 U4308 ( .A1(n6953), .A2(n5577), .ZN(n7203) );
  OR3_X1 U4309 ( .A1(n6421), .A2(n5581), .A3(n7296), .ZN(n7196) );
  OR2_X1 U4310 ( .A1(n6421), .A2(n7305), .ZN(n7215) );
  AND2_X1 U4311 ( .A1(n5027), .A2(n3694), .ZN(n5028) );
  NAND2_X1 U4312 ( .A1(n6880), .A2(n6310), .ZN(n6876) );
  INV_X1 U4313 ( .A(n6479), .ZN(n6482) );
  INV_X1 U4314 ( .A(n6755), .ZN(n6784) );
  NAND2_X1 U4315 ( .A1(n5206), .A2(n5226), .ZN(n5492) );
  INV_X1 U4316 ( .A(n6552), .ZN(n6558) );
  NAND2_X1 U4317 ( .A1(n7241), .A2(n4785), .ZN(n6906) );
  AND2_X1 U4318 ( .A1(n5012), .A2(n5011), .ZN(n5013) );
  AND2_X1 U4319 ( .A1(n6630), .A2(n4987), .ZN(n6628) );
  NAND2_X1 U4320 ( .A1(n4976), .A2(n4953), .ZN(n7023) );
  INV_X1 U4321 ( .A(n7065), .ZN(n7029) );
  INV_X1 U4322 ( .A(n6693), .ZN(n7465) );
  INV_X1 U4323 ( .A(n6700), .ZN(n7488) );
  INV_X1 U4324 ( .A(n6731), .ZN(n7652) );
  INV_X1 U4325 ( .A(n7591), .ZN(n6112) );
  INV_X1 U4326 ( .A(n5426), .ZN(n6273) );
  CLKBUF_X1 U4327 ( .A(n6837), .Z(n6826) );
  AOI22_X1 U4328 ( .A1(n3901), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4329 ( .A1(n3670), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3784) );
  NOR2_X4 U4330 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5104) );
  AOI22_X1 U4331 ( .A1(n3669), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3783) );
  AND2_X2 U4332 ( .A1(n5071), .A2(n6671), .ZN(n3961) );
  AOI22_X1 U4333 ( .A1(n3961), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4334 ( .A1(n4009), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3789) );
  AND2_X4 U4335 ( .A1(n5104), .A2(n6671), .ZN(n3909) );
  AOI22_X1 U4336 ( .A1(n3658), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3787) );
  NAND2_X1 U4337 ( .A1(n4009), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3793) );
  NAND2_X1 U4338 ( .A1(n3909), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3792)
         );
  NAND2_X1 U4339 ( .A1(n3793), .A2(n3792), .ZN(n3797) );
  NAND2_X1 U4340 ( .A1(n4003), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U4341 ( .A1(n3666), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3794) );
  NAND2_X1 U4342 ( .A1(n3795), .A2(n3794), .ZN(n3796) );
  NOR2_X1 U4343 ( .A1(n3797), .A2(n3796), .ZN(n3805) );
  NAND2_X1 U4344 ( .A1(n3900), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3799) );
  NAND2_X1 U4345 ( .A1(n3901), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3798) );
  NAND2_X1 U4346 ( .A1(n3799), .A2(n3798), .ZN(n3803) );
  NAND2_X1 U4347 ( .A1(n3961), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3801)
         );
  NAND2_X1 U4348 ( .A1(n3673), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3800)
         );
  NAND2_X1 U4349 ( .A1(n3801), .A2(n3800), .ZN(n3802) );
  NOR2_X1 U4350 ( .A1(n3803), .A2(n3802), .ZN(n3804) );
  NAND2_X1 U4351 ( .A1(n3805), .A2(n3804), .ZN(n3817) );
  NAND2_X1 U4352 ( .A1(n3660), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3809) );
  NAND2_X1 U4353 ( .A1(n3911), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3808) );
  NAND2_X1 U4354 ( .A1(n3912), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3807) );
  NAND2_X1 U4355 ( .A1(n3910), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3806) );
  NAND2_X1 U4356 ( .A1(n3671), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3813)
         );
  NAND2_X1 U4357 ( .A1(n4063), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3812)
         );
  NAND2_X1 U4358 ( .A1(n3665), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3811) );
  NAND2_X1 U4359 ( .A1(n3651), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3810)
         );
  NAND2_X1 U4360 ( .A1(n3926), .A2(n3923), .ZN(n3828) );
  AOI22_X1 U4361 ( .A1(n4003), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4362 ( .A1(n3660), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4363 ( .A1(n3670), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4364 ( .A1(n3961), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4365 ( .A1(n4009), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3652), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4366 ( .A1(n3901), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4367 ( .A1(n3911), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4368 ( .A1(n3669), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3822) );
  NAND2_X4 U4369 ( .A1(n3827), .A2(n3826), .ZN(n6233) );
  NAND2_X1 U4370 ( .A1(n3828), .A2(n6233), .ZN(n3918) );
  NAND2_X1 U4371 ( .A1(n3910), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3831) );
  NAND2_X1 U4372 ( .A1(n3911), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3830) );
  NAND2_X1 U4373 ( .A1(n3912), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3829) );
  NAND3_X1 U4374 ( .A1(n3831), .A2(n3830), .A3(n3829), .ZN(n3832) );
  NAND2_X1 U4375 ( .A1(n4009), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3836) );
  NAND2_X1 U4376 ( .A1(n4003), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3835) );
  NAND2_X1 U4377 ( .A1(n3667), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U4378 ( .A1(n3909), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3833)
         );
  NAND2_X1 U4379 ( .A1(n3900), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3840) );
  NAND2_X1 U4380 ( .A1(n3901), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4381 ( .A1(n3961), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3838)
         );
  NAND2_X1 U4382 ( .A1(n4065), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3837)
         );
  NAND2_X1 U4383 ( .A1(n4063), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3844)
         );
  NAND2_X1 U4384 ( .A1(n3671), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3843)
         );
  NAND2_X1 U4385 ( .A1(n3665), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U4386 ( .A1(n3651), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3841)
         );
  INV_X1 U4387 ( .A(n3938), .ZN(n3887) );
  NAND2_X1 U4388 ( .A1(n4009), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3852) );
  NAND2_X1 U4389 ( .A1(n4003), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3851) );
  NAND2_X1 U4390 ( .A1(n3652), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3850) );
  NAND2_X1 U4391 ( .A1(n3909), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3849)
         );
  NAND2_X1 U4392 ( .A1(n3900), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3856) );
  NAND2_X1 U4393 ( .A1(n3901), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3855) );
  NAND2_X1 U4394 ( .A1(n3961), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3854)
         );
  NAND2_X1 U4395 ( .A1(n3673), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3853)
         );
  NAND2_X1 U4396 ( .A1(n3668), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3860)
         );
  NAND2_X1 U4397 ( .A1(n3670), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3859)
         );
  NAND2_X1 U4398 ( .A1(n3664), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3858) );
  NAND2_X1 U4399 ( .A1(n3675), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3857)
         );
  NAND2_X1 U4400 ( .A1(n3660), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3864) );
  NAND2_X1 U4401 ( .A1(n3658), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4402 ( .A1(n3912), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3862) );
  NAND2_X1 U4403 ( .A1(n3910), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3861) );
  NAND4_X4 U4404 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3983)
         );
  NAND2_X1 U4405 ( .A1(n3900), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3872) );
  NAND2_X1 U4406 ( .A1(n3901), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4407 ( .A1(n3961), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3870)
         );
  NAND2_X1 U4408 ( .A1(n3672), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3869)
         );
  NAND2_X1 U4409 ( .A1(n4003), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3876) );
  NAND2_X1 U4410 ( .A1(n3666), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U4411 ( .A1(n3910), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3874) );
  NAND2_X1 U4412 ( .A1(n3909), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3873)
         );
  NAND2_X1 U4413 ( .A1(n3668), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3880)
         );
  NAND2_X1 U4414 ( .A1(n3670), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3879)
         );
  NAND2_X1 U4415 ( .A1(n3664), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3878) );
  NAND2_X1 U4416 ( .A1(n3651), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3877)
         );
  NAND2_X1 U4417 ( .A1(n4009), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3886) );
  NAND2_X1 U4418 ( .A1(n3912), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3885) );
  NAND2_X1 U4419 ( .A1(n3661), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3884) );
  NAND2_X1 U4420 ( .A1(n3887), .A2(n4017), .ZN(n3899) );
  AOI22_X1 U4421 ( .A1(n4003), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4009), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4422 ( .A1(n4063), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3671), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4423 ( .A1(n3911), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4424 ( .A1(n3901), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4425 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3897)
         );
  AOI22_X1 U4426 ( .A1(n3665), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4427 ( .A1(n3900), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3961), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4428 ( .A1(n3661), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4429 ( .A1(n3666), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3892) );
  NAND4_X1 U4430 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3896)
         );
  AOI22_X1 U4431 ( .A1(n3901), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3900), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4432 ( .A1(n3669), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4433 ( .A1(n3671), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4434 ( .A1(n3961), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4435 ( .A1(n4009), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3652), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4436 ( .A1(n4003), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4437 ( .A1(n3911), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3914) );
  INV_X1 U4438 ( .A(n3918), .ZN(n3919) );
  NAND2_X1 U4439 ( .A1(n7343), .A2(STATE_REG_1__SCAN_IN), .ZN(n7339) );
  NAND2_X1 U4440 ( .A1(n7334), .A2(STATE_REG_2__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4441 ( .A1(n7339), .A2(n3922), .ZN(n4813) );
  OAI21_X1 U4442 ( .B1(n5226), .B2(n4813), .A(n3981), .ZN(n3924) );
  OAI22_X1 U4443 ( .A1(n3939), .A2(n3925), .B1(n3984), .B2(n4018), .ZN(n3927)
         );
  NAND2_X1 U4444 ( .A1(n3927), .A2(n3980), .ZN(n3929) );
  NAND2_X1 U4445 ( .A1(n3938), .A2(n3928), .ZN(n3990) );
  NAND2_X1 U4446 ( .A1(n3929), .A2(n3990), .ZN(n3930) );
  AOI21_X1 U4447 ( .B1(n5146), .B2(n4044), .A(n5226), .ZN(n3944) );
  NAND2_X1 U4448 ( .A1(n3930), .A2(n3944), .ZN(n3931) );
  NAND2_X1 U4449 ( .A1(n3931), .A2(n4963), .ZN(n3954) );
  NAND2_X1 U4450 ( .A1(n3932), .A2(n3954), .ZN(n3933) );
  NAND2_X1 U4451 ( .A1(n3933), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U4452 ( .A1(n4269), .A2(n5146), .ZN(n3934) );
  NAND2_X1 U4453 ( .A1(n4055), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3937) );
  NOR2_X1 U4454 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7294) );
  MUX2_X1 U4455 ( .A(n4286), .B(n4784), .S(n7394), .Z(n3936) );
  INV_X1 U4456 ( .A(n3959), .ZN(n3957) );
  NAND2_X1 U4457 ( .A1(n3938), .A2(n5146), .ZN(n4938) );
  INV_X1 U4458 ( .A(n3939), .ZN(n3941) );
  NOR2_X1 U4459 ( .A1(n3981), .A2(n3925), .ZN(n3940) );
  NAND2_X1 U4460 ( .A1(n3941), .A2(n3940), .ZN(n4479) );
  NAND2_X1 U4461 ( .A1(n4938), .A2(n4479), .ZN(n3943) );
  AOI21_X1 U4462 ( .B1(n3943), .B2(n4044), .A(n3942), .ZN(n3952) );
  INV_X1 U4463 ( .A(n3944), .ZN(n3945) );
  NAND2_X1 U4464 ( .A1(n3945), .A2(n3980), .ZN(n3948) );
  AND2_X1 U4465 ( .A1(n7294), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3946) );
  OAI21_X1 U4466 ( .B1(n4799), .B2(n3939), .A(n3946), .ZN(n3947) );
  AOI21_X1 U4467 ( .B1(n3983), .B2(n3948), .A(n3947), .ZN(n3950) );
  NAND2_X1 U4468 ( .A1(n3950), .A2(n3949), .ZN(n3951) );
  NOR2_X1 U4469 ( .A1(n3952), .A2(n3951), .ZN(n3955) );
  INV_X1 U4470 ( .A(n4288), .ZN(n4239) );
  NOR2_X1 U4471 ( .A1(n4239), .A2(n3942), .ZN(n3953) );
  NAND2_X1 U4472 ( .A1(n3955), .A2(n4975), .ZN(n3958) );
  NAND2_X1 U4473 ( .A1(n3957), .A2(n3956), .ZN(n3960) );
  NAND2_X1 U4474 ( .A1(n3960), .A2(n4053), .ZN(n4292) );
  INV_X1 U4475 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3974) );
  INV_X1 U4476 ( .A(n4061), .ZN(n3972) );
  AOI22_X1 U4477 ( .A1(n3660), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4478 ( .A1(n3961), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4479 ( .A1(n3652), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4480 ( .A1(n4754), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4481 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3971)
         );
  AOI22_X1 U4482 ( .A1(n3669), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3670), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4483 ( .A1(n3901), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4484 ( .A1(n4753), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4485 ( .A1(n3665), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4486 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  NAND2_X1 U4487 ( .A1(n3972), .A2(n4080), .ZN(n3973) );
  OAI211_X1 U4488 ( .C1(n4252), .C2(n3974), .A(n4062), .B(n3973), .ZN(n3975)
         );
  INV_X1 U4489 ( .A(n3975), .ZN(n3976) );
  NAND2_X1 U4490 ( .A1(n4055), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3995) );
  INV_X1 U4491 ( .A(n3977), .ZN(n3979) );
  AND2_X1 U4492 ( .A1(n3981), .A2(n3925), .ZN(n3978) );
  INV_X1 U4493 ( .A(n4813), .ZN(n3987) );
  NOR2_X1 U4494 ( .A1(n3983), .A2(n5226), .ZN(n6328) );
  INV_X1 U4495 ( .A(n5142), .ZN(n3986) );
  NAND2_X1 U4496 ( .A1(n3986), .A2(n3985), .ZN(n4949) );
  NOR2_X1 U4497 ( .A1(n4799), .A2(n5226), .ZN(n3991) );
  NAND2_X1 U4498 ( .A1(n4800), .A2(n3991), .ZN(n5074) );
  INV_X1 U4499 ( .A(n4784), .ZN(n4090) );
  XNOR2_X1 U4500 ( .A(n7394), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5382)
         );
  INV_X1 U4501 ( .A(n4286), .ZN(n4089) );
  AND2_X1 U4502 ( .A1(n4089), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3994)
         );
  NAND3_X1 U4503 ( .A1(n3995), .A2(n3996), .A3(n3997), .ZN(n4051) );
  INV_X1 U4504 ( .A(n3996), .ZN(n3999) );
  INV_X1 U4505 ( .A(n3997), .ZN(n3998) );
  NAND2_X1 U4506 ( .A1(n3999), .A2(n3774), .ZN(n4000) );
  AOI22_X1 U4507 ( .A1(n3911), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4508 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4754), .B1(n3901), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4509 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3671), .B1(n4756), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4510 ( .A1(n3661), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4511 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4015)
         );
  AOI22_X1 U4512 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3664), .B1(n3961), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4513 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3668), .B1(n3653), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4514 ( .A1(n4753), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4515 ( .A1(n3909), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4516 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4014)
         );
  XNOR2_X1 U4517 ( .A(n4016), .B(n4081), .ZN(n4020) );
  NAND3_X1 U4518 ( .A1(n3980), .A2(n4018), .A3(n4044), .ZN(n4019) );
  AOI21_X1 U4519 ( .B1(n4020), .B2(n4017), .A(n4019), .ZN(n4021) );
  INV_X1 U4520 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4034) );
  AOI21_X1 U4521 ( .B1(n4963), .B2(n4081), .A(n7313), .ZN(n4033) );
  AOI22_X1 U4522 ( .A1(n4755), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4523 ( .A1(n3668), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4524 ( .A1(n3670), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4024) );
  INV_X1 U4525 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4526 ( .A1(n3961), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U4527 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4032)
         );
  AOI22_X1 U4528 ( .A1(n4753), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4529 ( .A1(n3661), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4530 ( .A1(n3658), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4531 ( .A1(n4754), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4027) );
  NAND4_X1 U4532 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4031)
         );
  NAND2_X1 U4533 ( .A1(n3925), .A2(n4206), .ZN(n4203) );
  OAI211_X1 U4534 ( .C1(n4252), .C2(n4034), .A(n4033), .B(n4203), .ZN(n4039)
         );
  INV_X1 U4535 ( .A(n4062), .ZN(n4037) );
  INV_X1 U4536 ( .A(n4206), .ZN(n4035) );
  XNOR2_X1 U4537 ( .A(n4035), .B(n4081), .ZN(n4036) );
  NAND2_X1 U4538 ( .A1(n4037), .A2(n4036), .ZN(n4038) );
  NOR2_X1 U4539 ( .A1(n4039), .A2(n4038), .ZN(n4041) );
  AND2_X1 U4540 ( .A1(n4039), .A2(n4038), .ZN(n4040) );
  NAND2_X1 U4541 ( .A1(n5161), .A2(n4259), .ZN(n4047) );
  NAND2_X1 U4542 ( .A1(n4963), .A2(n4044), .ZN(n4082) );
  OAI21_X1 U4543 ( .B1(n4957), .B2(n4081), .A(n4082), .ZN(n4045) );
  INV_X1 U4544 ( .A(n4045), .ZN(n4046) );
  NAND2_X1 U4545 ( .A1(n4047), .A2(n4046), .ZN(n5125) );
  AND2_X1 U4546 ( .A1(n5125), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5269)
         );
  OAI21_X1 U4547 ( .B1(n5271), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n5269), 
        .ZN(n4049) );
  NAND2_X1 U4548 ( .A1(n5271), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4048)
         );
  NAND2_X1 U4549 ( .A1(n4049), .A2(n4048), .ZN(n4085) );
  NAND2_X1 U4550 ( .A1(n4085), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6894)
         );
  INV_X1 U4551 ( .A(n4050), .ZN(n4054) );
  INV_X1 U4552 ( .A(n4051), .ZN(n4052) );
  AOI21_X2 U4553 ( .B1(n4054), .B2(n4053), .A(n4052), .ZN(n4059) );
  NAND2_X1 U4554 ( .A1(n4055), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4057) );
  NAND2_X1 U4555 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7433) );
  XNOR2_X1 U4556 ( .A(n7433), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5168)
         );
  AOI22_X1 U4557 ( .A1(n4090), .A2(n5168), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4089), .ZN(n4056) );
  NAND2_X1 U4558 ( .A1(n4057), .A2(n4056), .ZN(n4058) );
  OR2_X1 U4559 ( .A1(n4059), .A2(n4058), .ZN(n4060) );
  AOI22_X1 U4560 ( .A1(n4755), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4561 ( .A1(n3663), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U4562 ( .A1(n3671), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U4563 ( .A1(n3961), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4066) );
  NAND4_X1 U4564 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4075)
         );
  AOI22_X1 U4565 ( .A1(n4753), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3652), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4566 ( .A1(n4004), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4567 ( .A1(n3658), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4568 ( .A1(n4754), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4070) );
  NAND4_X1 U4569 ( .A1(n4073), .A2(n4072), .A3(n4071), .A4(n4070), .ZN(n4074)
         );
  AOI22_X1 U4570 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n4269), .B1(n4280), 
        .B2(n4105), .ZN(n4076) );
  OAI21_X2 U4571 ( .B1(n5163), .B2(STATE2_REG_0__SCAN_IN), .A(n4076), .ZN(
        n4079) );
  NAND2_X2 U4572 ( .A1(n4079), .A2(n4078), .ZN(n4114) );
  AND2_X2 U4573 ( .A1(n4114), .A2(n5159), .ZN(n4289) );
  NAND2_X1 U4574 ( .A1(n4081), .A2(n4080), .ZN(n4107) );
  XNOR2_X1 U4575 ( .A(n4107), .B(n4105), .ZN(n4083) );
  OAI21_X1 U4576 ( .B1(n4083), .B2(n4957), .A(n4082), .ZN(n4084) );
  INV_X1 U4577 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4111) );
  NAND2_X1 U4578 ( .A1(n4055), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4092) );
  NOR3_X1 U4579 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6251), .A3(n7448), 
        .ZN(n7414) );
  NAND2_X1 U4580 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7414), .ZN(n7408) );
  NAND2_X1 U4581 ( .A1(n7268), .A2(n7408), .ZN(n4088) );
  NAND3_X1 U4582 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5424) );
  NOR2_X1 U4583 ( .A1(n7394), .A2(n5424), .ZN(n5426) );
  AOI22_X1 U4584 ( .A1(n4090), .A2(n5285), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4089), .ZN(n4091) );
  NAND2_X1 U4585 ( .A1(n5110), .A2(n7313), .ZN(n4104) );
  AOI22_X1 U4586 ( .A1(n3660), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U4587 ( .A1(n3663), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3670), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U4588 ( .A1(n4753), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3652), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U4589 ( .A1(n3665), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4093) );
  NAND4_X1 U4590 ( .A1(n4096), .A2(n4095), .A3(n4094), .A4(n4093), .ZN(n4102)
         );
  AOI22_X1 U4591 ( .A1(n4755), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U4592 ( .A1(n4761), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U4593 ( .A1(n4762), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U4594 ( .A1(n4754), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4097) );
  NAND4_X1 U4595 ( .A1(n4100), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4101)
         );
  AOI22_X1 U4596 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n4269), .B1(n4280), 
        .B2(n4133), .ZN(n4103) );
  XNOR2_X2 U4597 ( .A(n4115), .B(n4114), .ZN(n5112) );
  INV_X1 U4598 ( .A(n4105), .ZN(n4106) );
  NAND2_X1 U4599 ( .A1(n4107), .A2(n4106), .ZN(n4134) );
  INV_X1 U4600 ( .A(n4133), .ZN(n4108) );
  XNOR2_X1 U4601 ( .A(n4134), .B(n4108), .ZN(n4109) );
  AND2_X1 U4602 ( .A1(n4109), .A2(n4017), .ZN(n4110) );
  AOI21_X1 U4603 ( .B1(n5112), .B2(n4259), .A(n4110), .ZN(n5177) );
  NAND2_X1 U4604 ( .A1(n5174), .A2(n5177), .ZN(n4113) );
  NAND2_X1 U4605 ( .A1(n4112), .A2(n4111), .ZN(n5175) );
  NAND2_X1 U4606 ( .A1(n4269), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U4607 ( .A1(n4755), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U4608 ( .A1(n3663), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U4609 ( .A1(n3671), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U4610 ( .A1(n4761), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4116) );
  NAND4_X1 U4611 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(n4125)
         );
  AOI22_X1 U4612 ( .A1(n4753), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3652), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U4613 ( .A1(n3661), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U4614 ( .A1(n3911), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U4615 ( .A1(n4754), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4120) );
  NAND4_X1 U4616 ( .A1(n4123), .A2(n4122), .A3(n4121), .A4(n4120), .ZN(n4124)
         );
  NAND2_X1 U4617 ( .A1(n4280), .A2(n4137), .ZN(n4126) );
  NAND2_X1 U4618 ( .A1(n4129), .A2(n4130), .ZN(n4131) );
  NAND2_X1 U4619 ( .A1(n4156), .A2(n4131), .ZN(n4324) );
  INV_X1 U4620 ( .A(n4324), .ZN(n4132) );
  NAND2_X1 U4621 ( .A1(n4134), .A2(n4133), .ZN(n4136) );
  INV_X1 U4622 ( .A(n4136), .ZN(n4138) );
  INV_X1 U4623 ( .A(n4137), .ZN(n4135) );
  OR2_X1 U4624 ( .A1(n4136), .A2(n4135), .ZN(n4181) );
  OAI211_X1 U4625 ( .C1(n4138), .C2(n4137), .A(n4017), .B(n4181), .ZN(n4139)
         );
  NAND2_X1 U4626 ( .A1(n4141), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4142)
         );
  OAI21_X1 U4627 ( .B1(n5221), .B2(n5222), .A(n4142), .ZN(n5319) );
  INV_X1 U4628 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U4629 ( .A1(n4004), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U4630 ( .A1(n3663), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3671), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U4631 ( .A1(n4756), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U4632 ( .A1(n4755), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4143) );
  NAND4_X1 U4633 ( .A1(n4146), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(n4152)
         );
  AOI22_X1 U4634 ( .A1(n4754), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U4635 ( .A1(n3664), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U4636 ( .A1(n4753), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U4637 ( .A1(n3909), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U4638 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4151)
         );
  NAND2_X1 U4639 ( .A1(n4280), .A2(n4182), .ZN(n4153) );
  OAI21_X1 U4640 ( .B1(n4154), .B2(n4252), .A(n4153), .ZN(n4175) );
  INV_X1 U4641 ( .A(n4175), .ZN(n4155) );
  NAND2_X1 U4642 ( .A1(n4156), .A2(n4155), .ZN(n4157) );
  INV_X1 U4643 ( .A(n4156), .ZN(n4178) );
  NAND2_X1 U4644 ( .A1(n4178), .A2(n4175), .ZN(n4180) );
  NAND2_X1 U4645 ( .A1(n4157), .A2(n4180), .ZN(n4325) );
  INV_X1 U4646 ( .A(n4259), .ZN(n4202) );
  XNOR2_X1 U4647 ( .A(n4181), .B(n4182), .ZN(n4158) );
  NAND2_X1 U4648 ( .A1(n4158), .A2(n4017), .ZN(n4159) );
  INV_X1 U4649 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5320) );
  XNOR2_X1 U4650 ( .A(n4160), .B(n5320), .ZN(n5318) );
  NAND2_X1 U4651 ( .A1(n5319), .A2(n5318), .ZN(n4162) );
  NAND2_X1 U4652 ( .A1(n4160), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4161)
         );
  NAND2_X1 U4653 ( .A1(n4162), .A2(n4161), .ZN(n5434) );
  NAND2_X1 U4654 ( .A1(n4269), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U4655 ( .A1(n4755), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U4656 ( .A1(n3663), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4657 ( .A1(n3670), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4658 ( .A1(n4761), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4163) );
  NAND4_X1 U4659 ( .A1(n4166), .A2(n4165), .A3(n4164), .A4(n4163), .ZN(n4172)
         );
  AOI22_X1 U4660 ( .A1(n4753), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U4661 ( .A1(n3660), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U4662 ( .A1(n3911), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4663 ( .A1(n4754), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U4664 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4171)
         );
  NAND2_X1 U4665 ( .A1(n4280), .A2(n4194), .ZN(n4173) );
  NAND2_X1 U4666 ( .A1(n4180), .A2(n4179), .ZN(n4348) );
  NAND3_X1 U4667 ( .A1(n4191), .A2(n4348), .A3(n4259), .ZN(n4186) );
  INV_X1 U4668 ( .A(n4181), .ZN(n4183) );
  NAND2_X1 U4669 ( .A1(n4183), .A2(n4182), .ZN(n4193) );
  XNOR2_X1 U4670 ( .A(n4193), .B(n4194), .ZN(n4184) );
  NAND2_X1 U4671 ( .A1(n4184), .A2(n4017), .ZN(n4185) );
  NAND2_X1 U4672 ( .A1(n4186), .A2(n4185), .ZN(n4187) );
  OR2_X1 U4673 ( .A1(n4187), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5436)
         );
  NAND2_X1 U4674 ( .A1(n5434), .A2(n5436), .ZN(n4188) );
  NAND2_X1 U4675 ( .A1(n4187), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5435)
         );
  NAND2_X1 U4676 ( .A1(n4188), .A2(n5435), .ZN(n6911) );
  NAND2_X1 U4677 ( .A1(n4280), .A2(n4206), .ZN(n4189) );
  OAI21_X1 U4678 ( .B1(n4022), .B2(n4252), .A(n4189), .ZN(n4190) );
  INV_X1 U4679 ( .A(n4339), .ZN(n4192) );
  OR2_X1 U4680 ( .A1(n4192), .A2(n4202), .ZN(n4198) );
  INV_X1 U4681 ( .A(n4193), .ZN(n4195) );
  NAND2_X1 U4682 ( .A1(n4195), .A2(n4194), .ZN(n4205) );
  XNOR2_X1 U4683 ( .A(n4205), .B(n4206), .ZN(n4196) );
  NAND2_X1 U4684 ( .A1(n4196), .A2(n4017), .ZN(n4197) );
  NAND2_X1 U4685 ( .A1(n4198), .A2(n4197), .ZN(n4200) );
  INV_X1 U4686 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4199) );
  XNOR2_X1 U4687 ( .A(n4200), .B(n4199), .ZN(n6910) );
  NAND2_X1 U4688 ( .A1(n6911), .A2(n6910), .ZN(n6913) );
  NAND2_X1 U4689 ( .A1(n4200), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4201)
         );
  NAND2_X1 U4690 ( .A1(n6913), .A2(n4201), .ZN(n5546) );
  NOR2_X1 U4691 ( .A1(n4203), .A2(n4202), .ZN(n4204) );
  INV_X1 U4692 ( .A(n4205), .ZN(n4207) );
  NAND3_X1 U4693 ( .A1(n4207), .A2(n4017), .A3(n4206), .ZN(n4208) );
  NAND2_X1 U4694 ( .A1(n4221), .A2(n4208), .ZN(n4210) );
  INV_X1 U4695 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4209) );
  XNOR2_X1 U4696 ( .A(n4210), .B(n4209), .ZN(n5545) );
  NAND2_X1 U4697 ( .A1(n5546), .A2(n5545), .ZN(n5544) );
  NAND2_X1 U4698 ( .A1(n4210), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4211)
         );
  XNOR2_X1 U4699 ( .A(n3650), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5995)
         );
  INV_X1 U4700 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7040) );
  OR2_X1 U4701 ( .A1(n3650), .A2(n7040), .ZN(n4213) );
  INV_X1 U4702 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4215) );
  INV_X1 U4703 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4214) );
  INV_X1 U4704 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U4705 ( .A1(n4216), .A2(n6155), .ZN(n4218) );
  NAND2_X1 U4706 ( .A1(n3650), .A2(n4214), .ZN(n4217) );
  XNOR2_X1 U4707 ( .A(n3650), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6178)
         );
  INV_X1 U4708 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4219) );
  INV_X1 U4709 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6662) );
  NOR2_X1 U4710 ( .A1(n3650), .A2(n6662), .ZN(n6567) );
  INV_X1 U4711 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4872) );
  NOR2_X1 U4712 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4220) );
  AND2_X1 U4713 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6644) );
  NAND2_X1 U4714 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U4715 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4988) );
  NOR2_X1 U4716 ( .A1(n6622), .A2(n4988), .ZN(n5006) );
  AND2_X1 U4717 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U4718 ( .A1(n5006), .A2(n6647), .ZN(n4222) );
  AND2_X1 U4719 ( .A1(n3650), .A2(n4222), .ZN(n4226) );
  INV_X1 U4720 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6629) );
  INV_X1 U4721 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6536) );
  INV_X1 U4722 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6627) );
  INV_X1 U4723 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4991) );
  NAND4_X1 U4724 ( .A1(n6629), .A2(n6536), .A3(n6627), .A4(n4991), .ZN(n4223)
         );
  INV_X1 U4725 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4883) );
  INV_X1 U4726 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U4727 ( .A1(n4883), .A2(n6545), .ZN(n6645) );
  NOR2_X1 U4728 ( .A1(n4223), .A2(n6645), .ZN(n4224) );
  INV_X1 U4729 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6934) );
  NOR2_X1 U4730 ( .A1(n3650), .A2(n6934), .ZN(n4228) );
  NAND2_X1 U4731 ( .A1(n3650), .A2(n6934), .ZN(n4227) );
  INV_X1 U4732 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U4733 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5008) );
  INV_X1 U4734 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6586) );
  NOR2_X1 U4735 ( .A1(n5008), .A2(n6586), .ZN(n5004) );
  NOR2_X1 U4736 ( .A1(n3650), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6498)
         );
  AOI21_X1 U4737 ( .B1(n4997), .B2(n5004), .A(n6498), .ZN(n4231) );
  INV_X1 U4738 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U4739 ( .A1(n6507), .A2(n6612), .ZN(n6221) );
  NOR2_X1 U4740 ( .A1(n6221), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4230)
         );
  NAND2_X1 U4741 ( .A1(n4229), .A2(n4230), .ZN(n4998) );
  XNOR2_X1 U4742 ( .A(n4232), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6582)
         );
  INV_X1 U4743 ( .A(n4280), .ZN(n4235) );
  XNOR2_X1 U4744 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4248) );
  NAND2_X1 U4745 ( .A1(n7394), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4234) );
  XNOR2_X1 U4746 ( .A(n4248), .B(n4247), .ZN(n4803) );
  NAND2_X1 U4747 ( .A1(n4269), .A2(n4803), .ZN(n4233) );
  OAI211_X1 U4748 ( .C1(n4235), .C2(n3942), .A(n4233), .B(n4018), .ZN(n4242)
         );
  INV_X1 U4749 ( .A(n4242), .ZN(n4246) );
  OAI21_X1 U4750 ( .B1(n7313), .B2(n4803), .A(n4271), .ZN(n4243) );
  INV_X1 U4751 ( .A(n4243), .ZN(n4245) );
  OAI21_X1 U4752 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7394), .A(n4234), 
        .ZN(n4236) );
  NOR2_X1 U4753 ( .A1(n4235), .A2(n4236), .ZN(n4241) );
  INV_X1 U4754 ( .A(n6328), .ZN(n5571) );
  OAI21_X1 U4755 ( .B1(n3981), .B2(n5226), .A(n5571), .ZN(n4261) );
  INV_X1 U4756 ( .A(n4236), .ZN(n4238) );
  AOI21_X1 U4757 ( .B1(n4239), .B2(n4238), .A(n4237), .ZN(n4240) );
  OAI222_X1 U4758 ( .A1(n4243), .A2(n4242), .B1(n4283), .B2(n4241), .C1(n4261), 
        .C2(n4240), .ZN(n4244) );
  OAI21_X1 U4759 ( .B1(n4246), .B2(n4245), .A(n4244), .ZN(n4263) );
  NAND2_X1 U4760 ( .A1(n4248), .A2(n4247), .ZN(n4250) );
  NAND2_X1 U4761 ( .A1(n7448), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4249) );
  NAND2_X1 U4762 ( .A1(n4250), .A2(n4249), .ZN(n4256) );
  XNOR2_X1 U4763 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4255) );
  XNOR2_X1 U4764 ( .A(n4256), .B(n4255), .ZN(n4802) );
  INV_X1 U4765 ( .A(n4802), .ZN(n4253) );
  INV_X1 U4766 ( .A(n4261), .ZN(n4251) );
  NAND2_X1 U4767 ( .A1(n4280), .A2(n4253), .ZN(n4254) );
  OAI211_X1 U4768 ( .C1(n4253), .C2(n4252), .A(n4251), .B(n4254), .ZN(n4262)
         );
  INV_X1 U4769 ( .A(n4254), .ZN(n4260) );
  NAND2_X1 U4770 ( .A1(n4256), .A2(n4255), .ZN(n4258) );
  NAND2_X1 U4771 ( .A1(n6251), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4257) );
  XNOR2_X1 U4772 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4264) );
  XNOR2_X1 U4773 ( .A(n4265), .B(n4264), .ZN(n4801) );
  AOI222_X1 U4774 ( .A1(n4263), .A2(n4262), .B1(n4261), .B2(n4260), .C1(n4801), 
        .C2(n4259), .ZN(n4273) );
  INV_X1 U4775 ( .A(n4801), .ZN(n4270) );
  NAND2_X1 U4776 ( .A1(n4265), .A2(n4264), .ZN(n4267) );
  NAND2_X1 U4777 ( .A1(n7268), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U4778 ( .A1(n4267), .A2(n4266), .ZN(n4277) );
  AOI21_X1 U4779 ( .B1(n4270), .B2(n4806), .A(n4269), .ZN(n4272) );
  OAI22_X1 U4780 ( .A1(n4273), .A2(n4272), .B1(n4271), .B2(n4806), .ZN(n4274)
         );
  AOI21_X1 U4781 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7313), .A(n4274), 
        .ZN(n4282) );
  NAND2_X1 U4782 ( .A1(n4275), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U4783 ( .A1(n4277), .A2(n4276), .ZN(n4278) );
  NAND2_X1 U4784 ( .A1(n4280), .A2(n4805), .ZN(n4281) );
  NAND2_X1 U4785 ( .A1(n4282), .A2(n4281), .ZN(n4285) );
  NAND2_X1 U4786 ( .A1(n4479), .A2(n4963), .ZN(n4287) );
  AND2_X1 U4787 ( .A1(n4962), .A2(n4287), .ZN(n4939) );
  NAND2_X1 U4788 ( .A1(n4289), .A2(n4468), .ZN(n4290) );
  NAND2_X1 U4789 ( .A1(n7295), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4643) );
  NAND2_X1 U4790 ( .A1(n4291), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U4791 ( .A1(n3985), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4321) );
  INV_X1 U4792 ( .A(n4468), .ZN(n4425) );
  NOR2_X4 U4793 ( .A1(n6233), .A2(n7295), .ZN(n4794) );
  AOI22_X1 U4794 ( .A1(n4794), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n7295), .ZN(n4293) );
  NAND2_X1 U4795 ( .A1(n7295), .A2(n7330), .ZN(n4317) );
  AOI22_X1 U4796 ( .A1(n4794), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n7295), .ZN(n4298) );
  NAND2_X1 U4797 ( .A1(n5087), .A2(n5088), .ZN(n4307) );
  INV_X1 U4798 ( .A(n4321), .ZN(n4301) );
  NAND2_X1 U4799 ( .A1(n4301), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4306) );
  INV_X1 U4800 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4303) );
  OAI21_X1 U4801 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4311), .ZN(n7085) );
  NAND2_X1 U4802 ( .A1(n4777), .A2(n7085), .ZN(n4302) );
  OAI21_X1 U4803 ( .B1(n4303), .B2(n4643), .A(n4302), .ZN(n4304) );
  AOI21_X1 U4804 ( .B1(n4794), .B2(EAX_REG_2__SCAN_IN), .A(n4304), .ZN(n4305)
         );
  AND2_X1 U4805 ( .A1(n4306), .A2(n4305), .ZN(n5089) );
  NAND2_X1 U4806 ( .A1(n4307), .A2(n5089), .ZN(n4309) );
  NAND2_X1 U4807 ( .A1(n4309), .A2(n4308), .ZN(n5086) );
  INV_X1 U4808 ( .A(n4311), .ZN(n4313) );
  INV_X1 U4809 ( .A(n4318), .ZN(n4312) );
  OAI21_X1 U4810 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n4313), .A(n4312), 
        .ZN(n6008) );
  AOI22_X1 U4811 ( .A1(n4777), .A2(n6008), .B1(n4793), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U4812 ( .A1(n4794), .A2(EAX_REG_3__SCAN_IN), .ZN(n4314) );
  OAI211_X1 U4813 ( .C1(n4321), .C2(n4310), .A(n4315), .B(n4314), .ZN(n4316)
         );
  AOI21_X1 U4814 ( .B1(n5112), .B2(n4468), .A(n4316), .ZN(n5132) );
  OAI21_X1 U4815 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n4318), .A(n4327), 
        .ZN(n7096) );
  OAI21_X1 U4816 ( .B1(n7330), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7295), 
        .ZN(n4320) );
  NAND2_X1 U4817 ( .A1(n4794), .A2(EAX_REG_4__SCAN_IN), .ZN(n4319) );
  OAI211_X1 U4818 ( .C1(n4321), .C2(n7250), .A(n4320), .B(n4319), .ZN(n4322)
         );
  OAI21_X1 U4819 ( .B1(n4317), .B2(n7096), .A(n4322), .ZN(n4323) );
  OAI21_X1 U4820 ( .B1(n4324), .B2(n4425), .A(n4323), .ZN(n5151) );
  NAND2_X1 U4821 ( .A1(n5131), .A2(n5151), .ZN(n5149) );
  INV_X1 U4822 ( .A(n5149), .ZN(n4334) );
  INV_X1 U4823 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4330) );
  INV_X1 U4824 ( .A(n4335), .ZN(n4341) );
  INV_X1 U4825 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n7106) );
  NAND2_X1 U4826 ( .A1(n7106), .A2(n4327), .ZN(n4328) );
  NAND2_X1 U4827 ( .A1(n4341), .A2(n4328), .ZN(n7119) );
  AOI22_X1 U4828 ( .A1(n7119), .A2(n4777), .B1(n4793), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4329) );
  OAI21_X1 U4829 ( .B1(n4751), .B2(n4330), .A(n4329), .ZN(n4331) );
  INV_X1 U4830 ( .A(n5256), .ZN(n4333) );
  NAND2_X1 U4831 ( .A1(n4334), .A2(n4333), .ZN(n5254) );
  INV_X1 U4832 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4337) );
  OAI21_X1 U4833 ( .B1(n4340), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4367), 
        .ZN(n7141) );
  AOI22_X1 U4834 ( .A1(n7141), .A2(n4777), .B1(n4793), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4336) );
  OAI21_X1 U4835 ( .B1(n4751), .B2(n4337), .A(n4336), .ZN(n4338) );
  AOI21_X1 U4836 ( .B1(n4339), .B2(n4468), .A(n4338), .ZN(n5535) );
  INV_X1 U4837 ( .A(n5535), .ZN(n4350) );
  INV_X1 U4838 ( .A(n4340), .ZN(n4343) );
  INV_X1 U4839 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U4840 ( .A1(n4341), .A2(n4344), .ZN(n4342) );
  NAND2_X1 U4841 ( .A1(n4343), .A2(n4342), .ZN(n7128) );
  INV_X1 U4842 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4345) );
  OAI22_X1 U4843 ( .A1(n4751), .A2(n4345), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4344), .ZN(n4346) );
  MUX2_X1 U4844 ( .A(n7128), .B(n4346), .S(n4317), .Z(n4347) );
  INV_X1 U4845 ( .A(n5533), .ZN(n4349) );
  NAND2_X1 U4846 ( .A1(n4350), .A2(n4349), .ZN(n4351) );
  AOI22_X1 U4847 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4753), .B1(n3911), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4355) );
  AOI22_X1 U4848 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3663), .B1(n3671), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4354) );
  AOI22_X1 U4849 ( .A1(n3652), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4353) );
  AOI22_X1 U4850 ( .A1(n3661), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4352) );
  NAND4_X1 U4851 ( .A1(n4355), .A2(n4354), .A3(n4353), .A4(n4352), .ZN(n4361)
         );
  AOI22_X1 U4852 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3651), .B1(n3665), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U4853 ( .A1(n4754), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U4854 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n4755), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4357) );
  AOI22_X1 U4855 ( .A1(n4761), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4356) );
  NAND4_X1 U4856 ( .A1(n4359), .A2(n4358), .A3(n4357), .A4(n4356), .ZN(n4360)
         );
  OAI21_X1 U4857 ( .B1(n4361), .B2(n4360), .A(n4468), .ZN(n4366) );
  NAND2_X1 U4858 ( .A1(n4794), .A2(EAX_REG_8__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U4859 ( .A1(n4793), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4364)
         );
  INV_X1 U4860 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4362) );
  XNOR2_X1 U4861 ( .A(n4367), .B(n4362), .ZN(n5983) );
  NAND2_X1 U4862 ( .A1(n5983), .A2(n4777), .ZN(n4363) );
  NAND4_X1 U4863 ( .A1(n4366), .A2(n4365), .A3(n4364), .A4(n4363), .ZN(n5526)
         );
  XOR2_X1 U4864 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4381), .Z(n5588) );
  AOI22_X1 U4865 ( .A1(n4754), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4371) );
  AOI22_X1 U4866 ( .A1(n4756), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4370) );
  AOI22_X1 U4867 ( .A1(n3665), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U4868 ( .A1(n4755), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4368) );
  NAND4_X1 U4869 ( .A1(n4371), .A2(n4370), .A3(n4369), .A4(n4368), .ZN(n4377)
         );
  AOI22_X1 U4870 ( .A1(n3663), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3671), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4375) );
  AOI22_X1 U4871 ( .A1(n3661), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4374) );
  AOI22_X1 U4872 ( .A1(n3658), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U4873 ( .A1(n3652), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4372) );
  NAND4_X1 U4874 ( .A1(n4375), .A2(n4374), .A3(n4373), .A4(n4372), .ZN(n4376)
         );
  OR2_X1 U4875 ( .A1(n4377), .A2(n4376), .ZN(n4378) );
  AOI22_X1 U4876 ( .A1(n4468), .A2(n4378), .B1(n4793), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U4877 ( .A1(n4794), .A2(EAX_REG_9__SCAN_IN), .ZN(n4379) );
  OAI211_X1 U4878 ( .C1(n5588), .C2(n4317), .A(n4380), .B(n4379), .ZN(n5539)
         );
  XNOR2_X1 U4879 ( .A(n4397), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6135)
         );
  AOI22_X1 U4880 ( .A1(n3911), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U4881 ( .A1(n4755), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4384) );
  AOI22_X1 U4882 ( .A1(n3664), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U4883 ( .A1(n4754), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4382) );
  NAND4_X1 U4884 ( .A1(n4385), .A2(n4384), .A3(n4383), .A4(n4382), .ZN(n4391)
         );
  AOI22_X1 U4885 ( .A1(n3663), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3671), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4389) );
  AOI22_X1 U4886 ( .A1(n3660), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4388) );
  AOI22_X1 U4887 ( .A1(n3652), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U4888 ( .A1(n4761), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4386) );
  NAND4_X1 U4889 ( .A1(n4389), .A2(n4388), .A3(n4387), .A4(n4386), .ZN(n4390)
         );
  OAI21_X1 U4890 ( .B1(n4391), .B2(n4390), .A(n4468), .ZN(n4394) );
  NAND2_X1 U4891 ( .A1(n4794), .A2(EAX_REG_10__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U4892 ( .A1(n4793), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4392)
         );
  NAND3_X1 U4893 ( .A1(n4394), .A2(n4393), .A3(n4392), .ZN(n4395) );
  AOI21_X1 U4894 ( .B1(n6135), .B2(n4777), .A(n4395), .ZN(n6021) );
  XOR2_X1 U4895 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4422), .Z(n6047) );
  INV_X1 U4896 ( .A(n6047), .ZN(n6089) );
  AOI22_X1 U4897 ( .A1(n3660), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U4898 ( .A1(n4755), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4400) );
  AOI22_X1 U4899 ( .A1(n4754), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4399) );
  AOI22_X1 U4900 ( .A1(n4761), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4398) );
  NAND4_X1 U4901 ( .A1(n4401), .A2(n4400), .A3(n4399), .A4(n4398), .ZN(n4407)
         );
  AOI22_X1 U4902 ( .A1(n4753), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U4903 ( .A1(n3663), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4404) );
  AOI22_X1 U4904 ( .A1(n3670), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4403) );
  AOI22_X1 U4905 ( .A1(n4762), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4402) );
  NAND4_X1 U4906 ( .A1(n4405), .A2(n4404), .A3(n4403), .A4(n4402), .ZN(n4406)
         );
  OAI21_X1 U4907 ( .B1(n4407), .B2(n4406), .A(n4468), .ZN(n4410) );
  NAND2_X1 U4908 ( .A1(n4794), .A2(EAX_REG_11__SCAN_IN), .ZN(n4409) );
  NAND2_X1 U4909 ( .A1(n4793), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4408)
         );
  NAND3_X1 U4910 ( .A1(n4410), .A2(n4409), .A3(n4408), .ZN(n4411) );
  AOI21_X1 U4911 ( .B1(n6089), .B2(n4777), .A(n4411), .ZN(n6038) );
  AOI22_X1 U4912 ( .A1(n4004), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4913 ( .A1(n4754), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4755), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U4914 ( .A1(n4753), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U4915 ( .A1(n3651), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4412) );
  NAND4_X1 U4916 ( .A1(n4415), .A2(n4414), .A3(n4413), .A4(n4412), .ZN(n4421)
         );
  AOI22_X1 U4917 ( .A1(n3663), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3671), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4419) );
  AOI22_X1 U4918 ( .A1(n4761), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U4919 ( .A1(n3666), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4417) );
  AOI22_X1 U4920 ( .A1(n4756), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4416) );
  NAND4_X1 U4921 ( .A1(n4419), .A2(n4418), .A3(n4417), .A4(n4416), .ZN(n4420)
         );
  NOR2_X1 U4922 ( .A1(n4421), .A2(n4420), .ZN(n4426) );
  XNOR2_X1 U4923 ( .A(n4438), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6171)
         );
  NAND2_X1 U4924 ( .A1(n6171), .A2(n4777), .ZN(n4424) );
  AOI22_X1 U4925 ( .A1(n4794), .A2(EAX_REG_12__SCAN_IN), .B1(n4793), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4423) );
  OAI211_X1 U4926 ( .C1(n4426), .C2(n4425), .A(n4424), .B(n4423), .ZN(n6072)
         );
  AOI22_X1 U4927 ( .A1(n3660), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U4928 ( .A1(n4754), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4429) );
  AOI22_X1 U4929 ( .A1(n3663), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U4930 ( .A1(n4756), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4427) );
  NAND4_X1 U4931 ( .A1(n4430), .A2(n4429), .A3(n4428), .A4(n4427), .ZN(n4436)
         );
  AOI22_X1 U4932 ( .A1(n4755), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4434) );
  AOI22_X1 U4933 ( .A1(n3670), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U4934 ( .A1(n4762), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U4935 ( .A1(n3667), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4431) );
  NAND4_X1 U4936 ( .A1(n4434), .A2(n4433), .A3(n4432), .A4(n4431), .ZN(n4435)
         );
  OR2_X1 U4937 ( .A1(n4436), .A2(n4435), .ZN(n4437) );
  NAND2_X1 U4938 ( .A1(n4468), .A2(n4437), .ZN(n4440) );
  XNOR2_X1 U4939 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4455), .ZN(n6181)
         );
  OAI22_X1 U4940 ( .A1(n4317), .A2(n6181), .B1(n4643), .B2(n6179), .ZN(n4439)
         );
  AOI21_X1 U4941 ( .B1(n4794), .B2(EAX_REG_13__SCAN_IN), .A(n4439), .ZN(n6143)
         );
  INV_X1 U4942 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4443) );
  INV_X1 U4943 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4442) );
  OAI22_X1 U4944 ( .A1(n4751), .A2(n4443), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4442), .ZN(n4444) );
  NAND2_X1 U4945 ( .A1(n4444), .A2(n4317), .ZN(n4458) );
  AOI22_X1 U4946 ( .A1(n4754), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U4947 ( .A1(n3663), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4447) );
  AOI22_X1 U4948 ( .A1(n3661), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4446) );
  AOI22_X1 U4949 ( .A1(n4761), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4445) );
  NAND4_X1 U4950 ( .A1(n4448), .A2(n4447), .A3(n4446), .A4(n4445), .ZN(n4454)
         );
  AOI22_X1 U4951 ( .A1(n4755), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4452) );
  AOI22_X1 U4952 ( .A1(n3671), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4451) );
  AOI22_X1 U4953 ( .A1(n4753), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4450) );
  AOI22_X1 U4954 ( .A1(n3652), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4449) );
  NAND4_X1 U4955 ( .A1(n4452), .A2(n4451), .A3(n4450), .A4(n4449), .ZN(n4453)
         );
  OR2_X1 U4956 ( .A1(n4454), .A2(n4453), .ZN(n4456) );
  XNOR2_X1 U4957 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4459), .ZN(n6204)
         );
  AOI22_X1 U4958 ( .A1(n4468), .A2(n4456), .B1(n4777), .B2(n6204), .ZN(n4457)
         );
  NAND2_X1 U4959 ( .A1(n4458), .A2(n4457), .ZN(n6189) );
  NAND2_X1 U4960 ( .A1(n6186), .A2(n6189), .ZN(n6187) );
  INV_X1 U4961 ( .A(n6187), .ZN(n4477) );
  XOR2_X1 U4962 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4478), .Z(n7146) );
  INV_X1 U4963 ( .A(n7146), .ZN(n4475) );
  AOI22_X1 U4964 ( .A1(n3660), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4463) );
  AOI22_X1 U4965 ( .A1(n4761), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4462) );
  AOI22_X1 U4966 ( .A1(n4754), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4461) );
  AOI22_X1 U4967 ( .A1(n4755), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4460) );
  NAND4_X1 U4968 ( .A1(n4463), .A2(n4462), .A3(n4461), .A4(n4460), .ZN(n4470)
         );
  AOI22_X1 U4969 ( .A1(n3663), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4467) );
  AOI22_X1 U4970 ( .A1(n3671), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4466) );
  AOI22_X1 U4971 ( .A1(n4753), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4465) );
  AOI22_X1 U4972 ( .A1(n3667), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4464) );
  NAND4_X1 U4973 ( .A1(n4467), .A2(n4466), .A3(n4465), .A4(n4464), .ZN(n4469)
         );
  OAI21_X1 U4974 ( .B1(n4470), .B2(n4469), .A(n4468), .ZN(n4473) );
  NAND2_X1 U4975 ( .A1(n4794), .A2(EAX_REG_15__SCAN_IN), .ZN(n4472) );
  NAND2_X1 U4976 ( .A1(n4793), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4471)
         );
  NAND3_X1 U4977 ( .A1(n4473), .A2(n4472), .A3(n4471), .ZN(n4474) );
  AOI21_X1 U4978 ( .B1(n4475), .B2(n4777), .A(n4474), .ZN(n6211) );
  NAND2_X1 U4979 ( .A1(n4477), .A2(n4476), .ZN(n6210) );
  INV_X1 U4980 ( .A(n6210), .ZN(n4494) );
  XNOR2_X1 U4981 ( .A(n4496), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n7160)
         );
  INV_X1 U4982 ( .A(n7160), .ZN(n6563) );
  AOI22_X1 U4983 ( .A1(n3660), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4483) );
  AOI22_X1 U4984 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4761), .B1(n4756), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U4985 ( .A1(n4753), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4481) );
  AOI22_X1 U4986 ( .A1(n4754), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4480) );
  NAND4_X1 U4987 ( .A1(n4483), .A2(n4482), .A3(n4481), .A4(n4480), .ZN(n4489)
         );
  AOI22_X1 U4988 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n3663), .B1(n3664), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4487) );
  AOI22_X1 U4989 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3670), .B1(n3675), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4486) );
  AOI22_X1 U4990 ( .A1(n3666), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4485) );
  AOI22_X1 U4991 ( .A1(n4755), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4484) );
  NAND4_X1 U4992 ( .A1(n4487), .A2(n4486), .A3(n4485), .A4(n4484), .ZN(n4488)
         );
  NOR2_X1 U4993 ( .A1(n4489), .A2(n4488), .ZN(n4491) );
  AOI22_X1 U4994 ( .A1(n4794), .A2(EAX_REG_16__SCAN_IN), .B1(n4793), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4490) );
  OAI21_X1 U4995 ( .B1(n4727), .B2(n4491), .A(n4490), .ZN(n4492) );
  AOI21_X1 U4996 ( .B1(n6563), .B2(n4777), .A(n4492), .ZN(n6470) );
  OR2_X1 U4997 ( .A1(n4497), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4498)
         );
  NAND2_X1 U4998 ( .A1(n4498), .A2(n4529), .ZN(n7173) );
  AOI22_X1 U4999 ( .A1(n3660), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4502) );
  AOI22_X1 U5000 ( .A1(n4754), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5001 ( .A1(n4761), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5002 ( .A1(n4756), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4499) );
  NAND4_X1 U5003 ( .A1(n4502), .A2(n4501), .A3(n4500), .A4(n4499), .ZN(n4508)
         );
  AOI22_X1 U5004 ( .A1(n4755), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3663), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5005 ( .A1(n3670), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4505) );
  AOI22_X1 U5006 ( .A1(n4762), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U5007 ( .A1(n3666), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4503) );
  NAND4_X1 U5008 ( .A1(n4506), .A2(n4505), .A3(n4504), .A4(n4503), .ZN(n4507)
         );
  NOR2_X1 U5009 ( .A1(n4508), .A2(n4507), .ZN(n4511) );
  OAI21_X1 U5010 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n7330), .A(n7295), 
        .ZN(n4510) );
  NAND2_X1 U5011 ( .A1(n4794), .A2(EAX_REG_17__SCAN_IN), .ZN(n4509) );
  OAI211_X1 U5012 ( .C1(n4727), .C2(n4511), .A(n4510), .B(n4509), .ZN(n4512)
         );
  OAI21_X1 U5013 ( .B1(n7173), .B2(n4317), .A(n4512), .ZN(n6462) );
  AOI22_X1 U5014 ( .A1(n4754), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4516) );
  AOI22_X1 U5015 ( .A1(n3911), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5016 ( .A1(n4756), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U5017 ( .A1(n3651), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4513) );
  NAND4_X1 U5018 ( .A1(n4516), .A2(n4515), .A3(n4514), .A4(n4513), .ZN(n4524)
         );
  AOI22_X1 U5019 ( .A1(n4753), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4755), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4522) );
  AOI21_X1 U5020 ( .B1(n4762), .B2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n4777), 
        .ZN(n4518) );
  NAND2_X1 U5021 ( .A1(n3670), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4517)
         );
  AND2_X1 U5022 ( .A1(n4518), .A2(n4517), .ZN(n4521) );
  AOI22_X1 U5023 ( .A1(n3661), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3652), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4520) );
  AOI22_X1 U5024 ( .A1(n3663), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4519) );
  NAND4_X1 U5025 ( .A1(n4522), .A2(n4521), .A3(n4520), .A4(n4519), .ZN(n4523)
         );
  NAND2_X1 U5026 ( .A1(n4727), .A2(n4317), .ZN(n4595) );
  OAI21_X1 U5027 ( .B1(n4524), .B2(n4523), .A(n4595), .ZN(n4527) );
  AOI22_X1 U5028 ( .A1(n4794), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n7295), .ZN(n4526) );
  XNOR2_X1 U5029 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4529), .ZN(n6556)
         );
  AOI21_X1 U5030 ( .B1(n4527), .B2(n4526), .A(n4525), .ZN(n6406) );
  OR2_X1 U5031 ( .A1(n4530), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4531)
         );
  NAND2_X1 U5032 ( .A1(n4531), .A2(n4565), .ZN(n7188) );
  AOI22_X1 U5033 ( .A1(n3658), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5034 ( .A1(n3663), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3671), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4534) );
  AOI22_X1 U5035 ( .A1(n4761), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4533) );
  AOI22_X1 U5036 ( .A1(n4755), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4532) );
  NAND4_X1 U5037 ( .A1(n4535), .A2(n4534), .A3(n4533), .A4(n4532), .ZN(n4541)
         );
  AOI22_X1 U5038 ( .A1(n4754), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5039 ( .A1(n3652), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5040 ( .A1(n4004), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4537) );
  AOI22_X1 U5041 ( .A1(n3651), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4536) );
  NAND4_X1 U5042 ( .A1(n4539), .A2(n4538), .A3(n4537), .A4(n4536), .ZN(n4540)
         );
  NOR2_X1 U5043 ( .A1(n4541), .A2(n4540), .ZN(n4542) );
  NOR2_X1 U5044 ( .A1(n4727), .A2(n4542), .ZN(n4546) );
  INV_X1 U5045 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4544) );
  NAND2_X1 U5046 ( .A1(n7295), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4543)
         );
  OAI211_X1 U5047 ( .C1(n4751), .C2(n4544), .A(n4317), .B(n4543), .ZN(n4545)
         );
  OAI22_X1 U5048 ( .A1(n7188), .A2(n4317), .B1(n4546), .B2(n4545), .ZN(n6870)
         );
  AOI22_X1 U5049 ( .A1(n3652), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4550) );
  AOI22_X1 U5050 ( .A1(n4755), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4549) );
  AOI22_X1 U5051 ( .A1(n4753), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4548) );
  AOI22_X1 U5052 ( .A1(n4754), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4547) );
  NAND4_X1 U5053 ( .A1(n4550), .A2(n4549), .A3(n4548), .A4(n4547), .ZN(n4558)
         );
  NAND2_X1 U5054 ( .A1(n3911), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4552) );
  NAND2_X1 U5055 ( .A1(n3675), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4551)
         );
  AND3_X1 U5056 ( .A1(n4552), .A2(n4551), .A3(n4317), .ZN(n4556) );
  AOI22_X1 U5057 ( .A1(n3660), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4555) );
  AOI22_X1 U5058 ( .A1(n3670), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4554) );
  AOI22_X1 U5059 ( .A1(n3663), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4553) );
  NAND4_X1 U5060 ( .A1(n4556), .A2(n4555), .A3(n4554), .A4(n4553), .ZN(n4557)
         );
  OAI21_X1 U5061 ( .B1(n4558), .B2(n4557), .A(n4595), .ZN(n4560) );
  AOI22_X1 U5062 ( .A1(n4794), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n7295), .ZN(n4559) );
  NAND2_X1 U5063 ( .A1(n4560), .A2(n4559), .ZN(n4562) );
  XNOR2_X1 U5064 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4565), .ZN(n7200)
         );
  NAND2_X1 U5065 ( .A1(n7200), .A2(n4777), .ZN(n4561) );
  NAND2_X1 U5066 ( .A1(n4562), .A2(n4561), .ZN(n6454) );
  INV_X1 U5067 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4564) );
  INV_X1 U5068 ( .A(n4604), .ZN(n4568) );
  OR2_X1 U5069 ( .A1(n4566), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4567)
         );
  NAND2_X1 U5070 ( .A1(n4568), .A2(n4567), .ZN(n7213) );
  AOI22_X1 U5071 ( .A1(n3661), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4572) );
  AOI22_X1 U5072 ( .A1(n3663), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5073 ( .A1(n3652), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5074 ( .A1(n4754), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4569) );
  NAND4_X1 U5075 ( .A1(n4572), .A2(n4571), .A3(n4570), .A4(n4569), .ZN(n4578)
         );
  AOI22_X1 U5076 ( .A1(n4755), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5077 ( .A1(n3670), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4575) );
  AOI22_X1 U5078 ( .A1(n4753), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4574) );
  AOI22_X1 U5079 ( .A1(n4761), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4573) );
  NAND4_X1 U5080 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n4577)
         );
  NOR2_X1 U5081 ( .A1(n4578), .A2(n4577), .ZN(n4582) );
  NAND2_X1 U5082 ( .A1(n7295), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4579)
         );
  NAND2_X1 U5083 ( .A1(n4317), .A2(n4579), .ZN(n4580) );
  AOI21_X1 U5084 ( .B1(n4794), .B2(EAX_REG_21__SCAN_IN), .A(n4580), .ZN(n4581)
         );
  OAI21_X1 U5085 ( .B1(n4727), .B2(n4582), .A(n4581), .ZN(n4583) );
  INV_X1 U5086 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6539) );
  XNOR2_X1 U5087 ( .A(n4604), .B(n6539), .ZN(n6542) );
  NAND2_X1 U5088 ( .A1(n6542), .A2(n4777), .ZN(n4601) );
  AOI22_X1 U5089 ( .A1(n4753), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3671), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U5090 ( .A1(n4756), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5091 ( .A1(n3665), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U5092 ( .A1(n3652), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4585) );
  NAND4_X1 U5093 ( .A1(n4588), .A2(n4587), .A3(n4586), .A4(n4585), .ZN(n4597)
         );
  NAND2_X1 U5094 ( .A1(n3663), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4590) );
  NAND2_X1 U5095 ( .A1(n3658), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4589) );
  AND3_X1 U5096 ( .A1(n4590), .A2(n4589), .A3(n4317), .ZN(n4594) );
  AOI22_X1 U5097 ( .A1(n4755), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4593) );
  AOI22_X1 U5098 ( .A1(n3660), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4592) );
  AOI22_X1 U5099 ( .A1(n4754), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4591) );
  NAND4_X1 U5100 ( .A1(n4594), .A2(n4593), .A3(n4592), .A4(n4591), .ZN(n4596)
         );
  OAI21_X1 U5101 ( .B1(n4597), .B2(n4596), .A(n4595), .ZN(n4599) );
  AOI22_X1 U5102 ( .A1(n4794), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n7295), .ZN(n4598) );
  NAND2_X1 U5103 ( .A1(n4599), .A2(n4598), .ZN(n4600) );
  NAND2_X1 U5104 ( .A1(n4601), .A2(n4600), .ZN(n6392) );
  AND2_X1 U5105 ( .A1(n4605), .A2(n7216), .ZN(n4606) );
  OR2_X1 U5106 ( .A1(n4606), .A2(n4649), .ZN(n7223) );
  AOI22_X1 U5107 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4755), .B1(n4756), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4610) );
  AOI22_X1 U5108 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3663), .B1(n3664), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4609) );
  AOI22_X1 U5109 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3670), .B1(n3653), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4608) );
  AOI22_X1 U5110 ( .A1(n4761), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4607) );
  NAND4_X1 U5111 ( .A1(n4610), .A2(n4609), .A3(n4608), .A4(n4607), .ZN(n4616)
         );
  AOI22_X1 U5112 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4753), .B1(n3652), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4614) );
  AOI22_X1 U5113 ( .A1(n3660), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4613) );
  AOI22_X1 U5114 ( .A1(n3658), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4612) );
  AOI22_X1 U5115 ( .A1(n4754), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4611) );
  NAND4_X1 U5116 ( .A1(n4614), .A2(n4613), .A3(n4612), .A4(n4611), .ZN(n4615)
         );
  OR2_X1 U5117 ( .A1(n4616), .A2(n4615), .ZN(n4628) );
  AOI22_X1 U5118 ( .A1(n4755), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4620) );
  AOI22_X1 U5119 ( .A1(n3663), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4619) );
  AOI22_X1 U5120 ( .A1(n3670), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4618) );
  AOI22_X1 U5121 ( .A1(n4761), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4617) );
  NAND4_X1 U5122 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n4626)
         );
  AOI22_X1 U5123 ( .A1(n4753), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3652), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4624) );
  AOI22_X1 U5124 ( .A1(n3660), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5125 ( .A1(n3658), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4622) );
  AOI22_X1 U5126 ( .A1(n4754), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4621) );
  NAND4_X1 U5127 ( .A1(n4624), .A2(n4623), .A3(n4622), .A4(n4621), .ZN(n4625)
         );
  OR2_X1 U5128 ( .A1(n4626), .A2(n4625), .ZN(n4627) );
  NAND2_X1 U5129 ( .A1(n4627), .A2(n4628), .ZN(n4663) );
  OAI21_X1 U5130 ( .B1(n4628), .B2(n4627), .A(n4663), .ZN(n4631) );
  OAI21_X1 U5131 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7216), .A(n4317), .ZN(
        n4629) );
  AOI21_X1 U5132 ( .B1(n4794), .B2(EAX_REG_23__SCAN_IN), .A(n4629), .ZN(n4630)
         );
  OAI21_X1 U5133 ( .B1(n4727), .B2(n4631), .A(n4630), .ZN(n4632) );
  OAI21_X1 U5134 ( .B1(n7223), .B2(n4317), .A(n4632), .ZN(n6439) );
  XNOR2_X1 U5135 ( .A(n4649), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6523)
         );
  NAND2_X1 U5136 ( .A1(n6523), .A2(n4777), .ZN(n4648) );
  INV_X1 U5137 ( .A(n4727), .ZN(n4774) );
  AOI22_X1 U5138 ( .A1(n4754), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4755), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5139 ( .A1(n4756), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U5140 ( .A1(n3665), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4634) );
  AOI22_X1 U5141 ( .A1(n3666), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4633) );
  NAND4_X1 U5142 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), .ZN(n4642)
         );
  AOI22_X1 U5143 ( .A1(n3661), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5144 ( .A1(n3663), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3670), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5145 ( .A1(n4753), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4638) );
  AOI22_X1 U5146 ( .A1(n3909), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4637) );
  NAND4_X1 U5147 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4641)
         );
  OR2_X1 U5148 ( .A1(n4642), .A2(n4641), .ZN(n4662) );
  XNOR2_X1 U5149 ( .A(n4663), .B(n4662), .ZN(n4646) );
  INV_X1 U5150 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4644) );
  INV_X1 U5151 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6383) );
  OAI22_X1 U5152 ( .A1(n4751), .A2(n4644), .B1(n4643), .B2(n6383), .ZN(n4645)
         );
  AOI21_X1 U5153 ( .B1(n4774), .B2(n4646), .A(n4645), .ZN(n4647) );
  NAND2_X1 U5154 ( .A1(n4648), .A2(n4647), .ZN(n6381) );
  OR2_X1 U5155 ( .A1(n4650), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4651)
         );
  NAND2_X1 U5156 ( .A1(n4651), .A2(n4691), .ZN(n7240) );
  AOI22_X1 U5157 ( .A1(n4755), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4756), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5158 ( .A1(n3663), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5159 ( .A1(n3671), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4653) );
  AOI22_X1 U5160 ( .A1(n4761), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4652) );
  NAND4_X1 U5161 ( .A1(n4655), .A2(n4654), .A3(n4653), .A4(n4652), .ZN(n4661)
         );
  AOI22_X1 U5162 ( .A1(n4753), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3652), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5163 ( .A1(n3661), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5164 ( .A1(n3911), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5165 ( .A1(n4754), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4656) );
  NAND4_X1 U5166 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4660)
         );
  OR2_X1 U5167 ( .A1(n4661), .A2(n4660), .ZN(n4681) );
  INV_X1 U5168 ( .A(n4662), .ZN(n4664) );
  NOR2_X1 U5169 ( .A1(n4664), .A2(n4663), .ZN(n4682) );
  XNOR2_X1 U5170 ( .A(n4681), .B(n4682), .ZN(n4668) );
  NAND2_X1 U5171 ( .A1(n7295), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4665)
         );
  NAND2_X1 U5172 ( .A1(n4317), .A2(n4665), .ZN(n4666) );
  AOI21_X1 U5173 ( .B1(n4794), .B2(EAX_REG_25__SCAN_IN), .A(n4666), .ZN(n4667)
         );
  OAI21_X1 U5174 ( .B1(n4727), .B2(n4668), .A(n4667), .ZN(n4669) );
  AOI22_X1 U5175 ( .A1(n4756), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5176 ( .A1(n3663), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4673) );
  AOI22_X1 U5177 ( .A1(n3911), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U5178 ( .A1(n4754), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4671) );
  NAND4_X1 U5179 ( .A1(n4674), .A2(n4673), .A3(n4672), .A4(n4671), .ZN(n4680)
         );
  AOI22_X1 U5180 ( .A1(n4753), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4678) );
  AOI22_X1 U5181 ( .A1(n3670), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4677) );
  AOI22_X1 U5182 ( .A1(n3660), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5183 ( .A1(n4755), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4675) );
  NAND4_X1 U5184 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4679)
         );
  NOR2_X1 U5185 ( .A1(n4680), .A2(n4679), .ZN(n4697) );
  NAND2_X1 U5186 ( .A1(n4682), .A2(n4681), .ZN(n4696) );
  XOR2_X1 U5187 ( .A(n4697), .B(n4696), .Z(n4683) );
  NAND2_X1 U5188 ( .A1(n4683), .A2(n4774), .ZN(n4686) );
  INV_X1 U5189 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6517) );
  OAI21_X1 U5190 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6517), .A(n4317), .ZN(
        n4684) );
  AOI21_X1 U5191 ( .B1(n4794), .B2(EAX_REG_26__SCAN_IN), .A(n4684), .ZN(n4685)
         );
  NAND2_X1 U5192 ( .A1(n4686), .A2(n4685), .ZN(n4688) );
  XNOR2_X1 U5193 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4691), .ZN(n6515)
         );
  NAND2_X1 U5194 ( .A1(n4777), .A2(n6515), .ZN(n4687) );
  NAND2_X1 U5195 ( .A1(n4688), .A2(n4687), .ZN(n6366) );
  NAND2_X2 U5196 ( .A1(n4690), .A2(n4689), .ZN(n6351) );
  INV_X1 U5197 ( .A(n4691), .ZN(n4692) );
  INV_X1 U5198 ( .A(n4693), .ZN(n4694) );
  INV_X1 U5199 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U5200 ( .A1(n4694), .A2(n6357), .ZN(n4695) );
  NAND2_X1 U5201 ( .A1(n4713), .A2(n4695), .ZN(n6510) );
  NOR2_X1 U5202 ( .A1(n4697), .A2(n4696), .ZN(n4715) );
  AOI22_X1 U5203 ( .A1(n3660), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5204 ( .A1(n4754), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4700) );
  AOI22_X1 U5205 ( .A1(n4756), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4699) );
  AOI22_X1 U5206 ( .A1(n3663), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4698) );
  NAND4_X1 U5207 ( .A1(n4701), .A2(n4700), .A3(n4699), .A4(n4698), .ZN(n4707)
         );
  AOI22_X1 U5208 ( .A1(n3671), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4705) );
  AOI22_X1 U5209 ( .A1(n4762), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5210 ( .A1(n4753), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4703) );
  AOI22_X1 U5211 ( .A1(n4755), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4702) );
  NAND4_X1 U5212 ( .A1(n4705), .A2(n4704), .A3(n4703), .A4(n4702), .ZN(n4706)
         );
  OR2_X1 U5213 ( .A1(n4707), .A2(n4706), .ZN(n4716) );
  XNOR2_X1 U5214 ( .A(n4715), .B(n4716), .ZN(n4710) );
  AOI21_X1 U5215 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n7295), .A(n4777), 
        .ZN(n4709) );
  NAND2_X1 U5216 ( .A1(n4794), .A2(EAX_REG_27__SCAN_IN), .ZN(n4708) );
  OAI211_X1 U5217 ( .C1(n4710), .C2(n4727), .A(n4709), .B(n4708), .ZN(n4711)
         );
  OAI21_X1 U5218 ( .B1(n4317), .B2(n6510), .A(n4711), .ZN(n6353) );
  INV_X1 U5219 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U5220 ( .A1(n4713), .A2(n6225), .ZN(n4714) );
  OAI21_X1 U5221 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6225), .A(n4317), .ZN(
        n4730) );
  NAND2_X1 U5222 ( .A1(n4716), .A2(n4715), .ZN(n4770) );
  AOI22_X1 U5223 ( .A1(n3671), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4720) );
  AOI22_X1 U5224 ( .A1(n4754), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4719) );
  AOI22_X1 U5225 ( .A1(n4004), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4718) );
  AOI22_X1 U5226 ( .A1(n4756), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4717) );
  NAND4_X1 U5227 ( .A1(n4720), .A2(n4719), .A3(n4718), .A4(n4717), .ZN(n4726)
         );
  AOI22_X1 U5228 ( .A1(n3658), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4724) );
  AOI22_X1 U5229 ( .A1(n4755), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3961), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4723) );
  AOI22_X1 U5230 ( .A1(n3663), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U5231 ( .A1(n3652), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4721) );
  NAND4_X1 U5232 ( .A1(n4724), .A2(n4723), .A3(n4722), .A4(n4721), .ZN(n4725)
         );
  NOR2_X1 U5233 ( .A1(n4726), .A2(n4725), .ZN(n4769) );
  XNOR2_X1 U5234 ( .A(n4770), .B(n4769), .ZN(n4728) );
  NOR2_X1 U5235 ( .A1(n4728), .A2(n4727), .ZN(n4729) );
  AOI211_X1 U5236 ( .C1(n4794), .C2(EAX_REG_28__SCAN_IN), .A(n4730), .B(n4729), 
        .ZN(n4731) );
  INV_X1 U5237 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4733) );
  NAND2_X1 U5238 ( .A1(n4734), .A2(n4733), .ZN(n4735) );
  NAND2_X1 U5239 ( .A1(n4811), .A2(n4735), .ZN(n6502) );
  INV_X1 U5240 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4750) );
  NOR2_X1 U5241 ( .A1(n4770), .A2(n4769), .ZN(n4746) );
  AOI22_X1 U5242 ( .A1(n4004), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4739) );
  AOI22_X1 U5243 ( .A1(n3671), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3651), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4738) );
  AOI22_X1 U5244 ( .A1(n3666), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4737) );
  AOI22_X1 U5245 ( .A1(n4755), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4065), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4736) );
  NAND4_X1 U5246 ( .A1(n4739), .A2(n4738), .A3(n4737), .A4(n4736), .ZN(n4745)
         );
  AOI22_X1 U5247 ( .A1(n4756), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4743) );
  AOI22_X1 U5248 ( .A1(n3663), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3665), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4742) );
  AOI22_X1 U5249 ( .A1(n4753), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4741) );
  AOI22_X1 U5250 ( .A1(n4754), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4740) );
  NAND4_X1 U5251 ( .A1(n4743), .A2(n4742), .A3(n4741), .A4(n4740), .ZN(n4744)
         );
  NOR2_X1 U5252 ( .A1(n4745), .A2(n4744), .ZN(n4771) );
  XNOR2_X1 U5253 ( .A(n4746), .B(n4771), .ZN(n4747) );
  NAND2_X1 U5254 ( .A1(n4747), .A2(n4774), .ZN(n4749) );
  AOI21_X1 U5255 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n7295), .A(n4777), 
        .ZN(n4748) );
  OAI211_X1 U5256 ( .C1(n4751), .C2(n4750), .A(n4749), .B(n4748), .ZN(n4752)
         );
  OAI21_X1 U5257 ( .B1(n4317), .B2(n6502), .A(n4752), .ZN(n6340) );
  AOI22_X1 U5258 ( .A1(n4754), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4753), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4760) );
  AOI22_X1 U5259 ( .A1(n3670), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3653), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4759) );
  AOI22_X1 U5260 ( .A1(n4755), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4758) );
  AOI22_X1 U5261 ( .A1(n4756), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4757) );
  NAND4_X1 U5262 ( .A1(n4760), .A2(n4759), .A3(n4758), .A4(n4757), .ZN(n4768)
         );
  AOI22_X1 U5263 ( .A1(n3667), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4761), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4766) );
  AOI22_X1 U5264 ( .A1(n3663), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3664), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5265 ( .A1(n3658), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4762), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5266 ( .A1(n3660), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4763) );
  NAND4_X1 U5267 ( .A1(n4766), .A2(n4765), .A3(n4764), .A4(n4763), .ZN(n4767)
         );
  NOR2_X1 U5268 ( .A1(n4768), .A2(n4767), .ZN(n4773) );
  NOR3_X1 U5269 ( .A1(n4771), .A2(n4770), .A3(n4769), .ZN(n4772) );
  XNOR2_X1 U5270 ( .A(n4773), .B(n4772), .ZN(n4775) );
  NAND2_X1 U5271 ( .A1(n4775), .A2(n4774), .ZN(n4780) );
  INV_X1 U5272 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4810) );
  AOI21_X1 U5273 ( .B1(n4810), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4776) );
  AOI21_X1 U5274 ( .B1(n4794), .B2(EAX_REG_30__SCAN_IN), .A(n4776), .ZN(n4779)
         );
  XNOR2_X1 U5275 ( .A(n4811), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6331)
         );
  AND2_X1 U5276 ( .A1(n6331), .A2(n4777), .ZN(n4778) );
  NAND2_X1 U5277 ( .A1(n7313), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5370) );
  INV_X1 U5278 ( .A(n5370), .ZN(n4782) );
  NAND2_X1 U5279 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4782), .ZN(n6952) );
  INV_X1 U5280 ( .A(n6952), .ZN(n4783) );
  NAND2_X1 U5281 ( .A1(n7457), .A2(n4783), .ZN(n6914) );
  INV_X2 U5282 ( .A(n6914), .ZN(n6937) );
  AND2_X1 U5283 ( .A1(n7445), .A2(n4784), .ZN(n6954) );
  OR2_X1 U5284 ( .A1(n6954), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4785) );
  NAND2_X1 U5285 ( .A1(n7313), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4787) );
  NAND2_X1 U5286 ( .A1(n7330), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4786) );
  NAND2_X1 U5287 ( .A1(n4787), .A2(n4786), .ZN(n6884) );
  NAND2_X1 U5288 ( .A1(n6901), .A2(n6331), .ZN(n4788) );
  AND2_X1 U5289 ( .A1(n7457), .A2(n7296), .ZN(n5049) );
  NAND2_X1 U5290 ( .A1(n7059), .A2(REIP_REG_30__SCAN_IN), .ZN(n6577) );
  OAI211_X1 U5291 ( .C1(n4810), .C2(n6906), .A(n4788), .B(n6577), .ZN(n4789)
         );
  AOI21_X1 U5292 ( .B1(n6479), .B2(n6937), .A(n4789), .ZN(n4790) );
  OAI21_X1 U5293 ( .B1(n6582), .B2(n7241), .A(n4790), .ZN(U2956) );
  AOI22_X1 U5294 ( .A1(n4794), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4793), .ZN(n4795) );
  INV_X1 U5295 ( .A(n4795), .ZN(n4796) );
  INV_X1 U5296 ( .A(n4799), .ZN(n4967) );
  NOR3_X1 U5297 ( .A1(n4803), .A2(n4802), .A3(n4801), .ZN(n4804) );
  OR2_X1 U5298 ( .A1(n4805), .A2(n4804), .ZN(n4807) );
  NOR2_X1 U5299 ( .A1(n6323), .A2(n6317), .ZN(n6326) );
  NAND2_X1 U5300 ( .A1(n6326), .A2(n7292), .ZN(n5048) );
  NAND2_X1 U5301 ( .A1(n7295), .A2(n7296), .ZN(n7314) );
  NOR3_X1 U5302 ( .A1(n7313), .A2(n7305), .A3(n7314), .ZN(n7310) );
  NOR2_X1 U5303 ( .A1(n4317), .A2(n5370), .ZN(n7301) );
  OR2_X1 U5304 ( .A1(n7059), .A2(n7301), .ZN(n4808) );
  NOR2_X1 U5305 ( .A1(n7310), .A2(n4808), .ZN(n4809) );
  INV_X1 U5306 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U5307 ( .A1(n6313), .A2(n7236), .ZN(n4925) );
  NAND2_X1 U5308 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .ZN(
        n4826) );
  INV_X1 U5309 ( .A(n4826), .ZN(n4822) );
  NAND2_X1 U5310 ( .A1(n4813), .A2(n7345), .ZN(n6950) );
  NOR2_X1 U5311 ( .A1(n5226), .A2(n5364), .ZN(n4931) );
  NOR2_X1 U5312 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n5573) );
  NAND2_X1 U5313 ( .A1(n3983), .A2(n5573), .ZN(n4814) );
  NAND2_X1 U5314 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4821) );
  INV_X1 U5315 ( .A(n6421), .ZN(n7114) );
  AND2_X1 U5316 ( .A1(n7192), .A2(n7114), .ZN(n6407) );
  INV_X1 U5317 ( .A(n6407), .ZN(n5586) );
  NAND3_X1 U5318 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        REIP_REG_22__SCAN_IN), .ZN(n4815) );
  NAND2_X1 U5319 ( .A1(n5586), .A2(n4815), .ZN(n4817) );
  INV_X1 U5320 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7190) );
  INV_X1 U5321 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6812) );
  NAND3_X1 U5322 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_14__SCAN_IN), .ZN(n6195) );
  NAND3_X1 U5323 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6014) );
  INV_X1 U5324 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7086) );
  INV_X1 U5325 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6791) );
  NOR3_X1 U5326 ( .A1(n6014), .A2(n7086), .A3(n6791), .ZN(n7115) );
  NAND4_X1 U5327 ( .A1(n7115), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .A4(REIP_REG_8__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U5328 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n6032) );
  NOR2_X1 U5329 ( .A1(n6030), .A2(n6032), .ZN(n6049) );
  NAND2_X1 U5330 ( .A1(n6049), .A2(REIP_REG_11__SCAN_IN), .ZN(n6194) );
  NOR2_X1 U5331 ( .A1(n6195), .A2(n6194), .ZN(n7142) );
  NAND4_X1 U5332 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n7142), .ZN(n6413) );
  NOR2_X1 U5333 ( .A1(n6812), .A2(n6413), .ZN(n7177) );
  NAND2_X1 U5334 ( .A1(REIP_REG_19__SCAN_IN), .A2(n7177), .ZN(n7191) );
  NOR2_X1 U5335 ( .A1(n7190), .A2(n7191), .ZN(n4825) );
  INV_X1 U5336 ( .A(n4825), .ZN(n7208) );
  NAND2_X1 U5337 ( .A1(n7178), .A2(n7208), .ZN(n4816) );
  AND2_X1 U5338 ( .A1(n4816), .A2(n7114), .ZN(n7189) );
  INV_X1 U5339 ( .A(REIP_REG_24__SCAN_IN), .ZN(n7224) );
  INV_X1 U5340 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7232) );
  NOR2_X1 U5341 ( .A1(n7224), .A2(n7232), .ZN(n4818) );
  NAND2_X1 U5342 ( .A1(n4818), .A2(REIP_REG_26__SCAN_IN), .ZN(n4819) );
  NAND2_X1 U5343 ( .A1(n7178), .A2(n4819), .ZN(n4820) );
  NAND2_X1 U5344 ( .A1(n7225), .A2(n4820), .ZN(n6373) );
  AOI21_X1 U5345 ( .B1(n7178), .B2(n4821), .A(n6373), .ZN(n6342) );
  OAI21_X1 U5346 ( .B1(n4822), .B2(n7192), .A(n6342), .ZN(n6336) );
  INV_X1 U5347 ( .A(n5573), .ZN(n4921) );
  OR2_X1 U5348 ( .A1(n6950), .A2(n4921), .ZN(n7288) );
  AND2_X1 U5349 ( .A1(n4017), .A2(n7288), .ZN(n5576) );
  NAND2_X1 U5350 ( .A1(n5576), .A2(EBX_REG_31__SCAN_IN), .ZN(n4823) );
  OAI22_X1 U5351 ( .A1(n4824), .A2(n7215), .B1(n6953), .B2(n4823), .ZN(n4828)
         );
  INV_X1 U5352 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6819) );
  NAND3_X1 U5353 ( .A1(n7178), .A2(n4825), .A3(REIP_REG_21__SCAN_IN), .ZN(
        n6396) );
  NOR2_X1 U5354 ( .A1(n6819), .A2(n6396), .ZN(n7214) );
  NAND2_X1 U5355 ( .A1(REIP_REG_23__SCAN_IN), .A2(n7214), .ZN(n7226) );
  NOR3_X1 U5356 ( .A1(n7224), .A2(n7232), .A3(n7226), .ZN(n6372) );
  AND3_X1 U5357 ( .A1(n6372), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U5358 ( .A1(n6242), .A2(REIP_REG_28__SCAN_IN), .ZN(n6350) );
  NOR3_X1 U5359 ( .A1(n6350), .A2(REIP_REG_31__SCAN_IN), .A3(n4826), .ZN(n4827) );
  AOI211_X1 U5360 ( .C1(REIP_REG_31__SCAN_IN), .C2(n6336), .A(n4828), .B(n4827), .ZN(n4924) );
  INV_X1 U5361 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4831) );
  NAND2_X1 U5362 ( .A1(n5099), .A2(n4831), .ZN(n4830) );
  INV_X1 U5363 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U5364 ( .A1(n4909), .A2(n5268), .ZN(n4829) );
  NAND3_X1 U5365 ( .A1(n4830), .A2(n4916), .A3(n4829), .ZN(n4833) );
  NAND2_X1 U5366 ( .A1(n3659), .A2(n4831), .ZN(n4832) );
  NAND2_X1 U5367 ( .A1(n4833), .A2(n4832), .ZN(n4835) );
  NAND2_X1 U5368 ( .A1(n4909), .A2(EBX_REG_0__SCAN_IN), .ZN(n4834) );
  OAI21_X1 U5369 ( .B1(n3659), .B2(EBX_REG_0__SCAN_IN), .A(n4834), .ZN(n5122)
         );
  XNOR2_X1 U5370 ( .A(n4835), .B(n5122), .ZN(n5100) );
  NAND2_X1 U5371 ( .A1(n5102), .A2(n4835), .ZN(n5093) );
  INV_X1 U5372 ( .A(n4909), .ZN(n4893) );
  MUX2_X1 U5373 ( .A(n3659), .B(n4893), .S(EBX_REG_2__SCAN_IN), .Z(n4837) );
  AND2_X1 U5374 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4836)
         );
  NOR2_X1 U5375 ( .A1(n4837), .A2(n4836), .ZN(n5092) );
  MUX2_X1 U5376 ( .A(n4906), .B(n4916), .S(EBX_REG_3__SCAN_IN), .Z(n4839) );
  NAND2_X1 U5377 ( .A1(n5121), .A2(n4111), .ZN(n4838) );
  NAND2_X1 U5378 ( .A1(n4839), .A2(n4838), .ZN(n5134) );
  MUX2_X1 U5379 ( .A(n4916), .B(n4909), .S(EBX_REG_4__SCAN_IN), .Z(n4841) );
  NAND2_X1 U5380 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4840)
         );
  NAND2_X1 U5381 ( .A1(n4841), .A2(n4840), .ZN(n5153) );
  MUX2_X1 U5382 ( .A(n4906), .B(n4916), .S(EBX_REG_5__SCAN_IN), .Z(n4843) );
  NAND2_X1 U5383 ( .A1(n5121), .A2(n5320), .ZN(n4842) );
  NAND2_X1 U5384 ( .A1(n4843), .A2(n4842), .ZN(n5259) );
  INV_X1 U5385 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U5386 ( .A1(n4909), .A2(n5442), .ZN(n4845) );
  INV_X1 U5387 ( .A(EBX_REG_6__SCAN_IN), .ZN(n7121) );
  NAND2_X1 U5388 ( .A1(n5099), .A2(n7121), .ZN(n4844) );
  NAND3_X1 U5389 ( .A1(n4845), .A2(n4916), .A3(n4844), .ZN(n4847) );
  NAND2_X1 U5390 ( .A1(n3659), .A2(n7121), .ZN(n4846) );
  AND2_X1 U5391 ( .A1(n4847), .A2(n4846), .ZN(n5328) );
  INV_X1 U5392 ( .A(EBX_REG_7__SCAN_IN), .ZN(n7132) );
  NAND2_X1 U5393 ( .A1(n4881), .A2(n7132), .ZN(n4850) );
  NAND2_X1 U5394 ( .A1(n5099), .A2(n7132), .ZN(n4848) );
  OAI211_X1 U5395 ( .C1(n3659), .C2(n4199), .A(n4848), .B(n4909), .ZN(n4849)
         );
  NAND2_X1 U5396 ( .A1(n4850), .A2(n4849), .ZN(n6864) );
  MUX2_X1 U5397 ( .A(n4916), .B(n4909), .S(EBX_REG_8__SCAN_IN), .Z(n4852) );
  NAND2_X1 U5398 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4851)
         );
  NAND2_X1 U5399 ( .A1(n4852), .A2(n4851), .ZN(n5531) );
  INV_X1 U5400 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U5401 ( .A1(n4881), .A2(n4853), .ZN(n4856) );
  NAND2_X1 U5402 ( .A1(n5099), .A2(n4853), .ZN(n4854) );
  OAI211_X1 U5403 ( .C1(n3659), .C2(n7040), .A(n4854), .B(n4909), .ZN(n4855)
         );
  NAND2_X1 U5404 ( .A1(n4856), .A2(n4855), .ZN(n5541) );
  MUX2_X1 U5405 ( .A(n3659), .B(n4893), .S(EBX_REG_10__SCAN_IN), .Z(n4859) );
  AND2_X1 U5406 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4858)
         );
  NOR2_X1 U5407 ( .A1(n4859), .A2(n4858), .ZN(n6022) );
  MUX2_X1 U5408 ( .A(n4881), .B(n3659), .S(EBX_REG_11__SCAN_IN), .Z(n4861) );
  INV_X1 U5409 ( .A(n5121), .ZN(n4918) );
  NOR2_X1 U5410 ( .A1(n4918), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4860)
         );
  NOR2_X1 U5411 ( .A1(n4861), .A2(n4860), .ZN(n6039) );
  MUX2_X1 U5412 ( .A(n4916), .B(n4909), .S(EBX_REG_12__SCAN_IN), .Z(n4863) );
  NAND2_X1 U5413 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U5414 ( .A1(n4863), .A2(n4862), .ZN(n6074) );
  MUX2_X1 U5415 ( .A(n4906), .B(n4916), .S(EBX_REG_13__SCAN_IN), .Z(n4866) );
  INV_X1 U5416 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4864) );
  NAND2_X1 U5417 ( .A1(n5121), .A2(n4864), .ZN(n4865) );
  NAND2_X1 U5418 ( .A1(n4866), .A2(n4865), .ZN(n6145) );
  MUX2_X1 U5419 ( .A(n4906), .B(n4916), .S(EBX_REG_15__SCAN_IN), .Z(n4868) );
  NAND2_X1 U5420 ( .A1(n5121), .A2(n6662), .ZN(n4867) );
  AND2_X1 U5421 ( .A1(n4868), .A2(n4867), .ZN(n6213) );
  MUX2_X1 U5422 ( .A(n4916), .B(n4909), .S(EBX_REG_14__SCAN_IN), .Z(n4870) );
  NAND2_X1 U5423 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U5424 ( .A1(n4870), .A2(n4869), .ZN(n6214) );
  NAND2_X1 U5425 ( .A1(n6213), .A2(n6214), .ZN(n4871) );
  NAND2_X1 U5426 ( .A1(n4909), .A2(n4872), .ZN(n4874) );
  INV_X1 U5427 ( .A(EBX_REG_16__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U5428 ( .A1(n5099), .A2(n7163), .ZN(n4873) );
  NAND3_X1 U5429 ( .A1(n4874), .A2(n4916), .A3(n4873), .ZN(n4876) );
  NAND2_X1 U5430 ( .A1(n3659), .A2(n7163), .ZN(n4875) );
  NAND2_X1 U5431 ( .A1(n4876), .A2(n4875), .ZN(n6471) );
  MUX2_X1 U5432 ( .A(n4906), .B(n4916), .S(EBX_REG_17__SCAN_IN), .Z(n4878) );
  INV_X1 U5433 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U5434 ( .A1(n5121), .A2(n7055), .ZN(n4877) );
  MUX2_X1 U5435 ( .A(n3659), .B(n4893), .S(EBX_REG_18__SCAN_IN), .Z(n4880) );
  AND2_X1 U5436 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4879)
         );
  NOR2_X1 U5437 ( .A1(n4880), .A2(n4879), .ZN(n5034) );
  INV_X1 U5438 ( .A(EBX_REG_19__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U5439 ( .A1(n4881), .A2(n7181), .ZN(n4885) );
  NAND2_X1 U5440 ( .A1(n5099), .A2(n7181), .ZN(n4882) );
  OAI211_X1 U5441 ( .C1(n3659), .C2(n4883), .A(n4882), .B(n4909), .ZN(n4884)
         );
  NAND2_X1 U5442 ( .A1(n4885), .A2(n4884), .ZN(n6872) );
  NAND2_X1 U5443 ( .A1(n4909), .A2(n6545), .ZN(n4887) );
  INV_X1 U5444 ( .A(EBX_REG_20__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U5445 ( .A1(n5099), .A2(n7204), .ZN(n4886) );
  NAND3_X1 U5446 ( .A1(n4887), .A2(n4916), .A3(n4886), .ZN(n4889) );
  NAND2_X1 U5447 ( .A1(n3659), .A2(n7204), .ZN(n4888) );
  NAND2_X1 U5448 ( .A1(n4889), .A2(n4888), .ZN(n6455) );
  MUX2_X1 U5449 ( .A(n4906), .B(n4916), .S(EBX_REG_21__SCAN_IN), .Z(n4891) );
  NAND2_X1 U5450 ( .A1(n5121), .A2(n6629), .ZN(n4890) );
  NAND2_X1 U5451 ( .A1(n4891), .A2(n4890), .ZN(n6450) );
  MUX2_X1 U5452 ( .A(n3659), .B(n4893), .S(EBX_REG_22__SCAN_IN), .Z(n4895) );
  AND2_X1 U5453 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4894)
         );
  NOR2_X1 U5454 ( .A1(n4895), .A2(n4894), .ZN(n6394) );
  MUX2_X1 U5455 ( .A(n4906), .B(n4916), .S(EBX_REG_23__SCAN_IN), .Z(n4897) );
  NAND2_X1 U5456 ( .A1(n5121), .A2(n6627), .ZN(n4896) );
  NAND2_X1 U5457 ( .A1(n4897), .A2(n4896), .ZN(n6443) );
  MUX2_X1 U5458 ( .A(n4916), .B(n4909), .S(EBX_REG_24__SCAN_IN), .Z(n4899) );
  NAND2_X1 U5459 ( .A1(n3989), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U5460 ( .A1(n4899), .A2(n4898), .ZN(n4955) );
  MUX2_X1 U5461 ( .A(n4906), .B(n4916), .S(EBX_REG_25__SCAN_IN), .Z(n4901) );
  NAND2_X1 U5462 ( .A1(n5121), .A2(n6934), .ZN(n4900) );
  AND2_X1 U5463 ( .A1(n4901), .A2(n4900), .ZN(n6434) );
  NAND2_X1 U5464 ( .A1(n4909), .A2(n6612), .ZN(n4903) );
  INV_X1 U5465 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U5466 ( .A1(n5099), .A2(n6370), .ZN(n4902) );
  NAND3_X1 U5467 ( .A1(n4903), .A2(n4916), .A3(n4902), .ZN(n4905) );
  NAND2_X1 U5468 ( .A1(n3659), .A2(n6370), .ZN(n4904) );
  AND2_X1 U5469 ( .A1(n4905), .A2(n4904), .ZN(n6368) );
  MUX2_X1 U5470 ( .A(n4906), .B(n4916), .S(EBX_REG_27__SCAN_IN), .Z(n4908) );
  NAND2_X1 U5471 ( .A1(n5121), .A2(n6507), .ZN(n4907) );
  NAND2_X1 U5472 ( .A1(n4908), .A2(n4907), .ZN(n6354) );
  INV_X1 U5473 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U5474 ( .A1(n4909), .A2(n6593), .ZN(n4910) );
  OAI211_X1 U5475 ( .C1(EBX_REG_28__SCAN_IN), .C2(n3989), .A(n4910), .B(n4916), 
        .ZN(n4912) );
  INV_X1 U5476 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U5477 ( .A1(n3659), .A2(n6232), .ZN(n4911) );
  NAND2_X1 U5478 ( .A1(n4912), .A2(n4911), .ZN(n6230) );
  NOR2_X1 U5479 ( .A1(n3989), .A2(EBX_REG_29__SCAN_IN), .ZN(n4913) );
  AOI21_X1 U5480 ( .B1(n5121), .B2(n6586), .A(n4913), .ZN(n5024) );
  INV_X1 U5481 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6428) );
  AND2_X1 U5482 ( .A1(n3659), .A2(n6428), .ZN(n4915) );
  AOI21_X1 U5483 ( .B1(n5024), .B2(n4916), .A(n4915), .ZN(n6346) );
  OAI22_X1 U5484 ( .A1(n4918), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n3989), .ZN(n5025) );
  NOR2_X1 U5485 ( .A1(n6346), .A2(n5025), .ZN(n4917) );
  AOI21_X1 U5486 ( .B1(n6345), .B2(n6428), .A(n4916), .ZN(n5023) );
  OAI22_X1 U5487 ( .A1(n4918), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3989), .ZN(n4919) );
  XNOR2_X1 U5488 ( .A(n4920), .B(n4919), .ZN(n6427) );
  NAND2_X1 U5489 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4921), .ZN(n4922) );
  NAND3_X1 U5490 ( .A1(n4925), .A2(n4924), .A3(n4923), .ZN(U2796) );
  XNOR2_X1 U5491 ( .A(n3650), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6923)
         );
  NOR2_X1 U5492 ( .A1(n3650), .A2(n6545), .ZN(n4926) );
  XNOR2_X1 U5493 ( .A(n3650), .B(n6629), .ZN(n6929) );
  NOR2_X1 U5494 ( .A1(n6928), .A2(n6929), .ZN(n6927) );
  NAND3_X1 U5495 ( .A1(n3650), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4928) );
  NAND3_X1 U5496 ( .A1(n6629), .A2(n6545), .A3(n6536), .ZN(n4927) );
  OR3_X1 U5497 ( .A1(n6922), .A2(n3650), .A3(n4927), .ZN(n6532) );
  OAI22_X1 U5498 ( .A1(n6538), .A2(n4928), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6532), .ZN(n4929) );
  XNOR2_X1 U5499 ( .A(n4929), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6526)
         );
  NOR2_X1 U5500 ( .A1(READY_N), .A2(n6317), .ZN(n5058) );
  INV_X1 U5501 ( .A(n5058), .ZN(n4930) );
  AOI21_X1 U5502 ( .B1(n5226), .B2(n6950), .A(n4930), .ZN(n4935) );
  OR2_X1 U5503 ( .A1(n4931), .A2(READY_N), .ZN(n4932) );
  OR2_X1 U5504 ( .A1(n6325), .A2(n4932), .ZN(n5061) );
  NOR2_X1 U5505 ( .A1(n5061), .A2(n4933), .ZN(n4934) );
  MUX2_X1 U5506 ( .A(n4935), .B(n4934), .S(n3980), .Z(n4942) );
  NOR2_X1 U5507 ( .A1(n5079), .A2(n3942), .ZN(n4972) );
  NAND2_X1 U5508 ( .A1(n6325), .A2(n4972), .ZN(n4940) );
  NAND2_X1 U5509 ( .A1(n5146), .A2(n3983), .ZN(n4936) );
  NAND2_X1 U5510 ( .A1(n4957), .A2(n4936), .ZN(n4937) );
  NAND2_X1 U5511 ( .A1(n4938), .A2(n4937), .ZN(n4965) );
  NAND2_X1 U5512 ( .A1(n4939), .A2(n4965), .ZN(n4948) );
  NAND2_X1 U5513 ( .A1(n4948), .A2(n6323), .ZN(n5065) );
  NAND2_X1 U5514 ( .A1(n4940), .A2(n5065), .ZN(n4941) );
  OAI21_X1 U5515 ( .B1(n4942), .B2(n4941), .A(n7292), .ZN(n4945) );
  AOI21_X1 U5516 ( .B1(n3984), .B2(n3983), .A(n5239), .ZN(n4943) );
  NAND2_X1 U5517 ( .A1(n5367), .A2(n4943), .ZN(n4944) );
  INV_X1 U5518 ( .A(n4946), .ZN(n4952) );
  INV_X1 U5519 ( .A(n4947), .ZN(n7273) );
  INV_X1 U5520 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U5521 ( .A1(n4950), .A2(n5246), .ZN(n4951) );
  NAND4_X1 U5522 ( .A1(n4952), .A2(n7273), .A3(n6319), .A4(n4951), .ZN(n4953)
         );
  NOR2_X1 U5523 ( .A1(n6441), .A2(n4955), .ZN(n4956) );
  OR2_X1 U5524 ( .A1(n4954), .A2(n4956), .ZN(n6437) );
  NAND2_X1 U5525 ( .A1(n3985), .A2(n3925), .ZN(n4958) );
  OR2_X1 U5526 ( .A1(n5142), .A2(n4958), .ZN(n4959) );
  AND2_X1 U5527 ( .A1(n7289), .A2(n4959), .ZN(n4960) );
  NOR2_X2 U5528 ( .A1(n4983), .A2(n4960), .ZN(n7065) );
  NAND2_X1 U5529 ( .A1(n7183), .A2(REIP_REG_24__SCAN_IN), .ZN(n6522) );
  OAI21_X1 U5530 ( .B1(n6437), .B2(n7029), .A(n6522), .ZN(n4961) );
  INV_X1 U5531 ( .A(n4961), .ZN(n4996) );
  INV_X1 U5532 ( .A(n6974), .ZN(n4970) );
  OR2_X1 U5533 ( .A1(n4962), .A2(n5121), .ZN(n4973) );
  NAND2_X1 U5534 ( .A1(n4963), .A2(n5226), .ZN(n5580) );
  OR2_X1 U5535 ( .A1(n5580), .A2(n5239), .ZN(n5064) );
  OAI21_X1 U5536 ( .B1(n3984), .B2(n3983), .A(n5239), .ZN(n4964) );
  AND4_X1 U5537 ( .A1(n4973), .A2(n4965), .A3(n5064), .A4(n4964), .ZN(n4966)
         );
  NAND2_X1 U5538 ( .A1(n4975), .A2(n4966), .ZN(n5076) );
  NAND2_X1 U5539 ( .A1(n6245), .A2(n4967), .ZN(n6680) );
  OAI21_X1 U5540 ( .B1(n5142), .B2(n3939), .A(n6680), .ZN(n4968) );
  NOR2_X1 U5541 ( .A1(n5076), .A2(n4968), .ZN(n4969) );
  NOR2_X1 U5542 ( .A1(n4983), .A2(n4969), .ZN(n5128) );
  NAND2_X1 U5543 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5128), .ZN(n5041)
         );
  NAND2_X1 U5544 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U5545 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5314) );
  INV_X1 U5546 ( .A(n5314), .ZN(n5322) );
  NAND3_X1 U5547 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n5322), .ZN(n7004) );
  NOR2_X1 U5548 ( .A1(n7022), .A2(n7004), .ZN(n7026) );
  NAND3_X1 U5549 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n7026), .ZN(n6160) );
  NOR3_X1 U5550 ( .A1(n4086), .A2(n5268), .A3(n6160), .ZN(n5044) );
  INV_X1 U5551 ( .A(n5044), .ZN(n5042) );
  NAND3_X1 U5552 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6973) );
  NOR2_X1 U5553 ( .A1(n4219), .A2(n6973), .ZN(n6652) );
  NAND3_X1 U5554 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6652), .ZN(n4977) );
  NOR2_X1 U5555 ( .A1(n5042), .A2(n4977), .ZN(n5031) );
  NAND2_X1 U5556 ( .A1(n6644), .A2(n5031), .ZN(n6638) );
  INV_X1 U5557 ( .A(n6638), .ZN(n4971) );
  NAND2_X1 U5558 ( .A1(n4971), .A2(n6647), .ZN(n4984) );
  AND2_X1 U5559 ( .A1(n4973), .A2(n4972), .ZN(n4974) );
  NOR2_X1 U5560 ( .A1(n7055), .A2(n4977), .ZN(n5045) );
  AOI21_X1 U5561 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5313) );
  NOR2_X1 U5562 ( .A1(n5313), .A2(n6160), .ZN(n5040) );
  NAND2_X1 U5563 ( .A1(n5045), .A2(n5040), .ZN(n5030) );
  NAND2_X1 U5564 ( .A1(n6647), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4978) );
  NOR2_X1 U5565 ( .A1(n5030), .A2(n4978), .ZN(n4982) );
  INV_X1 U5566 ( .A(n4982), .ZN(n4979) );
  OR2_X1 U5567 ( .A1(n5316), .A2(n4979), .ZN(n4980) );
  INV_X1 U5568 ( .A(n6622), .ZN(n6529) );
  OR2_X1 U5569 ( .A1(n7064), .A2(n6529), .ZN(n6630) );
  OR2_X1 U5570 ( .A1(n5316), .A2(n4982), .ZN(n4986) );
  OR2_X1 U5571 ( .A1(n6974), .A2(n5128), .ZN(n6639) );
  INV_X1 U5572 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5120) );
  AOI22_X1 U5573 ( .A1(n7105), .A2(n4983), .B1(n5120), .B2(n5128), .ZN(n5127)
         );
  INV_X1 U5574 ( .A(n5127), .ZN(n5311) );
  AOI21_X1 U5575 ( .B1(n6639), .B2(n4984), .A(n5311), .ZN(n4985) );
  NAND2_X1 U5576 ( .A1(n4986), .A2(n4985), .ZN(n7060) );
  INV_X1 U5577 ( .A(n7060), .ZN(n4987) );
  NAND2_X1 U5578 ( .A1(n6992), .A2(n5316), .ZN(n4989) );
  NAND2_X1 U5579 ( .A1(n4989), .A2(n4988), .ZN(n4990) );
  NAND2_X1 U5580 ( .A1(n6628), .A2(n4990), .ZN(n7069) );
  INV_X1 U5581 ( .A(n7069), .ZN(n4995) );
  NAND2_X1 U5582 ( .A1(n6529), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4992) );
  OAI21_X1 U5583 ( .B1(n7064), .B2(n4992), .A(n4991), .ZN(n4993) );
  INV_X1 U5584 ( .A(n4993), .ZN(n4994) );
  OAI21_X1 U5585 ( .B1(n6526), .B2(n7023), .A(n3770), .ZN(U2994) );
  NAND2_X1 U5586 ( .A1(n4997), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U5587 ( .A1(n6223), .A2(n3776), .ZN(n5001) );
  INV_X1 U5588 ( .A(n4998), .ZN(n4999) );
  INV_X1 U5589 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U5590 ( .A1(n4999), .A2(n3777), .ZN(n5000) );
  NAND2_X1 U5591 ( .A1(n5001), .A2(n5000), .ZN(n5002) );
  XNOR2_X1 U5592 ( .A(n5002), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5018)
         );
  INV_X1 U5593 ( .A(n6427), .ZN(n5003) );
  NAND2_X1 U5594 ( .A1(n5003), .A2(n7065), .ZN(n5012) );
  INV_X1 U5595 ( .A(n6639), .ZN(n5032) );
  NAND2_X1 U5596 ( .A1(n5032), .A2(n5316), .ZN(n7021) );
  INV_X1 U5597 ( .A(n7021), .ZN(n5272) );
  INV_X1 U5598 ( .A(n5004), .ZN(n5005) );
  AND2_X1 U5599 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6610) );
  OAI21_X1 U5600 ( .B1(n5272), .B2(n6610), .A(n4995), .ZN(n6607) );
  AOI21_X1 U5601 ( .B1(n7021), .B2(n5005), .A(n6607), .ZN(n6584) );
  OAI21_X1 U5602 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5272), .A(n6584), 
        .ZN(n5010) );
  INV_X1 U5603 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6836) );
  NOR2_X1 U5604 ( .A1(n7105), .A2(n6836), .ZN(n5014) );
  INV_X1 U5605 ( .A(n5006), .ZN(n5007) );
  NOR2_X1 U5606 ( .A1(n7064), .A2(n5007), .ZN(n7070) );
  NAND2_X1 U5607 ( .A1(n7070), .A2(n6610), .ZN(n6597) );
  OR2_X1 U5608 ( .A1(n6597), .A2(n5008), .ZN(n6585) );
  NOR4_X1 U5609 ( .A1(n6585), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6586), 
        .A4(n6578), .ZN(n5009) );
  AOI211_X1 U5610 ( .C1(n5010), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5014), .B(n5009), .ZN(n5011) );
  OAI21_X1 U5611 ( .B1(n5018), .B2(n7023), .A(n5013), .ZN(U2987) );
  AOI21_X1 U5612 ( .B1(n6932), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5014), 
        .ZN(n5015) );
  OAI21_X1 U5613 ( .B1(n5018), .B2(n7241), .A(n5017), .ZN(U2955) );
  NAND2_X1 U5614 ( .A1(n6325), .A2(n6254), .ZN(n5066) );
  INV_X1 U5615 ( .A(n6233), .ZN(n6310) );
  NAND3_X1 U5616 ( .A1(n6310), .A2(n3925), .A3(n3926), .ZN(n5141) );
  INV_X1 U5617 ( .A(n5141), .ZN(n5020) );
  NAND3_X1 U5618 ( .A1(n5020), .A2(n5019), .A3(n5099), .ZN(n5021) );
  NAND2_X1 U5619 ( .A1(n5066), .A2(n5021), .ZN(n5022) );
  NAND2_X1 U5620 ( .A1(n6880), .A2(n6233), .ZN(n6478) );
  NAND2_X1 U5621 ( .A1(n6479), .A2(n6878), .ZN(n5029) );
  XNOR2_X1 U5622 ( .A(n5026), .B(n5025), .ZN(n6574) );
  INV_X1 U5623 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U5624 ( .A1(n5029), .A2(n5028), .ZN(U2829) );
  AOI21_X1 U5625 ( .B1(n6995), .B2(n5030), .A(n5311), .ZN(n6642) );
  OAI21_X1 U5626 ( .B1(n5032), .B2(n5031), .A(n6642), .ZN(n7054) );
  INV_X1 U5627 ( .A(n7054), .ZN(n5033) );
  OAI21_X1 U5628 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6992), .A(n5033), 
        .ZN(n5039) );
  AOI21_X1 U5629 ( .B1(n5034), .B2(n6466), .A(n3704), .ZN(n6410) );
  NOR2_X1 U5630 ( .A1(n5035), .A2(n4212), .ZN(n6530) );
  NOR3_X1 U5631 ( .A1(n5036), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n3650), 
        .ZN(n5037) );
  AOI21_X1 U5632 ( .B1(n6530), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5037), 
        .ZN(n5038) );
  AOI222_X1 U5633 ( .A1(n5039), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n7065), .B2(n6410), .C1(n6552), .C2(n7066), .ZN(n5047) );
  INV_X1 U5634 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6640) );
  INV_X1 U5635 ( .A(n5040), .ZN(n5043) );
  OAI22_X1 U5636 ( .A1(n5316), .A2(n5043), .B1(n5042), .B2(n5041), .ZN(n6983)
         );
  AOI21_X1 U5637 ( .B1(n6974), .B2(n5044), .A(n6983), .ZN(n6981) );
  INV_X1 U5638 ( .A(n6981), .ZN(n6161) );
  NAND3_X1 U5639 ( .A1(n5045), .A2(n6640), .A3(n6161), .ZN(n5046) );
  NAND3_X1 U5640 ( .A1(n5047), .A2(n5046), .A3(n3773), .ZN(U3000) );
  INV_X1 U5641 ( .A(n5048), .ZN(n5054) );
  INV_X1 U5642 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n5052) );
  INV_X1 U5643 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U5644 ( .A1(n5140), .A2(n5050), .ZN(n5055) );
  INV_X1 U5645 ( .A(n5055), .ZN(n5051) );
  OAI21_X1 U5646 ( .B1(n5054), .B2(n5052), .A(n5051), .ZN(U2788) );
  INV_X1 U5647 ( .A(n6953), .ZN(n5057) );
  INV_X1 U5648 ( .A(n5580), .ZN(n5053) );
  OR2_X1 U5649 ( .A1(n5053), .A2(n4017), .ZN(n6330) );
  NOR3_X1 U5650 ( .A1(n5055), .A2(n5054), .A3(READREQUEST_REG_SCAN_IN), .ZN(
        n5056) );
  AOI21_X1 U5651 ( .B1(n5057), .B2(n6330), .A(n5056), .ZN(U3474) );
  NAND2_X1 U5652 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n7313), .ZN(n7304) );
  INV_X1 U5653 ( .A(n7304), .ZN(n5070) );
  OR2_X1 U5654 ( .A1(n6325), .A2(n6319), .ZN(n5060) );
  INV_X1 U5655 ( .A(n5074), .ZN(n7245) );
  NAND2_X1 U5656 ( .A1(n7245), .A2(n5058), .ZN(n5059) );
  NAND2_X1 U5657 ( .A1(n5060), .A2(n5059), .ZN(n5144) );
  INV_X1 U5658 ( .A(n5144), .ZN(n5069) );
  INV_X1 U5659 ( .A(n5061), .ZN(n5063) );
  NAND2_X1 U5660 ( .A1(n7257), .A2(n5364), .ZN(n5365) );
  NAND2_X1 U5661 ( .A1(n5365), .A2(n4798), .ZN(n5062) );
  NAND2_X1 U5662 ( .A1(n5063), .A2(n5062), .ZN(n5068) );
  AND3_X1 U5663 ( .A1(n5066), .A2(n5065), .A3(n5064), .ZN(n5067) );
  NAND2_X1 U5664 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n7306) );
  OR2_X1 U5665 ( .A1(n7313), .A2(n7306), .ZN(n7303) );
  INV_X1 U5666 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7242) );
  OAI22_X1 U5667 ( .A1(n7271), .A2(n7318), .B1(n7303), .B2(n7242), .ZN(n7248)
         );
  NOR2_X1 U5668 ( .A1(n5072), .A2(n5071), .ZN(n5081) );
  NAND3_X1 U5669 ( .A1(n5074), .A2(n4933), .A3(n5142), .ZN(n5075) );
  OR2_X1 U5670 ( .A1(n5076), .A2(n5075), .ZN(n6688) );
  INV_X1 U5671 ( .A(n6688), .ZN(n5077) );
  OR2_X1 U5672 ( .A1(n5073), .A2(n5077), .ZN(n5078) );
  NAND2_X1 U5673 ( .A1(n7257), .A2(n4297), .ZN(n6675) );
  OAI211_X1 U5674 ( .C1(n5081), .C2(n5079), .A(n5078), .B(n6675), .ZN(n7258)
         );
  INV_X1 U5675 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5080) );
  AOI22_X1 U5676 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5080), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5268), .ZN(n6262) );
  NAND2_X1 U5677 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6261) );
  INV_X1 U5678 ( .A(n6261), .ZN(n5083) );
  INV_X1 U5679 ( .A(n5081), .ZN(n5082) );
  AOI222_X1 U5680 ( .A1(n7258), .A2(n7294), .B1(n6262), .B2(n5083), .C1(n5082), 
        .C2(n6689), .ZN(n5085) );
  NAND2_X1 U5681 ( .A1(n7244), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5084) );
  OAI21_X1 U5682 ( .B1(n7244), .B2(n5085), .A(n5084), .ZN(U3460) );
  INV_X1 U5683 ( .A(n5087), .ZN(n5090) );
  INV_X1 U5684 ( .A(n5088), .ZN(n5096) );
  NAND3_X1 U5685 ( .A1(n5090), .A2(n5089), .A3(n5096), .ZN(n5091) );
  AND2_X1 U5686 ( .A1(n5086), .A2(n5091), .ZN(n7077) );
  INV_X1 U5687 ( .A(n7077), .ZN(n5332) );
  INV_X1 U5688 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U5689 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  NAND2_X1 U5690 ( .A1(n5135), .A2(n5094), .ZN(n7079) );
  OAI222_X1 U5691 ( .A1(n5332), .A2(n6478), .B1(n5095), .B2(n6880), .C1(n7079), 
        .C2(n6876), .ZN(U2857) );
  OAI21_X1 U5692 ( .B1(n5098), .B2(n5097), .A(n5096), .ZN(n6888) );
  OR2_X1 U5693 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  NAND2_X1 U5694 ( .A1(n5102), .A2(n5101), .ZN(n6422) );
  AOI22_X1 U5695 ( .A1(n6868), .A2(n6422), .B1(EBX_REG_1__SCAN_IN), .B2(n6475), 
        .ZN(n5103) );
  OAI21_X1 U5696 ( .B1(n6468), .B2(n6888), .A(n5103), .ZN(U2858) );
  INV_X1 U5697 ( .A(n6671), .ZN(n5105) );
  OAI21_X1 U5698 ( .B1(n5105), .B2(n5104), .A(n7250), .ZN(n5106) );
  NAND2_X1 U5699 ( .A1(n5106), .A2(n7242), .ZN(n7308) );
  NAND2_X1 U5700 ( .A1(n7308), .A2(n7242), .ZN(n5108) );
  INV_X1 U5701 ( .A(n7303), .ZN(n5107) );
  NAND2_X1 U5702 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  NAND2_X1 U5703 ( .A1(n5419), .A2(n5109), .ZN(n7328) );
  INV_X1 U5704 ( .A(n3662), .ZN(n6005) );
  OAI21_X1 U5705 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7296), .A(n7328), .ZN(
        n7320) );
  NAND2_X1 U5706 ( .A1(n7328), .A2(n7457), .ZN(n7325) );
  INV_X1 U5707 ( .A(n5112), .ZN(n7431) );
  AOI21_X1 U5708 ( .B1(n3654), .B2(STATEBS16_REG_SCAN_IN), .A(n7431), .ZN(
        n5118) );
  INV_X1 U5709 ( .A(n4115), .ZN(n5113) );
  NAND2_X1 U5710 ( .A1(n3654), .A2(n5113), .ZN(n5162) );
  INV_X1 U5711 ( .A(n5162), .ZN(n5115) );
  AND2_X1 U5712 ( .A1(n4115), .A2(n5114), .ZN(n5116) );
  NAND2_X1 U5713 ( .A1(n3654), .A2(n5116), .ZN(n7369) );
  AOI21_X1 U5714 ( .B1(n7404), .B2(n7369), .A(n7330), .ZN(n5117) );
  NOR2_X1 U5715 ( .A1(n5118), .A2(n5117), .ZN(n5119) );
  OAI222_X1 U5716 ( .A1(n7328), .A2(n7268), .B1(n6005), .B2(n7320), .C1(n7325), 
        .C2(n5119), .ZN(U3462) );
  NAND2_X1 U5717 ( .A1(n5121), .A2(n5120), .ZN(n5123) );
  NAND2_X1 U5718 ( .A1(n5123), .A2(n5122), .ZN(n5578) );
  INV_X1 U5719 ( .A(n5269), .ZN(n5124) );
  OAI21_X1 U5720 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5125), .A(n5124), 
        .ZN(n6887) );
  INV_X1 U5721 ( .A(n6887), .ZN(n5126) );
  AND2_X1 U5722 ( .A1(n7183), .A2(REIP_REG_0__SCAN_IN), .ZN(n6882) );
  AOI21_X1 U5723 ( .B1(n7066), .B2(n5126), .A(n6882), .ZN(n5130) );
  OAI21_X1 U5724 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5316), .A(n5127), 
        .ZN(n5275) );
  OR2_X1 U5725 ( .A1(n6995), .A2(n5128), .ZN(n6971) );
  OAI22_X1 U5726 ( .A1(n6974), .A2(n5275), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6971), .ZN(n5129) );
  OAI211_X1 U5727 ( .C1(n7029), .C2(n5578), .A(n5130), .B(n5129), .ZN(U3018)
         );
  AND2_X1 U5728 ( .A1(n5132), .A2(n5086), .ZN(n5133) );
  OR2_X1 U5729 ( .A1(n5131), .A2(n5133), .ZN(n6018) );
  INV_X1 U5730 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6006) );
  AND2_X1 U5731 ( .A1(n5135), .A2(n5134), .ZN(n5136) );
  NOR2_X1 U5732 ( .A1(n5154), .A2(n5136), .ZN(n5201) );
  INV_X1 U5733 ( .A(n5201), .ZN(n6007) );
  OAI222_X1 U5734 ( .A1(n6018), .A2(n6478), .B1(n6006), .B2(n6880), .C1(n6007), 
        .C2(n6876), .ZN(U2856) );
  XOR2_X1 U5735 ( .A(n5138), .B(n5137), .Z(n6881) );
  INV_X1 U5736 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5139) );
  OAI222_X1 U5737 ( .A1(n5578), .A2(n6876), .B1(n6468), .B2(n6881), .C1(n5139), 
        .C2(n6880), .ZN(U2859) );
  NOR2_X1 U5738 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U5739 ( .A1(n5146), .A2(n6233), .ZN(n5147) );
  INV_X1 U5740 ( .A(n5147), .ZN(n5148) );
  INV_X1 U5741 ( .A(DATAI_0_), .ZN(n5214) );
  INV_X1 U5742 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6757) );
  OAI222_X1 U5743 ( .A1(n7352), .A2(n6881), .B1(n6219), .B2(n5214), .C1(n6311), 
        .C2(n6757), .ZN(U2891) );
  OAI21_X1 U5744 ( .B1(n5131), .B2(n5151), .A(n5150), .ZN(n7098) );
  INV_X1 U5745 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5156) );
  OR2_X1 U5746 ( .A1(n5154), .A2(n5153), .ZN(n5155) );
  NAND2_X1 U5747 ( .A1(n5152), .A2(n5155), .ZN(n7093) );
  OAI222_X1 U5748 ( .A1(n7098), .A2(n6478), .B1(n6880), .B2(n5156), .C1(n7093), 
        .C2(n6876), .ZN(U2855) );
  INV_X1 U5749 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6765) );
  INV_X1 U5750 ( .A(DATAI_4_), .ZN(n5247) );
  OAI222_X1 U5751 ( .A1(n7098), .A2(n7352), .B1(n6311), .B2(n6765), .C1(n6219), 
        .C2(n5247), .ZN(U2887) );
  NOR3_X1 U5752 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6251), .ZN(n7421) );
  INV_X1 U5753 ( .A(n7421), .ZN(n7425) );
  OR2_X1 U5754 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7425), .ZN(n6301)
         );
  NOR2_X1 U5755 ( .A1(n5159), .A2(n5114), .ZN(n6058) );
  INV_X1 U5756 ( .A(n6058), .ZN(n5160) );
  NOR2_X1 U5757 ( .A1(n5160), .A2(n5112), .ZN(n5380) );
  NAND2_X1 U5758 ( .A1(n5380), .A2(n5161), .ZN(n5167) );
  NAND2_X1 U5759 ( .A1(n7420), .A2(n7324), .ZN(n7422) );
  AOI21_X1 U5760 ( .B1(n5167), .B2(n7422), .A(n7330), .ZN(n5166) );
  INV_X1 U5761 ( .A(n5073), .ZN(n6420) );
  NOR2_X1 U5762 ( .A1(n5163), .A2(n6420), .ZN(n7417) );
  NOR2_X1 U5763 ( .A1(n7417), .A2(n7445), .ZN(n6060) );
  NOR2_X1 U5764 ( .A1(n6060), .A2(n6093), .ZN(n5165) );
  NOR2_X1 U5765 ( .A1(n3779), .A2(n7295), .ZN(n5336) );
  OR2_X1 U5766 ( .A1(n5168), .A2(n7295), .ZN(n5287) );
  NAND2_X1 U5767 ( .A1(n5280), .A2(n5287), .ZN(n6095) );
  AOI211_X1 U5768 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6301), .A(n5336), .B(
        n6095), .ZN(n5164) );
  NAND2_X1 U5769 ( .A1(n6295), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U5770 ( .A1(n6937), .A2(DATAI_30_), .ZN(n6108) );
  INV_X1 U5771 ( .A(n6108), .ZN(n7593) );
  NAND2_X1 U5772 ( .A1(n6937), .A2(DATAI_22_), .ZN(n5973) );
  NAND2_X1 U5773 ( .A1(n6103), .A2(n7417), .ZN(n5170) );
  NAND2_X1 U5774 ( .A1(n5168), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5279) );
  INV_X1 U5775 ( .A(n5279), .ZN(n6101) );
  NAND2_X1 U5776 ( .A1(n3779), .A2(n6101), .ZN(n5169) );
  NAND2_X1 U5777 ( .A1(DATAI_6_), .A2(n5280), .ZN(n7596) );
  OAI22_X1 U5778 ( .A1(n7422), .A2(n5973), .B1(n6296), .B2(n7596), .ZN(n5171)
         );
  AOI21_X1 U5779 ( .B1(n7593), .B2(n7637), .A(n5171), .ZN(n5172) );
  OAI211_X1 U5780 ( .C1(n6301), .C2(n6112), .A(n5173), .B(n5172), .ZN(U3058)
         );
  CLKBUF_X1 U5781 ( .A(n5174), .Z(n5176) );
  NAND2_X1 U5782 ( .A1(n5176), .A2(n5175), .ZN(n5178) );
  XNOR2_X1 U5783 ( .A(n5178), .B(n5177), .ZN(n5204) );
  INV_X1 U5784 ( .A(n6018), .ZN(n5181) );
  AND2_X1 U5785 ( .A1(n7183), .A2(REIP_REG_3__SCAN_IN), .ZN(n5200) );
  AOI21_X1 U5786 ( .B1(n6932), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5200), 
        .ZN(n5179) );
  OAI21_X1 U5787 ( .B1(n6008), .B2(n6940), .A(n5179), .ZN(n5180) );
  AOI21_X1 U5788 ( .B1(n5181), .B2(n6937), .A(n5180), .ZN(n5182) );
  OAI21_X1 U5789 ( .B1(n5204), .B2(n7241), .A(n5182), .ZN(U2983) );
  INV_X1 U5790 ( .A(DATAI_3_), .ZN(n5184) );
  INV_X1 U5791 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6763) );
  OAI222_X1 U5792 ( .A1(n5184), .A2(n6219), .B1(n6311), .B2(n6763), .C1(n7352), 
        .C2(n6018), .ZN(U2888) );
  INV_X1 U5793 ( .A(n7533), .ZN(n6117) );
  NAND2_X1 U5794 ( .A1(n6295), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U5795 ( .A1(n6937), .A2(DATAI_27_), .ZN(n6113) );
  INV_X1 U5796 ( .A(n6113), .ZN(n7535) );
  AND2_X1 U5797 ( .A1(n6937), .A2(DATAI_19_), .ZN(n7534) );
  INV_X1 U5798 ( .A(n7534), .ZN(n5428) );
  NOR2_X1 U5799 ( .A1(n5184), .A2(n5419), .ZN(n6066) );
  OAI22_X1 U5800 ( .A1(n7422), .A2(n5428), .B1(n6296), .B2(n7538), .ZN(n5185)
         );
  AOI21_X1 U5801 ( .B1(n7535), .B2(n7637), .A(n5185), .ZN(n5186) );
  OAI211_X1 U5802 ( .C1(n6301), .C2(n6117), .A(n5187), .B(n5186), .ZN(U3055)
         );
  OR2_X1 U5803 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5424), .ZN(n6280)
         );
  AOI21_X1 U5804 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n5382), .A(n7295), 
        .ZN(n5968) );
  AOI211_X1 U5805 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6280), .A(n5968), .B(
        n6095), .ZN(n5192) );
  NOR2_X1 U5806 ( .A1(n5163), .A2(n5073), .ZN(n7409) );
  NOR2_X1 U5807 ( .A1(n7409), .A2(n7445), .ZN(n6094) );
  NOR2_X2 U5808 ( .A1(n7369), .A2(n7324), .ZN(n7599) );
  AND2_X1 U5809 ( .A1(n4115), .A2(n5281), .ZN(n5188) );
  INV_X1 U5810 ( .A(n5421), .ZN(n5189) );
  NOR2_X1 U5811 ( .A1(n5189), .A2(n5161), .ZN(n5430) );
  OAI21_X1 U5812 ( .B1(n7599), .B2(n5430), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5190) );
  OAI21_X1 U5813 ( .B1(n6103), .B2(n6094), .A(n5190), .ZN(n5191) );
  NAND2_X1 U5814 ( .A1(n5192), .A2(n5191), .ZN(n6274) );
  NAND2_X1 U5815 ( .A1(n6274), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5195)
         );
  INV_X1 U5816 ( .A(n5382), .ZN(n5286) );
  NOR2_X1 U5817 ( .A1(n5286), .A2(n7268), .ZN(n5974) );
  AOI22_X1 U5818 ( .A1(n6093), .A2(n7409), .B1(n5974), .B2(n6101), .ZN(n6275)
         );
  OAI22_X1 U5819 ( .A1(n6276), .A2(n5973), .B1(n6275), .B2(n7596), .ZN(n5193)
         );
  AOI21_X1 U5820 ( .B1(n7593), .B2(n7599), .A(n5193), .ZN(n5194) );
  OAI211_X1 U5821 ( .C1(n6280), .C2(n6112), .A(n5195), .B(n5194), .ZN(U3138)
         );
  NAND2_X1 U5822 ( .A1(n6274), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5198)
         );
  OAI22_X1 U5823 ( .A1(n6276), .A2(n5428), .B1(n6275), .B2(n7538), .ZN(n5196)
         );
  AOI21_X1 U5824 ( .B1(n7535), .B2(n7599), .A(n5196), .ZN(n5197) );
  OAI211_X1 U5825 ( .C1(n6280), .C2(n6117), .A(n5198), .B(n5197), .ZN(U3135)
         );
  NAND2_X1 U5826 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5199) );
  AOI21_X1 U5827 ( .B1(n6639), .B2(n5199), .A(n5311), .ZN(n7002) );
  NAND2_X1 U5828 ( .A1(n6995), .A2(n5313), .ZN(n6997) );
  NAND2_X1 U5829 ( .A1(n7002), .A2(n6997), .ZN(n6159) );
  NOR2_X1 U5830 ( .A1(n6992), .A2(n5199), .ZN(n5321) );
  NOR2_X1 U5831 ( .A1(n6995), .A2(n5321), .ZN(n5441) );
  NOR2_X1 U5832 ( .A1(n5313), .A2(n5441), .ZN(n7025) );
  AOI22_X1 U5833 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n6159), .B1(n7025), 
        .B2(n4111), .ZN(n5203) );
  AOI21_X1 U5834 ( .B1(n7065), .B2(n5201), .A(n5200), .ZN(n5202) );
  OAI211_X1 U5835 ( .C1(n5204), .C2(n7023), .A(n5203), .B(n5202), .ZN(U3015)
         );
  NAND2_X1 U5836 ( .A1(n5475), .A2(DATAI_5_), .ZN(n5482) );
  AOI22_X1 U5837 ( .A1(n5487), .A2(EAX_REG_21__SCAN_IN), .B1(n5448), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U5838 ( .A1(n5482), .A2(n5207), .ZN(U2929) );
  NAND2_X1 U5839 ( .A1(n5475), .A2(DATAI_3_), .ZN(n5455) );
  AOI22_X1 U5840 ( .A1(n5487), .A2(EAX_REG_19__SCAN_IN), .B1(n5448), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U5841 ( .A1(n5455), .A2(n5208), .ZN(U2927) );
  NAND2_X1 U5842 ( .A1(n5475), .A2(DATAI_7_), .ZN(n5465) );
  AOI22_X1 U5843 ( .A1(n5487), .A2(EAX_REG_23__SCAN_IN), .B1(n5448), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U5844 ( .A1(n5465), .A2(n5209), .ZN(U2931) );
  NAND2_X1 U5845 ( .A1(n5475), .A2(DATAI_6_), .ZN(n5467) );
  AOI22_X1 U5846 ( .A1(n5487), .A2(EAX_REG_22__SCAN_IN), .B1(n5448), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U5847 ( .A1(n5467), .A2(n5210), .ZN(U2930) );
  NAND2_X1 U5848 ( .A1(n5475), .A2(DATAI_2_), .ZN(n5457) );
  AOI22_X1 U5849 ( .A1(n5487), .A2(EAX_REG_18__SCAN_IN), .B1(n5448), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U5850 ( .A1(n5457), .A2(n5211), .ZN(U2926) );
  NAND2_X1 U5851 ( .A1(n5475), .A2(DATAI_4_), .ZN(n5453) );
  AOI22_X1 U5852 ( .A1(n5487), .A2(EAX_REG_20__SCAN_IN), .B1(n5448), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U5853 ( .A1(n5453), .A2(n5212), .ZN(U2928) );
  NAND2_X1 U5854 ( .A1(n5405), .A2(n3983), .ZN(n6107) );
  NAND2_X1 U5855 ( .A1(n6274), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5217)
         );
  NAND2_X1 U5856 ( .A1(n6937), .A2(DATAI_24_), .ZN(n6694) );
  INV_X1 U5857 ( .A(n6694), .ZN(n7462) );
  AND2_X1 U5858 ( .A1(n6937), .A2(DATAI_16_), .ZN(n7454) );
  INV_X1 U5859 ( .A(n7454), .ZN(n5511) );
  NOR2_X1 U5860 ( .A1(n5214), .A2(n5419), .ZN(n6693) );
  OAI22_X1 U5861 ( .A1(n6276), .A2(n5511), .B1(n6275), .B2(n7465), .ZN(n5215)
         );
  AOI21_X1 U5862 ( .B1(n7462), .B2(n7599), .A(n5215), .ZN(n5216) );
  OAI211_X1 U5863 ( .C1(n6107), .C2(n6280), .A(n5217), .B(n5216), .ZN(U3132)
         );
  NAND2_X1 U5864 ( .A1(n6295), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5220) );
  OAI22_X1 U5865 ( .A1(n7422), .A2(n5511), .B1(n6296), .B2(n7465), .ZN(n5218)
         );
  AOI21_X1 U5866 ( .B1(n7462), .B2(n7637), .A(n5218), .ZN(n5219) );
  OAI211_X1 U5867 ( .C1(n6107), .C2(n6301), .A(n5220), .B(n5219), .ZN(U3052)
         );
  XOR2_X1 U5868 ( .A(n5222), .B(n5221), .Z(n5263) );
  NAND2_X1 U5869 ( .A1(n5263), .A2(n6936), .ZN(n5225) );
  NOR2_X1 U5870 ( .A1(n7105), .A2(n7086), .ZN(n5262) );
  NOR2_X1 U5871 ( .A1(n6940), .A2(n7096), .ZN(n5223) );
  AOI211_X1 U5872 ( .C1(n6932), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5262), 
        .B(n5223), .ZN(n5224) );
  OAI211_X1 U5873 ( .C1(n6914), .C2(n7098), .A(n5225), .B(n5224), .ZN(U2982)
         );
  NAND2_X1 U5874 ( .A1(n5405), .A2(n5226), .ZN(n6701) );
  NAND2_X1 U5875 ( .A1(n6295), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U5876 ( .A1(n6937), .A2(DATAI_25_), .ZN(n6122) );
  INV_X1 U5877 ( .A(n6122), .ZN(n7485) );
  AND2_X1 U5878 ( .A1(n6937), .A2(DATAI_17_), .ZN(n7484) );
  INV_X1 U5879 ( .A(n7484), .ZN(n5518) );
  INV_X1 U5880 ( .A(DATAI_1_), .ZN(n5327) );
  NOR2_X1 U5881 ( .A1(n5327), .A2(n5419), .ZN(n6700) );
  OAI22_X1 U5882 ( .A1(n7422), .A2(n5518), .B1(n6296), .B2(n7488), .ZN(n5227)
         );
  AOI21_X1 U5883 ( .B1(n7485), .B2(n7637), .A(n5227), .ZN(n5228) );
  OAI211_X1 U5884 ( .C1(n6301), .C2(n6701), .A(n5229), .B(n5228), .ZN(U3053)
         );
  NAND2_X1 U5885 ( .A1(n6274), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5232)
         );
  OAI22_X1 U5886 ( .A1(n6276), .A2(n5518), .B1(n6275), .B2(n7488), .ZN(n5230)
         );
  AOI21_X1 U5887 ( .B1(n7485), .B2(n7599), .A(n5230), .ZN(n5231) );
  OAI211_X1 U5888 ( .C1(n6280), .C2(n6701), .A(n5232), .B(n5231), .ZN(U3133)
         );
  NAND2_X1 U5889 ( .A1(n5405), .A2(n6233), .ZN(n6732) );
  NAND2_X1 U5890 ( .A1(n6295), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U5891 ( .A1(n6937), .A2(DATAI_31_), .ZN(n6126) );
  INV_X1 U5892 ( .A(n6126), .ZN(n7648) );
  AND2_X1 U5893 ( .A1(n6937), .A2(DATAI_23_), .ZN(n7645) );
  INV_X1 U5894 ( .A(n7645), .ZN(n5522) );
  INV_X1 U5895 ( .A(DATAI_7_), .ZN(n5537) );
  NOR2_X1 U5896 ( .A1(n5537), .A2(n5419), .ZN(n6731) );
  OAI22_X1 U5897 ( .A1(n7422), .A2(n5522), .B1(n6296), .B2(n7652), .ZN(n5233)
         );
  AOI21_X1 U5898 ( .B1(n7648), .B2(n7637), .A(n5233), .ZN(n5234) );
  OAI211_X1 U5899 ( .C1(n6301), .C2(n6732), .A(n5235), .B(n5234), .ZN(U3059)
         );
  NAND2_X1 U5900 ( .A1(n6274), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5238)
         );
  OAI22_X1 U5901 ( .A1(n6276), .A2(n5522), .B1(n6275), .B2(n7652), .ZN(n5236)
         );
  AOI21_X1 U5902 ( .B1(n7648), .B2(n7599), .A(n5236), .ZN(n5237) );
  OAI211_X1 U5903 ( .C1(n6280), .C2(n6732), .A(n5238), .B(n5237), .ZN(U3139)
         );
  NAND2_X1 U5904 ( .A1(n5405), .A2(n5239), .ZN(n6707) );
  NAND2_X1 U5905 ( .A1(n6295), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5242) );
  AND2_X1 U5906 ( .A1(n6937), .A2(DATAI_26_), .ZN(n7508) );
  AND2_X1 U5907 ( .A1(n6937), .A2(DATAI_18_), .ZN(n7507) );
  INV_X1 U5908 ( .A(n7507), .ZN(n5503) );
  INV_X1 U5909 ( .A(DATAI_2_), .ZN(n5333) );
  NOR2_X1 U5910 ( .A1(n5333), .A2(n5419), .ZN(n6706) );
  OAI22_X1 U5911 ( .A1(n7422), .A2(n5503), .B1(n6296), .B2(n7511), .ZN(n5240)
         );
  AOI21_X1 U5912 ( .B1(n7508), .B2(n7637), .A(n5240), .ZN(n5241) );
  OAI211_X1 U5913 ( .C1(n6301), .C2(n6707), .A(n5242), .B(n5241), .ZN(U3054)
         );
  NAND2_X1 U5914 ( .A1(n6274), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5245)
         );
  OAI22_X1 U5915 ( .A1(n6276), .A2(n5503), .B1(n6275), .B2(n7511), .ZN(n5243)
         );
  AOI21_X1 U5916 ( .B1(n7508), .B2(n7599), .A(n5243), .ZN(n5244) );
  OAI211_X1 U5917 ( .C1(n6280), .C2(n6707), .A(n5245), .B(n5244), .ZN(U3134)
         );
  NAND2_X1 U5918 ( .A1(n5405), .A2(n5246), .ZN(n6713) );
  NAND2_X1 U5919 ( .A1(n6295), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5250) );
  AND2_X1 U5920 ( .A1(n6937), .A2(DATAI_28_), .ZN(n7555) );
  AND2_X1 U5921 ( .A1(n6937), .A2(DATAI_20_), .ZN(n7554) );
  INV_X1 U5922 ( .A(n7554), .ZN(n5507) );
  NOR2_X1 U5923 ( .A1(n5247), .A2(n5419), .ZN(n6712) );
  OAI22_X1 U5924 ( .A1(n7422), .A2(n5507), .B1(n6296), .B2(n7558), .ZN(n5248)
         );
  AOI21_X1 U5925 ( .B1(n7555), .B2(n7637), .A(n5248), .ZN(n5249) );
  OAI211_X1 U5926 ( .C1(n6301), .C2(n6713), .A(n5250), .B(n5249), .ZN(U3056)
         );
  NAND2_X1 U5927 ( .A1(n6274), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5253)
         );
  OAI22_X1 U5928 ( .A1(n6276), .A2(n5507), .B1(n6275), .B2(n7558), .ZN(n5251)
         );
  AOI21_X1 U5929 ( .B1(n7555), .B2(n7599), .A(n5251), .ZN(n5252) );
  OAI211_X1 U5930 ( .C1(n6280), .C2(n6713), .A(n5253), .B(n5252), .ZN(U3136)
         );
  NAND2_X1 U5931 ( .A1(n5150), .A2(n5256), .ZN(n5257) );
  AND2_X1 U5932 ( .A1(n5255), .A2(n5257), .ZN(n7113) );
  INV_X1 U5933 ( .A(n7113), .ZN(n5267) );
  INV_X1 U5934 ( .A(EBX_REG_5__SCAN_IN), .ZN(n7104) );
  NAND2_X1 U5935 ( .A1(n5152), .A2(n5259), .ZN(n5260) );
  NAND2_X1 U5936 ( .A1(n5258), .A2(n5260), .ZN(n7110) );
  OAI222_X1 U5937 ( .A1(n5267), .A2(n6468), .B1(n7104), .B2(n6880), .C1(n7110), 
        .C2(n6876), .ZN(U2854) );
  INV_X1 U5938 ( .A(n6159), .ZN(n7010) );
  INV_X1 U5939 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5266) );
  OAI211_X1 U5940 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n7025), .B(n5314), .ZN(n5265) );
  NOR2_X1 U5941 ( .A1(n7029), .A2(n7093), .ZN(n5261) );
  AOI211_X1 U5942 ( .C1(n5263), .C2(n7066), .A(n5262), .B(n5261), .ZN(n5264)
         );
  OAI211_X1 U5943 ( .C1(n7010), .C2(n5266), .A(n5265), .B(n5264), .ZN(U3014)
         );
  INV_X1 U5944 ( .A(DATAI_5_), .ZN(n5404) );
  OAI222_X1 U5945 ( .A1(n5404), .A2(n6219), .B1(n6311), .B2(n4330), .C1(n7352), 
        .C2(n5267), .ZN(U2886) );
  XNOR2_X1 U5946 ( .A(n5269), .B(n5268), .ZN(n5270) );
  XNOR2_X1 U5947 ( .A(n5271), .B(n5270), .ZN(n6893) );
  INV_X1 U5948 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6852) );
  NOR2_X1 U5949 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n6974), .ZN(n5273)
         );
  NOR3_X1 U5950 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5273), .A3(n5272), 
        .ZN(n5274) );
  AOI21_X1 U5951 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n5275), .A(n5274), 
        .ZN(n5276) );
  OAI21_X1 U5952 ( .B1(n7105), .B2(n6852), .A(n5276), .ZN(n5277) );
  AOI21_X1 U5953 ( .B1(n7065), .B2(n6422), .A(n5277), .ZN(n5278) );
  OAI21_X1 U5954 ( .B1(n6893), .B2(n7023), .A(n5278), .ZN(U3017) );
  NOR3_X1 U5955 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7268), .ZN(n7397) );
  INV_X1 U5956 ( .A(n7397), .ZN(n7398) );
  OR2_X1 U5957 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7398), .ZN(n6287)
         );
  AOI21_X1 U5958 ( .B1(n5285), .B2(n5286), .A(n7295), .ZN(n6056) );
  NAND2_X1 U5959 ( .A1(n5280), .A2(n5279), .ZN(n5967) );
  AOI211_X1 U5960 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6287), .A(n6056), .B(
        n5967), .ZN(n5284) );
  AND2_X1 U5961 ( .A1(n5163), .A2(n5073), .ZN(n7447) );
  NOR2_X1 U5962 ( .A1(n7447), .A2(n7445), .ZN(n5335) );
  NOR2_X1 U5963 ( .A1(n5111), .A2(n5281), .ZN(n5334) );
  NAND2_X1 U5964 ( .A1(n5334), .A2(n5112), .ZN(n7392) );
  OAI21_X1 U5965 ( .B1(n3771), .B2(n7625), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5282) );
  OAI21_X1 U5966 ( .B1(n6103), .B2(n5335), .A(n5282), .ZN(n5283) );
  NAND2_X1 U5967 ( .A1(n5284), .A2(n5283), .ZN(n6281) );
  NAND2_X1 U5968 ( .A1(n6281), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5292) );
  INV_X1 U5969 ( .A(n7508), .ZN(n6118) );
  NAND2_X1 U5970 ( .A1(n6093), .A2(n7447), .ZN(n5289) );
  AND2_X1 U5971 ( .A1(n5286), .A2(n5285), .ZN(n6063) );
  INV_X1 U5972 ( .A(n5287), .ZN(n5975) );
  NAND2_X1 U5973 ( .A1(n6063), .A2(n5975), .ZN(n5288) );
  OAI22_X1 U5974 ( .A1(n6283), .A2(n6118), .B1(n6282), .B2(n7511), .ZN(n5290)
         );
  AOI21_X1 U5975 ( .B1(n7507), .B2(n3771), .A(n5290), .ZN(n5291) );
  OAI211_X1 U5976 ( .C1(n6287), .C2(n6707), .A(n5292), .B(n5291), .ZN(U3086)
         );
  NAND2_X1 U5977 ( .A1(n6281), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5295) );
  OAI22_X1 U5978 ( .A1(n6283), .A2(n6694), .B1(n6282), .B2(n7465), .ZN(n5293)
         );
  AOI21_X1 U5979 ( .B1(n7454), .B2(n3771), .A(n5293), .ZN(n5294) );
  OAI211_X1 U5980 ( .C1(n6107), .C2(n6287), .A(n5295), .B(n5294), .ZN(U3084)
         );
  NAND2_X1 U5981 ( .A1(n6281), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5298) );
  OAI22_X1 U5982 ( .A1(n6283), .A2(n6122), .B1(n6282), .B2(n7488), .ZN(n5296)
         );
  AOI21_X1 U5983 ( .B1(n7484), .B2(n3771), .A(n5296), .ZN(n5297) );
  OAI211_X1 U5984 ( .C1(n6287), .C2(n6701), .A(n5298), .B(n5297), .ZN(U3085)
         );
  NAND2_X1 U5985 ( .A1(n6281), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5301) );
  INV_X1 U5986 ( .A(n5973), .ZN(n7592) );
  OAI22_X1 U5987 ( .A1(n6283), .A2(n6108), .B1(n6282), .B2(n7596), .ZN(n5299)
         );
  AOI21_X1 U5988 ( .B1(n7592), .B2(n3771), .A(n5299), .ZN(n5300) );
  OAI211_X1 U5989 ( .C1(n6287), .C2(n6112), .A(n5301), .B(n5300), .ZN(U3090)
         );
  NAND2_X1 U5990 ( .A1(n6281), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5304) );
  OAI22_X1 U5991 ( .A1(n6283), .A2(n6113), .B1(n6282), .B2(n7538), .ZN(n5302)
         );
  AOI21_X1 U5992 ( .B1(n7534), .B2(n3771), .A(n5302), .ZN(n5303) );
  OAI211_X1 U5993 ( .C1(n6287), .C2(n6117), .A(n5304), .B(n5303), .ZN(U3087)
         );
  NAND2_X1 U5994 ( .A1(n6281), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5307) );
  INV_X1 U5995 ( .A(n7555), .ZN(n6130) );
  OAI22_X1 U5996 ( .A1(n6283), .A2(n6130), .B1(n6282), .B2(n7558), .ZN(n5305)
         );
  AOI21_X1 U5997 ( .B1(n7554), .B2(n3771), .A(n5305), .ZN(n5306) );
  OAI211_X1 U5998 ( .C1(n6287), .C2(n6713), .A(n5307), .B(n5306), .ZN(U3088)
         );
  NAND2_X1 U5999 ( .A1(n6281), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5310) );
  OAI22_X1 U6000 ( .A1(n6283), .A2(n6126), .B1(n6282), .B2(n7652), .ZN(n5308)
         );
  AOI21_X1 U6001 ( .B1(n7645), .B2(n3771), .A(n5308), .ZN(n5309) );
  OAI211_X1 U6002 ( .C1(n6287), .C2(n6732), .A(n5310), .B(n5309), .ZN(U3091)
         );
  NOR3_X1 U6003 ( .A1(n5314), .A2(n5320), .A3(n5313), .ZN(n5439) );
  NOR2_X1 U6004 ( .A1(n5311), .A2(n7021), .ZN(n7009) );
  AOI21_X1 U6005 ( .B1(n7002), .B2(n5439), .A(n7009), .ZN(n5312) );
  INV_X1 U6006 ( .A(n5312), .ZN(n5443) );
  OR2_X1 U6007 ( .A1(n5314), .A2(n5313), .ZN(n5315) );
  OAI21_X1 U6008 ( .B1(n5316), .B2(n5315), .A(n5320), .ZN(n5317) );
  INV_X1 U6009 ( .A(n5317), .ZN(n5326) );
  XOR2_X1 U6010 ( .A(n5319), .B(n5318), .Z(n6903) );
  NAND3_X1 U6011 ( .A1(n5322), .A2(n5321), .A3(n5320), .ZN(n5323) );
  NAND2_X1 U6012 ( .A1(n7059), .A2(REIP_REG_5__SCAN_IN), .ZN(n6904) );
  OAI211_X1 U6013 ( .C1(n7029), .C2(n7110), .A(n5323), .B(n6904), .ZN(n5324)
         );
  AOI21_X1 U6014 ( .B1(n6903), .B2(n7066), .A(n5324), .ZN(n5325) );
  OAI21_X1 U6015 ( .B1(n5443), .B2(n5326), .A(n5325), .ZN(U3013) );
  INV_X1 U6016 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6759) );
  OAI222_X1 U6017 ( .A1(n6888), .A2(n7352), .B1(n6219), .B2(n5327), .C1(n6311), 
        .C2(n6759), .ZN(U2890) );
  XNOR2_X1 U6018 ( .A(n5255), .B(n4349), .ZN(n7126) );
  INV_X1 U6019 ( .A(n7126), .ZN(n5501) );
  NAND2_X1 U6020 ( .A1(n5258), .A2(n5328), .ZN(n5329) );
  NAND2_X1 U6021 ( .A1(n6865), .A2(n5329), .ZN(n7120) );
  INV_X1 U6022 ( .A(n7120), .ZN(n5330) );
  AOI22_X1 U6023 ( .A1(n6868), .A2(n5330), .B1(EBX_REG_6__SCAN_IN), .B2(n6475), 
        .ZN(n5331) );
  OAI21_X1 U6024 ( .B1(n5501), .B2(n6478), .A(n5331), .ZN(U2853) );
  INV_X1 U6025 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6761) );
  OAI222_X1 U6026 ( .A1(n6219), .A2(n5333), .B1(n6311), .B2(n6761), .C1(n7352), 
        .C2(n5332), .ZN(U2889) );
  NOR2_X1 U6027 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7449) );
  INV_X1 U6028 ( .A(n7449), .ZN(n7443) );
  OR3_X1 U6029 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n7443), .ZN(n6309) );
  NAND2_X1 U6030 ( .A1(n7431), .A2(n5334), .ZN(n7444) );
  AOI21_X1 U6031 ( .B1(n5340), .B2(n6305), .A(n7330), .ZN(n5339) );
  NOR2_X1 U6032 ( .A1(n5335), .A2(n6093), .ZN(n5338) );
  AOI211_X1 U6033 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6309), .A(n5336), .B(
        n5967), .ZN(n5337) );
  NAND2_X1 U6034 ( .A1(n6302), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6035 ( .A1(n6103), .A2(n7447), .ZN(n5342) );
  NAND2_X1 U6036 ( .A1(n3779), .A2(n5975), .ZN(n5341) );
  OAI22_X1 U6037 ( .A1(n6305), .A2(n6126), .B1(n6303), .B2(n7652), .ZN(n5343)
         );
  AOI21_X1 U6038 ( .B1(n7647), .B2(n7645), .A(n5343), .ZN(n5344) );
  OAI211_X1 U6039 ( .C1(n6309), .C2(n6732), .A(n5345), .B(n5344), .ZN(U3027)
         );
  NAND2_X1 U6040 ( .A1(n6302), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5348) );
  OAI22_X1 U6041 ( .A1(n6305), .A2(n6108), .B1(n6303), .B2(n7596), .ZN(n5346)
         );
  AOI21_X1 U6042 ( .B1(n7647), .B2(n7592), .A(n5346), .ZN(n5347) );
  OAI211_X1 U6043 ( .C1(n6309), .C2(n6112), .A(n5348), .B(n5347), .ZN(U3026)
         );
  NAND2_X1 U6044 ( .A1(n6302), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5351) );
  OAI22_X1 U6045 ( .A1(n6305), .A2(n6130), .B1(n6303), .B2(n7558), .ZN(n5349)
         );
  AOI21_X1 U6046 ( .B1(n7647), .B2(n7554), .A(n5349), .ZN(n5350) );
  OAI211_X1 U6047 ( .C1(n6309), .C2(n6713), .A(n5351), .B(n5350), .ZN(U3024)
         );
  NAND2_X1 U6048 ( .A1(n6302), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5354) );
  OAI22_X1 U6049 ( .A1(n6305), .A2(n6113), .B1(n6303), .B2(n7538), .ZN(n5352)
         );
  AOI21_X1 U6050 ( .B1(n7647), .B2(n7534), .A(n5352), .ZN(n5353) );
  OAI211_X1 U6051 ( .C1(n6309), .C2(n6117), .A(n5354), .B(n5353), .ZN(U3023)
         );
  NAND2_X1 U6052 ( .A1(n6302), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5357) );
  OAI22_X1 U6053 ( .A1(n6305), .A2(n6694), .B1(n6303), .B2(n7465), .ZN(n5355)
         );
  AOI21_X1 U6054 ( .B1(n7647), .B2(n7454), .A(n5355), .ZN(n5356) );
  OAI211_X1 U6055 ( .C1(n6107), .C2(n6309), .A(n5357), .B(n5356), .ZN(U3020)
         );
  NAND2_X1 U6056 ( .A1(n6302), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5360) );
  OAI22_X1 U6057 ( .A1(n6305), .A2(n6118), .B1(n6303), .B2(n7511), .ZN(n5358)
         );
  AOI21_X1 U6058 ( .B1(n7647), .B2(n7507), .A(n5358), .ZN(n5359) );
  OAI211_X1 U6059 ( .C1(n6309), .C2(n6707), .A(n5360), .B(n5359), .ZN(U3022)
         );
  NAND2_X1 U6060 ( .A1(n6302), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5363) );
  OAI22_X1 U6061 ( .A1(n6305), .A2(n6122), .B1(n6303), .B2(n7488), .ZN(n5361)
         );
  AOI21_X1 U6062 ( .B1(n7647), .B2(n7484), .A(n5361), .ZN(n5362) );
  OAI211_X1 U6063 ( .C1(n6309), .C2(n6701), .A(n5363), .B(n5362), .ZN(U3021)
         );
  INV_X1 U6064 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6065 ( .A1(n5487), .A2(n5364), .ZN(n5369) );
  INV_X1 U6066 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U6067 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  NAND2_X1 U6068 ( .A1(n6755), .A2(n3983), .ZN(n5568) );
  OR2_X1 U6069 ( .A1(n7295), .A2(n5370), .ZN(n6955) );
  INV_X2 U6070 ( .A(n6955), .ZN(n7285) );
  NOR2_X4 U6071 ( .A1(n7285), .A2(n6755), .ZN(n6767) );
  AOI22_X1 U6072 ( .A1(n7285), .A2(UWORD_REG_9__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5371) );
  OAI21_X1 U6073 ( .B1(n5372), .B2(n5568), .A(n5371), .ZN(U2898) );
  INV_X1 U6074 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5374) );
  AOI22_X1 U6075 ( .A1(n7285), .A2(UWORD_REG_7__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5373) );
  OAI21_X1 U6076 ( .B1(n5374), .B2(n5568), .A(n5373), .ZN(U2900) );
  INV_X1 U6077 ( .A(EAX_REG_21__SCAN_IN), .ZN(n5376) );
  AOI22_X1 U6078 ( .A1(n7285), .A2(UWORD_REG_5__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5375) );
  OAI21_X1 U6079 ( .B1(n5376), .B2(n5568), .A(n5375), .ZN(U2902) );
  INV_X1 U6080 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5378) );
  AOI22_X1 U6081 ( .A1(n7285), .A2(UWORD_REG_6__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5377) );
  OAI21_X1 U6082 ( .B1(n5378), .B2(n5568), .A(n5377), .ZN(U2901) );
  AOI22_X1 U6083 ( .A1(n7285), .A2(UWORD_REG_8__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5379) );
  OAI21_X1 U6084 ( .B1(n4644), .B2(n5568), .A(n5379), .ZN(U2899) );
  NAND2_X1 U6085 ( .A1(n5380), .A2(n7324), .ZN(n5493) );
  NOR2_X1 U6086 ( .A1(n7445), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5420) );
  AOI21_X1 U6087 ( .B1(n5493), .B2(n5495), .A(n5420), .ZN(n5381) );
  NAND2_X1 U6088 ( .A1(n5163), .A2(n6420), .ZN(n5966) );
  NOR2_X1 U6089 ( .A1(n3662), .A2(n5966), .ZN(n7434) );
  OAI21_X1 U6090 ( .B1(n5381), .B2(n7434), .A(n7305), .ZN(n5384) );
  NAND2_X1 U6091 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7449), .ZN(n7435) );
  NOR2_X1 U6092 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7435), .ZN(n5496)
         );
  INV_X1 U6093 ( .A(n5496), .ZN(n5414) );
  NAND2_X1 U6094 ( .A1(n5382), .A2(n7268), .ZN(n5385) );
  NAND2_X1 U6095 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5385), .ZN(n6098) );
  INV_X1 U6096 ( .A(n6098), .ZN(n5383) );
  AOI211_X2 U6097 ( .C1(n5384), .C2(n5414), .A(n5967), .B(n5383), .ZN(n5500)
         );
  INV_X1 U6098 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5391) );
  INV_X1 U6099 ( .A(n5385), .ZN(n6102) );
  NAND2_X1 U6100 ( .A1(n6102), .A2(n5975), .ZN(n5386) );
  OAI21_X1 U6101 ( .B1(n5387), .B2(n5966), .A(n5386), .ZN(n5494) );
  NOR2_X1 U6102 ( .A1(n5493), .A2(n5518), .ZN(n5389) );
  OAI22_X1 U6103 ( .A1(n5495), .A2(n6122), .B1(n6701), .B2(n5414), .ZN(n5388)
         );
  AOI211_X1 U6104 ( .C1(n6700), .C2(n5494), .A(n5389), .B(n5388), .ZN(n5390)
         );
  OAI21_X1 U6105 ( .B1(n5500), .B2(n5391), .A(n5390), .ZN(U3037) );
  INV_X1 U6106 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5395) );
  NOR2_X1 U6107 ( .A1(n5493), .A2(n5507), .ZN(n5393) );
  OAI22_X1 U6108 ( .A1(n5495), .A2(n6130), .B1(n6713), .B2(n5414), .ZN(n5392)
         );
  AOI211_X1 U6109 ( .C1(n6712), .C2(n5494), .A(n5393), .B(n5392), .ZN(n5394)
         );
  OAI21_X1 U6110 ( .B1(n5500), .B2(n5395), .A(n5394), .ZN(U3040) );
  INV_X1 U6111 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5399) );
  NOR2_X1 U6112 ( .A1(n5493), .A2(n5428), .ZN(n5397) );
  OAI22_X1 U6113 ( .A1(n6117), .A2(n5414), .B1(n6113), .B2(n5495), .ZN(n5396)
         );
  AOI211_X1 U6114 ( .C1(n6066), .C2(n5494), .A(n5397), .B(n5396), .ZN(n5398)
         );
  OAI21_X1 U6115 ( .B1(n5500), .B2(n5399), .A(n5398), .ZN(U3039) );
  INV_X1 U6116 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5403) );
  NOR2_X1 U6117 ( .A1(n5493), .A2(n5503), .ZN(n5401) );
  OAI22_X1 U6118 ( .A1(n5495), .A2(n6118), .B1(n6707), .B2(n5414), .ZN(n5400)
         );
  AOI211_X1 U6119 ( .C1(n6706), .C2(n5494), .A(n5401), .B(n5400), .ZN(n5402)
         );
  OAI21_X1 U6120 ( .B1(n5500), .B2(n5403), .A(n5402), .ZN(U3038) );
  INV_X1 U6121 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5409) );
  NOR2_X1 U6122 ( .A1(n5404), .A2(n5419), .ZN(n6718) );
  AND2_X1 U6123 ( .A1(n6937), .A2(DATAI_21_), .ZN(n7574) );
  INV_X1 U6124 ( .A(n7574), .ZN(n6297) );
  NOR2_X1 U6125 ( .A1(n5493), .A2(n6297), .ZN(n5407) );
  NAND2_X1 U6126 ( .A1(n6937), .A2(DATAI_29_), .ZN(n6304) );
  NAND2_X1 U6127 ( .A1(n5405), .A2(n4018), .ZN(n6719) );
  OAI22_X1 U6128 ( .A1(n5495), .A2(n6304), .B1(n6719), .B2(n5414), .ZN(n5406)
         );
  AOI211_X1 U6129 ( .C1(n6718), .C2(n5494), .A(n5407), .B(n5406), .ZN(n5408)
         );
  OAI21_X1 U6130 ( .B1(n5500), .B2(n5409), .A(n5408), .ZN(U3041) );
  INV_X1 U6131 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5413) );
  INV_X1 U6132 ( .A(n7596), .ZN(n6724) );
  NOR2_X1 U6133 ( .A1(n5493), .A2(n5973), .ZN(n5411) );
  OAI22_X1 U6134 ( .A1(n6112), .A2(n5414), .B1(n5495), .B2(n6108), .ZN(n5410)
         );
  AOI211_X1 U6135 ( .C1(n6724), .C2(n5494), .A(n5411), .B(n5410), .ZN(n5412)
         );
  OAI21_X1 U6136 ( .B1(n5500), .B2(n5413), .A(n5412), .ZN(U3042) );
  INV_X1 U6137 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5418) );
  NOR2_X1 U6138 ( .A1(n5493), .A2(n5522), .ZN(n5416) );
  OAI22_X1 U6139 ( .A1(n5495), .A2(n6126), .B1(n6732), .B2(n5414), .ZN(n5415)
         );
  AOI211_X1 U6140 ( .C1(n6731), .C2(n5494), .A(n5416), .B(n5415), .ZN(n5417)
         );
  OAI21_X1 U6141 ( .B1(n5500), .B2(n5418), .A(n5417), .ZN(U3043) );
  AND2_X1 U6142 ( .A1(n3662), .A2(n3739), .ZN(n7395) );
  AOI21_X1 U6143 ( .B1(n7395), .B2(n7409), .A(n5426), .ZN(n5425) );
  INV_X1 U6144 ( .A(n5420), .ZN(n7405) );
  OAI21_X1 U6145 ( .B1(n5421), .B2(n6914), .A(n7405), .ZN(n5422) );
  AOI22_X1 U6146 ( .A1(n5425), .A2(n5422), .B1(n5424), .B2(n7445), .ZN(n5423)
         );
  NAND2_X1 U6147 ( .A1(n7459), .A2(n5423), .ZN(n6268) );
  INV_X1 U6148 ( .A(n6268), .ZN(n5433) );
  INV_X1 U6149 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5432) );
  OAI22_X1 U6150 ( .A1(n5425), .A2(n7445), .B1(n5424), .B2(n7295), .ZN(n6270)
         );
  AOI22_X1 U6151 ( .A1(n5426), .A2(n7533), .B1(n6066), .B2(n6270), .ZN(n5427)
         );
  OAI21_X1 U6152 ( .B1(n6305), .B2(n5428), .A(n5427), .ZN(n5429) );
  AOI21_X1 U6153 ( .B1(n7535), .B2(n5430), .A(n5429), .ZN(n5431) );
  OAI21_X1 U6154 ( .B1(n5433), .B2(n5432), .A(n5431), .ZN(U3143) );
  NAND2_X1 U6155 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  XNOR2_X1 U6156 ( .A(n5434), .B(n5437), .ZN(n6907) );
  INV_X1 U6157 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5438) );
  OAI22_X1 U6158 ( .A1(n7029), .A2(n7120), .B1(n7105), .B2(n5438), .ZN(n5446)
         );
  INV_X1 U6160 ( .A(n5439), .ZN(n5440) );
  OAI33_X1 U6161 ( .A1(1'b0), .A2(n5443), .A3(n5442), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n5441), .B3(n5440), .ZN(n5445) );
  AOI211_X1 U6162 ( .C1(n7066), .C2(n6907), .A(n5446), .B(n5445), .ZN(n5447)
         );
  INV_X1 U6163 ( .A(n5447), .ZN(U3012) );
  NAND2_X1 U6164 ( .A1(n5475), .A2(DATAI_10_), .ZN(n5478) );
  AOI22_X1 U6165 ( .A1(n5487), .A2(EAX_REG_10__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6166 ( .A1(n5478), .A2(n5449), .ZN(U2949) );
  NAND2_X1 U6167 ( .A1(n5475), .A2(DATAI_1_), .ZN(n5459) );
  AOI22_X1 U6168 ( .A1(n5487), .A2(EAX_REG_17__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6169 ( .A1(n5459), .A2(n5450), .ZN(U2925) );
  NAND2_X1 U6170 ( .A1(n5475), .A2(DATAI_0_), .ZN(n5461) );
  AOI22_X1 U6171 ( .A1(n5487), .A2(EAX_REG_16__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6172 ( .A1(n5461), .A2(n5451), .ZN(U2924) );
  AOI22_X1 U6173 ( .A1(n5487), .A2(EAX_REG_4__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6174 ( .A1(n5453), .A2(n5452), .ZN(U2943) );
  AOI22_X1 U6175 ( .A1(n5487), .A2(EAX_REG_3__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6176 ( .A1(n5455), .A2(n5454), .ZN(U2942) );
  AOI22_X1 U6177 ( .A1(n5487), .A2(EAX_REG_2__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6178 ( .A1(n5457), .A2(n5456), .ZN(U2941) );
  AOI22_X1 U6179 ( .A1(n5487), .A2(EAX_REG_1__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6180 ( .A1(n5459), .A2(n5458), .ZN(U2940) );
  AOI22_X1 U6181 ( .A1(n5487), .A2(EAX_REG_0__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6182 ( .A1(n5461), .A2(n5460), .ZN(U2939) );
  NAND2_X1 U6183 ( .A1(n5475), .A2(DATAI_14_), .ZN(n5469) );
  AOI22_X1 U6184 ( .A1(n5487), .A2(EAX_REG_30__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6185 ( .A1(n5469), .A2(n5462), .ZN(U2938) );
  INV_X1 U6186 ( .A(DATAI_13_), .ZN(n6185) );
  OR2_X1 U6187 ( .A1(n5492), .A2(n6185), .ZN(n5471) );
  AOI22_X1 U6188 ( .A1(n5487), .A2(EAX_REG_29__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6189 ( .A1(n5471), .A2(n5463), .ZN(U2937) );
  AOI22_X1 U6190 ( .A1(n5487), .A2(EAX_REG_7__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6191 ( .A1(n5465), .A2(n5464), .ZN(U2946) );
  AOI22_X1 U6192 ( .A1(n5487), .A2(EAX_REG_6__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6193 ( .A1(n5467), .A2(n5466), .ZN(U2945) );
  AOI22_X1 U6194 ( .A1(n5487), .A2(EAX_REG_14__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6195 ( .A1(n5469), .A2(n5468), .ZN(U2953) );
  AOI22_X1 U6196 ( .A1(n5487), .A2(EAX_REG_13__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6197 ( .A1(n5471), .A2(n5470), .ZN(U2952) );
  NAND2_X1 U6198 ( .A1(n5475), .A2(DATAI_12_), .ZN(n5489) );
  AOI22_X1 U6199 ( .A1(n5487), .A2(EAX_REG_12__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6200 ( .A1(n5489), .A2(n5472), .ZN(U2951) );
  INV_X1 U6201 ( .A(DATAI_11_), .ZN(n6043) );
  OR2_X1 U6202 ( .A1(n5492), .A2(n6043), .ZN(n5484) );
  AOI22_X1 U6203 ( .A1(n5487), .A2(EAX_REG_11__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6204 ( .A1(n5484), .A2(n5473), .ZN(U2950) );
  NAND2_X1 U6205 ( .A1(n5475), .A2(DATAI_9_), .ZN(n5480) );
  AOI22_X1 U6206 ( .A1(n5487), .A2(EAX_REG_9__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6207 ( .A1(n5480), .A2(n5474), .ZN(U2948) );
  NAND2_X1 U6208 ( .A1(n5475), .A2(DATAI_8_), .ZN(n5486) );
  AOI22_X1 U6209 ( .A1(n5487), .A2(EAX_REG_8__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6210 ( .A1(n5486), .A2(n5476), .ZN(U2947) );
  AOI22_X1 U6211 ( .A1(n5487), .A2(EAX_REG_26__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6212 ( .A1(n5478), .A2(n5477), .ZN(U2934) );
  AOI22_X1 U6213 ( .A1(n5487), .A2(EAX_REG_25__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6214 ( .A1(n5480), .A2(n5479), .ZN(U2933) );
  AOI22_X1 U6215 ( .A1(n5487), .A2(EAX_REG_5__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U6216 ( .A1(n5482), .A2(n5481), .ZN(U2944) );
  AOI22_X1 U6217 ( .A1(n5487), .A2(EAX_REG_27__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U6218 ( .A1(n5484), .A2(n5483), .ZN(U2935) );
  AOI22_X1 U6219 ( .A1(n5487), .A2(EAX_REG_24__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U6220 ( .A1(n5486), .A2(n5485), .ZN(U2932) );
  AOI22_X1 U6221 ( .A1(n5487), .A2(EAX_REG_28__SCAN_IN), .B1(n5490), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6222 ( .A1(n5489), .A2(n5488), .ZN(U2936) );
  INV_X1 U6223 ( .A(DATAI_15_), .ZN(n6220) );
  AOI22_X1 U6224 ( .A1(n5487), .A2(EAX_REG_15__SCAN_IN), .B1(n5490), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n5491) );
  OAI21_X1 U6225 ( .B1(n5492), .B2(n6220), .A(n5491), .ZN(U2954) );
  INV_X1 U6226 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5499) );
  AOI22_X1 U6227 ( .A1(n7638), .A2(n7454), .B1(n6693), .B2(n5494), .ZN(n5498)
         );
  AOI22_X1 U6228 ( .A1(n7646), .A2(n7462), .B1(n7453), .B2(n5496), .ZN(n5497)
         );
  OAI211_X1 U6229 ( .C1(n5500), .C2(n5499), .A(n5498), .B(n5497), .ZN(U3036)
         );
  INV_X1 U6230 ( .A(DATAI_6_), .ZN(n5502) );
  OAI222_X1 U6231 ( .A1(n5502), .A2(n6219), .B1(n6311), .B2(n4345), .C1(n7352), 
        .C2(n5501), .ZN(U2885) );
  NAND2_X1 U6232 ( .A1(n6268), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5506)
         );
  OAI22_X1 U6233 ( .A1(n6276), .A2(n6118), .B1(n5503), .B2(n6305), .ZN(n5504)
         );
  AOI21_X1 U6234 ( .B1(n6706), .B2(n6270), .A(n5504), .ZN(n5505) );
  OAI211_X1 U6235 ( .C1(n6273), .C2(n6707), .A(n5506), .B(n5505), .ZN(U3142)
         );
  NAND2_X1 U6236 ( .A1(n6268), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5510)
         );
  OAI22_X1 U6237 ( .A1(n6276), .A2(n6130), .B1(n5507), .B2(n6305), .ZN(n5508)
         );
  AOI21_X1 U6238 ( .B1(n6712), .B2(n6270), .A(n5508), .ZN(n5509) );
  OAI211_X1 U6239 ( .C1(n6273), .C2(n6713), .A(n5510), .B(n5509), .ZN(U3144)
         );
  NAND2_X1 U6240 ( .A1(n6268), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5514)
         );
  OAI22_X1 U6241 ( .A1(n6276), .A2(n6694), .B1(n5511), .B2(n6305), .ZN(n5512)
         );
  AOI21_X1 U6242 ( .B1(n6693), .B2(n6270), .A(n5512), .ZN(n5513) );
  OAI211_X1 U6243 ( .C1(n6107), .C2(n6273), .A(n5514), .B(n5513), .ZN(U3140)
         );
  NAND2_X1 U6244 ( .A1(n6268), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5517)
         );
  OAI22_X1 U6245 ( .A1(n6276), .A2(n6108), .B1(n5973), .B2(n6305), .ZN(n5515)
         );
  AOI21_X1 U6246 ( .B1(n6724), .B2(n6270), .A(n5515), .ZN(n5516) );
  OAI211_X1 U6247 ( .C1(n6273), .C2(n6112), .A(n5517), .B(n5516), .ZN(U3146)
         );
  NAND2_X1 U6248 ( .A1(n6268), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5521)
         );
  OAI22_X1 U6249 ( .A1(n6276), .A2(n6122), .B1(n5518), .B2(n6305), .ZN(n5519)
         );
  AOI21_X1 U6250 ( .B1(n6700), .B2(n6270), .A(n5519), .ZN(n5520) );
  OAI211_X1 U6251 ( .C1(n6273), .C2(n6701), .A(n5521), .B(n5520), .ZN(U3141)
         );
  NAND2_X1 U6252 ( .A1(n6268), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5525)
         );
  OAI22_X1 U6253 ( .A1(n6276), .A2(n6126), .B1(n5522), .B2(n6305), .ZN(n5523)
         );
  AOI21_X1 U6254 ( .B1(n6731), .B2(n6270), .A(n5523), .ZN(n5524) );
  OAI211_X1 U6255 ( .C1(n6273), .C2(n6732), .A(n5525), .B(n5524), .ZN(U3147)
         );
  INV_X1 U6256 ( .A(n5526), .ZN(n5530) );
  INV_X1 U6257 ( .A(n5527), .ZN(n5529) );
  AOI21_X1 U6258 ( .B1(n5530), .B2(n5529), .A(n5528), .ZN(n5549) );
  INV_X1 U6259 ( .A(n5549), .ZN(n5993) );
  INV_X1 U6260 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5532) );
  XNOR2_X1 U6261 ( .A(n6867), .B(n5531), .ZN(n5987) );
  OAI222_X1 U6262 ( .A1(n6468), .A2(n5993), .B1(n5532), .B2(n6880), .C1(n6876), 
        .C2(n5987), .ZN(U2851) );
  OR2_X1 U6263 ( .A1(n5255), .A2(n5533), .ZN(n5534) );
  AND2_X1 U6264 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  OR2_X1 U6265 ( .A1(n5536), .A2(n5527), .ZN(n6915) );
  OAI222_X1 U6266 ( .A1(n5537), .A2(n6219), .B1(n6311), .B2(n4337), .C1(n7352), 
        .C2(n6915), .ZN(U2884) );
  OAI21_X1 U6267 ( .B1(n5528), .B2(n5539), .A(n5538), .ZN(n5997) );
  INV_X1 U6268 ( .A(n6023), .ZN(n5540) );
  AOI21_X1 U6269 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n7037) );
  AOI22_X1 U6270 ( .A1(n6868), .A2(n7037), .B1(EBX_REG_9__SCAN_IN), .B2(n6475), 
        .ZN(n5543) );
  OAI21_X1 U6271 ( .B1(n5997), .B2(n6478), .A(n5543), .ZN(U2850) );
  OAI21_X1 U6272 ( .B1(n5546), .B2(n5545), .A(n5544), .ZN(n7008) );
  NAND2_X1 U6273 ( .A1(n7059), .A2(REIP_REG_8__SCAN_IN), .ZN(n7005) );
  NAND2_X1 U6274 ( .A1(n6932), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5547)
         );
  OAI211_X1 U6275 ( .C1(n6940), .C2(n5983), .A(n7005), .B(n5547), .ZN(n5548)
         );
  AOI21_X1 U6276 ( .B1(n5549), .B2(n6937), .A(n5548), .ZN(n5550) );
  OAI21_X1 U6277 ( .B1(n7008), .B2(n7241), .A(n5550), .ZN(U2978) );
  INV_X1 U6278 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5552) );
  AOI22_X1 U6279 ( .A1(n7285), .A2(UWORD_REG_14__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5551) );
  OAI21_X1 U6280 ( .B1(n5552), .B2(n5568), .A(n5551), .ZN(U2893) );
  INV_X1 U6281 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5554) );
  AOI22_X1 U6282 ( .A1(n7285), .A2(UWORD_REG_11__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5553) );
  OAI21_X1 U6283 ( .B1(n5554), .B2(n5568), .A(n5553), .ZN(U2896) );
  INV_X1 U6284 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5556) );
  AOI22_X1 U6285 ( .A1(n7285), .A2(UWORD_REG_10__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5555) );
  OAI21_X1 U6286 ( .B1(n5556), .B2(n5568), .A(n5555), .ZN(U2897) );
  INV_X1 U6287 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5558) );
  AOI22_X1 U6288 ( .A1(n7285), .A2(UWORD_REG_4__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5557) );
  OAI21_X1 U6289 ( .B1(n5558), .B2(n5568), .A(n5557), .ZN(U2903) );
  AOI22_X1 U6290 ( .A1(n7285), .A2(UWORD_REG_3__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5559) );
  OAI21_X1 U6291 ( .B1(n4544), .B2(n5568), .A(n5559), .ZN(U2904) );
  INV_X1 U6292 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5561) );
  AOI22_X1 U6293 ( .A1(n7285), .A2(UWORD_REG_1__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5560) );
  OAI21_X1 U6294 ( .B1(n5561), .B2(n5568), .A(n5560), .ZN(U2906) );
  INV_X1 U6295 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5563) );
  AOI22_X1 U6296 ( .A1(n7285), .A2(UWORD_REG_0__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5562) );
  OAI21_X1 U6297 ( .B1(n5563), .B2(n5568), .A(n5562), .ZN(U2907) );
  AOI22_X1 U6298 ( .A1(n7285), .A2(UWORD_REG_13__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5564) );
  OAI21_X1 U6299 ( .B1(n4750), .B2(n5568), .A(n5564), .ZN(U2894) );
  INV_X1 U6300 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5566) );
  AOI22_X1 U6301 ( .A1(n7285), .A2(UWORD_REG_12__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5565) );
  OAI21_X1 U6302 ( .B1(n5566), .B2(n5568), .A(n5565), .ZN(U2895) );
  INV_X1 U6303 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5569) );
  AOI22_X1 U6304 ( .A1(n7285), .A2(UWORD_REG_2__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5567) );
  OAI21_X1 U6305 ( .B1(n5569), .B2(n5568), .A(n5567), .ZN(U2905) );
  INV_X1 U6306 ( .A(DATAI_8_), .ZN(n5570) );
  INV_X1 U6307 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6771) );
  OAI222_X1 U6308 ( .A1(n5570), .A2(n6219), .B1(n6311), .B2(n6771), .C1(n7352), 
        .C2(n5993), .ZN(U2883) );
  OR2_X1 U6309 ( .A1(n6953), .A2(n5571), .ZN(n5572) );
  NAND2_X1 U6310 ( .A1(n5572), .A2(n7196), .ZN(n7112) );
  NOR2_X1 U6311 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5573), .ZN(n5574) );
  AND2_X1 U6312 ( .A1(n3983), .A2(n5574), .ZN(n5575) );
  NOR2_X1 U6313 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  OAI22_X1 U6314 ( .A1(n5139), .A2(n7203), .B1(n7195), .B2(n5578), .ZN(n5579)
         );
  AOI21_X1 U6315 ( .B1(n5586), .B2(REIP_REG_0__SCAN_IN), .A(n5579), .ZN(n5585)
         );
  OR2_X1 U6316 ( .A1(n6953), .A2(n5580), .ZN(n7094) );
  INV_X1 U6317 ( .A(n7094), .ZN(n7074) );
  INV_X1 U6318 ( .A(n5581), .ZN(n5582) );
  NAND2_X1 U6319 ( .A1(n7215), .A2(n7239), .ZN(n5583) );
  AOI22_X1 U6320 ( .A1(n7074), .A2(n3739), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5583), .ZN(n5584) );
  OAI211_X1 U6321 ( .C1(n7097), .C2(n6881), .A(n5585), .B(n5584), .ZN(U2827)
         );
  OAI21_X1 U6322 ( .B1(n6421), .B2(n6030), .A(n5586), .ZN(n6027) );
  INV_X1 U6323 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6797) );
  AOI22_X1 U6324 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n7228), .B1(
        EBX_REG_9__SCAN_IN), .B2(n7227), .ZN(n5587) );
  OAI21_X1 U6325 ( .B1(n6027), .B2(n6797), .A(n5587), .ZN(n5592) );
  NOR3_X1 U6326 ( .A1(n7192), .A2(n6030), .A3(REIP_REG_9__SCAN_IN), .ZN(n5591)
         );
  INV_X1 U6327 ( .A(n5588), .ZN(n5999) );
  NAND2_X1 U6328 ( .A1(n7235), .A2(n7037), .ZN(n5589) );
  OAI211_X1 U6329 ( .C1(n7239), .C2(n5999), .A(n5589), .B(n7105), .ZN(n5590)
         );
  NOR3_X1 U6330 ( .A1(n5592), .A2(n5591), .A3(n5590), .ZN(n5593) );
  OAI21_X1 U6331 ( .B1(n5997), .B2(n7196), .A(n5593), .ZN(U2818) );
  INV_X1 U6332 ( .A(DATAI_9_), .ZN(n5594) );
  INV_X1 U6333 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6773) );
  OAI222_X1 U6334 ( .A1(n5594), .A2(n6219), .B1(n6311), .B2(n6773), .C1(n7352), 
        .C2(n5997), .ZN(U2882) );
  XOR2_X1 U6335 ( .A(DATAI_31_), .B(keyinput_128), .Z(n5598) );
  XOR2_X1 U6336 ( .A(DATAI_30_), .B(keyinput_129), .Z(n5597) );
  XNOR2_X1 U6337 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n5596) );
  XOR2_X1 U6338 ( .A(DATAI_29_), .B(keyinput_130), .Z(n5595) );
  AOI211_X1 U6339 ( .C1(n5598), .C2(n5597), .A(n5596), .B(n5595), .ZN(n5604)
         );
  XOR2_X1 U6340 ( .A(DATAI_27_), .B(keyinput_132), .Z(n5603) );
  XOR2_X1 U6341 ( .A(DATAI_25_), .B(keyinput_134), .Z(n5601) );
  XOR2_X1 U6342 ( .A(DATAI_26_), .B(keyinput_133), .Z(n5600) );
  XNOR2_X1 U6343 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n5599) );
  NOR3_X1 U6344 ( .A1(n5601), .A2(n5600), .A3(n5599), .ZN(n5602) );
  OAI21_X1 U6345 ( .B1(n5604), .B2(n5603), .A(n5602), .ZN(n5607) );
  XOR2_X1 U6346 ( .A(DATAI_23_), .B(keyinput_136), .Z(n5606) );
  XNOR2_X1 U6347 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n5605) );
  AOI21_X1 U6348 ( .B1(n5607), .B2(n5606), .A(n5605), .ZN(n5610) );
  XOR2_X1 U6349 ( .A(DATAI_21_), .B(keyinput_138), .Z(n5609) );
  XNOR2_X1 U6350 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n5608) );
  OAI21_X1 U6351 ( .B1(n5610), .B2(n5609), .A(n5608), .ZN(n5614) );
  XOR2_X1 U6352 ( .A(keyinput_140), .B(DATAI_19_), .Z(n5613) );
  XNOR2_X1 U6353 ( .A(keyinput_142), .B(DATAI_17_), .ZN(n5612) );
  XNOR2_X1 U6354 ( .A(keyinput_141), .B(DATAI_18_), .ZN(n5611) );
  NAND4_X1 U6355 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .ZN(n5617)
         );
  XNOR2_X1 U6356 ( .A(keyinput_143), .B(DATAI_16_), .ZN(n5616) );
  XOR2_X1 U6357 ( .A(keyinput_144), .B(DATAI_15_), .Z(n5615) );
  AOI21_X1 U6358 ( .B1(n5617), .B2(n5616), .A(n5615), .ZN(n5623) );
  XOR2_X1 U6359 ( .A(DATAI_14_), .B(keyinput_145), .Z(n5622) );
  XNOR2_X1 U6360 ( .A(DATAI_12_), .B(keyinput_147), .ZN(n5620) );
  XNOR2_X1 U6361 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n5619) );
  XNOR2_X1 U6362 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n5618) );
  NOR3_X1 U6363 ( .A1(n5620), .A2(n5619), .A3(n5618), .ZN(n5621) );
  OAI21_X1 U6364 ( .B1(n5623), .B2(n5622), .A(n5621), .ZN(n5626) );
  XOR2_X1 U6365 ( .A(keyinput_150), .B(DATAI_9_), .Z(n5625) );
  XNOR2_X1 U6366 ( .A(keyinput_149), .B(DATAI_10_), .ZN(n5624) );
  NAND3_X1 U6367 ( .A1(n5626), .A2(n5625), .A3(n5624), .ZN(n5633) );
  XOR2_X1 U6368 ( .A(keyinput_151), .B(DATAI_8_), .Z(n5632) );
  XOR2_X1 U6369 ( .A(keyinput_154), .B(DATAI_5_), .Z(n5630) );
  XOR2_X1 U6370 ( .A(keyinput_152), .B(DATAI_7_), .Z(n5629) );
  XOR2_X1 U6371 ( .A(keyinput_153), .B(DATAI_6_), .Z(n5628) );
  XNOR2_X1 U6372 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n5627) );
  NAND4_X1 U6373 ( .A1(n5630), .A2(n5629), .A3(n5628), .A4(n5627), .ZN(n5631)
         );
  AOI21_X1 U6374 ( .B1(n5633), .B2(n5632), .A(n5631), .ZN(n5636) );
  XOR2_X1 U6375 ( .A(keyinput_156), .B(DATAI_3_), .Z(n5635) );
  XNOR2_X1 U6376 ( .A(keyinput_157), .B(DATAI_2_), .ZN(n5634) );
  NOR3_X1 U6377 ( .A1(n5636), .A2(n5635), .A3(n5634), .ZN(n5639) );
  XNOR2_X1 U6378 ( .A(keyinput_158), .B(DATAI_1_), .ZN(n5638) );
  XNOR2_X1 U6379 ( .A(keyinput_159), .B(DATAI_0_), .ZN(n5637) );
  NOR3_X1 U6380 ( .A1(n5639), .A2(n5638), .A3(n5637), .ZN(n5645) );
  XOR2_X1 U6381 ( .A(keyinput_160), .B(MEMORYFETCH_REG_SCAN_IN), .Z(n5644) );
  INV_X1 U6382 ( .A(BS16_N), .ZN(n6738) );
  XNOR2_X1 U6383 ( .A(n6738), .B(keyinput_162), .ZN(n5642) );
  XNOR2_X1 U6384 ( .A(READY_N), .B(keyinput_163), .ZN(n5641) );
  XNOR2_X1 U6385 ( .A(keyinput_161), .B(NA_N), .ZN(n5640) );
  NOR3_X1 U6386 ( .A1(n5642), .A2(n5641), .A3(n5640), .ZN(n5643) );
  OAI21_X1 U6387 ( .B1(n5645), .B2(n5644), .A(n5643), .ZN(n5649) );
  XNOR2_X1 U6388 ( .A(keyinput_164), .B(HOLD), .ZN(n5648) );
  INV_X1 U6389 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6753) );
  XNOR2_X1 U6390 ( .A(n6753), .B(keyinput_166), .ZN(n5647) );
  XNOR2_X1 U6391 ( .A(keyinput_165), .B(READREQUEST_REG_SCAN_IN), .ZN(n5646)
         );
  AOI211_X1 U6392 ( .C1(n5649), .C2(n5648), .A(n5647), .B(n5646), .ZN(n5652)
         );
  INV_X1 U6393 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7351) );
  XNOR2_X1 U6394 ( .A(n7351), .B(keyinput_168), .ZN(n5651) );
  XNOR2_X1 U6395 ( .A(keyinput_167), .B(CODEFETCH_REG_SCAN_IN), .ZN(n5650) );
  NOR3_X1 U6396 ( .A1(n5652), .A2(n5651), .A3(n5650), .ZN(n5655) );
  XOR2_X1 U6397 ( .A(keyinput_170), .B(REQUESTPENDING_REG_SCAN_IN), .Z(n5654)
         );
  XNOR2_X1 U6398 ( .A(keyinput_169), .B(D_C_N_REG_SCAN_IN), .ZN(n5653) );
  NOR3_X1 U6399 ( .A1(n5655), .A2(n5654), .A3(n5653), .ZN(n5663) );
  XNOR2_X1 U6400 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_171), .ZN(n5662) );
  XNOR2_X1 U6401 ( .A(keyinput_173), .B(FLUSH_REG_SCAN_IN), .ZN(n5661) );
  XOR2_X1 U6402 ( .A(keyinput_176), .B(BYTEENABLE_REG_1__SCAN_IN), .Z(n5659)
         );
  XOR2_X1 U6403 ( .A(keyinput_175), .B(BYTEENABLE_REG_0__SCAN_IN), .Z(n5658)
         );
  INV_X1 U6404 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6946) );
  XNOR2_X1 U6405 ( .A(n6946), .B(keyinput_174), .ZN(n5657) );
  XNOR2_X1 U6406 ( .A(keyinput_172), .B(MORE_REG_SCAN_IN), .ZN(n5656) );
  NAND4_X1 U6407 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n5660)
         );
  NOR4_X1 U6408 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n5666)
         );
  XNOR2_X1 U6409 ( .A(keyinput_178), .B(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5665)
         );
  XNOR2_X1 U6410 ( .A(keyinput_177), .B(BYTEENABLE_REG_2__SCAN_IN), .ZN(n5664)
         );
  NOR3_X1 U6411 ( .A1(n5666), .A2(n5665), .A3(n5664), .ZN(n5669) );
  XNOR2_X1 U6412 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_179), .ZN(n5668) );
  XNOR2_X1 U6413 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_180), .ZN(n5667) );
  OAI21_X1 U6414 ( .B1(n5669), .B2(n5668), .A(n5667), .ZN(n5675) );
  OAI22_X1 U6415 ( .A1(n7232), .A2(keyinput_185), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_183), .ZN(n5670) );
  AOI221_X1 U6416 ( .B1(n7232), .B2(keyinput_185), .C1(keyinput_183), .C2(
        REIP_REG_27__SCAN_IN), .A(n5670), .ZN(n5674) );
  XOR2_X1 U6417 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_184), .Z(n5673) );
  INV_X1 U6418 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6829) );
  OAI22_X1 U6419 ( .A1(n6829), .A2(keyinput_182), .B1(REIP_REG_29__SCAN_IN), 
        .B2(keyinput_181), .ZN(n5671) );
  AOI221_X1 U6420 ( .B1(n6829), .B2(keyinput_182), .C1(keyinput_181), .C2(
        REIP_REG_29__SCAN_IN), .A(n5671), .ZN(n5672) );
  NAND4_X1 U6421 ( .A1(n5675), .A2(n5674), .A3(n5673), .A4(n5672), .ZN(n5678)
         );
  XOR2_X1 U6422 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_186), .Z(n5677) );
  INV_X1 U6423 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6527) );
  XNOR2_X1 U6424 ( .A(n6527), .B(keyinput_187), .ZN(n5676) );
  NAND3_X1 U6425 ( .A1(n5678), .A2(n5677), .A3(n5676), .ZN(n5681) );
  XOR2_X1 U6426 ( .A(keyinput_189), .B(REIP_REG_21__SCAN_IN), .Z(n5680) );
  XNOR2_X1 U6427 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_188), .ZN(n5679) );
  NAND3_X1 U6428 ( .A1(n5681), .A2(n5680), .A3(n5679), .ZN(n5686) );
  INV_X1 U6429 ( .A(keyinput_191), .ZN(n5682) );
  XNOR2_X1 U6430 ( .A(n5682), .B(REIP_REG_19__SCAN_IN), .ZN(n5685) );
  XNOR2_X1 U6431 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_192), .ZN(n5684) );
  XNOR2_X1 U6432 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_190), .ZN(n5683) );
  NAND4_X1 U6433 ( .A1(n5686), .A2(n5685), .A3(n5684), .A4(n5683), .ZN(n5689)
         );
  XOR2_X1 U6434 ( .A(keyinput_193), .B(REIP_REG_17__SCAN_IN), .Z(n5688) );
  XNOR2_X1 U6435 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_194), .ZN(n5687) );
  AOI21_X1 U6436 ( .B1(n5689), .B2(n5688), .A(n5687), .ZN(n5693) );
  INV_X1 U6437 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6838) );
  XNOR2_X1 U6438 ( .A(n6838), .B(keyinput_195), .ZN(n5692) );
  XNOR2_X1 U6439 ( .A(keyinput_196), .B(BE_N_REG_2__SCAN_IN), .ZN(n5691) );
  XNOR2_X1 U6440 ( .A(keyinput_197), .B(BE_N_REG_1__SCAN_IN), .ZN(n5690) );
  OAI211_X1 U6441 ( .C1(n5693), .C2(n5692), .A(n5691), .B(n5690), .ZN(n5696)
         );
  XNOR2_X1 U6442 ( .A(keyinput_198), .B(BE_N_REG_0__SCAN_IN), .ZN(n5695) );
  XNOR2_X1 U6443 ( .A(keyinput_199), .B(ADDRESS_REG_29__SCAN_IN), .ZN(n5694)
         );
  AOI21_X1 U6444 ( .B1(n5696), .B2(n5695), .A(n5694), .ZN(n5699) );
  INV_X1 U6445 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6832) );
  XNOR2_X1 U6446 ( .A(n6832), .B(keyinput_200), .ZN(n5698) );
  INV_X1 U6447 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6830) );
  XNOR2_X1 U6448 ( .A(n6830), .B(keyinput_201), .ZN(n5697) );
  OAI21_X1 U6449 ( .B1(n5699), .B2(n5698), .A(n5697), .ZN(n5703) );
  XNOR2_X1 U6450 ( .A(keyinput_202), .B(ADDRESS_REG_26__SCAN_IN), .ZN(n5702)
         );
  INV_X1 U6451 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6823) );
  XNOR2_X1 U6452 ( .A(n6823), .B(keyinput_203), .ZN(n5701) );
  XNOR2_X1 U6453 ( .A(keyinput_204), .B(ADDRESS_REG_24__SCAN_IN), .ZN(n5700)
         );
  AOI211_X1 U6454 ( .C1(n5703), .C2(n5702), .A(n5701), .B(n5700), .ZN(n5706)
         );
  INV_X1 U6455 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6821) );
  XNOR2_X1 U6456 ( .A(n6821), .B(keyinput_205), .ZN(n5705) );
  XNOR2_X1 U6457 ( .A(keyinput_206), .B(ADDRESS_REG_22__SCAN_IN), .ZN(n5704)
         );
  NOR3_X1 U6458 ( .A1(n5706), .A2(n5705), .A3(n5704), .ZN(n5709) );
  XNOR2_X1 U6459 ( .A(keyinput_207), .B(ADDRESS_REG_21__SCAN_IN), .ZN(n5708)
         );
  INV_X1 U6460 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6817) );
  XNOR2_X1 U6461 ( .A(n6817), .B(keyinput_208), .ZN(n5707) );
  OAI21_X1 U6462 ( .B1(n5709), .B2(n5708), .A(n5707), .ZN(n5712) );
  XNOR2_X1 U6463 ( .A(keyinput_209), .B(ADDRESS_REG_19__SCAN_IN), .ZN(n5711)
         );
  XNOR2_X1 U6464 ( .A(keyinput_210), .B(ADDRESS_REG_18__SCAN_IN), .ZN(n5710)
         );
  AOI21_X1 U6465 ( .B1(n5712), .B2(n5711), .A(n5710), .ZN(n5716) );
  INV_X1 U6466 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6813) );
  XNOR2_X1 U6467 ( .A(n6813), .B(keyinput_211), .ZN(n5715) );
  XNOR2_X1 U6468 ( .A(keyinput_213), .B(ADDRESS_REG_15__SCAN_IN), .ZN(n5714)
         );
  XNOR2_X1 U6469 ( .A(keyinput_212), .B(ADDRESS_REG_16__SCAN_IN), .ZN(n5713)
         );
  OAI211_X1 U6470 ( .C1(n5716), .C2(n5715), .A(n5714), .B(n5713), .ZN(n5719)
         );
  XNOR2_X1 U6471 ( .A(keyinput_214), .B(ADDRESS_REG_14__SCAN_IN), .ZN(n5718)
         );
  XNOR2_X1 U6472 ( .A(keyinput_215), .B(ADDRESS_REG_13__SCAN_IN), .ZN(n5717)
         );
  AOI21_X1 U6473 ( .B1(n5719), .B2(n5718), .A(n5717), .ZN(n5725) );
  INV_X1 U6474 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6805) );
  XNOR2_X1 U6475 ( .A(n6805), .B(keyinput_216), .ZN(n5724) );
  XNOR2_X1 U6476 ( .A(keyinput_217), .B(ADDRESS_REG_11__SCAN_IN), .ZN(n5722)
         );
  XNOR2_X1 U6477 ( .A(keyinput_219), .B(ADDRESS_REG_9__SCAN_IN), .ZN(n5721) );
  XNOR2_X1 U6478 ( .A(keyinput_218), .B(ADDRESS_REG_10__SCAN_IN), .ZN(n5720)
         );
  NOR3_X1 U6479 ( .A1(n5722), .A2(n5721), .A3(n5720), .ZN(n5723) );
  OAI21_X1 U6480 ( .B1(n5725), .B2(n5724), .A(n5723), .ZN(n5728) );
  XNOR2_X1 U6481 ( .A(keyinput_220), .B(ADDRESS_REG_8__SCAN_IN), .ZN(n5727) );
  INV_X1 U6482 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6796) );
  XNOR2_X1 U6483 ( .A(n6796), .B(keyinput_221), .ZN(n5726) );
  AOI21_X1 U6484 ( .B1(n5728), .B2(n5727), .A(n5726), .ZN(n5731) );
  INV_X1 U6485 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6794) );
  XNOR2_X1 U6486 ( .A(n6794), .B(keyinput_222), .ZN(n5730) );
  INV_X1 U6487 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6793) );
  XNOR2_X1 U6488 ( .A(n6793), .B(keyinput_223), .ZN(n5729) );
  OAI21_X1 U6489 ( .B1(n5731), .B2(n5730), .A(n5729), .ZN(n5733) );
  INV_X1 U6490 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6792) );
  XNOR2_X1 U6491 ( .A(n6792), .B(keyinput_224), .ZN(n5732) );
  NAND2_X1 U6492 ( .A1(n5733), .A2(n5732), .ZN(n5739) );
  INV_X1 U6493 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6790) );
  OAI22_X1 U6494 ( .A1(n6790), .A2(keyinput_225), .B1(ADDRESS_REG_0__SCAN_IN), 
        .B2(keyinput_228), .ZN(n5734) );
  AOI221_X1 U6495 ( .B1(n6790), .B2(keyinput_225), .C1(keyinput_228), .C2(
        ADDRESS_REG_0__SCAN_IN), .A(n5734), .ZN(n5738) );
  INV_X1 U6496 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6787) );
  XNOR2_X1 U6497 ( .A(n6787), .B(keyinput_227), .ZN(n5737) );
  OAI22_X1 U6498 ( .A1(STATE_REG_2__SCAN_IN), .A2(keyinput_229), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(keyinput_226), .ZN(n5735) );
  AOI221_X1 U6499 ( .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_229), .C1(
        keyinput_226), .C2(ADDRESS_REG_2__SCAN_IN), .A(n5735), .ZN(n5736) );
  NAND4_X1 U6500 ( .A1(n5739), .A2(n5738), .A3(n5737), .A4(n5736), .ZN(n5743)
         );
  XNOR2_X1 U6501 ( .A(n7334), .B(keyinput_230), .ZN(n5742) );
  XNOR2_X1 U6502 ( .A(n7345), .B(keyinput_231), .ZN(n5741) );
  XNOR2_X1 U6503 ( .A(keyinput_232), .B(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5740)
         );
  AOI211_X1 U6504 ( .C1(n5743), .C2(n5742), .A(n5741), .B(n5740), .ZN(n5746)
         );
  XNOR2_X1 U6505 ( .A(keyinput_233), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5745)
         );
  XOR2_X1 U6506 ( .A(keyinput_234), .B(DATAWIDTH_REG_2__SCAN_IN), .Z(n5744) );
  OAI21_X1 U6507 ( .B1(n5746), .B2(n5745), .A(n5744), .ZN(n5768) );
  INV_X1 U6508 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6742) );
  XNOR2_X1 U6509 ( .A(n6742), .B(keyinput_238), .ZN(n5750) );
  INV_X1 U6510 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6740) );
  XNOR2_X1 U6511 ( .A(n6740), .B(keyinput_235), .ZN(n5749) );
  XNOR2_X1 U6512 ( .A(keyinput_236), .B(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5748)
         );
  XNOR2_X1 U6513 ( .A(keyinput_237), .B(DATAWIDTH_REG_5__SCAN_IN), .ZN(n5747)
         );
  NOR4_X1 U6514 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n5767)
         );
  INV_X1 U6515 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6747) );
  INV_X1 U6516 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6748) );
  AOI22_X1 U6517 ( .A1(keyinput_245), .A2(n6747), .B1(n6748), .B2(keyinput_246), .ZN(n5762) );
  AOI22_X1 U6518 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput_242), .B1(
        DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_240), .ZN(n5761) );
  INV_X1 U6519 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6746) );
  AOI22_X1 U6520 ( .A1(n6746), .A2(keyinput_243), .B1(
        DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput_244), .ZN(n5760) );
  NAND2_X1 U6521 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(keyinput_248), .ZN(
        n5758) );
  NAND2_X1 U6522 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(keyinput_239), .ZN(n5757) );
  OAI22_X1 U6523 ( .A1(n6748), .A2(keyinput_246), .B1(DATAWIDTH_REG_7__SCAN_IN), .B2(keyinput_239), .ZN(n5752) );
  OAI22_X1 U6524 ( .A1(n6746), .A2(keyinput_243), .B1(n6747), .B2(keyinput_245), .ZN(n5751) );
  NOR2_X1 U6525 ( .A1(n5752), .A2(n5751), .ZN(n5756) );
  OAI22_X1 U6526 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput_242), .B1(
        DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_240), .ZN(n5754) );
  OAI22_X1 U6527 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(keyinput_248), .B1(
        DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput_244), .ZN(n5753) );
  NOR2_X1 U6528 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  AND4_X1 U6529 ( .A1(n5758), .A2(n5757), .A3(n5756), .A4(n5755), .ZN(n5759)
         );
  NAND4_X1 U6530 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n5766)
         );
  XNOR2_X1 U6531 ( .A(keyinput_247), .B(DATAWIDTH_REG_15__SCAN_IN), .ZN(n5764)
         );
  XNOR2_X1 U6532 ( .A(keyinput_241), .B(DATAWIDTH_REG_9__SCAN_IN), .ZN(n5763)
         );
  NAND2_X1 U6533 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  AOI211_X1 U6534 ( .C1(n5768), .C2(n5767), .A(n5766), .B(n5765), .ZN(n5778)
         );
  XOR2_X1 U6535 ( .A(keyinput_251), .B(DATAWIDTH_REG_19__SCAN_IN), .Z(n5772)
         );
  XOR2_X1 U6536 ( .A(keyinput_249), .B(DATAWIDTH_REG_17__SCAN_IN), .Z(n5771)
         );
  XOR2_X1 U6537 ( .A(keyinput_250), .B(DATAWIDTH_REG_18__SCAN_IN), .Z(n5770)
         );
  XOR2_X1 U6538 ( .A(keyinput_252), .B(DATAWIDTH_REG_20__SCAN_IN), .Z(n5769)
         );
  NAND4_X1 U6539 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n5777)
         );
  INV_X1 U6540 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6750) );
  XNOR2_X1 U6541 ( .A(n6750), .B(keyinput_255), .ZN(n5775) );
  XNOR2_X1 U6542 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_254), .ZN(n5774)
         );
  XNOR2_X1 U6543 ( .A(keyinput_253), .B(DATAWIDTH_REG_21__SCAN_IN), .ZN(n5773)
         );
  NOR3_X1 U6544 ( .A1(n5775), .A2(n5774), .A3(n5773), .ZN(n5776) );
  OAI21_X1 U6545 ( .B1(n5778), .B2(n5777), .A(n5776), .ZN(n5964) );
  XOR2_X1 U6546 ( .A(DATAI_31_), .B(keyinput_0), .Z(n5782) );
  XOR2_X1 U6547 ( .A(DATAI_30_), .B(keyinput_1), .Z(n5781) );
  XOR2_X1 U6548 ( .A(DATAI_29_), .B(keyinput_2), .Z(n5780) );
  XOR2_X1 U6549 ( .A(DATAI_28_), .B(keyinput_3), .Z(n5779) );
  AOI211_X1 U6550 ( .C1(n5782), .C2(n5781), .A(n5780), .B(n5779), .ZN(n5788)
         );
  XOR2_X1 U6551 ( .A(DATAI_27_), .B(keyinput_4), .Z(n5787) );
  XOR2_X1 U6552 ( .A(DATAI_25_), .B(keyinput_6), .Z(n5785) );
  XOR2_X1 U6553 ( .A(DATAI_26_), .B(keyinput_5), .Z(n5784) );
  XNOR2_X1 U6554 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n5783) );
  NOR3_X1 U6555 ( .A1(n5785), .A2(n5784), .A3(n5783), .ZN(n5786) );
  OAI21_X1 U6556 ( .B1(n5788), .B2(n5787), .A(n5786), .ZN(n5791) );
  XOR2_X1 U6557 ( .A(DATAI_23_), .B(keyinput_8), .Z(n5790) );
  XOR2_X1 U6558 ( .A(DATAI_22_), .B(keyinput_9), .Z(n5789) );
  AOI21_X1 U6559 ( .B1(n5791), .B2(n5790), .A(n5789), .ZN(n5794) );
  XNOR2_X1 U6560 ( .A(DATAI_21_), .B(keyinput_10), .ZN(n5793) );
  XOR2_X1 U6561 ( .A(DATAI_20_), .B(keyinput_11), .Z(n5792) );
  OAI21_X1 U6562 ( .B1(n5794), .B2(n5793), .A(n5792), .ZN(n5798) );
  XNOR2_X1 U6563 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n5797) );
  XNOR2_X1 U6564 ( .A(DATAI_17_), .B(keyinput_14), .ZN(n5796) );
  XNOR2_X1 U6565 ( .A(DATAI_18_), .B(keyinput_13), .ZN(n5795) );
  NAND4_X1 U6566 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n5801)
         );
  XOR2_X1 U6567 ( .A(DATAI_16_), .B(keyinput_15), .Z(n5800) );
  XOR2_X1 U6568 ( .A(DATAI_15_), .B(keyinput_16), .Z(n5799) );
  AOI21_X1 U6569 ( .B1(n5801), .B2(n5800), .A(n5799), .ZN(n5807) );
  XOR2_X1 U6570 ( .A(DATAI_14_), .B(keyinput_17), .Z(n5806) );
  XOR2_X1 U6571 ( .A(DATAI_12_), .B(keyinput_19), .Z(n5804) );
  XNOR2_X1 U6572 ( .A(DATAI_11_), .B(keyinput_20), .ZN(n5803) );
  XNOR2_X1 U6573 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n5802) );
  NOR3_X1 U6574 ( .A1(n5804), .A2(n5803), .A3(n5802), .ZN(n5805) );
  OAI21_X1 U6575 ( .B1(n5807), .B2(n5806), .A(n5805), .ZN(n5810) );
  XNOR2_X1 U6576 ( .A(DATAI_9_), .B(keyinput_22), .ZN(n5809) );
  XNOR2_X1 U6577 ( .A(DATAI_10_), .B(keyinput_21), .ZN(n5808) );
  NAND3_X1 U6578 ( .A1(n5810), .A2(n5809), .A3(n5808), .ZN(n5817) );
  XNOR2_X1 U6579 ( .A(DATAI_8_), .B(keyinput_23), .ZN(n5816) );
  XOR2_X1 U6580 ( .A(DATAI_4_), .B(keyinput_27), .Z(n5814) );
  XNOR2_X1 U6581 ( .A(DATAI_5_), .B(keyinput_26), .ZN(n5813) );
  XNOR2_X1 U6582 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n5812) );
  XNOR2_X1 U6583 ( .A(DATAI_7_), .B(keyinput_24), .ZN(n5811) );
  NAND4_X1 U6584 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n5815)
         );
  AOI21_X1 U6585 ( .B1(n5817), .B2(n5816), .A(n5815), .ZN(n5820) );
  XOR2_X1 U6586 ( .A(DATAI_3_), .B(keyinput_28), .Z(n5819) );
  XOR2_X1 U6587 ( .A(DATAI_2_), .B(keyinput_29), .Z(n5818) );
  NOR3_X1 U6588 ( .A1(n5820), .A2(n5819), .A3(n5818), .ZN(n5823) );
  XNOR2_X1 U6589 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n5822) );
  XNOR2_X1 U6590 ( .A(DATAI_0_), .B(keyinput_31), .ZN(n5821) );
  NOR3_X1 U6591 ( .A1(n5823), .A2(n5822), .A3(n5821), .ZN(n5829) );
  XNOR2_X1 U6592 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(keyinput_32), .ZN(n5828) );
  XNOR2_X1 U6593 ( .A(n6738), .B(keyinput_34), .ZN(n5826) );
  XNOR2_X1 U6594 ( .A(READY_N), .B(keyinput_35), .ZN(n5825) );
  XNOR2_X1 U6595 ( .A(NA_N), .B(keyinput_33), .ZN(n5824) );
  NOR3_X1 U6596 ( .A1(n5826), .A2(n5825), .A3(n5824), .ZN(n5827) );
  OAI21_X1 U6597 ( .B1(n5829), .B2(n5828), .A(n5827), .ZN(n5833) );
  XOR2_X1 U6598 ( .A(HOLD), .B(keyinput_36), .Z(n5832) );
  XNOR2_X1 U6599 ( .A(n6753), .B(keyinput_38), .ZN(n5831) );
  XNOR2_X1 U6600 ( .A(READREQUEST_REG_SCAN_IN), .B(keyinput_37), .ZN(n5830) );
  AOI211_X1 U6601 ( .C1(n5833), .C2(n5832), .A(n5831), .B(n5830), .ZN(n5836)
         );
  XOR2_X1 U6602 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_39), .Z(n5835) );
  XNOR2_X1 U6603 ( .A(n7351), .B(keyinput_40), .ZN(n5834) );
  NOR3_X1 U6604 ( .A1(n5836), .A2(n5835), .A3(n5834), .ZN(n5839) );
  XOR2_X1 U6605 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_42), .Z(n5838)
         );
  XNOR2_X1 U6606 ( .A(D_C_N_REG_SCAN_IN), .B(keyinput_41), .ZN(n5837) );
  NOR3_X1 U6607 ( .A1(n5839), .A2(n5838), .A3(n5837), .ZN(n5851) );
  XNOR2_X1 U6608 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(keyinput_48), .ZN(n5841)
         );
  XNOR2_X1 U6609 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_47), .ZN(n5840)
         );
  NOR2_X1 U6610 ( .A1(n5841), .A2(n5840), .ZN(n5847) );
  XNOR2_X1 U6611 ( .A(FLUSH_REG_SCAN_IN), .B(keyinput_45), .ZN(n5843) );
  XNOR2_X1 U6612 ( .A(MORE_REG_SCAN_IN), .B(keyinput_44), .ZN(n5842) );
  NOR2_X1 U6613 ( .A1(n5843), .A2(n5842), .ZN(n5846) );
  XNOR2_X1 U6614 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_43), .ZN(n5845) );
  XNOR2_X1 U6615 ( .A(W_R_N_REG_SCAN_IN), .B(keyinput_46), .ZN(n5844) );
  NAND4_X1 U6616 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n5850)
         );
  XNOR2_X1 U6617 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_50), .ZN(n5849)
         );
  XNOR2_X1 U6618 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_49), .ZN(n5848)
         );
  OAI211_X1 U6619 ( .C1(n5851), .C2(n5850), .A(n5849), .B(n5848), .ZN(n5854)
         );
  XNOR2_X1 U6620 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_51), .ZN(n5853) );
  XNOR2_X1 U6621 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_52), .ZN(n5852) );
  AOI21_X1 U6622 ( .B1(n5854), .B2(n5853), .A(n5852), .ZN(n5863) );
  INV_X1 U6623 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6831) );
  OAI22_X1 U6624 ( .A1(n6831), .A2(keyinput_53), .B1(n7232), .B2(keyinput_57), 
        .ZN(n5855) );
  AOI221_X1 U6625 ( .B1(n6831), .B2(keyinput_53), .C1(keyinput_57), .C2(n7232), 
        .A(n5855), .ZN(n5859) );
  XOR2_X1 U6626 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .Z(n5858) );
  INV_X1 U6627 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6828) );
  OAI22_X1 U6628 ( .A1(n6828), .A2(keyinput_55), .B1(REIP_REG_28__SCAN_IN), 
        .B2(keyinput_54), .ZN(n5856) );
  AOI221_X1 U6629 ( .B1(n6828), .B2(keyinput_55), .C1(keyinput_54), .C2(
        REIP_REG_28__SCAN_IN), .A(n5856), .ZN(n5857) );
  NAND3_X1 U6630 ( .A1(n5859), .A2(n5858), .A3(n5857), .ZN(n5862) );
  XOR2_X1 U6631 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .Z(n5861) );
  XNOR2_X1 U6632 ( .A(n6527), .B(keyinput_59), .ZN(n5860) );
  OAI211_X1 U6633 ( .C1(n5863), .C2(n5862), .A(n5861), .B(n5860), .ZN(n5866)
         );
  XOR2_X1 U6634 ( .A(REIP_REG_22__SCAN_IN), .B(keyinput_60), .Z(n5865) );
  XNOR2_X1 U6635 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_61), .ZN(n5864) );
  NAND3_X1 U6636 ( .A1(n5866), .A2(n5865), .A3(n5864), .ZN(n5870) );
  XOR2_X1 U6637 ( .A(REIP_REG_18__SCAN_IN), .B(keyinput_64), .Z(n5869) );
  XNOR2_X1 U6638 ( .A(REIP_REG_19__SCAN_IN), .B(keyinput_63), .ZN(n5868) );
  XNOR2_X1 U6639 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_62), .ZN(n5867) );
  NAND4_X1 U6640 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(n5873)
         );
  XOR2_X1 U6641 ( .A(REIP_REG_17__SCAN_IN), .B(keyinput_65), .Z(n5872) );
  XOR2_X1 U6642 ( .A(REIP_REG_16__SCAN_IN), .B(keyinput_66), .Z(n5871) );
  AOI21_X1 U6643 ( .B1(n5873), .B2(n5872), .A(n5871), .ZN(n5877) );
  XNOR2_X1 U6644 ( .A(BE_N_REG_3__SCAN_IN), .B(keyinput_67), .ZN(n5876) );
  INV_X1 U6645 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n6851) );
  XNOR2_X1 U6646 ( .A(n6851), .B(keyinput_68), .ZN(n5875) );
  XNOR2_X1 U6647 ( .A(BE_N_REG_1__SCAN_IN), .B(keyinput_69), .ZN(n5874) );
  OAI211_X1 U6648 ( .C1(n5877), .C2(n5876), .A(n5875), .B(n5874), .ZN(n5880)
         );
  XNOR2_X1 U6649 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_70), .ZN(n5879) );
  INV_X1 U6650 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6835) );
  XNOR2_X1 U6651 ( .A(n6835), .B(keyinput_71), .ZN(n5878) );
  AOI21_X1 U6652 ( .B1(n5880), .B2(n5879), .A(n5878), .ZN(n5883) );
  XNOR2_X1 U6653 ( .A(n6832), .B(keyinput_72), .ZN(n5882) );
  XNOR2_X1 U6654 ( .A(n6830), .B(keyinput_73), .ZN(n5881) );
  OAI21_X1 U6655 ( .B1(n5883), .B2(n5882), .A(n5881), .ZN(n5887) );
  XNOR2_X1 U6656 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_74), .ZN(n5886) );
  XNOR2_X1 U6657 ( .A(n6823), .B(keyinput_75), .ZN(n5885) );
  INV_X1 U6658 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6822) );
  XNOR2_X1 U6659 ( .A(n6822), .B(keyinput_76), .ZN(n5884) );
  AOI211_X1 U6660 ( .C1(n5887), .C2(n5886), .A(n5885), .B(n5884), .ZN(n5890)
         );
  XNOR2_X1 U6661 ( .A(n6821), .B(keyinput_77), .ZN(n5889) );
  INV_X1 U6662 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6820) );
  XNOR2_X1 U6663 ( .A(n6820), .B(keyinput_78), .ZN(n5888) );
  NOR3_X1 U6664 ( .A1(n5890), .A2(n5889), .A3(n5888), .ZN(n5893) );
  INV_X1 U6665 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6818) );
  XNOR2_X1 U6666 ( .A(n6818), .B(keyinput_79), .ZN(n5892) );
  XNOR2_X1 U6667 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_80), .ZN(n5891) );
  OAI21_X1 U6668 ( .B1(n5893), .B2(n5892), .A(n5891), .ZN(n5896) );
  XNOR2_X1 U6669 ( .A(ADDRESS_REG_19__SCAN_IN), .B(keyinput_81), .ZN(n5895) );
  INV_X1 U6670 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6814) );
  XNOR2_X1 U6671 ( .A(n6814), .B(keyinput_82), .ZN(n5894) );
  AOI21_X1 U6672 ( .B1(n5896), .B2(n5895), .A(n5894), .ZN(n5900) );
  XNOR2_X1 U6673 ( .A(n6813), .B(keyinput_83), .ZN(n5899) );
  INV_X1 U6674 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6810) );
  XNOR2_X1 U6675 ( .A(n6810), .B(keyinput_85), .ZN(n5898) );
  INV_X1 U6676 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6811) );
  XNOR2_X1 U6677 ( .A(n6811), .B(keyinput_84), .ZN(n5897) );
  OAI211_X1 U6678 ( .C1(n5900), .C2(n5899), .A(n5898), .B(n5897), .ZN(n5903)
         );
  INV_X1 U6679 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6808) );
  XNOR2_X1 U6680 ( .A(n6808), .B(keyinput_86), .ZN(n5902) );
  XNOR2_X1 U6681 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_87), .ZN(n5901) );
  AOI21_X1 U6682 ( .B1(n5903), .B2(n5902), .A(n5901), .ZN(n5909) );
  XNOR2_X1 U6683 ( .A(ADDRESS_REG_12__SCAN_IN), .B(keyinput_88), .ZN(n5908) );
  XOR2_X1 U6684 ( .A(ADDRESS_REG_9__SCAN_IN), .B(keyinput_91), .Z(n5906) );
  XNOR2_X1 U6685 ( .A(ADDRESS_REG_10__SCAN_IN), .B(keyinput_90), .ZN(n5905) );
  XNOR2_X1 U6686 ( .A(ADDRESS_REG_11__SCAN_IN), .B(keyinput_89), .ZN(n5904) );
  NOR3_X1 U6687 ( .A1(n5906), .A2(n5905), .A3(n5904), .ZN(n5907) );
  OAI21_X1 U6688 ( .B1(n5909), .B2(n5908), .A(n5907), .ZN(n5912) );
  XNOR2_X1 U6689 ( .A(ADDRESS_REG_8__SCAN_IN), .B(keyinput_92), .ZN(n5911) );
  XNOR2_X1 U6690 ( .A(ADDRESS_REG_7__SCAN_IN), .B(keyinput_93), .ZN(n5910) );
  AOI21_X1 U6691 ( .B1(n5912), .B2(n5911), .A(n5910), .ZN(n5915) );
  XNOR2_X1 U6692 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_94), .ZN(n5914) );
  XNOR2_X1 U6693 ( .A(n6793), .B(keyinput_95), .ZN(n5913) );
  OAI21_X1 U6694 ( .B1(n5915), .B2(n5914), .A(n5913), .ZN(n5924) );
  XNOR2_X1 U6695 ( .A(n6792), .B(keyinput_96), .ZN(n5923) );
  XOR2_X1 U6696 ( .A(ADDRESS_REG_3__SCAN_IN), .B(keyinput_97), .Z(n5918) );
  XNOR2_X1 U6697 ( .A(n7343), .B(keyinput_101), .ZN(n5917) );
  XNOR2_X1 U6698 ( .A(n6787), .B(keyinput_99), .ZN(n5916) );
  NOR3_X1 U6699 ( .A1(n5918), .A2(n5917), .A3(n5916), .ZN(n5921) );
  XNOR2_X1 U6700 ( .A(keyinput_100), .B(ADDRESS_REG_0__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U6701 ( .A(keyinput_98), .B(ADDRESS_REG_2__SCAN_IN), .ZN(n5919) );
  NAND3_X1 U6702 ( .A1(n5921), .A2(n5920), .A3(n5919), .ZN(n5922) );
  AOI21_X1 U6703 ( .B1(n5924), .B2(n5923), .A(n5922), .ZN(n5928) );
  XNOR2_X1 U6704 ( .A(n7334), .B(keyinput_102), .ZN(n5927) );
  XNOR2_X1 U6705 ( .A(DATAWIDTH_REG_0__SCAN_IN), .B(keyinput_104), .ZN(n5926)
         );
  XNOR2_X1 U6706 ( .A(STATE_REG_0__SCAN_IN), .B(keyinput_103), .ZN(n5925) );
  OAI211_X1 U6707 ( .C1(n5928), .C2(n5927), .A(n5926), .B(n5925), .ZN(n5931)
         );
  XOR2_X1 U6708 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_105), .Z(n5930) );
  XOR2_X1 U6709 ( .A(DATAWIDTH_REG_2__SCAN_IN), .B(keyinput_106), .Z(n5929) );
  AOI21_X1 U6710 ( .B1(n5931), .B2(n5930), .A(n5929), .ZN(n5951) );
  XOR2_X1 U6711 ( .A(DATAWIDTH_REG_4__SCAN_IN), .B(keyinput_108), .Z(n5935) );
  XNOR2_X1 U6712 ( .A(n6742), .B(keyinput_110), .ZN(n5934) );
  XNOR2_X1 U6713 ( .A(DATAWIDTH_REG_3__SCAN_IN), .B(keyinput_107), .ZN(n5933)
         );
  XNOR2_X1 U6714 ( .A(DATAWIDTH_REG_5__SCAN_IN), .B(keyinput_109), .ZN(n5932)
         );
  NAND4_X1 U6715 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n5950)
         );
  INV_X1 U6716 ( .A(keyinput_120), .ZN(n5936) );
  XNOR2_X1 U6717 ( .A(n5936), .B(DATAWIDTH_REG_16__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U6718 ( .A(DATAWIDTH_REG_11__SCAN_IN), .B(keyinput_115), .ZN(n5939)
         );
  XNOR2_X1 U6719 ( .A(DATAWIDTH_REG_14__SCAN_IN), .B(keyinput_118), .ZN(n5938)
         );
  XNOR2_X1 U6720 ( .A(DATAWIDTH_REG_15__SCAN_IN), .B(keyinput_119), .ZN(n5937)
         );
  NAND4_X1 U6721 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n5948)
         );
  XNOR2_X1 U6722 ( .A(DATAWIDTH_REG_9__SCAN_IN), .B(keyinput_113), .ZN(n5944)
         );
  XNOR2_X1 U6723 ( .A(DATAWIDTH_REG_7__SCAN_IN), .B(keyinput_111), .ZN(n5943)
         );
  XNOR2_X1 U6724 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_114), .ZN(n5942)
         );
  XNOR2_X1 U6725 ( .A(DATAWIDTH_REG_13__SCAN_IN), .B(keyinput_117), .ZN(n5941)
         );
  NAND4_X1 U6726 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n5947)
         );
  XNOR2_X1 U6727 ( .A(DATAWIDTH_REG_8__SCAN_IN), .B(keyinput_112), .ZN(n5946)
         );
  XNOR2_X1 U6728 ( .A(DATAWIDTH_REG_12__SCAN_IN), .B(keyinput_116), .ZN(n5945)
         );
  NOR4_X1 U6729 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n5949)
         );
  OAI21_X1 U6730 ( .B1(n5951), .B2(n5950), .A(n5949), .ZN(n5962) );
  XNOR2_X1 U6731 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_124), .ZN(n5955)
         );
  XNOR2_X1 U6732 ( .A(DATAWIDTH_REG_19__SCAN_IN), .B(keyinput_123), .ZN(n5954)
         );
  XNOR2_X1 U6733 ( .A(DATAWIDTH_REG_17__SCAN_IN), .B(keyinput_121), .ZN(n5953)
         );
  XNOR2_X1 U6734 ( .A(DATAWIDTH_REG_18__SCAN_IN), .B(keyinput_122), .ZN(n5952)
         );
  NOR4_X1 U6735 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n5961)
         );
  XNOR2_X1 U6736 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_125), .ZN(n5960)
         );
  INV_X1 U6737 ( .A(keyinput_127), .ZN(n5956) );
  XNOR2_X1 U6738 ( .A(n5956), .B(DATAWIDTH_REG_23__SCAN_IN), .ZN(n5958) );
  XNOR2_X1 U6739 ( .A(DATAWIDTH_REG_22__SCAN_IN), .B(keyinput_126), .ZN(n5957)
         );
  NAND2_X1 U6740 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  AOI211_X1 U6741 ( .C1(n5962), .C2(n5961), .A(n5960), .B(n5959), .ZN(n5963)
         );
  NAND2_X1 U6742 ( .A1(n5964), .A2(n5963), .ZN(n5982) );
  NAND3_X1 U6743 ( .A1(n5112), .A2(n7324), .A3(n6058), .ZN(n7385) );
  NAND2_X1 U6744 ( .A1(n7389), .A2(n7385), .ZN(n5965) );
  AOI21_X1 U6745 ( .B1(n5965), .B2(STATEBS16_REG_SCAN_IN), .A(n7445), .ZN(
        n5976) );
  NOR2_X1 U6746 ( .A1(n6005), .A2(n5966), .ZN(n7379) );
  INV_X1 U6747 ( .A(n7379), .ZN(n5971) );
  NOR3_X1 U6748 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7268), .A3(n7448), 
        .ZN(n7384) );
  NAND2_X1 U6749 ( .A1(n7384), .A2(n7394), .ZN(n5972) );
  AOI211_X1 U6750 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5972), .A(n5968), .B(
        n5967), .ZN(n5969) );
  INV_X1 U6751 ( .A(n5969), .ZN(n5970) );
  AOI21_X1 U6752 ( .B1(n5976), .B2(n5971), .A(n5970), .ZN(n7388) );
  INV_X1 U6753 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5980) );
  INV_X1 U6754 ( .A(n5972), .ZN(n7611) );
  OAI22_X1 U6755 ( .A1(n7389), .A2(n6108), .B1(n7385), .B2(n5973), .ZN(n5978)
         );
  AOI22_X1 U6756 ( .A1(n5976), .A2(n7379), .B1(n5975), .B2(n5974), .ZN(n7615)
         );
  NOR2_X1 U6757 ( .A1(n7615), .A2(n7596), .ZN(n5977) );
  AOI211_X1 U6758 ( .C1(n7591), .C2(n7611), .A(n5978), .B(n5977), .ZN(n5979)
         );
  OAI21_X1 U6759 ( .B1(n7388), .B2(n5980), .A(n5979), .ZN(n5981) );
  XNOR2_X1 U6760 ( .A(n5982), .B(n5981), .ZN(U3106) );
  INV_X1 U6761 ( .A(n5983), .ZN(n5986) );
  NAND2_X1 U6762 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n7137) );
  NOR2_X1 U6763 ( .A1(n7192), .A2(n6014), .ZN(n7087) );
  INV_X1 U6764 ( .A(n7087), .ZN(n5984) );
  NOR2_X1 U6765 ( .A1(n5984), .A2(n7086), .ZN(n7116) );
  NAND2_X1 U6766 ( .A1(REIP_REG_5__SCAN_IN), .A2(n7116), .ZN(n7134) );
  NOR3_X1 U6767 ( .A1(REIP_REG_8__SCAN_IN), .A2(n7137), .A3(n7134), .ZN(n5985)
         );
  AOI21_X1 U6768 ( .B1(n7199), .B2(n5986), .A(n5985), .ZN(n5992) );
  INV_X1 U6769 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6795) );
  AOI21_X1 U6770 ( .B1(n7228), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n7183), 
        .ZN(n5989) );
  INV_X1 U6771 ( .A(n5987), .ZN(n7007) );
  AOI22_X1 U6772 ( .A1(n7227), .A2(EBX_REG_8__SCAN_IN), .B1(n7235), .B2(n7007), 
        .ZN(n5988) );
  OAI211_X1 U6773 ( .C1(n6027), .C2(n6795), .A(n5989), .B(n5988), .ZN(n5990)
         );
  INV_X1 U6774 ( .A(n5990), .ZN(n5991) );
  OAI211_X1 U6775 ( .C1(n5993), .C2(n7196), .A(n5992), .B(n5991), .ZN(U2819)
         );
  OAI21_X1 U6776 ( .B1(n5996), .B2(n5995), .A(n3656), .ZN(n7035) );
  INV_X1 U6777 ( .A(n5997), .ZN(n6001) );
  AOI22_X1 U6778 ( .A1(n6932), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n7059), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5998) );
  OAI21_X1 U6779 ( .B1(n6940), .B2(n5999), .A(n5998), .ZN(n6000) );
  AOI21_X1 U6780 ( .B1(n6001), .B2(n6937), .A(n6000), .ZN(n6002) );
  OAI21_X1 U6781 ( .B1(n7035), .B2(n7241), .A(n6002), .ZN(U2977) );
  INV_X1 U6782 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6994) );
  NOR2_X1 U6783 ( .A1(n6852), .A2(n6994), .ZN(n6003) );
  NAND3_X1 U6784 ( .A1(n7178), .A2(n6003), .A3(n6014), .ZN(n6004) );
  OAI21_X1 U6785 ( .B1(n6005), .B2(n7094), .A(n6004), .ZN(n6013) );
  NOR2_X1 U6786 ( .A1(n7203), .A2(n6006), .ZN(n6012) );
  NOR2_X1 U6787 ( .A1(n7195), .A2(n6007), .ZN(n6011) );
  OAI22_X1 U6788 ( .A1(n6009), .A2(n7215), .B1(n7239), .B2(n6008), .ZN(n6010)
         );
  NOR4_X1 U6789 ( .A1(n6013), .A2(n6012), .A3(n6011), .A4(n6010), .ZN(n6017)
         );
  INV_X1 U6790 ( .A(n6014), .ZN(n6015) );
  OAI21_X1 U6791 ( .B1(n7192), .B2(n6015), .A(n7114), .ZN(n7088) );
  NAND2_X1 U6792 ( .A1(n7088), .A2(REIP_REG_3__SCAN_IN), .ZN(n6016) );
  OAI211_X1 U6793 ( .C1(n7097), .C2(n6018), .A(n6017), .B(n6016), .ZN(U2824)
         );
  INV_X1 U6794 ( .A(n6019), .ZN(n6020) );
  AOI21_X1 U6795 ( .B1(n6021), .B2(n5538), .A(n6020), .ZN(n6140) );
  INV_X1 U6796 ( .A(n6140), .ZN(n6044) );
  INV_X1 U6797 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6026) );
  AND2_X1 U6798 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  OR2_X1 U6799 ( .A1(n6024), .A2(n6040), .ZN(n7028) );
  OAI222_X1 U6800 ( .A1(n6044), .A2(n6478), .B1(n6880), .B2(n6026), .C1(n7028), 
        .C2(n6876), .ZN(U2849) );
  INV_X1 U6801 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6025) );
  OAI22_X1 U6802 ( .A1(n6025), .A2(n7215), .B1(n7239), .B2(n6135), .ZN(n6029)
         );
  INV_X1 U6803 ( .A(REIP_REG_10__SCAN_IN), .ZN(n7027) );
  OAI22_X1 U6804 ( .A1(n6027), .A2(n7027), .B1(n6026), .B2(n7203), .ZN(n6028)
         );
  OR3_X1 U6805 ( .A1(n6029), .A2(n7183), .A3(n6028), .ZN(n6035) );
  INV_X1 U6806 ( .A(n6030), .ZN(n6031) );
  OAI211_X1 U6807 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n6032), .B(n6031), .ZN(n6033) );
  OAI22_X1 U6808 ( .A1(n7195), .A2(n7028), .B1(n7192), .B2(n6033), .ZN(n6034)
         );
  AOI211_X1 U6809 ( .C1(n6140), .C2(n7236), .A(n6035), .B(n6034), .ZN(n6036)
         );
  INV_X1 U6810 ( .A(n6036), .ZN(U2817) );
  AOI21_X1 U6811 ( .B1(n6038), .B2(n6019), .A(n6037), .ZN(n6091) );
  INV_X1 U6812 ( .A(n6091), .ZN(n6055) );
  INV_X1 U6813 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6042) );
  NOR2_X1 U6814 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  OR2_X1 U6815 ( .A1(n6075), .A2(n6041), .ZN(n7042) );
  OAI222_X1 U6816 ( .A1(n6055), .A2(n6468), .B1(n6042), .B2(n6880), .C1(n6876), 
        .C2(n7042), .ZN(U2848) );
  INV_X1 U6817 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6777) );
  OAI222_X1 U6818 ( .A1(n6055), .A2(n7352), .B1(n6219), .B2(n6043), .C1(n6311), 
        .C2(n6777), .ZN(U2880) );
  INV_X1 U6819 ( .A(DATAI_10_), .ZN(n6045) );
  INV_X1 U6820 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6775) );
  OAI222_X1 U6821 ( .A1(n6045), .A2(n6219), .B1(n6311), .B2(n6775), .C1(n7352), 
        .C2(n6044), .ZN(U2881) );
  NOR2_X1 U6822 ( .A1(n6421), .A2(n6194), .ZN(n6046) );
  NOR2_X1 U6823 ( .A1(n6407), .A2(n6046), .ZN(n6147) );
  AOI21_X1 U6824 ( .B1(n7199), .B2(n6047), .A(n7183), .ZN(n6048) );
  OAI21_X1 U6825 ( .B1(n7195), .B2(n7042), .A(n6048), .ZN(n6053) );
  NAND2_X1 U6826 ( .A1(n7178), .A2(n6049), .ZN(n6051) );
  AOI22_X1 U6827 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n7228), .B1(
        EBX_REG_11__SCAN_IN), .B2(n7227), .ZN(n6050) );
  OAI21_X1 U6828 ( .B1(REIP_REG_11__SCAN_IN), .B2(n6051), .A(n6050), .ZN(n6052) );
  AOI211_X1 U6829 ( .C1(n6147), .C2(REIP_REG_11__SCAN_IN), .A(n6053), .B(n6052), .ZN(n6054) );
  OAI21_X1 U6830 ( .B1(n6055), .B2(n7196), .A(n6054), .ZN(U2816) );
  NOR3_X1 U6831 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6251), .A3(n7268), 
        .ZN(n7372) );
  INV_X1 U6832 ( .A(n7372), .ZN(n7373) );
  NOR2_X1 U6833 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7373), .ZN(n6733)
         );
  INV_X1 U6834 ( .A(n6733), .ZN(n6057) );
  AOI211_X1 U6835 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6057), .A(n6056), .B(
        n6095), .ZN(n6062) );
  OAI21_X1 U6836 ( .B1(n7597), .B2(n7604), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6059) );
  OAI21_X1 U6837 ( .B1(n6103), .B2(n6060), .A(n6059), .ZN(n6061) );
  NAND2_X1 U6838 ( .A1(n6062), .A2(n6061), .ZN(n6729) );
  INV_X1 U6839 ( .A(n7604), .ZN(n6695) );
  NAND2_X1 U6840 ( .A1(n6093), .A2(n7417), .ZN(n6065) );
  NAND2_X1 U6841 ( .A1(n6063), .A2(n6101), .ZN(n6064) );
  NAND2_X1 U6842 ( .A1(n6065), .A2(n6064), .ZN(n6730) );
  AOI22_X1 U6843 ( .A1(n7597), .A2(n7534), .B1(n6066), .B2(n6730), .ZN(n6068)
         );
  NAND2_X1 U6844 ( .A1(n7533), .A2(n6733), .ZN(n6067) );
  OAI211_X1 U6845 ( .C1(n6695), .C2(n6113), .A(n6068), .B(n6067), .ZN(n6069)
         );
  AOI21_X1 U6846 ( .B1(n6729), .B2(INSTQUEUE_REG_12__3__SCAN_IN), .A(n6069), 
        .ZN(n6070) );
  INV_X1 U6847 ( .A(n6070), .ZN(U3119) );
  OAI21_X1 U6848 ( .B1(n6037), .B2(n6072), .A(n6071), .ZN(n6176) );
  INV_X1 U6849 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6082) );
  AOI21_X1 U6850 ( .B1(n7228), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n7183), 
        .ZN(n6073) );
  OAI21_X1 U6851 ( .B1(n6082), .B2(n7203), .A(n6073), .ZN(n6080) );
  NOR2_X1 U6852 ( .A1(n7192), .A2(n6194), .ZN(n6193) );
  INV_X1 U6853 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6803) );
  OR2_X1 U6854 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  NAND2_X1 U6855 ( .A1(n6144), .A2(n6076), .ZN(n6164) );
  OAI22_X1 U6856 ( .A1(n7195), .A2(n6164), .B1(n6171), .B2(n7239), .ZN(n6077)
         );
  AOI21_X1 U6857 ( .B1(n6193), .B2(n6803), .A(n6077), .ZN(n6078) );
  INV_X1 U6858 ( .A(n6078), .ZN(n6079) );
  AOI211_X1 U6859 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6147), .A(n6080), .B(n6079), .ZN(n6081) );
  OAI21_X1 U6860 ( .B1(n6176), .B2(n7196), .A(n6081), .ZN(U2815) );
  OAI222_X1 U6861 ( .A1(n6164), .A2(n6876), .B1(n6880), .B2(n6082), .C1(n6176), 
        .C2(n6468), .ZN(U2847) );
  INV_X1 U6862 ( .A(DATAI_12_), .ZN(n6083) );
  INV_X1 U6863 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6779) );
  OAI222_X1 U6864 ( .A1(n6219), .A2(n6083), .B1(n6311), .B2(n6779), .C1(n7352), 
        .C2(n6176), .ZN(U2879) );
  XNOR2_X1 U6865 ( .A(n3650), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6136)
         );
  NAND2_X1 U6866 ( .A1(n6084), .A2(n6136), .ZN(n7032) );
  OAI21_X1 U6867 ( .B1(n4215), .B2(n3650), .A(n7032), .ZN(n6087) );
  INV_X1 U6868 ( .A(n6155), .ZN(n6085) );
  AOI21_X1 U6869 ( .B1(n3650), .B2(n6163), .A(n6085), .ZN(n6086) );
  NAND2_X1 U6870 ( .A1(n6087), .A2(n6086), .ZN(n6156) );
  OAI21_X1 U6871 ( .B1(n6087), .B2(n6086), .A(n6156), .ZN(n7046) );
  NAND2_X1 U6872 ( .A1(n7059), .A2(REIP_REG_11__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U6873 ( .A1(n6932), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6088)
         );
  OAI211_X1 U6874 ( .C1(n6940), .C2(n6089), .A(n7043), .B(n6088), .ZN(n6090)
         );
  AOI21_X1 U6875 ( .B1(n6091), .B2(n6937), .A(n6090), .ZN(n6092) );
  OAI21_X1 U6876 ( .B1(n7046), .B2(n7241), .A(n6092), .ZN(U2975) );
  AND2_X1 U6877 ( .A1(n7394), .A2(n7414), .ZN(n6100) );
  INV_X1 U6878 ( .A(n6100), .ZN(n6294) );
  NAND2_X1 U6879 ( .A1(n7420), .A2(n5161), .ZN(n6290) );
  OAI21_X1 U6880 ( .B1(n7630), .B2(n7622), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6097) );
  OR2_X1 U6881 ( .A1(n6094), .A2(n6093), .ZN(n6096) );
  AOI21_X1 U6882 ( .B1(n6097), .B2(n6096), .A(n6095), .ZN(n6099) );
  NAND2_X1 U6883 ( .A1(n6288), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6106) );
  AOI22_X1 U6884 ( .A1(n6103), .A2(n7409), .B1(n6102), .B2(n6101), .ZN(n6289)
         );
  OAI22_X1 U6885 ( .A1(n6290), .A2(n6694), .B1(n6289), .B2(n7465), .ZN(n6104)
         );
  AOI21_X1 U6886 ( .B1(n7454), .B2(n7622), .A(n6104), .ZN(n6105) );
  OAI211_X1 U6887 ( .C1(n6107), .C2(n6294), .A(n6106), .B(n6105), .ZN(U3068)
         );
  NAND2_X1 U6888 ( .A1(n6288), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6111) );
  OAI22_X1 U6889 ( .A1(n6290), .A2(n6108), .B1(n6289), .B2(n7596), .ZN(n6109)
         );
  AOI21_X1 U6890 ( .B1(n7592), .B2(n7622), .A(n6109), .ZN(n6110) );
  OAI211_X1 U6891 ( .C1(n6294), .C2(n6112), .A(n6111), .B(n6110), .ZN(U3074)
         );
  NAND2_X1 U6892 ( .A1(n6288), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6116) );
  OAI22_X1 U6893 ( .A1(n6290), .A2(n6113), .B1(n6289), .B2(n7538), .ZN(n6114)
         );
  AOI21_X1 U6894 ( .B1(n7622), .B2(n7534), .A(n6114), .ZN(n6115) );
  OAI211_X1 U6895 ( .C1(n6294), .C2(n6117), .A(n6116), .B(n6115), .ZN(U3071)
         );
  NAND2_X1 U6896 ( .A1(n6288), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6121) );
  OAI22_X1 U6897 ( .A1(n6290), .A2(n6118), .B1(n6289), .B2(n7511), .ZN(n6119)
         );
  AOI21_X1 U6898 ( .B1(n7622), .B2(n7507), .A(n6119), .ZN(n6120) );
  OAI211_X1 U6899 ( .C1(n6294), .C2(n6707), .A(n6121), .B(n6120), .ZN(U3070)
         );
  NAND2_X1 U6900 ( .A1(n6288), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6125) );
  OAI22_X1 U6901 ( .A1(n6290), .A2(n6122), .B1(n6289), .B2(n7488), .ZN(n6123)
         );
  AOI21_X1 U6902 ( .B1(n7622), .B2(n7484), .A(n6123), .ZN(n6124) );
  OAI211_X1 U6903 ( .C1(n6294), .C2(n6701), .A(n6125), .B(n6124), .ZN(U3069)
         );
  NAND2_X1 U6904 ( .A1(n6288), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6129) );
  OAI22_X1 U6905 ( .A1(n6290), .A2(n6126), .B1(n6289), .B2(n7652), .ZN(n6127)
         );
  AOI21_X1 U6906 ( .B1(n7622), .B2(n7645), .A(n6127), .ZN(n6128) );
  OAI211_X1 U6907 ( .C1(n6294), .C2(n6732), .A(n6129), .B(n6128), .ZN(U3075)
         );
  NAND2_X1 U6908 ( .A1(n6288), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6133) );
  OAI22_X1 U6909 ( .A1(n6290), .A2(n6130), .B1(n6289), .B2(n7558), .ZN(n6131)
         );
  AOI21_X1 U6910 ( .B1(n7622), .B2(n7554), .A(n6131), .ZN(n6132) );
  OAI211_X1 U6911 ( .C1(n6294), .C2(n6713), .A(n6133), .B(n6132), .ZN(U3072)
         );
  AOI22_X1 U6912 ( .A1(n6932), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n7183), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n6134) );
  OAI21_X1 U6913 ( .B1(n6135), .B2(n6940), .A(n6134), .ZN(n6139) );
  NOR2_X1 U6914 ( .A1(n6084), .A2(n6136), .ZN(n7024) );
  INV_X1 U6915 ( .A(n7032), .ZN(n6137) );
  NOR3_X1 U6916 ( .A1(n7024), .A2(n6137), .A3(n7241), .ZN(n6138) );
  AOI211_X1 U6917 ( .C1(n6937), .C2(n6140), .A(n6139), .B(n6138), .ZN(n6141)
         );
  INV_X1 U6918 ( .A(n6141), .ZN(U2976) );
  XNOR2_X1 U6919 ( .A(n6142), .B(n6143), .ZN(n6184) );
  INV_X1 U6920 ( .A(n6190), .ZN(n6215) );
  AOI21_X1 U6921 ( .B1(n6145), .B2(n6144), .A(n6215), .ZN(n6970) );
  AOI21_X1 U6922 ( .B1(n7199), .B2(n6181), .A(n7183), .ZN(n6146) );
  OAI21_X1 U6923 ( .B1(n6179), .B2(n7215), .A(n6146), .ZN(n6152) );
  AOI22_X1 U6924 ( .A1(EBX_REG_13__SCAN_IN), .A2(n7227), .B1(
        REIP_REG_13__SCAN_IN), .B2(n6147), .ZN(n6150) );
  NAND2_X1 U6925 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n6148) );
  OAI211_X1 U6926 ( .C1(REIP_REG_13__SCAN_IN), .C2(REIP_REG_12__SCAN_IN), .A(
        n6193), .B(n6148), .ZN(n6149) );
  NAND2_X1 U6927 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  AOI211_X1 U6928 ( .C1(n6970), .C2(n7235), .A(n6152), .B(n6151), .ZN(n6153)
         );
  OAI21_X1 U6929 ( .B1(n6184), .B2(n7196), .A(n6153), .ZN(U2814) );
  AOI22_X1 U6930 ( .A1(n6970), .A2(n6868), .B1(EBX_REG_13__SCAN_IN), .B2(n6475), .ZN(n6154) );
  OAI21_X1 U6931 ( .B1(n6184), .B2(n6468), .A(n6154), .ZN(U2846) );
  NAND2_X1 U6932 ( .A1(n6156), .A2(n6155), .ZN(n6158) );
  XNOR2_X1 U6933 ( .A(n3650), .B(n4214), .ZN(n6157) );
  XNOR2_X1 U6934 ( .A(n6158), .B(n6157), .ZN(n6170) );
  INV_X1 U6935 ( .A(n6170), .ZN(n6169) );
  NOR2_X1 U6936 ( .A1(n6160), .A2(n6159), .ZN(n6976) );
  NOR2_X1 U6937 ( .A1(n7009), .A2(n6976), .ZN(n7047) );
  INV_X1 U6938 ( .A(n7047), .ZN(n6162) );
  NAND2_X1 U6939 ( .A1(n6163), .A2(n6161), .ZN(n7049) );
  AOI21_X1 U6940 ( .B1(n6162), .B2(n7049), .A(n4214), .ZN(n6167) );
  AND2_X1 U6941 ( .A1(n7183), .A2(REIP_REG_12__SCAN_IN), .ZN(n6173) );
  NOR3_X1 U6942 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6981), .A3(n6163), 
        .ZN(n6166) );
  NOR2_X1 U6943 ( .A1(n7029), .A2(n6164), .ZN(n6165) );
  NOR4_X1 U6944 ( .A1(n6167), .A2(n6173), .A3(n6166), .A4(n6165), .ZN(n6168)
         );
  OAI21_X1 U6945 ( .B1(n6169), .B2(n7023), .A(n6168), .ZN(U3006) );
  NAND2_X1 U6946 ( .A1(n6170), .A2(n6936), .ZN(n6175) );
  NOR2_X1 U6947 ( .A1(n6940), .A2(n6171), .ZN(n6172) );
  AOI211_X1 U6948 ( .C1(n6932), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6173), 
        .B(n6172), .ZN(n6174) );
  OAI211_X1 U6949 ( .C1(n6914), .C2(n6176), .A(n6175), .B(n6174), .ZN(U2974)
         );
  XNOR2_X1 U6950 ( .A(n6177), .B(n6178), .ZN(n6977) );
  NAND2_X1 U6951 ( .A1(n6977), .A2(n6936), .ZN(n6183) );
  NAND2_X1 U6952 ( .A1(n7059), .A2(REIP_REG_13__SCAN_IN), .ZN(n6968) );
  OAI21_X1 U6953 ( .B1(n6906), .B2(n6179), .A(n6968), .ZN(n6180) );
  AOI21_X1 U6954 ( .B1(n6901), .B2(n6181), .A(n6180), .ZN(n6182) );
  OAI211_X1 U6955 ( .C1(n6184), .C2(n6914), .A(n6183), .B(n6182), .ZN(U2973)
         );
  INV_X1 U6956 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6781) );
  OAI222_X1 U6957 ( .A1(n6311), .A2(n6781), .B1(n6219), .B2(n6185), .C1(n7352), 
        .C2(n6184), .ZN(U2878) );
  OAI21_X1 U6958 ( .B1(n6186), .B2(n6189), .A(n6188), .ZN(n6208) );
  XNOR2_X1 U6959 ( .A(n6190), .B(n6214), .ZN(n6986) );
  AOI22_X1 U6960 ( .A1(n6986), .A2(n6868), .B1(EBX_REG_14__SCAN_IN), .B2(n6475), .ZN(n6191) );
  OAI21_X1 U6961 ( .B1(n6208), .B2(n6478), .A(n6191), .ZN(U2845) );
  NAND2_X1 U6962 ( .A1(n7228), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6192)
         );
  OAI211_X1 U6963 ( .C1(n7239), .C2(n6204), .A(n6192), .B(n7105), .ZN(n6199)
         );
  NAND3_X1 U6964 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        n6193), .ZN(n6197) );
  NOR3_X1 U6965 ( .A1(n6421), .A2(n6195), .A3(n6194), .ZN(n6408) );
  NOR2_X1 U6966 ( .A1(n6407), .A2(n6408), .ZN(n7153) );
  AOI22_X1 U6967 ( .A1(EBX_REG_14__SCAN_IN), .A2(n7227), .B1(
        REIP_REG_14__SCAN_IN), .B2(n7153), .ZN(n6196) );
  OAI21_X1 U6968 ( .B1(REIP_REG_14__SCAN_IN), .B2(n6197), .A(n6196), .ZN(n6198) );
  AOI211_X1 U6969 ( .C1(n7235), .C2(n6986), .A(n6199), .B(n6198), .ZN(n6200)
         );
  OAI21_X1 U6970 ( .B1(n6208), .B2(n7196), .A(n6200), .ZN(U2813) );
  NOR2_X1 U6971 ( .A1(n3688), .A2(n6202), .ZN(n6203) );
  XNOR2_X1 U6972 ( .A(n6201), .B(n6203), .ZN(n6988) );
  NAND2_X1 U6973 ( .A1(n6988), .A2(n6936), .ZN(n6207) );
  AND2_X1 U6974 ( .A1(n7183), .A2(REIP_REG_14__SCAN_IN), .ZN(n6985) );
  NOR2_X1 U6975 ( .A1(n6940), .A2(n6204), .ZN(n6205) );
  AOI211_X1 U6976 ( .C1(n6932), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6985), 
        .B(n6205), .ZN(n6206) );
  OAI211_X1 U6977 ( .C1(n6914), .C2(n6208), .A(n6207), .B(n6206), .ZN(U2972)
         );
  INV_X1 U6978 ( .A(DATAI_14_), .ZN(n6209) );
  OAI222_X1 U6979 ( .A1(n6219), .A2(n6209), .B1(n6311), .B2(n4443), .C1(n7352), 
        .C2(n6208), .ZN(U2877) );
  NAND2_X1 U6980 ( .A1(n6188), .A2(n6211), .ZN(n6212) );
  AND2_X1 U6981 ( .A1(n6210), .A2(n6212), .ZN(n7145) );
  INV_X1 U6982 ( .A(n7145), .ZN(n6218) );
  INV_X1 U6983 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6217) );
  AOI21_X1 U6984 ( .B1(n6215), .B2(n6214), .A(n6213), .ZN(n6216) );
  OR2_X1 U6985 ( .A1(n6216), .A2(n6472), .ZN(n7143) );
  OAI222_X1 U6986 ( .A1(n6218), .A2(n6468), .B1(n6217), .B2(n6880), .C1(n6876), 
        .C2(n7143), .ZN(U2844) );
  INV_X1 U6987 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6785) );
  OAI222_X1 U6988 ( .A1(n6220), .A2(n6219), .B1(n6311), .B2(n6785), .C1(n7352), 
        .C2(n6218), .ZN(U2876) );
  INV_X1 U6989 ( .A(n6221), .ZN(n6224) );
  NOR3_X1 U6990 ( .A1(n6222), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n3650), 
        .ZN(n6506) );
  NAND2_X1 U6991 ( .A1(n7059), .A2(REIP_REG_28__SCAN_IN), .ZN(n6594) );
  OAI21_X1 U6992 ( .B1(n6906), .B2(n6225), .A(n6594), .ZN(n6228) );
  NAND2_X2 U6993 ( .A1(n6339), .A2(n3681), .ZN(n6244) );
  NOR2_X1 U6994 ( .A1(n6244), .A2(n6914), .ZN(n6227) );
  AOI211_X2 U6995 ( .C1(n6901), .C2(n6237), .A(n6228), .B(n6227), .ZN(n6229)
         );
  OAI21_X1 U6996 ( .B1(n6601), .B2(n7241), .A(n6229), .ZN(U2958) );
  NOR2_X1 U6997 ( .A1(n6355), .A2(n6230), .ZN(n6231) );
  OR2_X1 U6998 ( .A1(n6345), .A2(n6231), .ZN(n6592) );
  AND2_X1 U6999 ( .A1(n6311), .A2(n3985), .ZN(n7512) );
  AOI22_X1 U7000 ( .A1(n7512), .A2(DATAI_28_), .B1(n7515), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6236) );
  AND2_X1 U7001 ( .A1(n3981), .A2(n6233), .ZN(n6234) );
  NAND2_X1 U7002 ( .A1(n7516), .A2(DATAI_12_), .ZN(n6235) );
  OAI211_X1 U7003 ( .C1(n6244), .C2(n7352), .A(n6236), .B(n6235), .ZN(U2863)
         );
  AOI22_X1 U7004 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n7228), .B1(n7199), 
        .B2(n6237), .ZN(n6239) );
  NAND2_X1 U7005 ( .A1(n7227), .A2(EBX_REG_28__SCAN_IN), .ZN(n6238) );
  OAI211_X1 U7006 ( .C1(n6342), .C2(n6829), .A(n6239), .B(n6238), .ZN(n6241)
         );
  NOR2_X1 U7007 ( .A1(n6592), .A2(n7195), .ZN(n6240) );
  AOI211_X1 U7008 ( .C1(n6242), .C2(n6829), .A(n6241), .B(n6240), .ZN(n6243)
         );
  OAI21_X1 U7009 ( .B1(n6244), .B2(n7196), .A(n6243), .ZN(U2799) );
  AOI21_X1 U7010 ( .B1(n7257), .B2(n7294), .A(n7244), .ZN(n6248) );
  AOI22_X1 U7011 ( .A1(n3739), .A2(n6688), .B1(n6245), .B2(n3781), .ZN(n7255)
         );
  OAI21_X1 U7012 ( .B1(n7255), .B2(STATE2_REG_3__SCAN_IN), .A(n7296), .ZN(
        n6246) );
  AOI22_X1 U7013 ( .A1(n6246), .A2(n6261), .B1(n6689), .B2(n3781), .ZN(n6247)
         );
  OAI22_X1 U7014 ( .A1(n6248), .A2(n3781), .B1(n7244), .B2(n6247), .ZN(U3461)
         );
  OR2_X1 U7015 ( .A1(n5114), .A2(n7330), .ZN(n6249) );
  NOR2_X1 U7016 ( .A1(n3654), .A2(n6249), .ZN(n7432) );
  AOI21_X1 U7017 ( .B1(n3654), .B2(n6249), .A(n7432), .ZN(n6250) );
  OAI222_X1 U7018 ( .A1(n7328), .A2(n6251), .B1(n7325), .B2(n6250), .C1(n5163), 
        .C2(n7320), .ZN(U3463) );
  INV_X1 U7019 ( .A(n6252), .ZN(n6253) );
  AOI21_X1 U7020 ( .B1(n6689), .B2(n6253), .A(n7244), .ZN(n6267) );
  INV_X1 U7021 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6266) );
  INV_X1 U7022 ( .A(n5163), .ZN(n7075) );
  XNOR2_X1 U7023 ( .A(n6252), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6258)
         );
  INV_X1 U7024 ( .A(n6254), .ZN(n6318) );
  NAND2_X1 U7025 ( .A1(n6318), .A2(n6319), .ZN(n6674) );
  NAND2_X1 U7026 ( .A1(n6674), .A2(n6258), .ZN(n6257) );
  NAND2_X1 U7027 ( .A1(n7257), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6255) );
  MUX2_X1 U7028 ( .A(n6675), .B(n6255), .S(n6266), .Z(n6256) );
  OAI211_X1 U7029 ( .C1(n6680), .C2(n6258), .A(n6257), .B(n6256), .ZN(n6259)
         );
  AOI21_X1 U7030 ( .B1(n7075), .B2(n6688), .A(n6259), .ZN(n7263) );
  INV_X1 U7031 ( .A(n7263), .ZN(n6264) );
  NAND3_X1 U7032 ( .A1(n6252), .A2(n6689), .A3(n6266), .ZN(n6260) );
  OAI21_X1 U7033 ( .B1(n6262), .B2(n6261), .A(n6260), .ZN(n6263) );
  AOI21_X1 U7034 ( .B1(n6264), .B2(n7294), .A(n6263), .ZN(n6265) );
  OAI22_X1 U7035 ( .A1(n6267), .A2(n6266), .B1(n7244), .B2(n6265), .ZN(U3459)
         );
  NAND2_X1 U7036 ( .A1(n6268), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6272)
         );
  OAI22_X1 U7037 ( .A1(n6276), .A2(n6304), .B1(n6297), .B2(n6305), .ZN(n6269)
         );
  AOI21_X1 U7038 ( .B1(n6718), .B2(n6270), .A(n6269), .ZN(n6271) );
  OAI211_X1 U7039 ( .C1(n6273), .C2(n6719), .A(n6272), .B(n6271), .ZN(U3145)
         );
  NAND2_X1 U7040 ( .A1(n6274), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6279)
         );
  INV_X1 U7041 ( .A(n6304), .ZN(n7575) );
  OAI22_X1 U7042 ( .A1(n6276), .A2(n6297), .B1(n6275), .B2(n7578), .ZN(n6277)
         );
  AOI21_X1 U7043 ( .B1(n7575), .B2(n7599), .A(n6277), .ZN(n6278) );
  OAI211_X1 U7044 ( .C1(n6280), .C2(n6719), .A(n6279), .B(n6278), .ZN(U3137)
         );
  NAND2_X1 U7045 ( .A1(n6281), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6286) );
  OAI22_X1 U7046 ( .A1(n6283), .A2(n6304), .B1(n6282), .B2(n7578), .ZN(n6284)
         );
  AOI21_X1 U7047 ( .B1(n7574), .B2(n3771), .A(n6284), .ZN(n6285) );
  OAI211_X1 U7048 ( .C1(n6287), .C2(n6719), .A(n6286), .B(n6285), .ZN(U3089)
         );
  NAND2_X1 U7049 ( .A1(n6288), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6293) );
  OAI22_X1 U7050 ( .A1(n6290), .A2(n6304), .B1(n6289), .B2(n7578), .ZN(n6291)
         );
  AOI21_X1 U7051 ( .B1(n7622), .B2(n7574), .A(n6291), .ZN(n6292) );
  OAI211_X1 U7052 ( .C1(n6294), .C2(n6719), .A(n6293), .B(n6292), .ZN(U3073)
         );
  NAND2_X1 U7053 ( .A1(n6295), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6300) );
  OAI22_X1 U7054 ( .A1(n7422), .A2(n6297), .B1(n6296), .B2(n7578), .ZN(n6298)
         );
  AOI21_X1 U7055 ( .B1(n7575), .B2(n7637), .A(n6298), .ZN(n6299) );
  OAI211_X1 U7056 ( .C1(n6301), .C2(n6719), .A(n6300), .B(n6299), .ZN(U3057)
         );
  NAND2_X1 U7057 ( .A1(n6302), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6308) );
  OAI22_X1 U7058 ( .A1(n6305), .A2(n6304), .B1(n6303), .B2(n7578), .ZN(n6306)
         );
  AOI21_X1 U7059 ( .B1(n7647), .B2(n7574), .A(n6306), .ZN(n6307) );
  OAI211_X1 U7060 ( .C1(n6309), .C2(n6719), .A(n6308), .B(n6307), .ZN(U3025)
         );
  AND2_X1 U7061 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  NAND2_X1 U7062 ( .A1(n6313), .A2(n6312), .ZN(n6315) );
  AOI22_X1 U7063 ( .A1(n7512), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7515), .ZN(n6314) );
  NAND2_X1 U7064 ( .A1(n6315), .A2(n6314), .ZN(U2860) );
  XNOR2_X1 U7065 ( .A(n5114), .B(n7330), .ZN(n6316) );
  OAI222_X1 U7066 ( .A1(n6316), .A2(n7325), .B1(n5073), .B2(n7320), .C1(n7448), 
        .C2(n7328), .ZN(U3464) );
  INV_X1 U7067 ( .A(n6317), .ZN(n6324) );
  OR2_X1 U7068 ( .A1(n6325), .A2(n6318), .ZN(n6322) );
  NAND3_X1 U7069 ( .A1(n7273), .A2(n4798), .A3(n6319), .ZN(n6320) );
  NAND2_X1 U7070 ( .A1(n6325), .A2(n6320), .ZN(n6321) );
  OAI211_X1 U7071 ( .C1(n6324), .C2(n6323), .A(n6322), .B(n6321), .ZN(n7276)
         );
  INV_X1 U7072 ( .A(n6325), .ZN(n6329) );
  OAI22_X1 U7073 ( .A1(n6329), .A2(n6328), .B1(n6327), .B2(n6326), .ZN(n6941)
         );
  AOI21_X1 U7074 ( .B1(n6330), .B2(n6950), .A(READY_N), .ZN(n6957) );
  NOR2_X1 U7075 ( .A1(n6941), .A2(n6957), .ZN(n7272) );
  NOR2_X1 U7076 ( .A1(n7272), .A2(n7318), .ZN(n7243) );
  MUX2_X1 U7077 ( .A(MORE_REG_SCAN_IN), .B(n7276), .S(n7243), .Z(U3471) );
  NAND2_X1 U7078 ( .A1(n6479), .A2(n7236), .ZN(n6338) );
  AOI22_X1 U7079 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n7228), .B1(n7199), 
        .B2(n6331), .ZN(n6332) );
  OAI21_X1 U7080 ( .B1(n6333), .B2(n7203), .A(n6332), .ZN(n6335) );
  NOR3_X1 U7081 ( .A1(n6350), .A2(REIP_REG_30__SCAN_IN), .A3(n6831), .ZN(n6334) );
  AOI211_X1 U7082 ( .C1(REIP_REG_30__SCAN_IN), .C2(n6336), .A(n6335), .B(n6334), .ZN(n6337) );
  OAI211_X1 U7083 ( .C1(n6574), .C2(n7195), .A(n6338), .B(n6337), .ZN(U2797)
         );
  NAND2_X1 U7084 ( .A1(n6504), .A2(n7236), .ZN(n6349) );
  INV_X1 U7085 ( .A(n6342), .ZN(n6348) );
  INV_X1 U7086 ( .A(n6502), .ZN(n6343) );
  AOI22_X1 U7087 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n7228), .B1(n7199), 
        .B2(n6343), .ZN(n6344) );
  OAI21_X1 U7088 ( .B1(n7203), .B2(n6428), .A(n6344), .ZN(n6347) );
  AOI21_X1 U7089 ( .B1(n6353), .B2(n6351), .A(n6352), .ZN(n6512) );
  INV_X1 U7090 ( .A(n6512), .ZN(n6488) );
  AND2_X1 U7091 ( .A1(n3717), .A2(n6354), .ZN(n6356) );
  OR2_X1 U7092 ( .A1(n6356), .A2(n6355), .ZN(n6605) );
  OAI22_X1 U7093 ( .A1(n6357), .A2(n7215), .B1(n7239), .B2(n6510), .ZN(n6358)
         );
  AOI21_X1 U7094 ( .B1(n7227), .B2(EBX_REG_27__SCAN_IN), .A(n6358), .ZN(n6360)
         );
  NAND2_X1 U7095 ( .A1(n6373), .A2(REIP_REG_27__SCAN_IN), .ZN(n6359) );
  OAI211_X1 U7096 ( .C1(n6605), .C2(n7195), .A(n6360), .B(n6359), .ZN(n6361)
         );
  INV_X1 U7097 ( .A(n6361), .ZN(n6363) );
  NAND3_X1 U7098 ( .A1(n6372), .A2(REIP_REG_26__SCAN_IN), .A3(n6828), .ZN(
        n6362) );
  OAI211_X1 U7099 ( .C1(n6488), .C2(n7196), .A(n6363), .B(n6362), .ZN(U2800)
         );
  NAND2_X1 U7100 ( .A1(n6365), .A2(n6366), .ZN(n6367) );
  NAND2_X1 U7101 ( .A1(n3682), .A2(n6368), .ZN(n6369) );
  NAND2_X1 U7102 ( .A1(n3717), .A2(n6369), .ZN(n6617) );
  OAI22_X1 U7103 ( .A1(n6517), .A2(n7215), .B1(n6370), .B2(n7203), .ZN(n6371)
         );
  AOI21_X1 U7104 ( .B1(n7199), .B2(n6515), .A(n6371), .ZN(n6376) );
  OR2_X1 U7105 ( .A1(n6372), .A2(REIP_REG_26__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U7106 ( .A1(n6374), .A2(n6373), .ZN(n6375) );
  OAI211_X1 U7107 ( .C1(n6617), .C2(n7195), .A(n6376), .B(n6375), .ZN(n6377)
         );
  AOI21_X1 U7108 ( .B1(n7514), .B2(n7236), .A(n6377), .ZN(n6378) );
  INV_X1 U7109 ( .A(n6378), .ZN(U2801) );
  NOR2_X1 U7110 ( .A1(n6380), .A2(n6381), .ZN(n6382) );
  OR2_X1 U7111 ( .A1(n6379), .A2(n6382), .ZN(n6520) );
  NOR2_X1 U7112 ( .A1(n6437), .A2(n7195), .ZN(n6387) );
  NOR2_X1 U7113 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7226), .ZN(n6386) );
  INV_X1 U7114 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6438) );
  OAI22_X1 U7115 ( .A1(n7225), .A2(n7224), .B1(n6438), .B2(n7203), .ZN(n6385)
         );
  OAI22_X1 U7116 ( .A1(n6383), .A2(n7215), .B1(n7239), .B2(n6523), .ZN(n6384)
         );
  NOR4_X1 U7117 ( .A1(n6387), .A2(n6386), .A3(n6385), .A4(n6384), .ZN(n6388)
         );
  OAI21_X1 U7118 ( .B1(n6520), .B2(n7196), .A(n6388), .ZN(U2803) );
  NAND2_X1 U7119 ( .A1(n6391), .A2(n6392), .ZN(n6393) );
  NAND2_X1 U7120 ( .A1(n6389), .A2(n6393), .ZN(n7362) );
  NAND2_X1 U7121 ( .A1(n4892), .A2(n6394), .ZN(n6395) );
  NAND2_X1 U7122 ( .A1(n6442), .A2(n6395), .ZN(n6632) );
  INV_X1 U7123 ( .A(n6632), .ZN(n6402) );
  INV_X1 U7124 ( .A(n6542), .ZN(n6400) );
  INV_X1 U7125 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U7126 ( .A1(n7178), .A2(n6816), .ZN(n7207) );
  AOI21_X1 U7127 ( .B1(n7189), .B2(n7207), .A(n6819), .ZN(n6398) );
  INV_X1 U7128 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6445) );
  OAI22_X1 U7129 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6396), .B1(n6445), .B2(
        n7203), .ZN(n6397) );
  AOI211_X1 U7130 ( .C1(n7228), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n6398), 
        .B(n6397), .ZN(n6399) );
  OAI21_X1 U7131 ( .B1(n6400), .B2(n7239), .A(n6399), .ZN(n6401) );
  AOI21_X1 U7132 ( .B1(n6402), .B2(n7235), .A(n6401), .ZN(n6403) );
  OAI21_X1 U7133 ( .B1(n7362), .B2(n7196), .A(n6403), .ZN(U2805) );
  OAI21_X1 U7134 ( .B1(n6404), .B2(n6406), .A(n6405), .ZN(n6553) );
  INV_X1 U7135 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7164) );
  INV_X1 U7136 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7166) );
  INV_X1 U7137 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6809) );
  NOR3_X1 U7138 ( .A1(n7164), .A2(n7166), .A3(n6809), .ZN(n6409) );
  AOI21_X1 U7139 ( .B1(n6409), .B2(n6408), .A(n6407), .ZN(n7174) );
  INV_X1 U7140 ( .A(n6410), .ZN(n6459) );
  INV_X1 U7141 ( .A(n6556), .ZN(n6411) );
  OR2_X1 U7142 ( .A1(n7239), .A2(n6411), .ZN(n6412) );
  OAI211_X1 U7143 ( .C1(n7215), .C2(n4528), .A(n6412), .B(n7105), .ZN(n6414)
         );
  NOR3_X1 U7144 ( .A1(n7192), .A2(REIP_REG_18__SCAN_IN), .A3(n6413), .ZN(n7175) );
  AOI211_X1 U7145 ( .C1(n7227), .C2(EBX_REG_18__SCAN_IN), .A(n6414), .B(n7175), 
        .ZN(n6415) );
  OAI21_X1 U7146 ( .B1(n7195), .B2(n6459), .A(n6415), .ZN(n6416) );
  AOI21_X1 U7147 ( .B1(REIP_REG_18__SCAN_IN), .B2(n7174), .A(n6416), .ZN(n6417) );
  OAI21_X1 U7148 ( .B1(n6553), .B2(n7196), .A(n6417), .ZN(U2809) );
  INV_X1 U7149 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6889) );
  OAI22_X1 U7150 ( .A1(n6889), .A2(n7215), .B1(n7239), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6419) );
  NOR2_X1 U7151 ( .A1(n7097), .A2(n6888), .ZN(n6418) );
  AOI211_X1 U7152 ( .C1(n6420), .C2(n7074), .A(n6419), .B(n6418), .ZN(n6425)
         );
  AOI22_X1 U7153 ( .A1(EBX_REG_1__SCAN_IN), .A2(n7227), .B1(n6421), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U7154 ( .A1(n7235), .A2(n6422), .ZN(n6423) );
  NAND2_X1 U7155 ( .A1(n7178), .A2(n6852), .ZN(n7073) );
  NAND4_X1 U7156 ( .A1(n6425), .A2(n6424), .A3(n6423), .A4(n7073), .ZN(U2826)
         );
  INV_X1 U7157 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6426) );
  OAI22_X1 U7158 ( .A1(n6427), .A2(n6876), .B1(n6880), .B2(n6426), .ZN(U2828)
         );
  OAI222_X1 U7159 ( .A1(n6485), .A2(n6468), .B1(n6428), .B2(n6880), .C1(n6876), 
        .C2(n6583), .ZN(U2830) );
  INV_X1 U7160 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6429) );
  OAI222_X1 U7161 ( .A1(n6876), .A2(n6605), .B1(n6429), .B2(n6880), .C1(n6488), 
        .C2(n6468), .ZN(U2832) );
  INV_X1 U7162 ( .A(n7514), .ZN(n6432) );
  INV_X1 U7163 ( .A(n6617), .ZN(n6430) );
  AOI22_X1 U7164 ( .A1(n6430), .A2(n6868), .B1(EBX_REG_26__SCAN_IN), .B2(n6475), .ZN(n6431) );
  OAI21_X1 U7165 ( .B1(n6432), .B2(n6478), .A(n6431), .ZN(U2833) );
  OAI21_X1 U7166 ( .B1(n6379), .B2(n6433), .A(n6365), .ZN(n6933) );
  OR2_X1 U7167 ( .A1(n4954), .A2(n6434), .ZN(n6435) );
  AND2_X1 U7168 ( .A1(n3682), .A2(n6435), .ZN(n7234) );
  AOI22_X1 U7169 ( .A1(n7234), .A2(n6868), .B1(EBX_REG_25__SCAN_IN), .B2(n6475), .ZN(n6436) );
  OAI21_X1 U7170 ( .B1(n6933), .B2(n6478), .A(n6436), .ZN(U2834) );
  OAI222_X1 U7171 ( .A1(n6468), .A2(n6520), .B1(n6880), .B2(n6438), .C1(n6437), 
        .C2(n6876), .ZN(U2835) );
  AND2_X1 U7172 ( .A1(n6389), .A2(n6439), .ZN(n6440) );
  OR2_X1 U7173 ( .A1(n6440), .A2(n6380), .ZN(n7219) );
  AOI21_X1 U7174 ( .B1(n6443), .B2(n6442), .A(n6441), .ZN(n7220) );
  AOI22_X1 U7175 ( .A1(n7220), .A2(n6868), .B1(EBX_REG_23__SCAN_IN), .B2(n6475), .ZN(n6444) );
  OAI21_X1 U7176 ( .B1(n7219), .B2(n6478), .A(n6444), .ZN(U2836) );
  OAI222_X1 U7177 ( .A1(n6632), .A2(n6876), .B1(n6880), .B2(n6445), .C1(n7362), 
        .C2(n6468), .ZN(U2837) );
  OR2_X1 U7178 ( .A1(n6447), .A2(n6448), .ZN(n6449) );
  AND2_X1 U7179 ( .A1(n6391), .A2(n6449), .ZN(n7359) );
  INV_X1 U7180 ( .A(n7359), .ZN(n6453) );
  NAND2_X1 U7181 ( .A1(n3680), .A2(n6450), .ZN(n6451) );
  AND2_X1 U7182 ( .A1(n4892), .A2(n6451), .ZN(n7210) );
  AOI22_X1 U7183 ( .A1(n7210), .A2(n6868), .B1(EBX_REG_21__SCAN_IN), .B2(n6475), .ZN(n6452) );
  OAI21_X1 U7184 ( .B1(n6453), .B2(n6478), .A(n6452), .ZN(U2838) );
  AOI21_X1 U7185 ( .B1(n6454), .B2(n3684), .A(n6447), .ZN(n6550) );
  OR2_X1 U7186 ( .A1(n6875), .A2(n6455), .ZN(n6456) );
  NAND2_X1 U7187 ( .A1(n3680), .A2(n6456), .ZN(n7194) );
  OAI22_X1 U7188 ( .A1(n7194), .A2(n6876), .B1(n7204), .B2(n6880), .ZN(n6457)
         );
  AOI21_X1 U7189 ( .B1(n6550), .B2(n6878), .A(n6457), .ZN(n6458) );
  INV_X1 U7190 ( .A(n6458), .ZN(U2839) );
  INV_X1 U7191 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6460) );
  OAI222_X1 U7192 ( .A1(n6553), .A2(n6468), .B1(n6880), .B2(n6460), .C1(n6459), 
        .C2(n6876), .ZN(U2841) );
  AND2_X1 U7193 ( .A1(n6461), .A2(n6462), .ZN(n6463) );
  NOR2_X1 U7194 ( .A1(n6404), .A2(n6463), .ZN(n7353) );
  INV_X1 U7195 ( .A(n7353), .ZN(n6469) );
  OR2_X1 U7196 ( .A1(n6474), .A2(n6464), .ZN(n6465) );
  AND2_X1 U7197 ( .A1(n6466), .A2(n6465), .ZN(n7170) );
  AOI22_X1 U7198 ( .A1(n7170), .A2(n6868), .B1(EBX_REG_17__SCAN_IN), .B2(n6475), .ZN(n6467) );
  OAI21_X1 U7199 ( .B1(n6469), .B2(n6468), .A(n6467), .ZN(U2842) );
  AOI21_X1 U7200 ( .B1(n6470), .B2(n6210), .A(n3757), .ZN(n6565) );
  INV_X1 U7201 ( .A(n6565), .ZN(n7158) );
  NOR2_X1 U7202 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  OR2_X1 U7203 ( .A1(n6474), .A2(n6473), .ZN(n7157) );
  INV_X1 U7204 ( .A(n7157), .ZN(n6476) );
  AOI22_X1 U7205 ( .A1(n6476), .A2(n6868), .B1(EBX_REG_16__SCAN_IN), .B2(n6475), .ZN(n6477) );
  OAI21_X1 U7206 ( .B1(n7158), .B2(n6478), .A(n6477), .ZN(U2843) );
  AOI22_X1 U7207 ( .A1(n7512), .A2(DATAI_30_), .B1(n7515), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U7208 ( .A1(n7516), .A2(DATAI_14_), .ZN(n6480) );
  OAI211_X1 U7209 ( .C1(n6482), .C2(n7352), .A(n6481), .B(n6480), .ZN(U2861)
         );
  AOI22_X1 U7210 ( .A1(n7512), .A2(DATAI_29_), .B1(n7515), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U7211 ( .A1(n7516), .A2(DATAI_13_), .ZN(n6483) );
  OAI211_X1 U7212 ( .C1(n6485), .C2(n7352), .A(n6484), .B(n6483), .ZN(U2862)
         );
  AOI22_X1 U7213 ( .A1(n7512), .A2(DATAI_27_), .B1(n7515), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7214 ( .A1(n7516), .A2(DATAI_11_), .ZN(n6486) );
  OAI211_X1 U7215 ( .C1(n6488), .C2(n7352), .A(n6487), .B(n6486), .ZN(U2864)
         );
  INV_X1 U7216 ( .A(n6550), .ZN(n7197) );
  AOI22_X1 U7217 ( .A1(n7512), .A2(DATAI_20_), .B1(n7515), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U7218 ( .A1(n7516), .A2(DATAI_4_), .ZN(n6489) );
  OAI211_X1 U7219 ( .C1(n7197), .C2(n7352), .A(n6490), .B(n6489), .ZN(U2871)
         );
  AOI22_X1 U7220 ( .A1(n7512), .A2(DATAI_18_), .B1(n7515), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U7221 ( .A1(n7516), .A2(DATAI_2_), .ZN(n6491) );
  OAI211_X1 U7222 ( .C1(n6553), .C2(n7352), .A(n6492), .B(n6491), .ZN(U2873)
         );
  AOI22_X1 U7223 ( .A1(n7512), .A2(DATAI_16_), .B1(n7515), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U7224 ( .A1(n7516), .A2(DATAI_0_), .ZN(n6493) );
  OAI211_X1 U7225 ( .C1(n7158), .C2(n7352), .A(n6494), .B(n6493), .ZN(U2875)
         );
  NOR2_X1 U7226 ( .A1(n6495), .A2(n6593), .ZN(n6497) );
  AOI21_X1 U7227 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n3650), .A(n6498), 
        .ZN(n6499) );
  XNOR2_X1 U7228 ( .A(n6500), .B(n6499), .ZN(n6591) );
  NOR2_X1 U7229 ( .A1(n7105), .A2(n6831), .ZN(n6588) );
  AOI21_X1 U7230 ( .B1(n6932), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6588), 
        .ZN(n6501) );
  OAI21_X1 U7231 ( .B1(n6502), .B2(n6940), .A(n6501), .ZN(n6503) );
  OAI21_X1 U7232 ( .B1(n7241), .B2(n6591), .A(n6505), .ZN(U2957) );
  OAI22_X1 U7233 ( .A1(n4997), .A2(n6506), .B1(n3650), .B2(n6612), .ZN(n6508)
         );
  XNOR2_X1 U7234 ( .A(n6508), .B(n6507), .ZN(n6609) );
  NAND2_X1 U7235 ( .A1(n7183), .A2(REIP_REG_27__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7236 ( .A1(n6932), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6509)
         );
  OAI211_X1 U7237 ( .C1(n6940), .C2(n6510), .A(n6604), .B(n6509), .ZN(n6511)
         );
  AOI21_X1 U7238 ( .B1(n6512), .B2(n6937), .A(n6511), .ZN(n6513) );
  OAI21_X1 U7239 ( .B1(n7241), .B2(n6609), .A(n6513), .ZN(U2959) );
  XNOR2_X1 U7240 ( .A(n3650), .B(n6612), .ZN(n6514) );
  XNOR2_X1 U7241 ( .A(n4229), .B(n6514), .ZN(n6620) );
  NAND2_X1 U7242 ( .A1(n6901), .A2(n6515), .ZN(n6516) );
  NAND2_X1 U7243 ( .A1(n7183), .A2(REIP_REG_26__SCAN_IN), .ZN(n6616) );
  OAI211_X1 U7244 ( .C1(n6906), .C2(n6517), .A(n6516), .B(n6616), .ZN(n6518)
         );
  AOI21_X1 U7245 ( .B1(n7514), .B2(n6937), .A(n6518), .ZN(n6519) );
  OAI21_X1 U7246 ( .B1(n7241), .B2(n6620), .A(n6519), .ZN(U2960) );
  INV_X1 U7247 ( .A(n6520), .ZN(n7466) );
  NAND2_X1 U7248 ( .A1(n6932), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6521)
         );
  OAI211_X1 U7249 ( .C1(n6523), .C2(n6940), .A(n6522), .B(n6521), .ZN(n6524)
         );
  AOI21_X1 U7250 ( .B1(n7466), .B2(n6937), .A(n6524), .ZN(n6525) );
  OAI21_X1 U7251 ( .B1(n6526), .B2(n7241), .A(n6525), .ZN(U2962) );
  NOR2_X1 U7252 ( .A1(n7105), .A2(n6527), .ZN(n6624) );
  NOR2_X1 U7253 ( .A1(n6940), .A2(n7223), .ZN(n6528) );
  AOI211_X1 U7254 ( .C1(n6932), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6624), 
        .B(n6528), .ZN(n6535) );
  NAND4_X1 U7255 ( .A1(n6530), .A2(n6647), .A3(n6529), .A4(n6644), .ZN(n6531)
         );
  NAND2_X1 U7256 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  XNOR2_X1 U7257 ( .A(n6533), .B(n6627), .ZN(n6621) );
  NAND2_X1 U7258 ( .A1(n6621), .A2(n6936), .ZN(n6534) );
  OAI211_X1 U7259 ( .C1(n7219), .C2(n6914), .A(n6535), .B(n6534), .ZN(U2963)
         );
  XNOR2_X1 U7260 ( .A(n3650), .B(n6536), .ZN(n6537) );
  XNOR2_X1 U7261 ( .A(n6538), .B(n6537), .ZN(n6637) );
  NAND2_X1 U7262 ( .A1(n7059), .A2(REIP_REG_22__SCAN_IN), .ZN(n6631) );
  OAI21_X1 U7263 ( .B1(n6906), .B2(n6539), .A(n6631), .ZN(n6541) );
  NOR2_X1 U7264 ( .A1(n7362), .A2(n6914), .ZN(n6540) );
  AOI211_X1 U7265 ( .C1(n6901), .C2(n6542), .A(n6541), .B(n6540), .ZN(n6543)
         );
  OAI21_X1 U7266 ( .B1(n6637), .B2(n7241), .A(n6543), .ZN(U2964) );
  NAND2_X1 U7267 ( .A1(n6922), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6544) );
  MUX2_X1 U7268 ( .A(n6922), .B(n6544), .S(n3650), .Z(n6546) );
  XNOR2_X1 U7269 ( .A(n6546), .B(n6545), .ZN(n6651) );
  INV_X1 U7270 ( .A(n7200), .ZN(n6548) );
  NAND2_X1 U7271 ( .A1(n6932), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6547)
         );
  NAND2_X1 U7272 ( .A1(n7059), .A2(REIP_REG_20__SCAN_IN), .ZN(n6643) );
  OAI211_X1 U7273 ( .C1(n6940), .C2(n6548), .A(n6547), .B(n6643), .ZN(n6549)
         );
  AOI21_X1 U7274 ( .B1(n6550), .B2(n6937), .A(n6549), .ZN(n6551) );
  OAI21_X1 U7275 ( .B1(n6651), .B2(n7241), .A(n6551), .ZN(U2966) );
  OAI22_X1 U7276 ( .A1(n6906), .A2(n4528), .B1(n7105), .B2(n6812), .ZN(n6555)
         );
  NOR2_X1 U7277 ( .A1(n6553), .A2(n6914), .ZN(n6554) );
  AOI211_X1 U7278 ( .C1(n6901), .C2(n6556), .A(n6555), .B(n6554), .ZN(n6557)
         );
  OAI21_X1 U7279 ( .B1(n6558), .B2(n7241), .A(n6557), .ZN(U2968) );
  NAND2_X1 U7280 ( .A1(n3778), .A2(n6560), .ZN(n6561) );
  XNOR2_X1 U7281 ( .A(n6559), .B(n6561), .ZN(n6661) );
  NAND2_X1 U7282 ( .A1(n6932), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6562)
         );
  NAND2_X1 U7283 ( .A1(n7059), .A2(REIP_REG_16__SCAN_IN), .ZN(n6657) );
  OAI211_X1 U7284 ( .C1(n6940), .C2(n6563), .A(n6562), .B(n6657), .ZN(n6564)
         );
  AOI21_X1 U7285 ( .B1(n6565), .B2(n6937), .A(n6564), .ZN(n6566) );
  OAI21_X1 U7286 ( .B1(n7241), .B2(n6661), .A(n6566), .ZN(U2970) );
  NOR2_X1 U7287 ( .A1(n6567), .A2(n3693), .ZN(n6568) );
  XNOR2_X1 U7288 ( .A(n6569), .B(n6568), .ZN(n6669) );
  INV_X1 U7289 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U7290 ( .A1(n7059), .A2(REIP_REG_15__SCAN_IN), .ZN(n6664) );
  OAI21_X1 U7291 ( .B1(n6906), .B2(n6570), .A(n6664), .ZN(n6571) );
  AOI21_X1 U7292 ( .B1(n6901), .B2(n7146), .A(n6571), .ZN(n6573) );
  NAND2_X1 U7293 ( .A1(n7145), .A2(n6937), .ZN(n6572) );
  OAI211_X1 U7294 ( .C1(n6669), .C2(n7241), .A(n6573), .B(n6572), .ZN(U2971)
         );
  INV_X1 U7295 ( .A(n6574), .ZN(n6580) );
  INV_X1 U7296 ( .A(n6585), .ZN(n6575) );
  NAND3_X1 U7297 ( .A1(n6575), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n6578), .ZN(n6576) );
  OAI211_X1 U7298 ( .C1(n6584), .C2(n6578), .A(n6577), .B(n6576), .ZN(n6579)
         );
  AOI21_X1 U7299 ( .B1(n6580), .B2(n7065), .A(n6579), .ZN(n6581) );
  OAI21_X1 U7300 ( .B1(n6582), .B2(n7023), .A(n6581), .ZN(U2988) );
  INV_X1 U7301 ( .A(n6583), .ZN(n6589) );
  AOI21_X1 U7302 ( .B1(n6586), .B2(n6585), .A(n6584), .ZN(n6587) );
  AOI211_X1 U7303 ( .C1(n6589), .C2(n7065), .A(n6588), .B(n6587), .ZN(n6590)
         );
  OAI21_X1 U7304 ( .B1(n6591), .B2(n7023), .A(n6590), .ZN(U2989) );
  INV_X1 U7305 ( .A(n6592), .ZN(n6599) );
  NAND2_X1 U7306 ( .A1(n6593), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6596) );
  NOR2_X1 U7307 ( .A1(n6597), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6602)
         );
  OAI21_X1 U7308 ( .B1(n6607), .B2(n6602), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n6595) );
  OAI211_X1 U7309 ( .C1(n6597), .C2(n6596), .A(n6595), .B(n6594), .ZN(n6598)
         );
  AOI21_X1 U7310 ( .B1(n6599), .B2(n7065), .A(n6598), .ZN(n6600) );
  INV_X1 U7311 ( .A(n6602), .ZN(n6603) );
  OAI211_X1 U7312 ( .C1(n6605), .C2(n7029), .A(n6604), .B(n6603), .ZN(n6606)
         );
  AOI21_X1 U7313 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6607), .A(n6606), 
        .ZN(n6608) );
  OAI21_X1 U7314 ( .B1(n6609), .B2(n7023), .A(n6608), .ZN(U2991) );
  INV_X1 U7315 ( .A(n6610), .ZN(n6614) );
  INV_X1 U7316 ( .A(n7070), .ZN(n6611) );
  AOI21_X1 U7317 ( .B1(n6612), .B2(n6934), .A(n6611), .ZN(n6613) );
  NAND2_X1 U7318 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  OAI211_X1 U7319 ( .C1(n6617), .C2(n7029), .A(n6616), .B(n6615), .ZN(n6618)
         );
  AOI21_X1 U7320 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n7069), .A(n6618), 
        .ZN(n6619) );
  OAI21_X1 U7321 ( .B1(n6620), .B2(n7023), .A(n6619), .ZN(U2992) );
  NAND2_X1 U7322 ( .A1(n6621), .A2(n7066), .ZN(n6626) );
  NOR3_X1 U7323 ( .A1(n7064), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n6622), 
        .ZN(n6623) );
  AOI211_X1 U7324 ( .C1(n7220), .C2(n7065), .A(n6624), .B(n6623), .ZN(n6625)
         );
  OAI211_X1 U7325 ( .C1(n6628), .C2(n6627), .A(n6626), .B(n6625), .ZN(U2995)
         );
  INV_X1 U7326 ( .A(n6628), .ZN(n6635) );
  NOR2_X1 U7327 ( .A1(n6630), .A2(n6629), .ZN(n6634) );
  OAI21_X1 U7328 ( .B1(n6632), .B2(n7029), .A(n6631), .ZN(n6633) );
  AOI211_X1 U7329 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n6635), .A(n6634), .B(n6633), .ZN(n6636) );
  OAI21_X1 U7330 ( .B1(n6637), .B2(n7023), .A(n6636), .ZN(U2996) );
  AOI22_X1 U7331 ( .A1(n6995), .A2(n6640), .B1(n6639), .B2(n6638), .ZN(n6641)
         );
  NAND2_X1 U7332 ( .A1(n6642), .A2(n6641), .ZN(n6962) );
  OAI21_X1 U7333 ( .B1(n7194), .B2(n7029), .A(n6643), .ZN(n6649) );
  NAND2_X1 U7334 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U7335 ( .A1(n6981), .A2(n6973), .ZN(n6987) );
  NAND2_X1 U7336 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6987), .ZN(n6653) );
  NOR2_X1 U7337 ( .A1(n6655), .A2(n6653), .ZN(n7056) );
  NAND2_X1 U7338 ( .A1(n6644), .A2(n7056), .ZN(n6967) );
  INV_X1 U7339 ( .A(n6645), .ZN(n6646) );
  NOR3_X1 U7340 ( .A1(n6967), .A2(n6647), .A3(n6646), .ZN(n6648) );
  AOI211_X1 U7341 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n6962), .A(n6649), .B(n6648), .ZN(n6650) );
  OAI21_X1 U7342 ( .B1(n6651), .B2(n7023), .A(n6650), .ZN(U2998) );
  AOI21_X1 U7343 ( .B1(n6652), .B2(n6976), .A(n7009), .ZN(n6667) );
  INV_X1 U7344 ( .A(n6653), .ZN(n6663) );
  OAI21_X1 U7345 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6663), .ZN(n6654) );
  INV_X1 U7346 ( .A(n6654), .ZN(n6656) );
  NAND2_X1 U7347 ( .A1(n6656), .A2(n6655), .ZN(n6658) );
  OAI211_X1 U7348 ( .C1(n7029), .C2(n7157), .A(n6658), .B(n6657), .ZN(n6659)
         );
  AOI21_X1 U7349 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n6667), .A(n6659), 
        .ZN(n6660) );
  OAI21_X1 U7350 ( .B1(n6661), .B2(n7023), .A(n6660), .ZN(U3002) );
  NAND2_X1 U7351 ( .A1(n6663), .A2(n6662), .ZN(n6665) );
  OAI211_X1 U7352 ( .C1(n7029), .C2(n7143), .A(n6665), .B(n6664), .ZN(n6666)
         );
  AOI21_X1 U7353 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6667), .A(n6666), 
        .ZN(n6668) );
  OAI21_X1 U7354 ( .B1(n6669), .B2(n7023), .A(n6668), .ZN(U3003) );
  MUX2_X1 U7355 ( .A(n6670), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6252), 
        .Z(n6672) );
  NOR2_X1 U7356 ( .A1(n6672), .A2(n6671), .ZN(n6673) );
  NAND2_X1 U7357 ( .A1(n6674), .A2(n6673), .ZN(n6686) );
  INV_X1 U7358 ( .A(n6675), .ZN(n6684) );
  AOI21_X1 U7359 ( .B1(n6676), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n6677), 
        .ZN(n6681) );
  INV_X1 U7360 ( .A(n6677), .ZN(n6678) );
  OAI21_X1 U7361 ( .B1(n6252), .B2(n4310), .A(n6678), .ZN(n6679) );
  NOR2_X1 U7362 ( .A1(n6679), .A2(n4004), .ZN(n6690) );
  OAI22_X1 U7363 ( .A1(n6682), .A2(n6681), .B1(n6690), .B2(n6680), .ZN(n6683)
         );
  AOI21_X1 U7364 ( .B1(n6684), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n6683), 
        .ZN(n6685) );
  NAND2_X1 U7365 ( .A1(n6686), .A2(n6685), .ZN(n6687) );
  AOI21_X1 U7366 ( .B1(n3662), .B2(n6688), .A(n6687), .ZN(n7252) );
  INV_X1 U7367 ( .A(n7294), .ZN(n6691) );
  INV_X1 U7368 ( .A(n6689), .ZN(n7315) );
  OAI22_X1 U7369 ( .A1(n7252), .A2(n6691), .B1(n6690), .B2(n7315), .ZN(n6692)
         );
  MUX2_X1 U7370 ( .A(n6692), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n7244), 
        .Z(U3456) );
  NAND2_X1 U7371 ( .A1(n6729), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6699)
         );
  AOI22_X1 U7372 ( .A1(n7597), .A2(n7454), .B1(n6693), .B2(n6730), .ZN(n6698)
         );
  NAND2_X1 U7373 ( .A1(n7453), .A2(n6733), .ZN(n6697) );
  OR2_X1 U7374 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  NAND4_X1 U7375 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(U3116)
         );
  NAND2_X1 U7376 ( .A1(n6729), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6705)
         );
  AOI22_X1 U7377 ( .A1(n7597), .A2(n7484), .B1(n6700), .B2(n6730), .ZN(n6704)
         );
  NAND2_X1 U7378 ( .A1(n7483), .A2(n6733), .ZN(n6703) );
  NAND2_X1 U7379 ( .A1(n7604), .A2(n7485), .ZN(n6702) );
  NAND4_X1 U7380 ( .A1(n6705), .A2(n6704), .A3(n6703), .A4(n6702), .ZN(U3117)
         );
  NAND2_X1 U7381 ( .A1(n6729), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6711)
         );
  AOI22_X1 U7382 ( .A1(n7597), .A2(n7507), .B1(n6706), .B2(n6730), .ZN(n6710)
         );
  NAND2_X1 U7383 ( .A1(n7506), .A2(n6733), .ZN(n6709) );
  NAND2_X1 U7384 ( .A1(n7604), .A2(n7508), .ZN(n6708) );
  NAND4_X1 U7385 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(U3118)
         );
  NAND2_X1 U7386 ( .A1(n6729), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6717)
         );
  AOI22_X1 U7387 ( .A1(n7597), .A2(n7554), .B1(n6712), .B2(n6730), .ZN(n6716)
         );
  NAND2_X1 U7388 ( .A1(n7553), .A2(n6733), .ZN(n6715) );
  NAND2_X1 U7389 ( .A1(n7604), .A2(n7555), .ZN(n6714) );
  NAND4_X1 U7390 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(U3120)
         );
  NAND2_X1 U7391 ( .A1(n6729), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6723)
         );
  AOI22_X1 U7392 ( .A1(n7597), .A2(n7574), .B1(n6718), .B2(n6730), .ZN(n6722)
         );
  NAND2_X1 U7393 ( .A1(n7573), .A2(n6733), .ZN(n6721) );
  NAND2_X1 U7394 ( .A1(n7604), .A2(n7575), .ZN(n6720) );
  NAND4_X1 U7395 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(U3121)
         );
  NAND2_X1 U7396 ( .A1(n6729), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6728)
         );
  AOI22_X1 U7397 ( .A1(n7597), .A2(n7592), .B1(n6724), .B2(n6730), .ZN(n6727)
         );
  NAND2_X1 U7398 ( .A1(n7591), .A2(n6733), .ZN(n6726) );
  NAND2_X1 U7399 ( .A1(n7604), .A2(n7593), .ZN(n6725) );
  NAND4_X1 U7400 ( .A1(n6728), .A2(n6727), .A3(n6726), .A4(n6725), .ZN(U3122)
         );
  NAND2_X1 U7401 ( .A1(n6729), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6737)
         );
  AOI22_X1 U7402 ( .A1(n7597), .A2(n7645), .B1(n6731), .B2(n6730), .ZN(n6736)
         );
  NAND2_X1 U7403 ( .A1(n7644), .A2(n6733), .ZN(n6735) );
  NAND2_X1 U7404 ( .A1(n7604), .A2(n7648), .ZN(n6734) );
  NAND4_X1 U7405 ( .A1(n6737), .A2(n6736), .A3(n6735), .A4(n6734), .ZN(U3123)
         );
  INV_X1 U7406 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6739) );
  AND2_X1 U7407 ( .A1(STATE_REG_0__SCAN_IN), .A2(n7339), .ZN(n6754) );
  NOR2_X2 U7408 ( .A1(n6947), .A2(n6754), .ZN(n7333) );
  NAND2_X1 U7409 ( .A1(n7343), .A2(n7345), .ZN(n6945) );
  AOI21_X1 U7410 ( .B1(n6738), .B2(n6945), .A(n6751), .ZN(n7329) );
  AOI21_X1 U7411 ( .B1(n6739), .B2(n6751), .A(n7329), .ZN(U3451) );
  AND2_X1 U7412 ( .A1(n6751), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  NOR2_X1 U7413 ( .A1(n7333), .A2(n6740), .ZN(U3179) );
  AND2_X1 U7414 ( .A1(n6751), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  INV_X1 U7415 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6741) );
  NOR2_X1 U7416 ( .A1(n7333), .A2(n6741), .ZN(U3177) );
  NOR2_X1 U7417 ( .A1(n7333), .A2(n6742), .ZN(U3176) );
  INV_X1 U7418 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6743) );
  NOR2_X1 U7419 ( .A1(n7333), .A2(n6743), .ZN(U3175) );
  AND2_X1 U7420 ( .A1(n6751), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  INV_X1 U7421 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6744) );
  NOR2_X1 U7422 ( .A1(n7333), .A2(n6744), .ZN(U3173) );
  INV_X1 U7423 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6745) );
  NOR2_X1 U7424 ( .A1(n7333), .A2(n6745), .ZN(U3172) );
  NOR2_X1 U7425 ( .A1(n7333), .A2(n6746), .ZN(U3171) );
  AND2_X1 U7426 ( .A1(n6751), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  NOR2_X1 U7427 ( .A1(n7333), .A2(n6747), .ZN(U3169) );
  NOR2_X1 U7428 ( .A1(n7333), .A2(n6748), .ZN(U3168) );
  INV_X1 U7429 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6749) );
  NOR2_X1 U7430 ( .A1(n7333), .A2(n6749), .ZN(U3167) );
  AND2_X1 U7431 ( .A1(n6751), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  AND2_X1 U7432 ( .A1(n6751), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  AND2_X1 U7433 ( .A1(n6751), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  AND2_X1 U7434 ( .A1(n6751), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U7435 ( .A1(n6751), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U7436 ( .A1(n6751), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  AND2_X1 U7437 ( .A1(n6751), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  NOR2_X1 U7438 ( .A1(n7333), .A2(n6750), .ZN(U3159) );
  AND2_X1 U7439 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6751), .ZN(U3158) );
  AND2_X1 U7440 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6751), .ZN(U3157) );
  AND2_X1 U7441 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6751), .ZN(U3156) );
  AND2_X1 U7442 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6751), .ZN(U3155) );
  AND2_X1 U7443 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6751), .ZN(U3154) );
  AND2_X1 U7444 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6751), .ZN(U3153) );
  AND2_X1 U7445 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6751), .ZN(U3152) );
  AND2_X1 U7446 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6751), .ZN(U3151) );
  INV_X1 U7447 ( .A(n7328), .ZN(n6752) );
  AND2_X1 U7448 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6752), .ZN(U3019)
         );
  AND2_X1 U7449 ( .A1(n6767), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U7450 ( .B1(n6754), .B2(n6753), .A(n6947), .ZN(U2789) );
  AOI22_X1 U7451 ( .A1(n7285), .A2(LWORD_REG_0__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6756) );
  OAI21_X1 U7452 ( .B1(n6757), .B2(n6784), .A(n6756), .ZN(U2923) );
  AOI22_X1 U7453 ( .A1(n7285), .A2(LWORD_REG_1__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6758) );
  OAI21_X1 U7454 ( .B1(n6759), .B2(n6784), .A(n6758), .ZN(U2922) );
  AOI22_X1 U7455 ( .A1(n7285), .A2(LWORD_REG_2__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6760) );
  OAI21_X1 U7456 ( .B1(n6761), .B2(n6784), .A(n6760), .ZN(U2921) );
  AOI22_X1 U7457 ( .A1(n7285), .A2(LWORD_REG_3__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6762) );
  OAI21_X1 U7458 ( .B1(n6763), .B2(n6784), .A(n6762), .ZN(U2920) );
  AOI22_X1 U7459 ( .A1(n7285), .A2(LWORD_REG_4__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6764) );
  OAI21_X1 U7460 ( .B1(n6765), .B2(n6784), .A(n6764), .ZN(U2919) );
  AOI22_X1 U7461 ( .A1(n7285), .A2(LWORD_REG_5__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6766) );
  OAI21_X1 U7462 ( .B1(n4330), .B2(n6784), .A(n6766), .ZN(U2918) );
  AOI22_X1 U7463 ( .A1(n7285), .A2(LWORD_REG_6__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6768) );
  OAI21_X1 U7464 ( .B1(n4345), .B2(n6784), .A(n6768), .ZN(U2917) );
  AOI22_X1 U7465 ( .A1(n7285), .A2(LWORD_REG_7__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6769) );
  OAI21_X1 U7466 ( .B1(n4337), .B2(n6784), .A(n6769), .ZN(U2916) );
  AOI22_X1 U7467 ( .A1(n7285), .A2(LWORD_REG_8__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6770) );
  OAI21_X1 U7468 ( .B1(n6771), .B2(n6784), .A(n6770), .ZN(U2915) );
  AOI22_X1 U7469 ( .A1(n7285), .A2(LWORD_REG_9__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6772) );
  OAI21_X1 U7470 ( .B1(n6773), .B2(n6784), .A(n6772), .ZN(U2914) );
  AOI22_X1 U7471 ( .A1(n7285), .A2(LWORD_REG_10__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6774) );
  OAI21_X1 U7472 ( .B1(n6775), .B2(n6784), .A(n6774), .ZN(U2913) );
  AOI22_X1 U7473 ( .A1(n7285), .A2(LWORD_REG_11__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6776) );
  OAI21_X1 U7474 ( .B1(n6777), .B2(n6784), .A(n6776), .ZN(U2912) );
  AOI22_X1 U7475 ( .A1(n7285), .A2(LWORD_REG_12__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6778) );
  OAI21_X1 U7476 ( .B1(n6779), .B2(n6784), .A(n6778), .ZN(U2911) );
  AOI22_X1 U7477 ( .A1(n7285), .A2(LWORD_REG_13__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6780) );
  OAI21_X1 U7478 ( .B1(n6781), .B2(n6784), .A(n6780), .ZN(U2910) );
  AOI22_X1 U7479 ( .A1(n7285), .A2(LWORD_REG_14__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6782) );
  OAI21_X1 U7480 ( .B1(n4443), .B2(n6784), .A(n6782), .ZN(U2909) );
  AOI22_X1 U7481 ( .A1(n7285), .A2(LWORD_REG_15__SCAN_IN), .B1(n6767), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6783) );
  OAI21_X1 U7482 ( .B1(n6785), .B2(n6784), .A(n6783), .ZN(U2908) );
  NAND2_X1 U7483 ( .A1(n6947), .A2(n7343), .ZN(n6837) );
  INV_X1 U7484 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U7485 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6947), .ZN(n6825) );
  CLKBUF_X1 U7486 ( .A(n6825), .Z(n6833) );
  OAI222_X1 U7487 ( .A1(n6837), .A2(n6994), .B1(n6786), .B2(n6947), .C1(n6852), 
        .C2(n6833), .ZN(U3184) );
  INV_X1 U7488 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6788) );
  OAI222_X1 U7489 ( .A1(n6837), .A2(n6788), .B1(n6787), .B2(n6947), .C1(n6994), 
        .C2(n6833), .ZN(U3185) );
  INV_X1 U7490 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6789) );
  OAI222_X1 U7491 ( .A1(n6837), .A2(n7086), .B1(n6789), .B2(n6947), .C1(n6788), 
        .C2(n6833), .ZN(U3186) );
  OAI222_X1 U7492 ( .A1(n6837), .A2(n6791), .B1(n6790), .B2(n6947), .C1(n7086), 
        .C2(n6833), .ZN(U3187) );
  OAI222_X1 U7493 ( .A1(n6837), .A2(n5438), .B1(n6792), .B2(n6947), .C1(n6791), 
        .C2(n6833), .ZN(U3188) );
  INV_X1 U7494 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7135) );
  OAI222_X1 U7495 ( .A1(n6837), .A2(n7135), .B1(n6793), .B2(n6947), .C1(n5438), 
        .C2(n6833), .ZN(U3189) );
  OAI222_X1 U7496 ( .A1(n6826), .A2(n6795), .B1(n6794), .B2(n6947), .C1(n7135), 
        .C2(n6833), .ZN(U3190) );
  OAI222_X1 U7497 ( .A1(n6826), .A2(n6797), .B1(n6796), .B2(n6947), .C1(n6795), 
        .C2(n6825), .ZN(U3191) );
  INV_X1 U7498 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6798) );
  OAI222_X1 U7499 ( .A1(n6826), .A2(n7027), .B1(n6798), .B2(n6947), .C1(n6797), 
        .C2(n6833), .ZN(U3192) );
  INV_X1 U7500 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6801) );
  INV_X1 U7501 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6799) );
  OAI222_X1 U7502 ( .A1(n6826), .A2(n6801), .B1(n6799), .B2(n6947), .C1(n7027), 
        .C2(n6833), .ZN(U3193) );
  INV_X1 U7503 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6800) );
  OAI222_X1 U7504 ( .A1(n6825), .A2(n6801), .B1(n6800), .B2(n6947), .C1(n6803), 
        .C2(n6826), .ZN(U3194) );
  INV_X1 U7505 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6802) );
  INV_X1 U7506 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6804) );
  OAI222_X1 U7507 ( .A1(n6825), .A2(n6803), .B1(n6802), .B2(n6947), .C1(n6804), 
        .C2(n6826), .ZN(U3195) );
  INV_X1 U7508 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6807) );
  OAI222_X1 U7509 ( .A1(n6826), .A2(n6807), .B1(n6805), .B2(n6947), .C1(n6804), 
        .C2(n6833), .ZN(U3196) );
  INV_X1 U7510 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6806) );
  OAI222_X1 U7511 ( .A1(n6825), .A2(n6807), .B1(n6806), .B2(n6947), .C1(n6809), 
        .C2(n6826), .ZN(U3197) );
  OAI222_X1 U7512 ( .A1(n6825), .A2(n6809), .B1(n6808), .B2(n6947), .C1(n7166), 
        .C2(n6826), .ZN(U3198) );
  OAI222_X1 U7513 ( .A1(n6825), .A2(n7166), .B1(n6810), .B2(n6947), .C1(n7164), 
        .C2(n6826), .ZN(U3199) );
  OAI222_X1 U7514 ( .A1(n6825), .A2(n7164), .B1(n6811), .B2(n6947), .C1(n6812), 
        .C2(n6826), .ZN(U3200) );
  INV_X1 U7515 ( .A(REIP_REG_19__SCAN_IN), .ZN(n7176) );
  OAI222_X1 U7516 ( .A1(n6826), .A2(n7176), .B1(n6813), .B2(n6947), .C1(n6812), 
        .C2(n6833), .ZN(U3201) );
  OAI222_X1 U7517 ( .A1(n6825), .A2(n7176), .B1(n6814), .B2(n6947), .C1(n7190), 
        .C2(n6826), .ZN(U3202) );
  INV_X1 U7518 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6815) );
  OAI222_X1 U7519 ( .A1(n6837), .A2(n6816), .B1(n6815), .B2(n6947), .C1(n7190), 
        .C2(n6833), .ZN(U3203) );
  OAI222_X1 U7520 ( .A1(n6837), .A2(n6819), .B1(n6817), .B2(n6947), .C1(n6816), 
        .C2(n6833), .ZN(U3204) );
  OAI222_X1 U7521 ( .A1(n6833), .A2(n6819), .B1(n6818), .B2(n6947), .C1(n6527), 
        .C2(n6826), .ZN(U3205) );
  OAI222_X1 U7522 ( .A1(n6825), .A2(n6527), .B1(n6820), .B2(n6947), .C1(n7224), 
        .C2(n6826), .ZN(U3206) );
  OAI222_X1 U7523 ( .A1(n6837), .A2(n7232), .B1(n6821), .B2(n6947), .C1(n7224), 
        .C2(n6833), .ZN(U3207) );
  INV_X1 U7524 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6824) );
  OAI222_X1 U7525 ( .A1(n6833), .A2(n7232), .B1(n6822), .B2(n6947), .C1(n6824), 
        .C2(n6826), .ZN(U3208) );
  OAI222_X1 U7526 ( .A1(n6825), .A2(n6824), .B1(n6823), .B2(n6947), .C1(n6828), 
        .C2(n6826), .ZN(U3209) );
  INV_X1 U7527 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6827) );
  OAI222_X1 U7528 ( .A1(n6833), .A2(n6828), .B1(n6827), .B2(n6947), .C1(n6829), 
        .C2(n6826), .ZN(U3210) );
  OAI222_X1 U7529 ( .A1(n6837), .A2(n6831), .B1(n6830), .B2(n6947), .C1(n6829), 
        .C2(n6833), .ZN(U3211) );
  INV_X1 U7530 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6834) );
  OAI222_X1 U7531 ( .A1(n6837), .A2(n6834), .B1(n6832), .B2(n6947), .C1(n6831), 
        .C2(n6833), .ZN(U3212) );
  OAI222_X1 U7532 ( .A1(n6837), .A2(n6836), .B1(n6835), .B2(n6947), .C1(n6834), 
        .C2(n6833), .ZN(U3213) );
  INV_X1 U7533 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6839) );
  AOI22_X1 U7534 ( .A1(n6947), .A2(n6839), .B1(n6838), .B2(n7350), .ZN(U3445)
         );
  AOI221_X1 U7535 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), 
        .C1(REIP_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6850) );
  NOR4_X1 U7536 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n6843) );
  NOR4_X1 U7537 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6842) );
  NOR4_X1 U7538 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(
        n6841) );
  NOR4_X1 U7539 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6840) );
  NAND4_X1 U7540 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n6849)
         );
  NOR4_X1 U7541 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6847)
         );
  AOI211_X1 U7542 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_9__SCAN_IN), .B(
        DATAWIDTH_REG_11__SCAN_IN), .ZN(n6846) );
  NOR4_X1 U7543 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6845) );
  NOR4_X1 U7544 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n6844) );
  NAND4_X1 U7545 ( .A1(n6847), .A2(n6846), .A3(n6845), .A4(n6844), .ZN(n6848)
         );
  NOR2_X1 U7546 ( .A1(n6849), .A2(n6848), .ZN(n6863) );
  MUX2_X1 U7547 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n6850), .S(n6863), .Z(
        U2795) );
  INV_X1 U7548 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6855) );
  AOI22_X1 U7549 ( .A1(n6947), .A2(n6855), .B1(n6851), .B2(n7350), .ZN(U3446)
         );
  AOI21_X1 U7550 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6853) );
  OAI221_X1 U7551 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6853), .C1(n6852), .C2(
        REIP_REG_0__SCAN_IN), .A(n6863), .ZN(n6854) );
  OAI21_X1 U7552 ( .B1(n6863), .B2(n6855), .A(n6854), .ZN(U3468) );
  INV_X1 U7553 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6859) );
  INV_X1 U7554 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U7555 ( .A1(n6947), .A2(n6859), .B1(n6856), .B2(n7350), .ZN(U3447)
         );
  NOR3_X1 U7556 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n6857) );
  OAI21_X1 U7557 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6857), .A(n6863), .ZN(n6858)
         );
  OAI21_X1 U7558 ( .B1(n6863), .B2(n6859), .A(n6858), .ZN(U2794) );
  INV_X1 U7559 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6862) );
  INV_X1 U7560 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7561 ( .A1(n6947), .A2(n6862), .B1(n6860), .B2(n7350), .ZN(U3448)
         );
  OAI21_X1 U7562 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .A(
        n6863), .ZN(n6861) );
  OAI21_X1 U7563 ( .B1(n6863), .B2(n6862), .A(n6861), .ZN(U3469) );
  INV_X1 U7564 ( .A(n6915), .ZN(n7136) );
  AND2_X1 U7565 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  NOR2_X1 U7566 ( .A1(n6867), .A2(n6866), .ZN(n7129) );
  AOI22_X1 U7567 ( .A1(n7136), .A2(n6878), .B1(n6868), .B2(n7129), .ZN(n6869)
         );
  OAI21_X1 U7568 ( .B1(n6880), .B2(n7132), .A(n6869), .ZN(U2852) );
  NAND2_X1 U7569 ( .A1(n6405), .A2(n6870), .ZN(n6871) );
  AND2_X1 U7570 ( .A1(n6873), .A2(n6872), .ZN(n6874) );
  OR2_X1 U7571 ( .A1(n6875), .A2(n6874), .ZN(n7184) );
  NOR2_X1 U7572 ( .A1(n7184), .A2(n6876), .ZN(n6877) );
  AOI21_X1 U7573 ( .B1(n7356), .B2(n6878), .A(n6877), .ZN(n6879) );
  OAI21_X1 U7574 ( .B1(n6880), .B2(n7181), .A(n6879), .ZN(U2840) );
  INV_X1 U7575 ( .A(n6881), .ZN(n6883) );
  AOI21_X1 U7576 ( .B1(n6883), .B2(n6937), .A(n6882), .ZN(n6886) );
  OAI21_X1 U7577 ( .B1(n6932), .B2(n6884), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6885) );
  OAI211_X1 U7578 ( .C1(n6887), .C2(n7241), .A(n6886), .B(n6885), .ZN(U2986)
         );
  AOI22_X1 U7579 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6932), .B1(n7059), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6892) );
  INV_X1 U7580 ( .A(n6888), .ZN(n6890) );
  AOI22_X1 U7581 ( .A1(n6937), .A2(n6890), .B1(n6901), .B2(n6889), .ZN(n6891)
         );
  OAI211_X1 U7582 ( .C1(n7241), .C2(n6893), .A(n6892), .B(n6891), .ZN(U2985)
         );
  AOI22_X1 U7583 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6932), .B1(n7183), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6900) );
  NAND2_X1 U7584 ( .A1(n6895), .A2(n6894), .ZN(n6898) );
  INV_X1 U7585 ( .A(n6896), .ZN(n6897) );
  XNOR2_X1 U7586 ( .A(n6898), .B(n6897), .ZN(n7000) );
  AOI22_X1 U7587 ( .A1(n6936), .A2(n7000), .B1(n7077), .B2(n6937), .ZN(n6899)
         );
  OAI211_X1 U7588 ( .C1(n6940), .C2(n7085), .A(n6900), .B(n6899), .ZN(U2984)
         );
  INV_X1 U7589 ( .A(n7119), .ZN(n6902) );
  AOI222_X1 U7590 ( .A1(n6903), .A2(n6936), .B1(n6902), .B2(n6901), .C1(n6937), 
        .C2(n7113), .ZN(n6905) );
  OAI211_X1 U7591 ( .C1(n6906), .C2(n7106), .A(n6905), .B(n6904), .ZN(U2981)
         );
  AOI22_X1 U7592 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6932), .B1(n7059), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7593 ( .A1(n6907), .A2(n6936), .B1(n6937), .B2(n7126), .ZN(n6908)
         );
  OAI211_X1 U7594 ( .C1(n6940), .C2(n7128), .A(n6909), .B(n6908), .ZN(U2980)
         );
  AOI22_X1 U7595 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6932), .B1(n7059), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6918) );
  OR2_X1 U7596 ( .A1(n6911), .A2(n6910), .ZN(n6912) );
  AND2_X1 U7597 ( .A1(n6913), .A2(n6912), .ZN(n7016) );
  NOR2_X1 U7598 ( .A1(n6915), .A2(n6914), .ZN(n6916) );
  AOI21_X1 U7599 ( .B1(n7016), .B2(n6936), .A(n6916), .ZN(n6917) );
  OAI211_X1 U7600 ( .C1(n6940), .C2(n7141), .A(n6918), .B(n6917), .ZN(U2979)
         );
  AOI22_X1 U7601 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6932), .B1(n7059), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n6921) );
  XNOR2_X1 U7602 ( .A(n3650), .B(n7055), .ZN(n6919) );
  XNOR2_X1 U7603 ( .A(n5036), .B(n6919), .ZN(n7052) );
  AOI22_X1 U7604 ( .A1(n7052), .A2(n6936), .B1(n6937), .B2(n7353), .ZN(n6920)
         );
  OAI211_X1 U7605 ( .C1(n6940), .C2(n7173), .A(n6921), .B(n6920), .ZN(U2969)
         );
  AOI22_X1 U7606 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6932), .B1(n7059), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n6926) );
  OAI21_X1 U7607 ( .B1(n6924), .B2(n6923), .A(n6922), .ZN(n6964) );
  AOI22_X1 U7608 ( .A1(n6964), .A2(n6936), .B1(n6937), .B2(n7356), .ZN(n6925)
         );
  OAI211_X1 U7609 ( .C1(n6940), .C2(n7188), .A(n6926), .B(n6925), .ZN(U2967)
         );
  AOI22_X1 U7610 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6932), .B1(n7183), 
        .B2(REIP_REG_21__SCAN_IN), .ZN(n6931) );
  AOI21_X1 U7611 ( .B1(n6929), .B2(n6928), .A(n6927), .ZN(n7061) );
  AOI22_X1 U7612 ( .A1(n7061), .A2(n6936), .B1(n6937), .B2(n7359), .ZN(n6930)
         );
  OAI211_X1 U7613 ( .C1(n6940), .C2(n7213), .A(n6931), .B(n6930), .ZN(U2965)
         );
  AOI22_X1 U7614 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6932), .B1(n7183), 
        .B2(REIP_REG_25__SCAN_IN), .ZN(n6939) );
  INV_X1 U7615 ( .A(n6933), .ZN(n7489) );
  XNOR2_X1 U7616 ( .A(n3650), .B(n6934), .ZN(n6935) );
  XNOR2_X1 U7617 ( .A(n6222), .B(n6935), .ZN(n7067) );
  AOI22_X1 U7618 ( .A1(n7489), .A2(n6937), .B1(n6936), .B2(n7067), .ZN(n6938)
         );
  OAI211_X1 U7619 ( .C1(n6940), .C2(n7240), .A(n6939), .B(n6938), .ZN(U2961)
         );
  INV_X1 U7620 ( .A(n7314), .ZN(n6959) );
  NAND2_X1 U7621 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6959), .ZN(n6943) );
  OAI21_X1 U7622 ( .B1(n6941), .B2(n7318), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6942) );
  OAI21_X1 U7623 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6943), .A(n6942), .ZN(
        U2790) );
  INV_X1 U7624 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6944) );
  OAI222_X1 U7625 ( .A1(n6947), .A2(n6945), .B1(n6947), .B2(n6944), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(n7350), .ZN(U2791) );
  AOI22_X1 U7626 ( .A1(n6947), .A2(READREQUEST_REG_SCAN_IN), .B1(n6946), .B2(
        n7350), .ZN(U3470) );
  NAND2_X1 U7627 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7348) );
  INV_X1 U7628 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7336) );
  NOR2_X1 U7629 ( .A1(n7345), .A2(n7336), .ZN(n7338) );
  INV_X1 U7630 ( .A(HOLD), .ZN(n7341) );
  NOR2_X1 U7631 ( .A1(n7334), .A2(n7341), .ZN(n6948) );
  OAI22_X1 U7632 ( .A1(n7338), .A2(n6948), .B1(n7343), .B2(n7341), .ZN(n6949)
         );
  NAND3_X1 U7633 ( .A1(n6950), .A2(n7348), .A3(n6949), .ZN(U3182) );
  NOR2_X1 U7634 ( .A1(READY_N), .A2(n7313), .ZN(n7293) );
  OAI211_X1 U7635 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n7293), .A(n7303), .B(
        n7314), .ZN(n6951) );
  NAND2_X1 U7636 ( .A1(n6952), .A2(n6951), .ZN(U3150) );
  OAI211_X1 U7637 ( .C1(READY_N), .C2(n6955), .A(n6954), .B(n6953), .ZN(n6961)
         );
  AOI21_X1 U7638 ( .B1(n4017), .B2(n7330), .A(n7295), .ZN(n6956) );
  AOI21_X1 U7639 ( .B1(n6957), .B2(n6956), .A(n7313), .ZN(n6958) );
  OAI21_X1 U7640 ( .B1(n6959), .B2(n6958), .A(n6961), .ZN(n6960) );
  OAI21_X1 U7641 ( .B1(n6961), .B2(n7336), .A(n6960), .ZN(U3472) );
  AOI22_X1 U7642 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6962), .B1(n7059), .B2(REIP_REG_19__SCAN_IN), .ZN(n6966) );
  INV_X1 U7643 ( .A(n7184), .ZN(n6963) );
  AOI22_X1 U7644 ( .A1(n6964), .A2(n7066), .B1(n7065), .B2(n6963), .ZN(n6965)
         );
  OAI211_X1 U7645 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6967), .A(n6966), .B(n6965), .ZN(U2999) );
  NAND2_X1 U7646 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6972) );
  NOR2_X1 U7647 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6972), .ZN(n6984)
         );
  INV_X1 U7648 ( .A(n6984), .ZN(n6980) );
  INV_X1 U7649 ( .A(n6968), .ZN(n6969) );
  AOI21_X1 U7650 ( .B1(n7065), .B2(n6970), .A(n6969), .ZN(n6979) );
  AOI22_X1 U7651 ( .A1(n6974), .A2(n6973), .B1(n6972), .B2(n6971), .ZN(n6975)
         );
  OAI21_X1 U7652 ( .B1(n7009), .B2(n6976), .A(n6975), .ZN(n6982) );
  AOI22_X1 U7653 ( .A1(n6977), .A2(n7066), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6982), .ZN(n6978) );
  OAI211_X1 U7654 ( .C1(n6981), .C2(n6980), .A(n6979), .B(n6978), .ZN(U3005)
         );
  AOI21_X1 U7655 ( .B1(n6984), .B2(n6983), .A(n6982), .ZN(n6991) );
  AOI21_X1 U7656 ( .B1(n7065), .B2(n6986), .A(n6985), .ZN(n6990) );
  AOI22_X1 U7657 ( .A1(n6988), .A2(n7066), .B1(n6987), .B2(n4219), .ZN(n6989)
         );
  OAI211_X1 U7658 ( .C1(n6991), .C2(n4219), .A(n6990), .B(n6989), .ZN(U3004)
         );
  INV_X1 U7659 ( .A(n6992), .ZN(n6993) );
  NAND2_X1 U7660 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6993), .ZN(n7003)
         );
  OAI22_X1 U7661 ( .A1(n7029), .A2(n7079), .B1(n6994), .B2(n7105), .ZN(n6999)
         );
  NAND4_X1 U7662 ( .A1(n6995), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A4(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6996) );
  NAND2_X1 U7663 ( .A1(n6997), .A2(n6996), .ZN(n6998) );
  AOI211_X1 U7664 ( .C1(n7066), .C2(n7000), .A(n6999), .B(n6998), .ZN(n7001)
         );
  OAI221_X1 U7665 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n7003), .C1(n4086), .C2(n7002), .A(n7001), .ZN(U3016) );
  INV_X1 U7666 ( .A(n7004), .ZN(n7011) );
  NAND2_X1 U7667 ( .A1(n7011), .A2(n7025), .ZN(n7019) );
  OAI21_X1 U7668 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n7022), .ZN(n7015) );
  INV_X1 U7669 ( .A(n7005), .ZN(n7006) );
  AOI21_X1 U7670 ( .B1(n7065), .B2(n7007), .A(n7006), .ZN(n7014) );
  INV_X1 U7671 ( .A(n7008), .ZN(n7012) );
  AOI21_X1 U7672 ( .B1(n7011), .B2(n7010), .A(n7009), .ZN(n7020) );
  AOI22_X1 U7673 ( .A1(n7066), .A2(n7012), .B1(n7020), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n7013) );
  OAI211_X1 U7674 ( .C1(n7019), .C2(n7015), .A(n7014), .B(n7013), .ZN(U3010)
         );
  AOI22_X1 U7675 ( .A1(n7065), .A2(n7129), .B1(n7059), .B2(REIP_REG_7__SCAN_IN), .ZN(n7018) );
  AOI22_X1 U7676 ( .A1(n7020), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .B1(n7066), 
        .B2(n7016), .ZN(n7017) );
  OAI211_X1 U7677 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n7019), .A(n7018), 
        .B(n7017), .ZN(U3011) );
  AOI21_X1 U7678 ( .B1(n7022), .B2(n7021), .A(n7020), .ZN(n7039) );
  NOR2_X1 U7679 ( .A1(n7024), .A2(n7023), .ZN(n7033) );
  NAND2_X1 U7680 ( .A1(n7026), .A2(n7025), .ZN(n7041) );
  AOI221_X1 U7681 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n4215), .C2(n7040), .A(n7041), 
        .ZN(n7031) );
  OAI22_X1 U7682 ( .A1(n7029), .A2(n7028), .B1(n7027), .B2(n7105), .ZN(n7030)
         );
  AOI211_X1 U7683 ( .C1(n7033), .C2(n7032), .A(n7031), .B(n7030), .ZN(n7034)
         );
  OAI21_X1 U7684 ( .B1(n7039), .B2(n4215), .A(n7034), .ZN(U3008) );
  INV_X1 U7685 ( .A(n7035), .ZN(n7036) );
  AOI222_X1 U7686 ( .A1(REIP_REG_9__SCAN_IN), .A2(n7183), .B1(n7065), .B2(
        n7037), .C1(n7066), .C2(n7036), .ZN(n7038) );
  OAI221_X1 U7687 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n7041), .C1(n7040), .C2(n7039), .A(n7038), .ZN(U3009) );
  INV_X1 U7688 ( .A(n7042), .ZN(n7045) );
  INV_X1 U7689 ( .A(n7043), .ZN(n7044) );
  AOI21_X1 U7690 ( .B1(n7065), .B2(n7045), .A(n7044), .ZN(n7051) );
  INV_X1 U7691 ( .A(n7046), .ZN(n7048) );
  AOI22_X1 U7692 ( .A1(n7048), .A2(n7066), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n7047), .ZN(n7050) );
  NAND3_X1 U7693 ( .A1(n7051), .A2(n7050), .A3(n7049), .ZN(U3007) );
  AOI22_X1 U7694 ( .A1(n7052), .A2(n7066), .B1(n7065), .B2(n7170), .ZN(n7058)
         );
  NOR2_X1 U7695 ( .A1(n7105), .A2(n7164), .ZN(n7053) );
  AOI221_X1 U7696 ( .B1(n7056), .B2(n7055), .C1(n7054), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n7053), .ZN(n7057) );
  NAND2_X1 U7697 ( .A1(n7058), .A2(n7057), .ZN(U3001) );
  AOI22_X1 U7698 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n7060), .B1(n7059), .B2(REIP_REG_21__SCAN_IN), .ZN(n7063) );
  AOI22_X1 U7699 ( .A1(n7061), .A2(n7066), .B1(n7065), .B2(n7210), .ZN(n7062)
         );
  OAI211_X1 U7700 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n7064), .A(n7063), .B(n7062), .ZN(U2997) );
  AOI22_X1 U7701 ( .A1(n7067), .A2(n7066), .B1(n7065), .B2(n7234), .ZN(n7072)
         );
  NOR2_X1 U7702 ( .A1(n7105), .A2(n7232), .ZN(n7068) );
  AOI221_X1 U7703 ( .B1(n7070), .B2(n6934), .C1(n7069), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n7068), .ZN(n7071) );
  NAND2_X1 U7704 ( .A1(n7072), .A2(n7071), .ZN(U2993) );
  NAND2_X1 U7705 ( .A1(n7073), .A2(n7114), .ZN(n7076) );
  AOI222_X1 U7706 ( .A1(n7076), .A2(REIP_REG_2__SCAN_IN), .B1(n7227), .B2(
        EBX_REG_2__SCAN_IN), .C1(n7075), .C2(n7074), .ZN(n7084) );
  NAND2_X1 U7707 ( .A1(n7112), .A2(n7077), .ZN(n7078) );
  OAI21_X1 U7708 ( .B1(n7079), .B2(n7195), .A(n7078), .ZN(n7082) );
  NAND2_X1 U7709 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6994), .ZN(n7080) );
  OAI22_X1 U7710 ( .A1(n7192), .A2(n7080), .B1(n4303), .B2(n7215), .ZN(n7081)
         );
  NOR2_X1 U7711 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  OAI211_X1 U7712 ( .C1(n7085), .C2(n7239), .A(n7084), .B(n7083), .ZN(U2825)
         );
  INV_X1 U7713 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n7103) );
  AOI221_X1 U7714 ( .B1(n7088), .B2(REIP_REG_4__SCAN_IN), .C1(n7087), .C2(
        n7086), .A(n7183), .ZN(n7102) );
  INV_X1 U7715 ( .A(n7089), .ZN(n7090) );
  NOR2_X1 U7716 ( .A1(n7091), .A2(n7090), .ZN(n7092) );
  XNOR2_X1 U7717 ( .A(n7092), .B(n7250), .ZN(n7246) );
  INV_X1 U7718 ( .A(n7246), .ZN(n7095) );
  OAI22_X1 U7719 ( .A1(n7095), .A2(n7094), .B1(n7195), .B2(n7093), .ZN(n7100)
         );
  OAI22_X1 U7720 ( .A1(n7098), .A2(n7097), .B1(n7096), .B2(n7239), .ZN(n7099)
         );
  AOI211_X1 U7721 ( .C1(EBX_REG_4__SCAN_IN), .C2(n7227), .A(n7100), .B(n7099), 
        .ZN(n7101) );
  OAI211_X1 U7722 ( .C1(n7103), .C2(n7215), .A(n7102), .B(n7101), .ZN(U2823)
         );
  OR2_X1 U7723 ( .A1(n7203), .A2(n7104), .ZN(n7109) );
  OAI21_X1 U7724 ( .B1(n7215), .B2(n7106), .A(n7105), .ZN(n7107) );
  INV_X1 U7725 ( .A(n7107), .ZN(n7108) );
  OAI211_X1 U7726 ( .C1(n7110), .C2(n7195), .A(n7109), .B(n7108), .ZN(n7111)
         );
  AOI21_X1 U7727 ( .B1(n7113), .B2(n7112), .A(n7111), .ZN(n7118) );
  OAI21_X1 U7728 ( .B1(n7192), .B2(n7115), .A(n7114), .ZN(n7130) );
  OAI21_X1 U7729 ( .B1(REIP_REG_5__SCAN_IN), .B2(n7116), .A(n7130), .ZN(n7117)
         );
  OAI211_X1 U7730 ( .C1(n7239), .C2(n7119), .A(n7118), .B(n7117), .ZN(U2822)
         );
  NAND2_X1 U7731 ( .A1(n7130), .A2(REIP_REG_6__SCAN_IN), .ZN(n7124) );
  OAI22_X1 U7732 ( .A1(n7121), .A2(n7203), .B1(n7120), .B2(n7195), .ZN(n7122)
         );
  AOI211_X1 U7733 ( .C1(n7228), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n7183), 
        .B(n7122), .ZN(n7123) );
  OAI211_X1 U7734 ( .C1(REIP_REG_6__SCAN_IN), .C2(n7134), .A(n7124), .B(n7123), 
        .ZN(n7125) );
  AOI21_X1 U7735 ( .B1(n7126), .B2(n7236), .A(n7125), .ZN(n7127) );
  OAI21_X1 U7736 ( .B1(n7128), .B2(n7239), .A(n7127), .ZN(U2821) );
  AOI22_X1 U7737 ( .A1(n7130), .A2(REIP_REG_7__SCAN_IN), .B1(n7235), .B2(n7129), .ZN(n7131) );
  OAI21_X1 U7738 ( .B1(n7132), .B2(n7203), .A(n7131), .ZN(n7133) );
  AOI211_X1 U7739 ( .C1(n7228), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n7183), 
        .B(n7133), .ZN(n7140) );
  AOI21_X1 U7740 ( .B1(n5438), .B2(n7135), .A(n7134), .ZN(n7138) );
  AOI22_X1 U7741 ( .A1(n7138), .A2(n7137), .B1(n7136), .B2(n7236), .ZN(n7139)
         );
  OAI211_X1 U7742 ( .C1(n7141), .C2(n7239), .A(n7140), .B(n7139), .ZN(U2820)
         );
  AOI22_X1 U7743 ( .A1(EBX_REG_15__SCAN_IN), .A2(n7227), .B1(
        REIP_REG_15__SCAN_IN), .B2(n7153), .ZN(n7150) );
  NAND2_X1 U7744 ( .A1(n7178), .A2(n7142), .ZN(n7151) );
  NOR2_X1 U7745 ( .A1(REIP_REG_15__SCAN_IN), .A2(n7151), .ZN(n7154) );
  AOI211_X1 U7746 ( .C1(n7228), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n7183), 
        .B(n7154), .ZN(n7149) );
  NOR2_X1 U7747 ( .A1(n7195), .A2(n7143), .ZN(n7144) );
  AOI21_X1 U7748 ( .B1(n7145), .B2(n7236), .A(n7144), .ZN(n7148) );
  NAND2_X1 U7749 ( .A1(n7146), .A2(n7199), .ZN(n7147) );
  NAND4_X1 U7750 ( .A1(n7150), .A2(n7149), .A3(n7148), .A4(n7147), .ZN(U2812)
         );
  INV_X1 U7751 ( .A(n7151), .ZN(n7152) );
  NAND2_X1 U7752 ( .A1(n7152), .A2(REIP_REG_15__SCAN_IN), .ZN(n7165) );
  OAI21_X1 U7753 ( .B1(n7154), .B2(n7153), .A(REIP_REG_16__SCAN_IN), .ZN(n7155) );
  OAI21_X1 U7754 ( .B1(REIP_REG_16__SCAN_IN), .B2(n7165), .A(n7155), .ZN(n7156) );
  AOI211_X1 U7755 ( .C1(n7228), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n7183), 
        .B(n7156), .ZN(n7162) );
  OAI22_X1 U7756 ( .A1(n7158), .A2(n7196), .B1(n7195), .B2(n7157), .ZN(n7159)
         );
  AOI21_X1 U7757 ( .B1(n7160), .B2(n7199), .A(n7159), .ZN(n7161) );
  OAI211_X1 U7758 ( .C1(n7163), .C2(n7203), .A(n7162), .B(n7161), .ZN(U2811)
         );
  OAI21_X1 U7759 ( .B1(n7166), .B2(n7165), .A(n7164), .ZN(n7169) );
  AOI22_X1 U7760 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n7228), .B1(
        EBX_REG_17__SCAN_IN), .B2(n7227), .ZN(n7167) );
  INV_X1 U7761 ( .A(n7167), .ZN(n7168) );
  AOI211_X1 U7762 ( .C1(n7174), .C2(n7169), .A(n7183), .B(n7168), .ZN(n7172)
         );
  AOI22_X1 U7763 ( .A1(n7353), .A2(n7236), .B1(n7235), .B2(n7170), .ZN(n7171)
         );
  OAI211_X1 U7764 ( .C1(n7173), .C2(n7239), .A(n7172), .B(n7171), .ZN(U2810)
         );
  OAI21_X1 U7765 ( .B1(n7175), .B2(n7174), .A(REIP_REG_19__SCAN_IN), .ZN(n7180) );
  NAND3_X1 U7766 ( .A1(n7178), .A2(n7177), .A3(n7176), .ZN(n7179) );
  OAI211_X1 U7767 ( .C1(n7203), .C2(n7181), .A(n7180), .B(n7179), .ZN(n7182)
         );
  AOI211_X1 U7768 ( .C1(n7228), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n7183), 
        .B(n7182), .ZN(n7187) );
  NOR2_X1 U7769 ( .A1(n7184), .A2(n7195), .ZN(n7185) );
  AOI21_X1 U7770 ( .B1(n7356), .B2(n7236), .A(n7185), .ZN(n7186) );
  OAI211_X1 U7771 ( .C1(n7188), .C2(n7239), .A(n7187), .B(n7186), .ZN(U2808)
         );
  INV_X1 U7772 ( .A(n7189), .ZN(n7205) );
  OAI21_X1 U7773 ( .B1(n7192), .B2(n7191), .A(n7190), .ZN(n7193) );
  AOI22_X1 U7774 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n7228), .B1(n7205), 
        .B2(n7193), .ZN(n7202) );
  OAI22_X1 U7775 ( .A1(n7197), .A2(n7196), .B1(n7195), .B2(n7194), .ZN(n7198)
         );
  AOI21_X1 U7776 ( .B1(n7200), .B2(n7199), .A(n7198), .ZN(n7201) );
  OAI211_X1 U7777 ( .C1(n7204), .C2(n7203), .A(n7202), .B(n7201), .ZN(U2807)
         );
  AOI22_X1 U7778 ( .A1(EBX_REG_21__SCAN_IN), .A2(n7227), .B1(
        REIP_REG_21__SCAN_IN), .B2(n7205), .ZN(n7206) );
  OAI21_X1 U7779 ( .B1(n7208), .B2(n7207), .A(n7206), .ZN(n7209) );
  AOI21_X1 U7780 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n7228), .A(n7209), 
        .ZN(n7212) );
  AOI22_X1 U7781 ( .A1(n7359), .A2(n7236), .B1(n7235), .B2(n7210), .ZN(n7211)
         );
  OAI211_X1 U7782 ( .C1(n7213), .C2(n7239), .A(n7212), .B(n7211), .ZN(U2806)
         );
  NOR2_X1 U7783 ( .A1(REIP_REG_23__SCAN_IN), .A2(n7214), .ZN(n7217) );
  INV_X1 U7784 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n7216) );
  OAI22_X1 U7785 ( .A1(n7225), .A2(n7217), .B1(n7216), .B2(n7215), .ZN(n7218)
         );
  AOI21_X1 U7786 ( .B1(EBX_REG_23__SCAN_IN), .B2(n7227), .A(n7218), .ZN(n7222)
         );
  INV_X1 U7787 ( .A(n7219), .ZN(n7366) );
  AOI22_X1 U7788 ( .A1(n7366), .A2(n7236), .B1(n7235), .B2(n7220), .ZN(n7221)
         );
  OAI211_X1 U7789 ( .C1(n7223), .C2(n7239), .A(n7222), .B(n7221), .ZN(U2804)
         );
  NOR2_X1 U7790 ( .A1(n7224), .A2(n7226), .ZN(n7233) );
  OAI21_X1 U7791 ( .B1(REIP_REG_24__SCAN_IN), .B2(n7226), .A(n7225), .ZN(n7231) );
  AOI22_X1 U7792 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n7228), .B1(
        EBX_REG_25__SCAN_IN), .B2(n7227), .ZN(n7229) );
  INV_X1 U7793 ( .A(n7229), .ZN(n7230) );
  AOI221_X1 U7794 ( .B1(n7233), .B2(n7232), .C1(n7231), .C2(
        REIP_REG_25__SCAN_IN), .A(n7230), .ZN(n7238) );
  AOI22_X1 U7795 ( .A1(n7489), .A2(n7236), .B1(n7235), .B2(n7234), .ZN(n7237)
         );
  OAI211_X1 U7796 ( .C1(n7240), .C2(n7239), .A(n7238), .B(n7237), .ZN(U2802)
         );
  OAI21_X1 U7797 ( .B1(n7243), .B2(n7242), .A(n7241), .ZN(U2793) );
  INV_X1 U7798 ( .A(n7244), .ZN(n7251) );
  NAND2_X1 U7799 ( .A1(n7246), .A2(n7245), .ZN(n7275) );
  INV_X1 U7800 ( .A(n7275), .ZN(n7247) );
  NAND3_X1 U7801 ( .A1(n7248), .A2(n7247), .A3(n7294), .ZN(n7249) );
  OAI21_X1 U7802 ( .B1(n7251), .B2(n7250), .A(n7249), .ZN(U3455) );
  OR2_X1 U7803 ( .A1(n7271), .A2(n7252), .ZN(n7254) );
  NAND2_X1 U7804 ( .A1(n7271), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n7253) );
  NAND2_X1 U7805 ( .A1(n7254), .A2(n7253), .ZN(n7281) );
  INV_X1 U7806 ( .A(n7255), .ZN(n7256) );
  AOI211_X1 U7807 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n7257), .A(n7394), .B(n7256), .ZN(n7259) );
  INV_X1 U7808 ( .A(n7259), .ZN(n7262) );
  INV_X1 U7809 ( .A(n7258), .ZN(n7260) );
  OAI22_X1 U7810 ( .A1(n7271), .A2(n7260), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n7259), .ZN(n7261) );
  OAI21_X1 U7811 ( .B1(n7262), .B2(n7448), .A(n7261), .ZN(n7266) );
  OR2_X1 U7812 ( .A1(n7271), .A2(n7263), .ZN(n7265) );
  NAND2_X1 U7813 ( .A1(n7271), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n7264) );
  AOI222_X1 U7814 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7266), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7270), .C1(n7266), .C2(n7270), 
        .ZN(n7267) );
  AOI222_X1 U7815 ( .A1(n7268), .A2(n7281), .B1(n7268), .B2(n7267), .C1(n7281), 
        .C2(n7267), .ZN(n7269) );
  OR2_X1 U7816 ( .A1(n7269), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7284)
         );
  INV_X1 U7817 ( .A(n7270), .ZN(n7282) );
  NAND2_X1 U7818 ( .A1(n7271), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7279) );
  OAI21_X1 U7819 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n7272), 
        .ZN(n7274) );
  NAND3_X1 U7820 ( .A1(n7275), .A2(n7274), .A3(n7273), .ZN(n7277) );
  NOR2_X1 U7821 ( .A1(n7277), .A2(n7276), .ZN(n7278) );
  NAND2_X1 U7822 ( .A1(n7279), .A2(n7278), .ZN(n7280) );
  AOI21_X1 U7823 ( .B1(n7282), .B2(n7281), .A(n7280), .ZN(n7283) );
  NAND2_X1 U7824 ( .A1(n7319), .A2(n7292), .ZN(n7287) );
  NAND2_X1 U7825 ( .A1(READY_N), .A2(n7285), .ZN(n7286) );
  NAND2_X1 U7826 ( .A1(n7287), .A2(n7286), .ZN(n7291) );
  OR2_X1 U7827 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  AOI21_X1 U7828 ( .B1(n7294), .B2(n7293), .A(n7292), .ZN(n7299) );
  AOI21_X1 U7829 ( .B1(READY_N), .B2(n7295), .A(n7302), .ZN(n7309) );
  NOR2_X1 U7830 ( .A1(n7309), .A2(n7296), .ZN(n7297) );
  OAI21_X1 U7831 ( .B1(n7302), .B2(STATE2_REG_0__SCAN_IN), .A(n7297), .ZN(
        n7298) );
  OAI21_X1 U7832 ( .B1(n7302), .B2(n7299), .A(n7298), .ZN(n7300) );
  OR2_X1 U7833 ( .A1(n7301), .A2(n7300), .ZN(U3149) );
  INV_X1 U7834 ( .A(n7302), .ZN(n7312) );
  OAI211_X1 U7835 ( .C1(n7305), .C2(n7312), .A(n7304), .B(n7303), .ZN(U3453)
         );
  INV_X1 U7836 ( .A(n7306), .ZN(n7307) );
  AND2_X1 U7837 ( .A1(n7308), .A2(n7307), .ZN(n7322) );
  INV_X1 U7838 ( .A(n7309), .ZN(n7311) );
  AOI221_X1 U7839 ( .B1(n7322), .B2(STATE2_REG_0__SCAN_IN), .C1(n7311), .C2(
        STATE2_REG_0__SCAN_IN), .A(n7310), .ZN(n7317) );
  OAI211_X1 U7840 ( .C1(n7315), .C2(n7314), .A(n7313), .B(n7312), .ZN(n7316)
         );
  OAI211_X1 U7841 ( .C1(n7319), .C2(n7318), .A(n7317), .B(n7316), .ZN(U3148)
         );
  NOR2_X1 U7842 ( .A1(n7407), .A2(n7320), .ZN(n7321) );
  AOI21_X1 U7843 ( .B1(n7328), .B2(n7322), .A(n7321), .ZN(n7323) );
  OAI21_X1 U7844 ( .B1(n7325), .B2(n7324), .A(n7323), .ZN(n7326) );
  INV_X1 U7845 ( .A(n7326), .ZN(n7327) );
  OAI21_X1 U7846 ( .B1(n7394), .B2(n7328), .A(n7327), .ZN(U3465) );
  INV_X1 U7847 ( .A(n7329), .ZN(n7331) );
  OAI21_X1 U7848 ( .B1(n7333), .B2(n7330), .A(n7331), .ZN(U2792) );
  INV_X1 U7849 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7332) );
  OAI21_X1 U7850 ( .B1(n7333), .B2(n7332), .A(n7331), .ZN(U3452) );
  OAI221_X1 U7851 ( .B1(n7343), .B2(NA_N), .C1(n7343), .C2(n7334), .A(n7345), 
        .ZN(n7344) );
  AOI21_X1 U7852 ( .B1(n7334), .B2(n7343), .A(n7341), .ZN(n7335) );
  OAI21_X1 U7853 ( .B1(n7336), .B2(n7335), .A(n7350), .ZN(n7337) );
  OAI211_X1 U7854 ( .C1(STATE_REG_2__SCAN_IN), .C2(n7348), .A(n7344), .B(n7337), .ZN(U3181) );
  INV_X1 U7855 ( .A(NA_N), .ZN(n7340) );
  AOI21_X1 U7856 ( .B1(n7338), .B2(n7340), .A(STATE_REG_2__SCAN_IN), .ZN(n7349) );
  AOI21_X1 U7857 ( .B1(READY_N), .B2(n7340), .A(n7339), .ZN(n7342) );
  AOI211_X1 U7858 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n7343), .A(n7342), 
        .B(n7341), .ZN(n7346) );
  OAI21_X1 U7859 ( .B1(n7346), .B2(n7345), .A(n7344), .ZN(n7347) );
  OAI21_X1 U7860 ( .B1(n7349), .B2(n7348), .A(n7347), .ZN(U3183) );
  AOI22_X1 U7861 ( .A1(n6947), .A2(n5052), .B1(n7351), .B2(n7350), .ZN(U3473)
         );
  AOI22_X1 U7862 ( .A1(n7353), .A2(n7513), .B1(n7512), .B2(DATAI_17_), .ZN(
        n7355) );
  AOI22_X1 U7863 ( .A1(n7516), .A2(DATAI_1_), .B1(n7515), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n7354) );
  NAND2_X1 U7864 ( .A1(n7355), .A2(n7354), .ZN(U2874) );
  AOI22_X1 U7865 ( .A1(n7356), .A2(n7513), .B1(n7512), .B2(DATAI_19_), .ZN(
        n7358) );
  AOI22_X1 U7866 ( .A1(n7516), .A2(DATAI_3_), .B1(n7515), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n7357) );
  NAND2_X1 U7867 ( .A1(n7358), .A2(n7357), .ZN(U2872) );
  AOI22_X1 U7868 ( .A1(n7359), .A2(n7513), .B1(n7512), .B2(DATAI_21_), .ZN(
        n7361) );
  AOI22_X1 U7869 ( .A1(n7516), .A2(DATAI_5_), .B1(n7515), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n7360) );
  NAND2_X1 U7870 ( .A1(n7361), .A2(n7360), .ZN(U2870) );
  INV_X1 U7871 ( .A(n7362), .ZN(n7363) );
  AOI22_X1 U7872 ( .A1(n7363), .A2(n7513), .B1(n7512), .B2(DATAI_22_), .ZN(
        n7365) );
  AOI22_X1 U7873 ( .A1(n7516), .A2(DATAI_6_), .B1(n7515), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n7364) );
  NAND2_X1 U7874 ( .A1(n7365), .A2(n7364), .ZN(U2869) );
  AOI22_X1 U7875 ( .A1(n7366), .A2(n7513), .B1(n7512), .B2(DATAI_23_), .ZN(
        n7368) );
  AOI22_X1 U7876 ( .A1(n7516), .A2(DATAI_7_), .B1(n7515), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n7367) );
  NAND2_X1 U7877 ( .A1(n7368), .A2(n7367), .ZN(U2868) );
  INV_X1 U7878 ( .A(n7369), .ZN(n7370) );
  OAI21_X1 U7879 ( .B1(n7370), .B2(n7445), .A(n7405), .ZN(n7374) );
  NOR2_X1 U7880 ( .A1(n7394), .A2(n7373), .ZN(n7598) );
  AOI21_X1 U7881 ( .B1(n7395), .B2(n7417), .A(n7598), .ZN(n7375) );
  INV_X1 U7882 ( .A(n7375), .ZN(n7371) );
  AOI22_X1 U7883 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7372), .B1(n7374), .B2(
        n7371), .ZN(n7603) );
  AOI22_X1 U7884 ( .A1(n7453), .A2(n7598), .B1(n7462), .B2(n7597), .ZN(n7378)
         );
  AOI22_X1 U7885 ( .A1(n7375), .A2(n7374), .B1(n7445), .B2(n7373), .ZN(n7376)
         );
  NAND2_X1 U7886 ( .A1(n7459), .A2(n7376), .ZN(n7600) );
  AOI22_X1 U7887 ( .A1(n7600), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n7454), 
        .B2(n7599), .ZN(n7377) );
  OAI211_X1 U7888 ( .C1(n7603), .C2(n7465), .A(n7378), .B(n7377), .ZN(U3124)
         );
  AOI21_X1 U7889 ( .B1(n7432), .B2(n5112), .A(n7445), .ZN(n7382) );
  AND2_X1 U7890 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7384), .ZN(n7605)
         );
  AOI21_X1 U7891 ( .B1(n7379), .B2(n3739), .A(n7605), .ZN(n7381) );
  INV_X1 U7892 ( .A(n7381), .ZN(n7380) );
  AOI22_X1 U7893 ( .A1(n7382), .A2(n7380), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7384), .ZN(n7609) );
  AOI22_X1 U7894 ( .A1(n7453), .A2(n7605), .B1(n7454), .B2(n7604), .ZN(n7387)
         );
  NAND2_X1 U7895 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  OAI211_X1 U7896 ( .C1(n7457), .C2(n7384), .A(n7383), .B(n7459), .ZN(n7606)
         );
  AOI22_X1 U7897 ( .A1(n7606), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n7610), 
        .B2(n7462), .ZN(n7386) );
  OAI211_X1 U7898 ( .C1(n7609), .C2(n7465), .A(n7387), .B(n7386), .ZN(U3108)
         );
  AOI22_X1 U7899 ( .A1(n7453), .A2(n7611), .B1(n7610), .B2(n7454), .ZN(n7391)
         );
  AOI22_X1 U7900 ( .A1(n7612), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n7617), 
        .B2(n7462), .ZN(n7390) );
  OAI211_X1 U7901 ( .C1(n7615), .C2(n7465), .A(n7391), .B(n7390), .ZN(U3100)
         );
  INV_X1 U7902 ( .A(n7392), .ZN(n7393) );
  OAI21_X1 U7903 ( .B1(n7393), .B2(n7445), .A(n7405), .ZN(n7399) );
  NOR2_X1 U7904 ( .A1(n7394), .A2(n7398), .ZN(n7616) );
  AOI21_X1 U7905 ( .B1(n7395), .B2(n7447), .A(n7616), .ZN(n7400) );
  INV_X1 U7906 ( .A(n7400), .ZN(n7396) );
  AOI22_X1 U7907 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7397), .B1(n7399), .B2(
        n7396), .ZN(n7621) );
  AOI22_X1 U7908 ( .A1(n3771), .A2(n7462), .B1(n7453), .B2(n7616), .ZN(n7403)
         );
  AOI22_X1 U7909 ( .A1(n7400), .A2(n7399), .B1(n7445), .B2(n7398), .ZN(n7401)
         );
  NAND2_X1 U7910 ( .A1(n7459), .A2(n7401), .ZN(n7618) );
  AOI22_X1 U7911 ( .A1(n7618), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n7617), 
        .B2(n7454), .ZN(n7402) );
  OAI211_X1 U7912 ( .C1(n7621), .C2(n7465), .A(n7403), .B(n7402), .ZN(U3092)
         );
  INV_X1 U7913 ( .A(n7404), .ZN(n7406) );
  OAI21_X1 U7914 ( .B1(n7406), .B2(n7445), .A(n7405), .ZN(n7412) );
  OR2_X1 U7915 ( .A1(n3662), .A2(n7407), .ZN(n7450) );
  INV_X1 U7916 ( .A(n7450), .ZN(n7418) );
  INV_X1 U7917 ( .A(n7408), .ZN(n7623) );
  AOI21_X1 U7918 ( .B1(n7418), .B2(n7409), .A(n7623), .ZN(n7411) );
  INV_X1 U7919 ( .A(n7411), .ZN(n7410) );
  AOI22_X1 U7920 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7414), .B1(n7412), .B2(
        n7410), .ZN(n7628) );
  AOI22_X1 U7921 ( .A1(n7453), .A2(n7623), .B1(n7622), .B2(n7462), .ZN(n7416)
         );
  NAND2_X1 U7922 ( .A1(n7412), .A2(n7411), .ZN(n7413) );
  OAI211_X1 U7923 ( .C1(n7457), .C2(n7414), .A(n7459), .B(n7413), .ZN(n7624)
         );
  AOI22_X1 U7924 ( .A1(n7625), .A2(n7454), .B1(INSTQUEUE_REG_7__0__SCAN_IN), 
        .B2(n7624), .ZN(n7415) );
  OAI211_X1 U7925 ( .C1(n7628), .C2(n7465), .A(n7416), .B(n7415), .ZN(U3076)
         );
  NAND2_X1 U7926 ( .A1(n7418), .A2(n7417), .ZN(n7419) );
  NAND2_X1 U7927 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7421), .ZN(n7423) );
  NAND2_X1 U7928 ( .A1(n7419), .A2(n7423), .ZN(n7427) );
  AOI21_X1 U7929 ( .B1(n7420), .B2(STATEBS16_REG_SCAN_IN), .A(n7445), .ZN(
        n7424) );
  AOI22_X1 U7930 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7421), .B1(n7427), .B2(
        n7424), .ZN(n7635) );
  INV_X1 U7931 ( .A(n7423), .ZN(n7629) );
  AOI22_X1 U7932 ( .A1(n7462), .A2(n7631), .B1(n7453), .B2(n7629), .ZN(n7430)
         );
  INV_X1 U7933 ( .A(n7424), .ZN(n7428) );
  NAND2_X1 U7934 ( .A1(n7445), .A2(n7425), .ZN(n7426) );
  OAI211_X1 U7935 ( .C1(n7428), .C2(n7427), .A(n7459), .B(n7426), .ZN(n7632)
         );
  AOI22_X1 U7936 ( .A1(n7632), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n7454), 
        .B2(n7630), .ZN(n7429) );
  OAI211_X1 U7937 ( .C1(n7635), .C2(n7465), .A(n7430), .B(n7429), .ZN(U3060)
         );
  AOI21_X1 U7938 ( .B1(n7432), .B2(n7431), .A(n7445), .ZN(n7438) );
  NOR2_X1 U7939 ( .A1(n7433), .A2(n7443), .ZN(n7636) );
  AOI21_X1 U7940 ( .B1(n7434), .B2(n3739), .A(n7636), .ZN(n7437) );
  INV_X1 U7941 ( .A(n7437), .ZN(n7436) );
  INV_X1 U7942 ( .A(n7435), .ZN(n7440) );
  AOI22_X1 U7943 ( .A1(n7438), .A2(n7436), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7440), .ZN(n7642) );
  AOI22_X1 U7944 ( .A1(n7637), .A2(n7454), .B1(n7453), .B2(n7636), .ZN(n7442)
         );
  NAND2_X1 U7945 ( .A1(n7438), .A2(n7437), .ZN(n7439) );
  OAI211_X1 U7946 ( .C1(n7457), .C2(n7440), .A(n7439), .B(n7459), .ZN(n7639)
         );
  AOI22_X1 U7947 ( .A1(n7639), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n7462), 
        .B2(n7638), .ZN(n7441) );
  OAI211_X1 U7948 ( .C1(n7642), .C2(n7465), .A(n7442), .B(n7441), .ZN(U3044)
         );
  NOR2_X1 U7949 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7443), .ZN(n7456)
         );
  INV_X1 U7950 ( .A(n7444), .ZN(n7446) );
  AOI21_X1 U7951 ( .B1(n7446), .B2(STATEBS16_REG_SCAN_IN), .A(n7445), .ZN(
        n7455) );
  INV_X1 U7952 ( .A(n7447), .ZN(n7451) );
  NAND3_X1 U7953 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7449), .A3(n7448), .ZN(n7452) );
  OAI21_X1 U7954 ( .B1(n7451), .B2(n7450), .A(n7452), .ZN(n7460) );
  AOI22_X1 U7955 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7456), .B1(n7455), .B2(
        n7460), .ZN(n7653) );
  INV_X1 U7956 ( .A(n7452), .ZN(n7643) );
  AOI22_X1 U7957 ( .A1(n7646), .A2(n7454), .B1(n7453), .B2(n7643), .ZN(n7464)
         );
  INV_X1 U7958 ( .A(n7455), .ZN(n7461) );
  OR2_X1 U7959 ( .A1(n7457), .A2(n7456), .ZN(n7458) );
  OAI211_X1 U7960 ( .C1(n7461), .C2(n7460), .A(n7459), .B(n7458), .ZN(n7649)
         );
  AOI22_X1 U7961 ( .A1(n7649), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n7462), 
        .B2(n7647), .ZN(n7463) );
  OAI211_X1 U7962 ( .C1(n7653), .C2(n7465), .A(n7464), .B(n7463), .ZN(U3028)
         );
  AOI22_X1 U7963 ( .A1(n7466), .A2(n7513), .B1(n7512), .B2(DATAI_24_), .ZN(
        n7468) );
  AOI22_X1 U7964 ( .A1(n7516), .A2(DATAI_8_), .B1(n7515), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n7467) );
  NAND2_X1 U7965 ( .A1(n7468), .A2(n7467), .ZN(U2867) );
  AOI22_X1 U7966 ( .A1(n7483), .A2(n7598), .B1(n7484), .B2(n7599), .ZN(n7470)
         );
  AOI22_X1 U7967 ( .A1(n7600), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n7485), 
        .B2(n7597), .ZN(n7469) );
  OAI211_X1 U7968 ( .C1(n7603), .C2(n7488), .A(n7470), .B(n7469), .ZN(U3125)
         );
  AOI22_X1 U7969 ( .A1(n7483), .A2(n7605), .B1(n7484), .B2(n7604), .ZN(n7472)
         );
  AOI22_X1 U7970 ( .A1(n7606), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n7610), 
        .B2(n7485), .ZN(n7471) );
  OAI211_X1 U7971 ( .C1(n7609), .C2(n7488), .A(n7472), .B(n7471), .ZN(U3109)
         );
  AOI22_X1 U7972 ( .A1(n7483), .A2(n7611), .B1(n7610), .B2(n7484), .ZN(n7474)
         );
  AOI22_X1 U7973 ( .A1(n7612), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n7617), 
        .B2(n7485), .ZN(n7473) );
  OAI211_X1 U7974 ( .C1(n7615), .C2(n7488), .A(n7474), .B(n7473), .ZN(U3101)
         );
  AOI22_X1 U7975 ( .A1(n3771), .A2(n7485), .B1(n7483), .B2(n7616), .ZN(n7476)
         );
  AOI22_X1 U7976 ( .A1(n7618), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n7617), 
        .B2(n7484), .ZN(n7475) );
  OAI211_X1 U7977 ( .C1(n7621), .C2(n7488), .A(n7476), .B(n7475), .ZN(U3093)
         );
  AOI22_X1 U7978 ( .A1(n7483), .A2(n7623), .B1(n7625), .B2(n7484), .ZN(n7478)
         );
  AOI22_X1 U7979 ( .A1(n7622), .A2(n7485), .B1(INSTQUEUE_REG_7__1__SCAN_IN), 
        .B2(n7624), .ZN(n7477) );
  OAI211_X1 U7980 ( .C1(n7628), .C2(n7488), .A(n7478), .B(n7477), .ZN(U3077)
         );
  AOI22_X1 U7981 ( .A1(n7485), .A2(n7631), .B1(n7483), .B2(n7629), .ZN(n7480)
         );
  AOI22_X1 U7982 ( .A1(n7632), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n7630), 
        .B2(n7484), .ZN(n7479) );
  OAI211_X1 U7983 ( .C1(n7635), .C2(n7488), .A(n7480), .B(n7479), .ZN(U3061)
         );
  AOI22_X1 U7984 ( .A1(n7638), .A2(n7485), .B1(n7483), .B2(n7636), .ZN(n7482)
         );
  AOI22_X1 U7985 ( .A1(n7639), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n7484), 
        .B2(n7637), .ZN(n7481) );
  OAI211_X1 U7986 ( .C1(n7642), .C2(n7488), .A(n7482), .B(n7481), .ZN(U3045)
         );
  AOI22_X1 U7987 ( .A1(n7646), .A2(n7484), .B1(n7483), .B2(n7643), .ZN(n7487)
         );
  AOI22_X1 U7988 ( .A1(n7649), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n7485), 
        .B2(n7647), .ZN(n7486) );
  OAI211_X1 U7989 ( .C1(n7653), .C2(n7488), .A(n7487), .B(n7486), .ZN(U3029)
         );
  AOI22_X1 U7990 ( .A1(n7489), .A2(n7513), .B1(n7512), .B2(DATAI_25_), .ZN(
        n7491) );
  AOI22_X1 U7991 ( .A1(n7516), .A2(DATAI_9_), .B1(n7515), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n7490) );
  NAND2_X1 U7992 ( .A1(n7491), .A2(n7490), .ZN(U2866) );
  AOI22_X1 U7993 ( .A1(n7506), .A2(n7598), .B1(n7508), .B2(n7597), .ZN(n7493)
         );
  AOI22_X1 U7994 ( .A1(n7600), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n7507), 
        .B2(n7599), .ZN(n7492) );
  OAI211_X1 U7995 ( .C1(n7603), .C2(n7511), .A(n7493), .B(n7492), .ZN(U3126)
         );
  AOI22_X1 U7996 ( .A1(n7506), .A2(n7605), .B1(n7610), .B2(n7508), .ZN(n7495)
         );
  AOI22_X1 U7997 ( .A1(n7606), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n7507), 
        .B2(n7604), .ZN(n7494) );
  OAI211_X1 U7998 ( .C1(n7609), .C2(n7511), .A(n7495), .B(n7494), .ZN(U3110)
         );
  AOI22_X1 U7999 ( .A1(n7506), .A2(n7611), .B1(n7610), .B2(n7507), .ZN(n7497)
         );
  AOI22_X1 U8000 ( .A1(n7612), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n7617), 
        .B2(n7508), .ZN(n7496) );
  OAI211_X1 U8001 ( .C1(n7615), .C2(n7511), .A(n7497), .B(n7496), .ZN(U3102)
         );
  AOI22_X1 U8002 ( .A1(n7617), .A2(n7507), .B1(n7506), .B2(n7616), .ZN(n7499)
         );
  AOI22_X1 U8003 ( .A1(n7618), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n7508), 
        .B2(n3771), .ZN(n7498) );
  OAI211_X1 U8004 ( .C1(n7621), .C2(n7511), .A(n7499), .B(n7498), .ZN(U3094)
         );
  AOI22_X1 U8005 ( .A1(n7506), .A2(n7623), .B1(n7625), .B2(n7507), .ZN(n7501)
         );
  AOI22_X1 U8006 ( .A1(n7622), .A2(n7508), .B1(INSTQUEUE_REG_7__2__SCAN_IN), 
        .B2(n7624), .ZN(n7500) );
  OAI211_X1 U8007 ( .C1(n7628), .C2(n7511), .A(n7501), .B(n7500), .ZN(U3078)
         );
  AOI22_X1 U8008 ( .A1(n7630), .A2(n7507), .B1(n7506), .B2(n7629), .ZN(n7503)
         );
  AOI22_X1 U8009 ( .A1(n7632), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n7508), 
        .B2(n7631), .ZN(n7502) );
  OAI211_X1 U8010 ( .C1(n7635), .C2(n7511), .A(n7503), .B(n7502), .ZN(U3062)
         );
  AOI22_X1 U8011 ( .A1(n7638), .A2(n7508), .B1(n7506), .B2(n7636), .ZN(n7505)
         );
  AOI22_X1 U8012 ( .A1(n7639), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n7507), 
        .B2(n7637), .ZN(n7504) );
  OAI211_X1 U8013 ( .C1(n7642), .C2(n7511), .A(n7505), .B(n7504), .ZN(U3046)
         );
  AOI22_X1 U8014 ( .A1(n7646), .A2(n7507), .B1(n7506), .B2(n7643), .ZN(n7510)
         );
  AOI22_X1 U8015 ( .A1(n7649), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n7508), 
        .B2(n7647), .ZN(n7509) );
  OAI211_X1 U8016 ( .C1(n7653), .C2(n7511), .A(n7510), .B(n7509), .ZN(U3030)
         );
  AOI22_X1 U8017 ( .A1(n7514), .A2(n7513), .B1(n7512), .B2(DATAI_26_), .ZN(
        n7518) );
  AOI22_X1 U8018 ( .A1(n7516), .A2(DATAI_10_), .B1(n7515), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n7517) );
  NAND2_X1 U8019 ( .A1(n7518), .A2(n7517), .ZN(U2865) );
  AOI22_X1 U8020 ( .A1(n7533), .A2(n7598), .B1(n7534), .B2(n7599), .ZN(n7520)
         );
  AOI22_X1 U8021 ( .A1(n7600), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n7535), 
        .B2(n7597), .ZN(n7519) );
  OAI211_X1 U8022 ( .C1(n7603), .C2(n7538), .A(n7520), .B(n7519), .ZN(U3127)
         );
  AOI22_X1 U8023 ( .A1(n7533), .A2(n7605), .B1(n7534), .B2(n7604), .ZN(n7522)
         );
  AOI22_X1 U8024 ( .A1(n7606), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n7610), 
        .B2(n7535), .ZN(n7521) );
  OAI211_X1 U8025 ( .C1(n7609), .C2(n7538), .A(n7522), .B(n7521), .ZN(U3111)
         );
  AOI22_X1 U8026 ( .A1(n7533), .A2(n7611), .B1(n7610), .B2(n7534), .ZN(n7524)
         );
  AOI22_X1 U8027 ( .A1(n7612), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n7617), 
        .B2(n7535), .ZN(n7523) );
  OAI211_X1 U8028 ( .C1(n7615), .C2(n7538), .A(n7524), .B(n7523), .ZN(U3103)
         );
  AOI22_X1 U8029 ( .A1(n3771), .A2(n7535), .B1(n7533), .B2(n7616), .ZN(n7526)
         );
  AOI22_X1 U8030 ( .A1(n7618), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n7617), 
        .B2(n7534), .ZN(n7525) );
  OAI211_X1 U8031 ( .C1(n7621), .C2(n7538), .A(n7526), .B(n7525), .ZN(U3095)
         );
  AOI22_X1 U8032 ( .A1(n7622), .A2(n7535), .B1(n7533), .B2(n7623), .ZN(n7528)
         );
  AOI22_X1 U8033 ( .A1(n7625), .A2(n7534), .B1(INSTQUEUE_REG_7__3__SCAN_IN), 
        .B2(n7624), .ZN(n7527) );
  OAI211_X1 U8034 ( .C1(n7628), .C2(n7538), .A(n7528), .B(n7527), .ZN(U3079)
         );
  AOI22_X1 U8035 ( .A1(n7631), .A2(n7535), .B1(n7533), .B2(n7629), .ZN(n7530)
         );
  AOI22_X1 U8036 ( .A1(n7632), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n7630), 
        .B2(n7534), .ZN(n7529) );
  OAI211_X1 U8037 ( .C1(n7635), .C2(n7538), .A(n7530), .B(n7529), .ZN(U3063)
         );
  AOI22_X1 U8038 ( .A1(n7638), .A2(n7535), .B1(n7533), .B2(n7636), .ZN(n7532)
         );
  AOI22_X1 U8039 ( .A1(n7639), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n7534), 
        .B2(n7637), .ZN(n7531) );
  OAI211_X1 U8040 ( .C1(n7642), .C2(n7538), .A(n7532), .B(n7531), .ZN(U3047)
         );
  AOI22_X1 U8041 ( .A1(n7646), .A2(n7534), .B1(n7533), .B2(n7643), .ZN(n7537)
         );
  AOI22_X1 U8042 ( .A1(n7649), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n7535), 
        .B2(n7647), .ZN(n7536) );
  OAI211_X1 U8043 ( .C1(n7653), .C2(n7538), .A(n7537), .B(n7536), .ZN(U3031)
         );
  AOI22_X1 U8044 ( .A1(n7553), .A2(n7598), .B1(n7554), .B2(n7599), .ZN(n7540)
         );
  AOI22_X1 U8045 ( .A1(n7600), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n7555), 
        .B2(n7597), .ZN(n7539) );
  OAI211_X1 U8046 ( .C1(n7603), .C2(n7558), .A(n7540), .B(n7539), .ZN(U3128)
         );
  AOI22_X1 U8047 ( .A1(n7553), .A2(n7605), .B1(n7554), .B2(n7604), .ZN(n7542)
         );
  AOI22_X1 U8048 ( .A1(n7606), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n7610), 
        .B2(n7555), .ZN(n7541) );
  OAI211_X1 U8049 ( .C1(n7609), .C2(n7558), .A(n7542), .B(n7541), .ZN(U3112)
         );
  AOI22_X1 U8050 ( .A1(n7553), .A2(n7611), .B1(n7610), .B2(n7554), .ZN(n7544)
         );
  AOI22_X1 U8051 ( .A1(n7612), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n7617), 
        .B2(n7555), .ZN(n7543) );
  OAI211_X1 U8052 ( .C1(n7615), .C2(n7558), .A(n7544), .B(n7543), .ZN(U3104)
         );
  AOI22_X1 U8053 ( .A1(n7617), .A2(n7554), .B1(n7553), .B2(n7616), .ZN(n7546)
         );
  AOI22_X1 U8054 ( .A1(n7618), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n7555), 
        .B2(n3771), .ZN(n7545) );
  OAI211_X1 U8055 ( .C1(n7621), .C2(n7558), .A(n7546), .B(n7545), .ZN(U3096)
         );
  AOI22_X1 U8056 ( .A1(n7553), .A2(n7623), .B1(n7622), .B2(n7555), .ZN(n7548)
         );
  AOI22_X1 U8057 ( .A1(n7625), .A2(n7554), .B1(INSTQUEUE_REG_7__4__SCAN_IN), 
        .B2(n7624), .ZN(n7547) );
  OAI211_X1 U8058 ( .C1(n7628), .C2(n7558), .A(n7548), .B(n7547), .ZN(U3080)
         );
  AOI22_X1 U8059 ( .A1(n7630), .A2(n7554), .B1(n7553), .B2(n7629), .ZN(n7550)
         );
  AOI22_X1 U8060 ( .A1(n7632), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n7555), 
        .B2(n7631), .ZN(n7549) );
  OAI211_X1 U8061 ( .C1(n7635), .C2(n7558), .A(n7550), .B(n7549), .ZN(U3064)
         );
  AOI22_X1 U8062 ( .A1(n7638), .A2(n7555), .B1(n7553), .B2(n7636), .ZN(n7552)
         );
  AOI22_X1 U8063 ( .A1(n7639), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n7554), 
        .B2(n7637), .ZN(n7551) );
  OAI211_X1 U8064 ( .C1(n7642), .C2(n7558), .A(n7552), .B(n7551), .ZN(U3048)
         );
  AOI22_X1 U8065 ( .A1(n7646), .A2(n7554), .B1(n7553), .B2(n7643), .ZN(n7557)
         );
  AOI22_X1 U8066 ( .A1(n7649), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n7555), 
        .B2(n7647), .ZN(n7556) );
  OAI211_X1 U8067 ( .C1(n7653), .C2(n7558), .A(n7557), .B(n7556), .ZN(U3032)
         );
  AOI22_X1 U8068 ( .A1(n7573), .A2(n7598), .B1(n7574), .B2(n7599), .ZN(n7560)
         );
  AOI22_X1 U8069 ( .A1(n7600), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n7575), 
        .B2(n7597), .ZN(n7559) );
  OAI211_X1 U8070 ( .C1(n7603), .C2(n7578), .A(n7560), .B(n7559), .ZN(U3129)
         );
  AOI22_X1 U8071 ( .A1(n7573), .A2(n7605), .B1(n7574), .B2(n7604), .ZN(n7562)
         );
  AOI22_X1 U8072 ( .A1(n7606), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n7610), 
        .B2(n7575), .ZN(n7561) );
  OAI211_X1 U8073 ( .C1(n7609), .C2(n7578), .A(n7562), .B(n7561), .ZN(U3113)
         );
  AOI22_X1 U8074 ( .A1(n7573), .A2(n7611), .B1(n7610), .B2(n7574), .ZN(n7564)
         );
  AOI22_X1 U8075 ( .A1(n7612), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n7617), 
        .B2(n7575), .ZN(n7563) );
  OAI211_X1 U8076 ( .C1(n7615), .C2(n7578), .A(n7564), .B(n7563), .ZN(U3105)
         );
  AOI22_X1 U8077 ( .A1(n3771), .A2(n7575), .B1(n7573), .B2(n7616), .ZN(n7566)
         );
  AOI22_X1 U8078 ( .A1(n7618), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n7617), 
        .B2(n7574), .ZN(n7565) );
  OAI211_X1 U8079 ( .C1(n7621), .C2(n7578), .A(n7566), .B(n7565), .ZN(U3097)
         );
  AOI22_X1 U8080 ( .A1(n7573), .A2(n7623), .B1(n7622), .B2(n7575), .ZN(n7568)
         );
  AOI22_X1 U8081 ( .A1(n7625), .A2(n7574), .B1(INSTQUEUE_REG_7__5__SCAN_IN), 
        .B2(n7624), .ZN(n7567) );
  OAI211_X1 U8082 ( .C1(n7628), .C2(n7578), .A(n7568), .B(n7567), .ZN(U3081)
         );
  AOI22_X1 U8083 ( .A1(n7575), .A2(n7631), .B1(n7573), .B2(n7629), .ZN(n7570)
         );
  AOI22_X1 U8084 ( .A1(n7632), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n7630), 
        .B2(n7574), .ZN(n7569) );
  OAI211_X1 U8085 ( .C1(n7635), .C2(n7578), .A(n7570), .B(n7569), .ZN(U3065)
         );
  AOI22_X1 U8086 ( .A1(n7638), .A2(n7575), .B1(n7573), .B2(n7636), .ZN(n7572)
         );
  AOI22_X1 U8087 ( .A1(n7639), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n7574), 
        .B2(n7637), .ZN(n7571) );
  OAI211_X1 U8088 ( .C1(n7642), .C2(n7578), .A(n7572), .B(n7571), .ZN(U3049)
         );
  AOI22_X1 U8089 ( .A1(n7646), .A2(n7574), .B1(n7573), .B2(n7643), .ZN(n7577)
         );
  AOI22_X1 U8090 ( .A1(n7649), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n7575), 
        .B2(n7647), .ZN(n7576) );
  OAI211_X1 U8091 ( .C1(n7653), .C2(n7578), .A(n7577), .B(n7576), .ZN(U3033)
         );
  AOI22_X1 U8092 ( .A1(n7591), .A2(n7598), .B1(n7599), .B2(n7592), .ZN(n7580)
         );
  AOI22_X1 U8093 ( .A1(n7600), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n7593), 
        .B2(n7597), .ZN(n7579) );
  OAI211_X1 U8094 ( .C1(n7603), .C2(n7596), .A(n7580), .B(n7579), .ZN(U3130)
         );
  AOI22_X1 U8095 ( .A1(n7591), .A2(n7605), .B1(n7610), .B2(n7593), .ZN(n7582)
         );
  AOI22_X1 U8096 ( .A1(n7606), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n7592), 
        .B2(n7604), .ZN(n7581) );
  OAI211_X1 U8097 ( .C1(n7609), .C2(n7596), .A(n7582), .B(n7581), .ZN(U3114)
         );
  AOI22_X1 U8098 ( .A1(n3771), .A2(n7593), .B1(n7591), .B2(n7616), .ZN(n7584)
         );
  AOI22_X1 U8099 ( .A1(n7618), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n7617), 
        .B2(n7592), .ZN(n7583) );
  OAI211_X1 U8100 ( .C1(n7621), .C2(n7596), .A(n7584), .B(n7583), .ZN(U3098)
         );
  AOI22_X1 U8101 ( .A1(n7625), .A2(n7592), .B1(n7591), .B2(n7623), .ZN(n7586)
         );
  AOI22_X1 U8102 ( .A1(n7622), .A2(n7593), .B1(INSTQUEUE_REG_7__6__SCAN_IN), 
        .B2(n7624), .ZN(n7585) );
  OAI211_X1 U8103 ( .C1(n7628), .C2(n7596), .A(n7586), .B(n7585), .ZN(U3082)
         );
  AOI22_X1 U8104 ( .A1(n7630), .A2(n7592), .B1(n7591), .B2(n7629), .ZN(n7588)
         );
  AOI22_X1 U8105 ( .A1(n7632), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n7593), 
        .B2(n7631), .ZN(n7587) );
  OAI211_X1 U8106 ( .C1(n7635), .C2(n7596), .A(n7588), .B(n7587), .ZN(U3066)
         );
  AOI22_X1 U8107 ( .A1(n7637), .A2(n7592), .B1(n7591), .B2(n7636), .ZN(n7590)
         );
  AOI22_X1 U8108 ( .A1(n7639), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n7593), 
        .B2(n7638), .ZN(n7589) );
  OAI211_X1 U8109 ( .C1(n7642), .C2(n7596), .A(n7590), .B(n7589), .ZN(U3050)
         );
  AOI22_X1 U8110 ( .A1(n7646), .A2(n7592), .B1(n7591), .B2(n7643), .ZN(n7595)
         );
  AOI22_X1 U8111 ( .A1(n7649), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n7593), 
        .B2(n7647), .ZN(n7594) );
  OAI211_X1 U8112 ( .C1(n7653), .C2(n7596), .A(n7595), .B(n7594), .ZN(U3034)
         );
  AOI22_X1 U8113 ( .A1(n7644), .A2(n7598), .B1(n7648), .B2(n7597), .ZN(n7602)
         );
  AOI22_X1 U8114 ( .A1(n7600), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n7645), 
        .B2(n7599), .ZN(n7601) );
  OAI211_X1 U8115 ( .C1(n7603), .C2(n7652), .A(n7602), .B(n7601), .ZN(U3131)
         );
  AOI22_X1 U8116 ( .A1(n7644), .A2(n7605), .B1(n7645), .B2(n7604), .ZN(n7608)
         );
  AOI22_X1 U8117 ( .A1(n7606), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n7610), 
        .B2(n7648), .ZN(n7607) );
  OAI211_X1 U8118 ( .C1(n7609), .C2(n7652), .A(n7608), .B(n7607), .ZN(U3115)
         );
  AOI22_X1 U8119 ( .A1(n7644), .A2(n7611), .B1(n7610), .B2(n7645), .ZN(n7614)
         );
  AOI22_X1 U8120 ( .A1(n7612), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n7617), 
        .B2(n7648), .ZN(n7613) );
  OAI211_X1 U8121 ( .C1(n7615), .C2(n7652), .A(n7614), .B(n7613), .ZN(U3107)
         );
  AOI22_X1 U8122 ( .A1(n3771), .A2(n7648), .B1(n7644), .B2(n7616), .ZN(n7620)
         );
  AOI22_X1 U8123 ( .A1(n7618), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n7617), 
        .B2(n7645), .ZN(n7619) );
  OAI211_X1 U8124 ( .C1(n7621), .C2(n7652), .A(n7620), .B(n7619), .ZN(U3099)
         );
  AOI22_X1 U8125 ( .A1(n7644), .A2(n7623), .B1(n7622), .B2(n7648), .ZN(n7627)
         );
  AOI22_X1 U8126 ( .A1(n7625), .A2(n7645), .B1(INSTQUEUE_REG_7__7__SCAN_IN), 
        .B2(n7624), .ZN(n7626) );
  OAI211_X1 U8127 ( .C1(n7628), .C2(n7652), .A(n7627), .B(n7626), .ZN(U3083)
         );
  AOI22_X1 U8128 ( .A1(n7630), .A2(n7645), .B1(n7644), .B2(n7629), .ZN(n7634)
         );
  AOI22_X1 U8129 ( .A1(n7632), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n7648), 
        .B2(n7631), .ZN(n7633) );
  OAI211_X1 U8130 ( .C1(n7635), .C2(n7652), .A(n7634), .B(n7633), .ZN(U3067)
         );
  AOI22_X1 U8131 ( .A1(n7637), .A2(n7645), .B1(n7644), .B2(n7636), .ZN(n7641)
         );
  AOI22_X1 U8132 ( .A1(n7639), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n7648), 
        .B2(n7638), .ZN(n7640) );
  OAI211_X1 U8133 ( .C1(n7642), .C2(n7652), .A(n7641), .B(n7640), .ZN(U3051)
         );
  AOI22_X1 U8134 ( .A1(n7646), .A2(n7645), .B1(n7644), .B2(n7643), .ZN(n7651)
         );
  AOI22_X1 U8135 ( .A1(n7649), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n7648), 
        .B2(n7647), .ZN(n7650) );
  OAI211_X1 U8136 ( .C1(n7653), .C2(n7652), .A(n7651), .B(n7650), .ZN(U3035)
         );
  CLKBUF_X1 U3698 ( .A(n3908), .Z(n3667) );
  CLKBUF_X1 U3709 ( .A(n3923), .Z(n3981) );
  CLKBUF_X2 U3724 ( .A(n4914), .Z(n3659) );
  CLKBUF_X1 U3728 ( .A(n5448), .Z(n5490) );
  CLKBUF_X1 U3791 ( .A(n5111), .Z(n3654) );
endmodule

