

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, 
        HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684;

  OAI21_X1 U3661 ( .B1(n6535), .B2(n6336), .A(n6335), .ZN(n6518) );
  NAND2_X1 U3662 ( .A1(n6271), .A2(n5825), .ZN(n6281) );
  INV_X1 U3663 ( .A(n6970), .ZN(n6962) );
  NAND2_X1 U3664 ( .A1(n5573), .A2(n5650), .ZN(n5649) );
  NOR2_X2 U3665 ( .A1(n5425), .A2(n4214), .ZN(n5573) );
  NAND2_X1 U3666 ( .A1(n5104), .A2(n3681), .ZN(n5425) );
  AND2_X1 U3667 ( .A1(n3712), .A2(n5599), .ZN(n3643) );
  INV_X2 U3668 ( .A(n6549), .ZN(n6526) );
  NAND2_X1 U3669 ( .A1(n4146), .A2(n4145), .ZN(n4719) );
  NOR2_X1 U3670 ( .A1(n4927), .A2(n4902), .ZN(n4930) );
  INV_X1 U3671 ( .A(n5112), .ZN(n5526) );
  BUF_X1 U3672 ( .A(n4666), .Z(n3665) );
  AND2_X1 U3673 ( .A1(n4658), .A2(n4657), .ZN(n3644) );
  NAND2_X1 U3674 ( .A1(n5579), .A2(n5672), .ZN(n5772) );
  NAND2_X2 U3675 ( .A1(n5125), .A2(n3664), .ZN(n5579) );
  CLKBUF_X1 U3676 ( .A(n3890), .Z(n6455) );
  AND3_X1 U3677 ( .A1(n3889), .A2(n3664), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4622) );
  NAND2_X1 U3678 ( .A1(n5129), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4003) );
  CLKBUF_X1 U3679 ( .A(n4185), .Z(n4565) );
  CLKBUF_X2 U3680 ( .A(n4515), .Z(n3678) );
  NAND4_X2 U3681 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3864)
         );
  AND4_X1 U3682 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3849)
         );
  AND2_X1 U3683 ( .A1(n5020), .A2(n4990), .ZN(n3877) );
  AND2_X1 U3684 ( .A1(n4992), .A2(n4989), .ZN(n3876) );
  AND2_X1 U3685 ( .A1(n4812), .A2(n4990), .ZN(n4515) );
  AND2_X2 U3686 ( .A1(n4992), .A2(n4812), .ZN(n3668) );
  AND2_X2 U3687 ( .A1(n5020), .A2(n3770), .ZN(n4381) );
  AND2_X2 U3688 ( .A1(n4992), .A2(n4812), .ZN(n3669) );
  BUF_X1 U3689 ( .A(n3867), .Z(n3674) );
  CLKBUF_X1 U3690 ( .A(n5262), .Z(n3628) );
  NOR2_X1 U3691 ( .A1(STATEBS16_REG_SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n5262) );
  NOR2_X1 U3692 ( .A1(n6423), .A2(n6414), .ZN(n3629) );
  AND2_X1 U3693 ( .A1(n5384), .A2(n5383), .ZN(n3630) );
  INV_X1 U3694 ( .A(n4929), .ZN(n3631) );
  NOR2_X1 U3695 ( .A1(n6423), .A2(n6414), .ZN(n6415) );
  NAND2_X1 U3696 ( .A1(n6440), .A2(n3697), .ZN(n6423) );
  AND2_X1 U3697 ( .A1(n5342), .A2(n5341), .ZN(n5384) );
  AND2_X2 U3698 ( .A1(n6954), .A2(n5335), .ZN(n3712) );
  NOR2_X1 U3700 ( .A1(n5103), .A2(n5102), .ZN(n3632) );
  INV_X1 U3701 ( .A(n6450), .ZN(n3633) );
  AND2_X1 U3702 ( .A1(n3634), .A2(n6451), .ZN(n3660) );
  NOR2_X1 U3703 ( .A1(n3661), .A2(n3633), .ZN(n3634) );
  NOR2_X1 U3705 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  NAND2_X1 U3706 ( .A1(n4142), .A2(n4141), .ZN(n5103) );
  OAI21_X1 U3707 ( .B1(n5649), .B2(n3702), .A(n3701), .ZN(n6451) );
  NAND2_X1 U3708 ( .A1(n3728), .A2(n3639), .ZN(n3636) );
  AND2_X1 U3709 ( .A1(n3636), .A2(n3637), .ZN(n4745) );
  OR2_X1 U3710 ( .A1(n3638), .A2(n4739), .ZN(n3637) );
  INV_X1 U3711 ( .A(n3738), .ZN(n3638) );
  AND2_X1 U3712 ( .A1(n3731), .A2(n3738), .ZN(n3639) );
  NAND2_X1 U3713 ( .A1(n6952), .A2(n3643), .ZN(n3640) );
  AND2_X2 U3714 ( .A1(n3640), .A2(n3641), .ZN(n5597) );
  OR2_X1 U3715 ( .A1(n3642), .A2(n3709), .ZN(n3641) );
  INV_X1 U3716 ( .A(n5599), .ZN(n3642) );
  CLKBUF_X2 U3717 ( .A(n3670), .Z(n4540) );
  AND2_X1 U3718 ( .A1(n3947), .A2(n3909), .ZN(n4659) );
  OR2_X1 U3719 ( .A1(n3885), .A2(n3898), .ZN(n4768) );
  AND2_X1 U3720 ( .A1(n5020), .A2(n4975), .ZN(n4535) );
  NAND2_X1 U3721 ( .A1(n4815), .A2(n6263), .ZN(n5763) );
  INV_X1 U3722 ( .A(n6263), .ZN(n4786) );
  NAND2_X1 U3723 ( .A1(n3890), .A2(n3888), .ZN(n3923) );
  INV_X2 U3724 ( .A(n3891), .ZN(n3947) );
  INV_X1 U3725 ( .A(n7339), .ZN(n7323) );
  XNOR2_X1 U3726 ( .A(n5774), .B(n5773), .ZN(n5803) );
  AND2_X4 U3728 ( .A1(n5020), .A2(n3770), .ZN(n3666) );
  INV_X1 U3729 ( .A(n4388), .ZN(n3645) );
  NAND2_X1 U3730 ( .A1(n4653), .A2(n3865), .ZN(n3904) );
  NAND2_X2 U3732 ( .A1(n3902), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3996) );
  XNOR2_X2 U3733 ( .A(n4016), .B(n4017), .ZN(n5303) );
  AOI21_X2 U3735 ( .B1(n3665), .B2(n4706), .A(n4665), .ZN(n6935) );
  NAND2_X1 U3738 ( .A1(n4678), .A2(n4913), .ZN(n4963) );
  INV_X4 U3739 ( .A(n6526), .ZN(n6668) );
  NAND3_X1 U3740 ( .A1(n3708), .A2(n6933), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n4912) );
  NAND2_X1 U3741 ( .A1(n4059), .A2(n4058), .ZN(n5524) );
  NAND2_X1 U3742 ( .A1(n3947), .A2(n5139), .ZN(n6261) );
  NAND2_X4 U3743 ( .A1(n3799), .A2(n3798), .ZN(n3891) );
  AND4_X1 U3744 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3883)
         );
  AND4_X1 U3745 ( .A1(n3817), .A2(n3816), .A3(n3815), .A4(n3814), .ZN(n3818)
         );
  AND4_X1 U3746 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3852)
         );
  BUF_X2 U3747 ( .A(n3877), .Z(n4497) );
  BUF_X2 U3748 ( .A(n3876), .Z(n4380) );
  BUF_X2 U3749 ( .A(n3836), .Z(n4533) );
  CLKBUF_X2 U3750 ( .A(n3875), .Z(n4564) );
  CLKBUF_X2 U3751 ( .A(n4535), .Z(n4559) );
  NAND2_X1 U3752 ( .A1(n3656), .A2(n6524), .ZN(n6558) );
  AOI21_X1 U3753 ( .B1(n6271), .B2(n6273), .A(n6272), .ZN(n6490) );
  OR2_X1 U3754 ( .A1(n6281), .A2(n6962), .ZN(n3756) );
  NOR2_X1 U3755 ( .A1(n6533), .A2(n6353), .ZN(n6546) );
  INV_X1 U3756 ( .A(n3707), .ZN(n6272) );
  XNOR2_X1 U3757 ( .A(n3707), .B(n3706), .ZN(n5775) );
  AND2_X1 U3758 ( .A1(n6400), .A2(n6352), .ZN(n6353) );
  OR2_X1 U3759 ( .A1(n6291), .A2(n5824), .ZN(n5825) );
  NAND2_X1 U3760 ( .A1(n6400), .A2(n6399), .ZN(n7442) );
  AND2_X1 U3761 ( .A1(n6290), .A2(n6289), .ZN(n3657) );
  AND2_X1 U3762 ( .A1(n6334), .A2(n6333), .ZN(n6535) );
  NOR2_X1 U3763 ( .A1(n6398), .A2(n6350), .ZN(n6533) );
  NOR2_X1 U3764 ( .A1(n6319), .A2(n6412), .ZN(n6413) );
  NOR2_X2 U3765 ( .A1(n6304), .A2(n6305), .ZN(n6290) );
  NAND2_X1 U3766 ( .A1(n3658), .A2(n3659), .ZN(n6304) );
  AND2_X2 U3767 ( .A1(n6410), .A2(n6411), .ZN(n6319) );
  AND2_X1 U3768 ( .A1(n6419), .A2(n6421), .ZN(n6410) );
  AND2_X1 U3769 ( .A1(n6419), .A2(n6421), .ZN(n3658) );
  INV_X1 U3770 ( .A(n3660), .ZN(n6435) );
  NOR2_X1 U3771 ( .A1(n3718), .A2(n3715), .ZN(n3714) );
  OAI21_X1 U3772 ( .B1(n5803), .B2(n7042), .A(n3699), .ZN(n5806) );
  NOR2_X1 U3773 ( .A1(n4734), .A2(n3720), .ZN(n3719) );
  XNOR2_X1 U3774 ( .A(n4719), .B(n4148), .ZN(n4707) );
  OAI21_X1 U3776 ( .B1(n4687), .B2(n4126), .A(n4125), .ZN(n4959) );
  XNOR2_X1 U3777 ( .A(n4685), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4964)
         );
  NAND2_X1 U3778 ( .A1(n4684), .A2(n4683), .ZN(n4685) );
  NAND2_X1 U3779 ( .A1(n4077), .A2(n4076), .ZN(n4969) );
  NAND2_X1 U3780 ( .A1(n4116), .A2(n4039), .ZN(n5112) );
  AND2_X1 U3781 ( .A1(n4781), .A2(n4780), .ZN(n4783) );
  NAND2_X1 U3782 ( .A1(n4038), .A2(n5042), .ZN(n4039) );
  NAND2_X1 U3783 ( .A1(n4054), .A2(n3748), .ZN(n4781) );
  NAND2_X1 U3784 ( .A1(n4036), .A2(n4035), .ZN(n5145) );
  AOI21_X1 U3785 ( .B1(n5303), .B2(n7400), .A(n4015), .ZN(n4071) );
  AND2_X1 U3786 ( .A1(n5675), .A2(n5674), .ZN(n5694) );
  NAND2_X2 U3787 ( .A1(n6927), .A2(n6455), .ZN(n6454) );
  MUX2_X1 U3788 ( .A(n3628), .B(n4777), .S(n4776), .Z(n4780) );
  NAND2_X1 U3789 ( .A1(n3630), .A2(n3680), .ZN(n5657) );
  AOI21_X1 U3790 ( .B1(n5524), .B2(n4061), .A(n7505), .ZN(n4777) );
  NOR2_X2 U3791 ( .A1(n5107), .A2(n5108), .ZN(n5342) );
  OR3_X2 U3792 ( .A1(n5031), .A2(n6921), .A3(n5036), .ZN(n5107) );
  NAND2_X1 U3793 ( .A1(n4024), .A2(n4023), .ZN(n4976) );
  OAI211_X1 U3794 ( .C1(n3915), .C2(n5778), .A(n3914), .B(n4820), .ZN(n3969)
         );
  NAND2_X1 U3795 ( .A1(n3913), .A2(n4717), .ZN(n4820) );
  AND4_X1 U3796 ( .A1(n3911), .A2(n3910), .A3(n3907), .A4(n5012), .ZN(n3914)
         );
  NOR2_X1 U3797 ( .A1(n4816), .A2(n4826), .ZN(n4640) );
  AND3_X1 U3798 ( .A1(n3961), .A2(n3960), .A3(n3959), .ZN(n3964) );
  NOR2_X1 U3799 ( .A1(n4768), .A2(n5125), .ZN(n3915) );
  NAND2_X1 U3800 ( .A1(n6263), .A2(n5672), .ZN(n5745) );
  AND2_X2 U3801 ( .A1(n5139), .A2(n3664), .ZN(n6995) );
  BUF_X4 U3802 ( .A(n4763), .Z(n5672) );
  INV_X1 U3803 ( .A(n6455), .ZN(n5717) );
  NAND2_X2 U3804 ( .A1(n3883), .A2(n3882), .ZN(n3887) );
  OR2_X1 U3805 ( .A1(n3958), .A2(n3957), .ZN(n4720) );
  OR2_X1 U3806 ( .A1(n3979), .A2(n3978), .ZN(n4660) );
  INV_X4 U3807 ( .A(n3889), .ZN(n5129) );
  OR2_X1 U3808 ( .A1(n3830), .A2(n3829), .ZN(n3890) );
  AND4_X1 U3809 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3863)
         );
  AND4_X1 U3810 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3778)
         );
  AND4_X1 U3811 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3851)
         );
  AND4_X1 U3812 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3808)
         );
  AND4_X1 U3813 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3809)
         );
  AND4_X1 U3814 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3798)
         );
  AND4_X1 U3815 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3775)
         );
  AND4_X1 U3816 ( .A1(n3769), .A2(n3768), .A3(n3767), .A4(n3766), .ZN(n3776)
         );
  AND4_X1 U3817 ( .A1(n3765), .A2(n3764), .A3(n3763), .A4(n3762), .ZN(n3777)
         );
  AND4_X1 U3818 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3850)
         );
  INV_X2 U3819 ( .A(n7376), .ZN(n6828) );
  BUF_X4 U3820 ( .A(n4369), .Z(n3673) );
  AND2_X1 U3821 ( .A1(n4515), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3820) );
  AND2_X2 U3822 ( .A1(n4992), .A2(n5020), .ZN(n3836) );
  AND2_X1 U3823 ( .A1(n3928), .A2(n3997), .ZN(n5529) );
  NOR2_X4 U3824 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5020) );
  AND2_X2 U3825 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4975) );
  INV_X1 U3826 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7496) );
  INV_X1 U3827 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5266) );
  INV_X1 U3828 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7502) );
  AOI21_X1 U3829 ( .B1(n4814), .B2(n7400), .A(n3946), .ZN(n3965) );
  OR2_X1 U3830 ( .A1(n6656), .A2(n7345), .ZN(n3646) );
  NAND2_X1 U3831 ( .A1(n3646), .A2(n6555), .ZN(U2964) );
  AOI211_X1 U3832 ( .C1(n6941), .C2(n7322), .A(n6554), .B(n6553), .ZN(n6555)
         );
  NAND2_X1 U3833 ( .A1(n3644), .A2(n3653), .ZN(n3647) );
  NAND2_X1 U3835 ( .A1(n3644), .A2(n3653), .ZN(n6711) );
  NAND2_X1 U3836 ( .A1(n6959), .A2(n6961), .ZN(n6960) );
  OAI22_X1 U3838 ( .A1(n6485), .A2(n4747), .B1(n5816), .B2(n4746), .ZN(n4748)
         );
  OAI21_X1 U3840 ( .B1(n3724), .B2(n3685), .A(n3722), .ZN(n6959) );
  NOR2_X2 U3841 ( .A1(n4745), .A2(n4744), .ZN(n6500) );
  NOR2_X2 U3842 ( .A1(n6523), .A2(n6565), .ZN(n6665) );
  NAND2_X1 U3843 ( .A1(n3679), .A2(n3654), .ZN(n3651) );
  AND2_X1 U3844 ( .A1(n3651), .A2(n3652), .ZN(n6710) );
  OR2_X1 U3845 ( .A1(n3653), .A2(n4657), .ZN(n3652) );
  INV_X1 U3846 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3653) );
  AND2_X1 U3847 ( .A1(n4706), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3654)
         );
  OR2_X1 U3848 ( .A1(n6558), .A2(n6557), .ZN(n3655) );
  OR2_X1 U3849 ( .A1(n6526), .A2(n6525), .ZN(n3656) );
  AND2_X1 U3850 ( .A1(n4490), .A2(n6411), .ZN(n3659) );
  AND2_X1 U3851 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  NAND2_X1 U3852 ( .A1(n4292), .A2(n4277), .ZN(n3661) );
  INV_X1 U3853 ( .A(n6375), .ZN(n6378) );
  INV_X2 U3854 ( .A(n6261), .ZN(n3921) );
  NAND2_X1 U3855 ( .A1(n4037), .A2(n5145), .ZN(n4116) );
  NAND2_X1 U3856 ( .A1(n3988), .A2(n3987), .ZN(n4050) );
  INV_X4 U3857 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6248) );
  INV_X2 U3858 ( .A(n3887), .ZN(n3900) );
  NAND2_X1 U3859 ( .A1(n3799), .A2(n3798), .ZN(n3664) );
  XNOR2_X1 U3860 ( .A(n4073), .B(n4072), .ZN(n4666) );
  INV_X1 U3861 ( .A(n3645), .ZN(n3676) );
  INV_X1 U3862 ( .A(n3645), .ZN(n3677) );
  INV_X2 U3864 ( .A(n3864), .ZN(n5139) );
  BUF_X1 U3865 ( .A(n3968), .Z(n3991) );
  AND3_X1 U3866 ( .A1(n3897), .A2(n3905), .A3(n3909), .ZN(n4792) );
  AND2_X2 U3867 ( .A1(n3831), .A2(n3890), .ZN(n3897) );
  NAND2_X4 U3868 ( .A1(n3819), .A2(n3818), .ZN(n3888) );
  NAND2_X2 U3869 ( .A1(n3683), .A2(n3863), .ZN(n3909) );
  AND2_X2 U3870 ( .A1(n4813), .A2(n4990), .ZN(n4388) );
  OAI222_X1 U3871 ( .A1(n6454), .A2(n6281), .B1(n6391), .B2(n6927), .C1(n6390), 
        .C2(n6916), .ZN(U2830) );
  INV_X2 U3872 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n7354) );
  AND2_X4 U3873 ( .A1(n6248), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4992)
         );
  INV_X2 U3874 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4994) );
  AND2_X2 U3875 ( .A1(n3770), .A2(n4989), .ZN(n3667) );
  AND2_X1 U3876 ( .A1(n4992), .A2(n4812), .ZN(n4393) );
  INV_X2 U3877 ( .A(n3886), .ZN(n4653) );
  AND2_X2 U3878 ( .A1(n3809), .A2(n3808), .ZN(n3886) );
  NAND2_X2 U3879 ( .A1(n3920), .A2(n5139), .ZN(n4821) );
  INV_X2 U3880 ( .A(n4759), .ZN(n3920) );
  NOR2_X2 U3881 ( .A1(n6428), .A2(n6429), .ZN(n6419) );
  AND2_X1 U3882 ( .A1(n4990), .A2(n4989), .ZN(n3670) );
  NOR2_X2 U3883 ( .A1(n4889), .A2(n4891), .ZN(n4890) );
  OR2_X1 U3884 ( .A1(n6306), .A2(n6290), .ZN(n7582) );
  BUF_X8 U3885 ( .A(n4369), .Z(n3672) );
  BUF_X8 U3886 ( .A(n3867), .Z(n3675) );
  AND2_X4 U3887 ( .A1(n3757), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4812)
         );
  OR2_X2 U3888 ( .A1(n4594), .A2(n4763), .ZN(n3907) );
  NAND2_X2 U3889 ( .A1(n3864), .A2(n3909), .ZN(n4763) );
  XNOR2_X2 U3890 ( .A(n3934), .B(n3990), .ZN(n4814) );
  AND2_X4 U3891 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4989) );
  AND2_X4 U3892 ( .A1(n4992), .A2(n4813), .ZN(n4185) );
  AND2_X4 U3893 ( .A1(n7354), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4813)
         );
  INV_X1 U3894 ( .A(n4116), .ZN(n4113) );
  NAND2_X1 U3895 ( .A1(n4884), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4525) );
  OR2_X1 U3896 ( .A1(n6668), .A2(n7139), .ZN(n4739) );
  INV_X1 U3897 ( .A(n4730), .ZN(n3715) );
  INV_X1 U3898 ( .A(n3719), .ZN(n3718) );
  AND2_X1 U3899 ( .A1(n6366), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U3900 ( .A1(n4637), .A2(n4636), .ZN(n6255) );
  NAND2_X1 U3901 ( .A1(n3657), .A2(n3688), .ZN(n3707) );
  INV_X1 U3902 ( .A(n6273), .ZN(n3705) );
  AND2_X1 U3903 ( .A1(n4489), .A2(n6320), .ZN(n4490) );
  INV_X1 U3904 ( .A(n4715), .ZN(n3710) );
  AND2_X1 U3905 ( .A1(n5266), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4638) );
  INV_X1 U3906 ( .A(n7337), .ZN(n7329) );
  AND2_X1 U3907 ( .A1(n7502), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4599)
         );
  OR2_X1 U3908 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  OR2_X1 U3909 ( .A1(n3945), .A2(n3944), .ZN(n4652) );
  INV_X1 U3910 ( .A(n4652), .ZN(n3948) );
  NAND2_X1 U3911 ( .A1(n3904), .A2(n3889), .ZN(n3905) );
  OR2_X1 U3912 ( .A1(n4627), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4756)
         );
  INV_X1 U3913 ( .A(n3916), .ZN(n4793) );
  OR2_X1 U3914 ( .A1(n6668), .A2(n3691), .ZN(n3682) );
  AND2_X1 U3915 ( .A1(n4488), .A2(n6365), .ZN(n6320) );
  AND2_X1 U3916 ( .A1(n6668), .A2(n4733), .ZN(n4734) );
  INV_X1 U3917 ( .A(n4732), .ZN(n3720) );
  INV_X1 U3918 ( .A(n4731), .ZN(n3717) );
  INV_X1 U3919 ( .A(n5745), .ZN(n5759) );
  NAND2_X1 U3920 ( .A1(n4050), .A2(n3989), .ZN(n4073) );
  NAND2_X1 U3921 ( .A1(n3967), .A2(n3969), .ZN(n3968) );
  OR2_X1 U3922 ( .A1(n3996), .A2(n6248), .ZN(n4001) );
  AOI22_X1 U3923 ( .A1(n4515), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3800) );
  NAND2_X1 U3924 ( .A1(n7460), .A2(n7400), .ZN(n4036) );
  NAND2_X1 U3925 ( .A1(n3904), .A2(n6455), .ZN(n4955) );
  NAND2_X1 U3926 ( .A1(n6334), .A2(n6351), .ZN(n6400) );
  AND2_X1 U3927 ( .A1(n4364), .A2(n4363), .ZN(n6411) );
  AND2_X1 U3928 ( .A1(n4342), .A2(n4341), .ZN(n6421) );
  NAND2_X1 U3929 ( .A1(n4171), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4184)
         );
  INV_X1 U3930 ( .A(n5028), .ZN(n4141) );
  AND2_X1 U3931 ( .A1(n4093), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4118)
         );
  AOI21_X1 U3932 ( .B1(n5526), .B2(n4270), .A(n4046), .ZN(n4920) );
  OAI211_X1 U3933 ( .C1(n4745), .C2(n4743), .A(n5815), .B(n4742), .ZN(n6485)
         );
  OAI21_X1 U3934 ( .B1(n4740), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n6526), 
        .ZN(n4742) );
  AND2_X1 U3935 ( .A1(n6415), .A2(n6367), .ZN(n6402) );
  OR2_X1 U3936 ( .A1(n6668), .A2(n5697), .ZN(n4731) );
  NOR2_X1 U3937 ( .A1(n3723), .A2(n3725), .ZN(n3722) );
  NAND2_X1 U3938 ( .A1(n3708), .A2(n6933), .ZN(n4677) );
  OR2_X1 U3939 ( .A1(n4863), .A2(n4862), .ZN(n4879) );
  NAND2_X1 U3940 ( .A1(n3727), .A2(n4055), .ZN(n4059) );
  OAI21_X1 U3941 ( .B1(n4062), .B2(STATE2_REG_0__SCAN_IN), .A(n4057), .ZN(
        n3727) );
  NOR2_X1 U3942 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5110), .ZN(n5388) );
  INV_X1 U3943 ( .A(n3909), .ZN(n5125) );
  INV_X1 U3944 ( .A(n7316), .ZN(n7151) );
  AND2_X1 U3945 ( .A1(n6366), .A2(n5267), .ZN(n7338) );
  AND2_X1 U3946 ( .A1(n6366), .A2(STATE2_REG_3__SCAN_IN), .ZN(n7335) );
  AND2_X1 U3947 ( .A1(n5776), .A2(n5265), .ZN(n7337) );
  INV_X1 U3948 ( .A(n6927), .ZN(n6426) );
  NAND2_X1 U3949 ( .A1(n5078), .A2(n4954), .ZN(n6479) );
  INV_X1 U3950 ( .A(n4583), .ZN(n3706) );
  NAND2_X1 U3951 ( .A1(n6965), .A2(n4645), .ZN(n6975) );
  NAND2_X1 U3952 ( .A1(n5771), .A2(n5770), .ZN(n5774) );
  OR2_X1 U3953 ( .A1(n6268), .A2(n4815), .ZN(n5771) );
  XNOR2_X1 U3954 ( .A(n3752), .B(n6483), .ZN(n3734) );
  INV_X1 U3955 ( .A(n6796), .ZN(n5045) );
  NAND2_X1 U3956 ( .A1(n5914), .A2(n3755), .ZN(n5918) );
  OAI21_X1 U3957 ( .B1(n3754), .B2(n5936), .A(n3743), .ZN(n5941) );
  OAI21_X1 U3958 ( .B1(n3744), .B2(n5962), .A(n5961), .ZN(n5965) );
  INV_X1 U3959 ( .A(n4635), .ZN(n4623) );
  NAND2_X1 U3960 ( .A1(n3875), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3787)
         );
  OR2_X1 U3961 ( .A1(n4112), .A2(n4111), .ZN(n4692) );
  OR2_X1 U3962 ( .A1(n4090), .A2(n4089), .ZN(n4689) );
  INV_X1 U3963 ( .A(n4622), .ZN(n4603) );
  AOI21_X1 U3964 ( .B1(n3675), .B2(INSTQUEUE_REG_6__7__SCAN_IN), .A(n3820), 
        .ZN(n3824) );
  NAND2_X1 U3965 ( .A1(n3897), .A2(n3899), .ZN(n4816) );
  AND2_X1 U3966 ( .A1(n3672), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U3967 ( .A1(n4388), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3813) );
  OR2_X1 U3968 ( .A1(n4034), .A2(n4033), .ZN(n4680) );
  AND2_X1 U3969 ( .A1(n4622), .A2(n4706), .ZN(n4635) );
  NOR2_X1 U3970 ( .A1(n4357), .A2(n7293), .ZN(n4358) );
  AND2_X1 U3971 ( .A1(n5377), .A2(n5352), .ZN(n3704) );
  OR2_X1 U3972 ( .A1(n4013), .A2(n4012), .ZN(n4669) );
  NAND2_X1 U3973 ( .A1(n6526), .A2(n4729), .ZN(n3726) );
  INV_X1 U3974 ( .A(n5702), .ZN(n3723) );
  NOR2_X1 U3975 ( .A1(n6526), .A2(n3753), .ZN(n3725) );
  OR2_X1 U3976 ( .A1(n6668), .A2(n4725), .ZN(n4726) );
  NAND2_X1 U3977 ( .A1(n3906), .A2(n3864), .ZN(n3911) );
  AND2_X2 U3978 ( .A1(n6248), .A2(n4994), .ZN(n4990) );
  AOI22_X1 U3979 ( .A1(n3935), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3671), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3804) );
  AND2_X1 U3980 ( .A1(n4758), .A2(n4757), .ZN(n6258) );
  CLKBUF_X1 U3981 ( .A(n4759), .Z(n4760) );
  AOI21_X1 U3982 ( .B1(n4707), .B2(n4270), .A(n4156), .ZN(n5102) );
  CLKBUF_X1 U3983 ( .A(n4822), .Z(n4823) );
  AND2_X1 U3984 ( .A1(n4795), .A2(n6264), .ZN(n6799) );
  NOR2_X1 U3985 ( .A1(n5260), .A2(READY_N), .ZN(n5047) );
  AND2_X1 U3986 ( .A1(n7505), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4582) );
  AND2_X1 U3987 ( .A1(n4555), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4646)
         );
  NOR2_X1 U3988 ( .A1(n4527), .A2(n6503), .ZN(n4528) );
  OR2_X1 U3989 ( .A1(n6496), .A2(n4581), .ZN(n4531) );
  AND2_X1 U3990 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4424), .ZN(n4425)
         );
  INV_X1 U3991 ( .A(n4434), .ZN(n4424) );
  NAND2_X1 U3992 ( .A1(n4425), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4527)
         );
  NAND2_X1 U3993 ( .A1(n6668), .A2(n3692), .ZN(n3731) );
  AND2_X1 U3994 ( .A1(n4467), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4437)
         );
  NOR2_X1 U3995 ( .A1(n4465), .A2(n6552), .ZN(n4467) );
  AND2_X1 U3996 ( .A1(n4487), .A2(n4486), .ZN(n6365) );
  AND2_X1 U3997 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4358), .ZN(n4485)
         );
  NOR2_X1 U3998 ( .A1(n4324), .A2(n7269), .ZN(n4325) );
  NAND2_X1 U3999 ( .A1(n4325), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4357)
         );
  OR2_X1 U4000 ( .A1(n4293), .A2(n7260), .ZN(n4324) );
  NOR2_X1 U4001 ( .A1(n4261), .A2(n7246), .ZN(n4278) );
  AOI21_X1 U4002 ( .B1(n5671), .B2(n3703), .A(n4248), .ZN(n3702) );
  NAND2_X1 U4003 ( .A1(n5649), .A2(n3689), .ZN(n3701) );
  NOR2_X1 U4004 ( .A1(n4244), .A2(n7223), .ZN(n4245) );
  NAND2_X1 U4005 ( .A1(n4215), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4244)
         );
  NOR2_X1 U4006 ( .A1(n4184), .A2(n5443), .ZN(n4201) );
  AND2_X1 U4007 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4149) );
  AOI21_X1 U4008 ( .B1(n4699), .B2(n4270), .A(n4140), .ZN(n5028) );
  AOI21_X1 U4009 ( .B1(n4679), .B2(n4270), .A(n4101), .ZN(n4891) );
  AND2_X1 U4010 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n4040), .ZN(n4093)
         );
  CLKBUF_X1 U4011 ( .A(n4889), .Z(n4918) );
  NAND2_X1 U4012 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4068) );
  NOR2_X1 U4013 ( .A1(n6294), .A2(n5817), .ZN(n6268) );
  XNOR2_X1 U4014 ( .A(n6668), .B(n6483), .ZN(n3733) );
  OR2_X2 U4015 ( .A1(n6309), .A2(n6296), .ZN(n6294) );
  XNOR2_X1 U4016 ( .A(n6526), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6494)
         );
  NAND2_X1 U4017 ( .A1(n6330), .A2(n6307), .ZN(n6309) );
  AND2_X1 U4018 ( .A1(n6668), .A2(n6623), .ZN(n4744) );
  NOR2_X2 U4019 ( .A1(n3696), .A2(n3690), .ZN(n6330) );
  NAND2_X1 U4020 ( .A1(n6402), .A2(n3694), .ZN(n6632) );
  NOR2_X1 U4021 ( .A1(n6356), .A2(n3695), .ZN(n3694) );
  INV_X1 U4022 ( .A(n6401), .ZN(n3695) );
  NOR2_X1 U4023 ( .A1(n7006), .A2(n6677), .ZN(n6650) );
  NOR2_X1 U4024 ( .A1(n6425), .A2(n3698), .ZN(n3697) );
  INV_X1 U4025 ( .A(n6431), .ZN(n3698) );
  AOI21_X1 U4026 ( .B1(n3719), .B2(n3717), .A(n3684), .ZN(n3716) );
  AND2_X1 U4027 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  AND2_X1 U4028 ( .A1(n5035), .A2(n5034), .ZN(n5036) );
  OR2_X1 U4029 ( .A1(n5031), .A2(n6921), .ZN(n6923) );
  NAND2_X1 U4030 ( .A1(n4703), .A2(n7047), .ZN(n6947) );
  XNOR2_X1 U4031 ( .A(n4696), .B(n7051), .ZN(n6940) );
  AND2_X1 U4032 ( .A1(n7063), .A2(n7038), .ZN(n5799) );
  AND2_X1 U4033 ( .A1(n5688), .A2(n5344), .ZN(n7019) );
  AND2_X1 U4034 ( .A1(n4877), .A2(n4876), .ZN(n7088) );
  OAI21_X1 U4035 ( .B1(n3996), .B2(n7354), .A(n3903), .ZN(n3967) );
  INV_X1 U4036 ( .A(n3908), .ZN(n4884) );
  INV_X1 U4037 ( .A(n6255), .ZN(n6262) );
  OR2_X1 U4038 ( .A1(n3996), .A2(n4994), .ZN(n4024) );
  NAND2_X1 U4039 ( .A1(n4018), .A2(n4017), .ZN(n4978) );
  NOR2_X1 U4040 ( .A1(n4847), .A2(n4953), .ZN(n5004) );
  OR2_X1 U4041 ( .A1(n5637), .A2(n7640), .ZN(n5527) );
  OR2_X1 U4042 ( .A1(n5146), .A2(n5042), .ZN(n5503) );
  AOI21_X1 U4043 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7502), .A(n5450), .ZN(
        n7513) );
  INV_X1 U4044 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U4045 ( .A1(n5260), .A2(n5259), .ZN(n6997) );
  INV_X1 U4046 ( .A(n7335), .ZN(n7294) );
  NAND2_X1 U4047 ( .A1(n5776), .A2(n5274), .ZN(n7316) );
  AND2_X1 U4048 ( .A1(n5776), .A2(n5282), .ZN(n7332) );
  INV_X1 U4049 ( .A(n6366), .ZN(n7268) );
  AND2_X1 U4050 ( .A1(n7325), .A2(n5268), .ZN(n7172) );
  INV_X1 U4051 ( .A(n6916), .ZN(n6924) );
  AND2_X1 U4052 ( .A1(n4775), .A2(n7397), .ZN(n6927) );
  INV_X1 U4053 ( .A(n6546), .ZN(n6473) );
  AND2_X1 U4054 ( .A1(n6479), .A2(n4955), .ZN(n7521) );
  AND2_X1 U4055 ( .A1(n3886), .A2(n6455), .ZN(n6456) );
  INV_X1 U4056 ( .A(n6479), .ZN(n7584) );
  NAND2_X1 U4057 ( .A1(n6479), .A2(n4956), .ZN(n6481) );
  INV_X1 U4058 ( .A(n7435), .ZN(n7286) );
  NAND2_X1 U4059 ( .A1(n5669), .A2(n5671), .ZN(n5670) );
  INV_X1 U4061 ( .A(n6965), .ZN(n6969) );
  INV_X1 U4062 ( .A(n7345), .ZN(n6971) );
  AND2_X1 U4063 ( .A1(n3700), .A2(n5804), .ZN(n3699) );
  OR2_X1 U4064 ( .A1(n5805), .A2(n5811), .ZN(n3700) );
  XNOR2_X1 U4065 ( .A(n6486), .B(n6600), .ZN(n6604) );
  OAI21_X1 U4066 ( .B1(n6485), .B2(n3736), .A(n6484), .ZN(n6486) );
  NOR2_X1 U4067 ( .A1(n6633), .A2(n5808), .ZN(n7140) );
  NAND2_X1 U4068 ( .A1(n5679), .A2(n4731), .ZN(n3721) );
  NAND2_X1 U4069 ( .A1(n4879), .A2(n4878), .ZN(n7042) );
  AND2_X1 U4070 ( .A1(n7019), .A2(n7063), .ZN(n7040) );
  AND2_X1 U4071 ( .A1(n4879), .A2(n4869), .ZN(n7133) );
  INV_X1 U4072 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7364) );
  AND2_X1 U4073 ( .A1(n5024), .A2(n5450), .ZN(n6796) );
  NOR2_X1 U4075 ( .A1(n7390), .A2(n6262), .ZN(n6721) );
  INV_X1 U4076 ( .A(n5418), .ZN(n7667) );
  AND2_X1 U4077 ( .A1(n7471), .A2(n3662), .ZN(n7652) );
  INV_X1 U4078 ( .A(n5409), .ZN(n7645) );
  NOR2_X1 U4079 ( .A1(n5387), .A2(n5139), .ZN(n7536) );
  NOR2_X1 U4080 ( .A1(n5387), .A2(n5125), .ZN(n7572) );
  NOR2_X1 U4081 ( .A1(n5387), .A2(n5129), .ZN(n7599) );
  NOR2_X1 U4082 ( .A1(n5387), .A2(n5717), .ZN(n7674) );
  INV_X1 U4083 ( .A(n7519), .ZN(n6740) );
  INV_X1 U4084 ( .A(n7535), .ZN(n7537) );
  INV_X1 U4085 ( .A(n7536), .ZN(n5619) );
  INV_X1 U4086 ( .A(n7554), .ZN(n5634) );
  INV_X1 U4087 ( .A(n7571), .ZN(n7573) );
  INV_X1 U4088 ( .A(n7598), .ZN(n7600) );
  INV_X1 U4089 ( .A(n7599), .ZN(n5628) );
  INV_X1 U4090 ( .A(n7616), .ZN(n7618) );
  INV_X1 U4091 ( .A(n7617), .ZN(n5625) );
  INV_X1 U4092 ( .A(n7637), .ZN(n6765) );
  INV_X1 U4093 ( .A(n7632), .ZN(n5622) );
  INV_X1 U4094 ( .A(n7671), .ZN(n7676) );
  INV_X1 U4095 ( .A(n7674), .ZN(n5616) );
  AND2_X1 U4096 ( .A1(n4638), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7397) );
  OAI21_X1 U4097 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7391) );
  NAND2_X1 U4098 ( .A1(n5775), .A2(n7338), .ZN(n5791) );
  OAI211_X1 U4099 ( .C1(n5827), .C2(n6975), .A(n5826), .B(n3756), .ZN(n5828)
         );
  NAND2_X1 U4100 ( .A1(n5333), .A2(n5335), .ZN(n5334) );
  AND2_X1 U4101 ( .A1(n5585), .A2(n5584), .ZN(n3680) );
  NAND2_X1 U4102 ( .A1(n6378), .A2(n4277), .ZN(n6377) );
  AND2_X1 U4103 ( .A1(n3704), .A2(n4200), .ZN(n3681) );
  AND4_X1 U4104 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3683)
         );
  XNOR2_X1 U4105 ( .A(n4116), .B(n4102), .ZN(n4679) );
  XNOR2_X1 U4106 ( .A(n5649), .B(n4248), .ZN(n5669) );
  NAND2_X1 U4107 ( .A1(n3657), .A2(n5824), .ZN(n6271) );
  OR2_X1 U4108 ( .A1(n6632), .A2(n5753), .ZN(n3696) );
  NAND2_X1 U4109 ( .A1(n4001), .A2(n4000), .ZN(n4017) );
  NOR2_X1 U4110 ( .A1(n6668), .A2(n4733), .ZN(n3684) );
  NAND2_X1 U4111 ( .A1(n6319), .A2(n6365), .ZN(n6398) );
  NAND2_X1 U4112 ( .A1(n4726), .A2(n3726), .ZN(n3685) );
  NAND2_X1 U4113 ( .A1(n3660), .A2(n4309), .ZN(n6428) );
  AND2_X1 U4114 ( .A1(n4724), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3686)
         );
  NAND2_X1 U4115 ( .A1(n3632), .A2(n3704), .ZN(n5376) );
  NAND2_X1 U4116 ( .A1(n6402), .A2(n6401), .ZN(n6354) );
  NAND2_X1 U4117 ( .A1(n6440), .A2(n6431), .ZN(n6422) );
  AND2_X1 U4118 ( .A1(n5597), .A2(n4726), .ZN(n3687) );
  AND2_X1 U4119 ( .A1(n3632), .A2(n5352), .ZN(n5353) );
  NAND2_X1 U4120 ( .A1(n3648), .A2(n4730), .ZN(n5679) );
  NAND2_X1 U4121 ( .A1(n3721), .A2(n4732), .ZN(n6583) );
  NAND2_X1 U4122 ( .A1(n6953), .A2(n4715), .ZN(n5333) );
  AND2_X1 U4123 ( .A1(n3705), .A2(n5824), .ZN(n3688) );
  AND2_X1 U4124 ( .A1(n4653), .A2(n3864), .ZN(n4706) );
  AND2_X1 U4125 ( .A1(n5671), .A2(n4248), .ZN(n3689) );
  NAND2_X1 U4126 ( .A1(n5384), .A2(n5383), .ZN(n5586) );
  INV_X1 U4127 ( .A(n5424), .ZN(n4200) );
  AND2_X1 U4128 ( .A1(n5758), .A2(n5757), .ZN(n3690) );
  AND4_X1 U4129 ( .A1(n6676), .A2(n6652), .A3(n5748), .A4(n6645), .ZN(n3691)
         );
  NAND2_X1 U4130 ( .A1(n3693), .A2(n4738), .ZN(n3692) );
  AND2_X1 U4131 ( .A1(n6525), .A2(n6651), .ZN(n3693) );
  INV_X1 U4132 ( .A(n3628), .ZN(n4581) );
  NOR3_X2 U4133 ( .A1(n7502), .A2(n7501), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n7666) );
  NOR3_X2 U4134 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n7501), .ZN(n7673) );
  NOR2_X2 U4135 ( .A1(n5657), .A2(n5656), .ZN(n5675) );
  INV_X1 U4136 ( .A(n3696), .ZN(n6338) );
  INV_X1 U4137 ( .A(n4248), .ZN(n3703) );
  NAND2_X1 U4138 ( .A1(n6932), .A2(n6935), .ZN(n3708) );
  NAND2_X1 U4139 ( .A1(n4668), .A2(n4897), .ZN(n6933) );
  NAND2_X1 U4140 ( .A1(n6952), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U4141 ( .A1(n3711), .A2(n3709), .ZN(n5596) );
  AOI21_X1 U4142 ( .B1(n3710), .B2(n5335), .A(n3686), .ZN(n3709) );
  NAND2_X1 U4143 ( .A1(n6952), .A2(n3712), .ZN(n3711) );
  NAND2_X1 U4144 ( .A1(n6960), .A2(n3714), .ZN(n3713) );
  NAND2_X1 U4145 ( .A1(n3713), .A2(n3716), .ZN(n6575) );
  INV_X1 U4146 ( .A(n5597), .ZN(n3724) );
  NAND2_X1 U4147 ( .A1(n4737), .A2(n4736), .ZN(n3729) );
  NAND2_X1 U4148 ( .A1(n4735), .A2(n6526), .ZN(n3730) );
  NAND2_X1 U4149 ( .A1(n3730), .A2(n3729), .ZN(n6523) );
  NAND2_X1 U4150 ( .A1(n3728), .A2(n3731), .ZN(n6515) );
  NAND3_X1 U4151 ( .A1(n3730), .A2(n3729), .A3(n3682), .ZN(n3728) );
  NAND2_X1 U4152 ( .A1(n6493), .A2(n3733), .ZN(n3732) );
  OAI21_X1 U4153 ( .B1(n6493), .B2(n3734), .A(n3732), .ZN(n5830) );
  OAI21_X1 U4154 ( .B1(n5830), .B2(n7055), .A(n5820), .ZN(U2989) );
  NAND2_X1 U4155 ( .A1(n6451), .A2(n6450), .ZN(n6375) );
  AND2_X1 U4156 ( .A1(n3665), .A2(n5175), .ZN(n5458) );
  INV_X1 U4157 ( .A(n4917), .ZN(n4079) );
  NAND2_X1 U4158 ( .A1(n4050), .A2(n4049), .ZN(n4651) );
  NAND4_X1 U4159 ( .A1(n3890), .A2(n3900), .A3(n3865), .A4(n3889), .ZN(n3908)
         );
  NAND2_X1 U4160 ( .A1(n3890), .A2(n3865), .ZN(n4060) );
  AOI22_X1 U4161 ( .A1(n3875), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3668), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4162 ( .A1(n3668), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3828) );
  INV_X1 U4163 ( .A(n3888), .ZN(n3865) );
  INV_X1 U4164 ( .A(n4098), .ZN(n4051) );
  OR2_X1 U4165 ( .A1(n6016), .A2(n6015), .ZN(n3735) );
  AND2_X1 U4166 ( .A1(n6526), .A2(n6483), .ZN(n3736) );
  OR2_X1 U4167 ( .A1(n6526), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3737)
         );
  OR2_X1 U4168 ( .A1(n6526), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3738)
         );
  NOR2_X1 U4169 ( .A1(n4115), .A2(n4114), .ZN(n3739) );
  AND3_X1 U4170 ( .A1(n5861), .A2(n5860), .A3(n5859), .ZN(n3740) );
  AND2_X1 U4171 ( .A1(n5884), .A2(n5883), .ZN(n3741) );
  NAND2_X1 U4172 ( .A1(keyinput_143), .A2(n5876), .ZN(n3742) );
  XOR2_X1 U4173 ( .A(n6906), .B(keyinput_176), .Z(n3743) );
  AND2_X1 U4174 ( .A1(n5959), .A2(n5958), .ZN(n3744) );
  AND2_X1 U4175 ( .A1(n4185), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3745) );
  AND2_X1 U4176 ( .A1(n4381), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3746) );
  AND2_X1 U4177 ( .A1(n3670), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3747) );
  AND2_X1 U4178 ( .A1(n4053), .A2(n4052), .ZN(n3748) );
  AND3_X1 U4179 ( .A1(n6010), .A2(n6009), .A3(n6008), .ZN(n3749) );
  AND3_X1 U4180 ( .A1(n7126), .A2(n6686), .A3(n6707), .ZN(n3750) );
  OR2_X1 U4181 ( .A1(n3931), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3751)
         );
  AND2_X1 U4182 ( .A1(n6668), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3752)
         );
  AND2_X1 U4183 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3753) );
  INV_X1 U4184 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5443) );
  AND2_X1 U4185 ( .A1(n5933), .A2(n5932), .ZN(n3754) );
  NAND2_X1 U4186 ( .A1(n4113), .A2(n3739), .ZN(n4143) );
  INV_X1 U4187 ( .A(n6376), .ZN(n4277) );
  AND2_X1 U4188 ( .A1(n5913), .A2(n5912), .ZN(n3755) );
  INV_X1 U4189 ( .A(keyinput_130), .ZN(n5840) );
  NAND2_X1 U4190 ( .A1(keyinput_129), .A2(DATAI_30_), .ZN(n5843) );
  OAI22_X1 U4191 ( .A1(n5853), .A2(keyinput_132), .B1(n5852), .B2(DATAI_27_), 
        .ZN(n5854) );
  INV_X1 U4192 ( .A(keyinput_133), .ZN(n5857) );
  XNOR2_X1 U4193 ( .A(n5857), .B(DATAI_26_), .ZN(n5860) );
  INV_X1 U4194 ( .A(keyinput_146), .ZN(n5881) );
  XNOR2_X1 U4195 ( .A(n5882), .B(n5881), .ZN(n5883) );
  NAND2_X1 U4196 ( .A1(n3742), .A2(n5878), .ZN(n5885) );
  NAND2_X1 U4197 ( .A1(n5885), .A2(n3741), .ZN(n5894) );
  NAND2_X1 U4198 ( .A1(keyinput_165), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5912)
         );
  INV_X1 U4199 ( .A(keyinput_168), .ZN(n5919) );
  NAND2_X1 U4200 ( .A1(M_IO_N_REG_SCAN_IN), .A2(n5919), .ZN(n5920) );
  OAI22_X1 U4201 ( .A1(n7373), .A2(n5930), .B1(FLUSH_REG_SCAN_IN), .B2(
        keyinput_173), .ZN(n5931) );
  INV_X1 U4202 ( .A(n5931), .ZN(n5932) );
  NAND2_X1 U4203 ( .A1(n6874), .A2(keyinput_183), .ZN(n5947) );
  OAI22_X1 U4204 ( .A1(n6868), .A2(n5951), .B1(REIP_REG_24__SCAN_IN), .B2(
        keyinput_186), .ZN(n5952) );
  OAI22_X1 U4205 ( .A1(n6867), .A2(keyinput_187), .B1(n5956), .B2(
        REIP_REG_23__SCAN_IN), .ZN(n5957) );
  INV_X1 U4206 ( .A(n5957), .ZN(n5958) );
  INV_X1 U4207 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U4208 ( .A(n5963), .B(keyinput_191), .ZN(n5964) );
  XNOR2_X1 U4209 ( .A(keyinput_199), .B(ADDRESS_REG_29__SCAN_IN), .ZN(n5976)
         );
  NOR3_X1 U4210 ( .A1(n5978), .A2(n5977), .A3(n5976), .ZN(n5980) );
  OR2_X1 U4211 ( .A1(n4596), .A2(n4611), .ZN(n4597) );
  INV_X1 U4212 ( .A(n6001), .ZN(n6002) );
  AND2_X1 U4213 ( .A1(n4609), .A2(n4608), .ZN(n4612) );
  INV_X1 U4214 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3868) );
  INV_X1 U4215 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4727) );
  OAI21_X1 U4216 ( .B1(n4116), .B2(n4115), .A(n4114), .ZN(n4117) );
  INV_X1 U4217 ( .A(n3923), .ZN(n3924) );
  AOI22_X1 U4218 ( .A1(n3673), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3874) );
  NAND2_X1 U4219 ( .A1(n4143), .A2(n4117), .ZN(n4687) );
  NAND2_X1 U4220 ( .A1(n3947), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4002) );
  AND4_X1 U4221 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3882)
         );
  NAND2_X1 U4222 ( .A1(n4388), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3835) );
  AND2_X1 U4223 ( .A1(n6036), .A2(n6035), .ZN(n6039) );
  NOR2_X1 U4224 ( .A1(n3747), .A2(n3782), .ZN(n3793) );
  NAND2_X1 U4225 ( .A1(n4003), .A2(n4002), .ZN(n4632) );
  OR2_X1 U4226 ( .A1(n4136), .A2(n4135), .ZN(n4709) );
  NAND2_X1 U4227 ( .A1(n3966), .A2(n3989), .ZN(n4048) );
  AOI21_X1 U4228 ( .B1(n3670), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n3858), 
        .ZN(n3860) );
  AND2_X1 U4229 ( .A1(n6039), .A2(n6038), .ZN(n6040) );
  OR2_X1 U4230 ( .A1(n4844), .A2(n3920), .ZN(n4854) );
  NOR2_X1 U4231 ( .A1(n6455), .A2(n7505), .ZN(n4063) );
  INV_X1 U4232 ( .A(n4063), .ZN(n4579) );
  INV_X1 U4233 ( .A(n4143), .ZN(n4146) );
  AND2_X1 U4234 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  INV_X1 U4235 ( .A(keyinput_248), .ZN(n6047) );
  INV_X1 U4236 ( .A(n6436), .ZN(n4309) );
  AND2_X1 U4237 ( .A1(n4854), .A2(n4825), .ZN(n4838) );
  AND2_X1 U4238 ( .A1(n4532), .A2(n4531), .ZN(n6289) );
  NAND2_X1 U4239 ( .A1(n4485), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4465)
         );
  INV_X1 U4240 ( .A(n6442), .ZN(n4292) );
  INV_X1 U4241 ( .A(n4579), .ZN(n4482) );
  OAI21_X1 U4242 ( .B1(n5570), .B2(n7390), .A(n5536), .ZN(n5565) );
  NAND2_X1 U4243 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6047), .ZN(n6048) );
  INV_X1 U4244 ( .A(n6995), .ZN(n5778) );
  NAND2_X1 U4245 ( .A1(n4245), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4261)
         );
  OR2_X1 U4246 ( .A1(n6997), .A2(n5263), .ZN(n6366) );
  INV_X1 U4247 ( .A(n6397), .ZN(n6351) );
  OR2_X1 U4248 ( .A1(n4861), .A2(n7380), .ZN(n5046) );
  NAND2_X1 U4249 ( .A1(n4437), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4434)
         );
  AND2_X1 U4250 ( .A1(n4201), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4215)
         );
  AND2_X1 U4251 ( .A1(n4150), .A2(n4149), .ZN(n4171) );
  INV_X1 U4252 ( .A(n6523), .ZN(n6540) );
  NAND2_X1 U4253 ( .A1(n4879), .A2(n6254), .ZN(n7063) );
  INV_X1 U4254 ( .A(n7659), .ZN(n5417) );
  INV_X1 U4255 ( .A(n5533), .ZN(n5227) );
  OR2_X1 U4256 ( .A1(n5302), .A2(n5301), .ZN(n5409) );
  OR2_X1 U4257 ( .A1(n7446), .A2(n3679), .ZN(n5605) );
  INV_X1 U4258 ( .A(n5637), .ZN(n5568) );
  AOI21_X1 U4259 ( .B1(n7393), .B2(n7388), .A(n6721), .ZN(n5110) );
  INV_X1 U4260 ( .A(n3662), .ZN(n5300) );
  OR3_X1 U4261 ( .A1(n7390), .A2(STATE2_REG_0__SCAN_IN), .A3(n5110), .ZN(n5387) );
  NAND2_X1 U4262 ( .A1(n4792), .A2(n3917), .ZN(n6260) );
  NOR2_X1 U4263 ( .A1(n7316), .A2(n5433), .ZN(n7218) );
  INV_X1 U4264 ( .A(n7279), .ZN(n7291) );
  NOR2_X1 U4265 ( .A1(n5368), .A2(n7268), .ZN(n7279) );
  AND2_X1 U4266 ( .A1(n6366), .A2(n5278), .ZN(n7339) );
  AND2_X1 U4267 ( .A1(n6479), .A2(n6456), .ZN(n7520) );
  INV_X1 U4269 ( .A(n5078), .ZN(n5065) );
  AND2_X1 U4270 ( .A1(n4118), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4150)
         );
  INV_X1 U4271 ( .A(n6975), .ZN(n6941) );
  NAND2_X1 U4272 ( .A1(n6255), .A2(n7397), .ZN(n4861) );
  INV_X1 U4273 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6483) );
  AOI21_X1 U4274 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n6526), .A(n6556), 
        .ZN(n6551) );
  NOR2_X1 U4275 ( .A1(n7119), .A2(n6700), .ZN(n7127) );
  NAND2_X1 U4276 ( .A1(n6689), .A2(n5696), .ZN(n7106) );
  INV_X1 U4277 ( .A(n7063), .ZN(n7087) );
  NOR2_X1 U4278 ( .A1(n7019), .A2(n6708), .ZN(n7068) );
  INV_X1 U4279 ( .A(n7042), .ZN(n7132) );
  NOR2_X1 U4280 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7383) );
  INV_X1 U4281 ( .A(n5488), .ZN(n7677) );
  AND2_X1 U4282 ( .A1(n5174), .A2(n3662), .ZN(n7680) );
  OAI211_X1 U4283 ( .C1(n5116), .C2(n5115), .A(n5306), .B(n5227), .ZN(n5416)
         );
  INV_X1 U4284 ( .A(n5410), .ZN(n7654) );
  OAI211_X1 U4285 ( .C1(n5308), .C2(n7390), .A(n5307), .B(n5306), .ZN(n5408)
         );
  OAI211_X1 U4286 ( .C1(n7390), .C2(n5230), .A(n5229), .B(n5228), .ZN(n5404)
         );
  AND2_X1 U4287 ( .A1(n5526), .A2(n5525), .ZN(n7640) );
  AND2_X1 U4288 ( .A1(n5458), .A2(n3662), .ZN(n6771) );
  INV_X1 U4289 ( .A(n7553), .ZN(n7555) );
  NOR2_X1 U4290 ( .A1(n5387), .A2(n3886), .ZN(n7617) );
  OR2_X1 U4291 ( .A1(n4861), .A2(n6260), .ZN(n5260) );
  INV_X1 U4292 ( .A(n7338), .ZN(n7325) );
  INV_X1 U4293 ( .A(n7332), .ZN(n7312) );
  NAND2_X1 U4294 ( .A1(n6927), .A2(n5717), .ZN(n6916) );
  INV_X2 U4295 ( .A(n7521), .ZN(n7581) );
  INV_X1 U4296 ( .A(n6799), .ZN(n6830) );
  NAND2_X1 U4297 ( .A1(n5047), .A2(n3864), .ZN(n5078) );
  NAND2_X1 U4298 ( .A1(n7345), .A2(n4642), .ZN(n6965) );
  OR2_X1 U4299 ( .A1(n4861), .A2(n4864), .ZN(n7345) );
  NAND2_X1 U4300 ( .A1(n5807), .A2(n7106), .ZN(n7119) );
  INV_X1 U4301 ( .A(n7133), .ZN(n7055) );
  INV_X1 U4302 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7363) );
  AOI21_X1 U4303 ( .B1(n5179), .B2(n5178), .A(n5177), .ZN(n7684) );
  INV_X1 U4304 ( .A(n7506), .ZN(n7672) );
  INV_X1 U4305 ( .A(n7474), .ZN(n7658) );
  INV_X1 U4306 ( .A(n7507), .ZN(n5642) );
  INV_X1 U4307 ( .A(n7572), .ZN(n5631) );
  INV_X1 U4308 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7400) );
  AOI211_X1 U4309 ( .C1(n6236), .C2(n6235), .A(n6234), .B(n6233), .ZN(n6239)
         );
  AND2_X4 U4310 ( .A1(n4994), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3770)
         );
  AND2_X4 U4311 ( .A1(n3770), .A2(n4813), .ZN(n3867) );
  NAND2_X1 U4312 ( .A1(n3675), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U4313 ( .A1(n4515), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3760) );
  AND2_X4 U4314 ( .A1(n3770), .A2(n4812), .ZN(n4369) );
  NAND2_X1 U4315 ( .A1(n3673), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3759) );
  AND2_X2 U4316 ( .A1(n4812), .A2(n4975), .ZN(n3935) );
  NAND2_X1 U4317 ( .A1(n3935), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3758)
         );
  NAND2_X1 U4318 ( .A1(n4185), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3765)
         );
  NAND2_X1 U4319 ( .A1(n3836), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3764) );
  AND2_X4 U4320 ( .A1(n3770), .A2(n4989), .ZN(n4451) );
  NAND2_X1 U4321 ( .A1(n4451), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4322 ( .A1(n3670), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3762) );
  NAND2_X1 U4323 ( .A1(n3668), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3769) );
  NAND2_X1 U4324 ( .A1(n3876), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3768)
         );
  NAND2_X1 U4325 ( .A1(n4388), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3767) );
  AND2_X4 U4326 ( .A1(n4989), .A2(n4975), .ZN(n4534) );
  NAND2_X1 U4327 ( .A1(n4534), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3766)
         );
  NAND2_X1 U4328 ( .A1(n4381), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3774) );
  AND2_X2 U4329 ( .A1(n4813), .A2(n4975), .ZN(n3875) );
  NAND2_X1 U4330 ( .A1(n3875), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3773)
         );
  NAND2_X1 U4331 ( .A1(n3877), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U4332 ( .A1(n4535), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3771)
         );
  NAND2_X1 U4333 ( .A1(n3935), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3781)
         );
  NAND2_X1 U4334 ( .A1(n3836), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3780) );
  NAND2_X1 U4335 ( .A1(n3672), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3779) );
  NAND3_X1 U4336 ( .A1(n3781), .A2(n3780), .A3(n3779), .ZN(n3782) );
  NAND2_X1 U4337 ( .A1(n4534), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3785)
         );
  NAND2_X1 U4338 ( .A1(n3876), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3784)
         );
  NAND2_X1 U4339 ( .A1(n3669), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3783) );
  NAND3_X1 U4340 ( .A1(n3785), .A2(n3784), .A3(n3783), .ZN(n3786) );
  NOR2_X1 U4341 ( .A1(n3746), .A2(n3786), .ZN(n3792) );
  NAND2_X1 U4342 ( .A1(n4535), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3789)
         );
  NAND2_X1 U4343 ( .A1(n3877), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3788) );
  NAND3_X1 U4344 ( .A1(n3789), .A2(n3788), .A3(n3787), .ZN(n3790) );
  NOR2_X1 U4345 ( .A1(n3745), .A2(n3790), .ZN(n3791) );
  AND3_X2 U4346 ( .A1(n3793), .A2(n3792), .A3(n3791), .ZN(n3799) );
  NAND2_X1 U4347 ( .A1(n4388), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3797) );
  NAND2_X1 U4348 ( .A1(n4515), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3796) );
  NAND2_X1 U4349 ( .A1(n3675), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U4350 ( .A1(n3667), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4351 ( .A1(n4451), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4352 ( .A1(n3666), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4353 ( .A1(n3836), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3670), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4354 ( .A1(n3669), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4355 ( .A1(n3876), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4535), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4356 ( .A1(n4185), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4357 ( .A1(n3935), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3670), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4358 ( .A1(n4515), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4359 ( .A1(n3673), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3810) );
  AND4_X2 U4360 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3819)
         );
  AOI22_X1 U4361 ( .A1(n3666), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4362 ( .A1(n4185), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4363 ( .A1(n4393), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4364 ( .A1(n3877), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4535), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3814) );
  NAND2_X1 U4365 ( .A1(n3886), .A2(n3888), .ZN(n3831) );
  AOI22_X1 U4366 ( .A1(n3672), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4367 ( .A1(n4388), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4368 ( .A1(n3935), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3670), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4369 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3830)
         );
  AOI22_X1 U4370 ( .A1(n4185), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4371 ( .A1(n4381), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4372 ( .A1(n3877), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4535), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4373 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3829)
         );
  NAND2_X1 U4374 ( .A1(n4515), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U4375 ( .A1(n3675), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3833) );
  NAND2_X1 U4376 ( .A1(n4451), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3832) );
  NAND2_X1 U4377 ( .A1(n3672), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3840) );
  NAND2_X1 U4378 ( .A1(n3836), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4379 ( .A1(n3935), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3838)
         );
  NAND2_X1 U4380 ( .A1(n3670), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4381 ( .A1(n3668), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3844) );
  NAND2_X1 U4382 ( .A1(n3876), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3843)
         );
  NAND2_X1 U4383 ( .A1(n3666), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3842) );
  NAND2_X1 U4384 ( .A1(n4534), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3841)
         );
  NAND2_X1 U4385 ( .A1(n4185), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3848)
         );
  NAND2_X1 U4386 ( .A1(n3875), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3847)
         );
  NAND2_X1 U4387 ( .A1(n3877), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3846) );
  NAND2_X1 U4388 ( .A1(n4535), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3845)
         );
  NAND4_X4 U4389 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3889)
         );
  NAND2_X2 U4390 ( .A1(n3897), .A2(n5129), .ZN(n3885) );
  INV_X1 U4391 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6988) );
  XNOR2_X1 U4392 ( .A(n6988), .B(STATE_REG_2__SCAN_IN), .ZN(n3853) );
  NOR2_X1 U4393 ( .A1(n3864), .A2(n3853), .ZN(n3926) );
  NAND2_X1 U4394 ( .A1(n4653), .A2(n5129), .ZN(n4594) );
  AOI22_X1 U4395 ( .A1(n3935), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4396 ( .A1(n4185), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4397 ( .A1(n3666), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4398 ( .A1(n4515), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3836), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4399 ( .A1(n4451), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3877), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4400 ( .A1(n3876), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4535), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3859) );
  OAI211_X1 U4401 ( .C1(n3926), .C2(n4653), .A(n3907), .B(n3905), .ZN(n3866)
         );
  AOI21_X1 U4402 ( .B1(n6995), .B2(n3885), .A(n3866), .ZN(n3901) );
  AOI22_X1 U4403 ( .A1(n4388), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3873) );
  INV_X1 U4404 ( .A(n3674), .ZN(n3869) );
  NOR2_X1 U4405 ( .A1(n3869), .A2(n3868), .ZN(n3870) );
  AOI21_X1 U4406 ( .B1(n4515), .B2(INSTQUEUE_REG_1__2__SCAN_IN), .A(n3870), 
        .ZN(n3872) );
  AOI22_X1 U4407 ( .A1(n3935), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3670), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4408 ( .A1(n4185), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4409 ( .A1(n3668), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3876), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4410 ( .A1(n4381), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4411 ( .A1(n3877), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4535), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3878) );
  NAND2_X1 U4412 ( .A1(n4060), .A2(n3887), .ZN(n3884) );
  NOR2_X2 U4413 ( .A1(n3885), .A2(n3884), .ZN(n3919) );
  INV_X1 U4414 ( .A(n3919), .ZN(n3896) );
  NAND2_X1 U4415 ( .A1(n3886), .A2(n3900), .ZN(n3916) );
  OAI211_X1 U4416 ( .C1(n3916), .C2(n3923), .A(n3908), .B(n3947), .ZN(n3892)
         );
  INV_X1 U4417 ( .A(n3892), .ZN(n3895) );
  NAND2_X1 U4418 ( .A1(n4659), .A2(n3904), .ZN(n3893) );
  NAND2_X1 U4419 ( .A1(n3947), .A2(n3864), .ZN(n5269) );
  NAND2_X1 U4420 ( .A1(n3893), .A2(n5269), .ZN(n3894) );
  AOI21_X2 U4421 ( .B1(n3896), .B2(n3895), .A(n3894), .ZN(n3912) );
  INV_X1 U4422 ( .A(n3904), .ZN(n3898) );
  NAND2_X1 U4423 ( .A1(n3898), .A2(n5129), .ZN(n3899) );
  NAND2_X1 U4424 ( .A1(n3900), .A2(n3909), .ZN(n4826) );
  NAND3_X1 U4425 ( .A1(n3901), .A2(n3912), .A3(n4640), .ZN(n3902) );
  NAND2_X1 U4426 ( .A1(n7383), .A2(n7400), .ZN(n4641) );
  MUX2_X1 U4427 ( .A(n4638), .B(n4641), .S(n7502), .Z(n3903) );
  INV_X1 U4428 ( .A(n4792), .ZN(n3906) );
  NAND2_X1 U4429 ( .A1(n7383), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6979) );
  AOI21_X1 U4430 ( .B1(n3887), .B2(n3891), .A(n6979), .ZN(n3910) );
  NOR2_X1 U4431 ( .A1(n3909), .A2(n3891), .ZN(n3918) );
  NAND2_X1 U4432 ( .A1(n4884), .A2(n3918), .ZN(n5012) );
  INV_X1 U4433 ( .A(n3912), .ZN(n3913) );
  NAND2_X1 U4434 ( .A1(n4706), .A2(n5129), .ZN(n4717) );
  INV_X1 U4435 ( .A(n3968), .ZN(n3934) );
  AND2_X1 U4436 ( .A1(n4793), .A2(n3664), .ZN(n3917) );
  NAND2_X1 U4437 ( .A1(n3919), .A2(n3918), .ZN(n4759) );
  NAND2_X1 U4438 ( .A1(n4793), .A2(n5125), .ZN(n4773) );
  INV_X1 U4439 ( .A(n4773), .ZN(n3922) );
  NAND2_X1 U4440 ( .A1(n3922), .A2(n3921), .ZN(n4822) );
  INV_X1 U4441 ( .A(n4822), .ZN(n3925) );
  NAND2_X1 U4442 ( .A1(n3925), .A2(n3924), .ZN(n4865) );
  OAI211_X1 U4443 ( .C1(n6260), .C2(n3926), .A(n4821), .B(n4865), .ZN(n3927)
         );
  NAND2_X1 U4444 ( .A1(n3927), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3929) );
  INV_X1 U4445 ( .A(n4641), .ZN(n4022) );
  NAND2_X1 U4446 ( .A1(n7496), .A2(n7502), .ZN(n3928) );
  NAND2_X1 U4447 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3997) );
  INV_X1 U4448 ( .A(n4638), .ZN(n3999) );
  AOI22_X1 U4449 ( .A1(n4022), .A2(n5529), .B1(n3999), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3930) );
  OAI211_X1 U4450 ( .C1(n3996), .C2(n3757), .A(n3929), .B(n3930), .ZN(n3993)
         );
  INV_X1 U4451 ( .A(n3929), .ZN(n3932) );
  INV_X1 U4452 ( .A(n3930), .ZN(n3931) );
  NAND2_X1 U4453 ( .A1(n3932), .A2(n3751), .ZN(n3933) );
  NAND2_X1 U4454 ( .A1(n3993), .A2(n3933), .ZN(n3990) );
  AOI22_X1 U4455 ( .A1(n3668), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3939) );
  BUF_X1 U4456 ( .A(n3935), .Z(n4558) );
  AOI22_X1 U4457 ( .A1(n4558), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4458 ( .A1(n3676), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4459 ( .A1(n4185), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4460 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3945)
         );
  AOI22_X1 U4461 ( .A1(n4533), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4462 ( .A1(n4564), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4463 ( .A1(n3672), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4464 ( .A1(n4380), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4465 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3944)
         );
  NOR2_X1 U4466 ( .A1(n4003), .A2(n3948), .ZN(n3946) );
  INV_X1 U4467 ( .A(n3965), .ZN(n3963) );
  OR2_X1 U4468 ( .A1(n4002), .A2(n3948), .ZN(n3961) );
  AOI22_X1 U4469 ( .A1(n3668), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4470 ( .A1(n3678), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4471 ( .A1(n3676), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4472 ( .A1(n3672), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3949) );
  NAND4_X1 U4473 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3958)
         );
  AOI22_X1 U4474 ( .A1(n4558), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4475 ( .A1(n4185), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4476 ( .A1(n4380), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4477 ( .A1(n4497), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4478 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3957)
         );
  OR2_X1 U4479 ( .A1(n4003), .A2(n4720), .ZN(n3960) );
  NAND2_X1 U4480 ( .A1(n4622), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3959) );
  INV_X1 U4481 ( .A(n3964), .ZN(n3962) );
  NAND2_X1 U4482 ( .A1(n3963), .A2(n3962), .ZN(n3966) );
  NAND2_X1 U4483 ( .A1(n3965), .A2(n3964), .ZN(n3989) );
  INV_X1 U4484 ( .A(n4048), .ZN(n3988) );
  OAI21_X1 U4485 ( .B1(n3967), .B2(n3969), .A(n3991), .ZN(n4062) );
  INV_X1 U4486 ( .A(n4720), .ZN(n3985) );
  AOI22_X1 U4487 ( .A1(n4380), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4488 ( .A1(n4558), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4489 ( .A1(n4533), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4490 ( .A1(n4565), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4491 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3979)
         );
  AOI22_X1 U4492 ( .A1(n3677), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4493 ( .A1(n4497), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4494 ( .A1(n3678), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4495 ( .A1(n3668), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U4496 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3978)
         );
  XNOR2_X1 U4497 ( .A(n3985), .B(n4660), .ZN(n3981) );
  INV_X1 U4498 ( .A(n4003), .ZN(n3980) );
  NAND2_X1 U4499 ( .A1(n3981), .A2(n3980), .ZN(n4057) );
  INV_X1 U4500 ( .A(n4660), .ZN(n3984) );
  NAND2_X1 U4501 ( .A1(n4622), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3983) );
  AOI21_X1 U4502 ( .B1(n5129), .B2(n4720), .A(n7400), .ZN(n3982) );
  OAI211_X1 U4503 ( .C1(n3984), .C2(n3891), .A(n3983), .B(n3982), .ZN(n4055)
         );
  OR2_X1 U4504 ( .A1(n4003), .A2(n3985), .ZN(n3986) );
  NAND2_X1 U4505 ( .A1(n4059), .A2(n3986), .ZN(n4047) );
  INV_X1 U4506 ( .A(n4047), .ZN(n3987) );
  INV_X1 U4507 ( .A(n3990), .ZN(n3992) );
  NAND2_X1 U4508 ( .A1(n3992), .A2(n3991), .ZN(n3995) );
  NAND2_X1 U4510 ( .A1(n3995), .A2(n3994), .ZN(n4016) );
  INV_X1 U4511 ( .A(n3997), .ZN(n7485) );
  AND2_X1 U4512 ( .A1(n7485), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5449)
         );
  INV_X1 U4513 ( .A(n5449), .ZN(n4019) );
  NAND2_X1 U4514 ( .A1(n3997), .A2(n7363), .ZN(n3998) );
  AND2_X1 U4515 ( .A1(n4019), .A2(n3998), .ZN(n5117) );
  AOI22_X1 U4516 ( .A1(n5117), .A2(n4022), .B1(n3999), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4000) );
  INV_X1 U4517 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n7560) );
  AOI22_X1 U4518 ( .A1(n3667), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4519 ( .A1(n3673), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4520 ( .A1(n3675), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3676), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4521 ( .A1(n4380), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4004) );
  NAND4_X1 U4522 ( .A1(n4007), .A2(n4006), .A3(n4005), .A4(n4004), .ZN(n4013)
         );
  AOI22_X1 U4523 ( .A1(n4565), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4524 ( .A1(n3668), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4525 ( .A1(n3935), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4526 ( .A1(n4381), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4008) );
  NAND4_X1 U4527 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4012)
         );
  NAND2_X1 U4528 ( .A1(n4632), .A2(n4669), .ZN(n4014) );
  OAI21_X1 U4529 ( .B1(n4603), .B2(n7560), .A(n4014), .ZN(n4015) );
  NOR2_X2 U4530 ( .A1(n4073), .A2(n4071), .ZN(n4037) );
  INV_X1 U4531 ( .A(n4016), .ZN(n4018) );
  NAND2_X1 U4532 ( .A1(n5449), .A2(n7364), .ZN(n7461) );
  NAND2_X1 U4533 ( .A1(n4019), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4020) );
  NAND2_X1 U4534 ( .A1(n7461), .A2(n4020), .ZN(n5195) );
  NOR2_X1 U4535 ( .A1(n4638), .A2(n7364), .ZN(n4021) );
  AOI21_X1 U4536 ( .B1(n5195), .B2(n4022), .A(n4021), .ZN(n4023) );
  XNOR2_X2 U4537 ( .A(n4978), .B(n4976), .ZN(n7460) );
  AOI22_X1 U4538 ( .A1(n3678), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4539 ( .A1(n3672), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4540 ( .A1(n3677), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4541 ( .A1(n3935), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4025) );
  NAND4_X1 U4542 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4034)
         );
  AOI22_X1 U4543 ( .A1(n3668), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4544 ( .A1(n4565), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4031) );
  INV_X1 U4545 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n7578) );
  AOI22_X1 U4546 ( .A1(n3666), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4547 ( .A1(n4497), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U4548 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4033)
         );
  AOI22_X1 U4549 ( .A1(n4632), .A2(n4680), .B1(n4622), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4035) );
  INV_X1 U4550 ( .A(n4037), .ZN(n4038) );
  INV_X1 U4551 ( .A(n5145), .ZN(n5042) );
  NOR2_X2 U4552 ( .A1(n3888), .A2(n7505), .ZN(n4270) );
  NAND2_X1 U4553 ( .A1(n3924), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4098) );
  INV_X1 U4554 ( .A(n4068), .ZN(n4040) );
  INV_X1 U4555 ( .A(n4093), .ZN(n4043) );
  INV_X1 U4556 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U4557 ( .A1(n4041), .A2(n4068), .ZN(n4042) );
  NAND2_X1 U4558 ( .A1(n4043), .A2(n4042), .ZN(n5290) );
  AOI22_X1 U4559 ( .A1(n5290), .A2(n3628), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U4560 ( .A1(n4482), .A2(EAX_REG_3__SCAN_IN), .ZN(n4044) );
  OAI211_X1 U4561 ( .C1(n4098), .C2(n4994), .A(n4045), .B(n4044), .ZN(n4046)
         );
  INV_X1 U4562 ( .A(n4920), .ZN(n4080) );
  NAND2_X1 U4563 ( .A1(n4048), .A2(n4047), .ZN(n4049) );
  NAND2_X1 U4564 ( .A1(n4651), .A2(n4270), .ZN(n4054) );
  AOI22_X1 U4565 ( .A1(n4063), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n7505), .ZN(n4053) );
  NAND2_X1 U4566 ( .A1(n4051), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4052) );
  INV_X1 U4567 ( .A(n4055), .ZN(n4056) );
  NAND2_X1 U4568 ( .A1(n4057), .A2(n4056), .ZN(n4058) );
  INV_X1 U4569 ( .A(n4060), .ZN(n4061) );
  INV_X1 U4570 ( .A(n4270), .ZN(n4126) );
  OR2_X1 U4571 ( .A1(n4062), .A2(n4126), .ZN(n4067) );
  AOI22_X1 U4572 ( .A1(n4063), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n7505), .ZN(n4065) );
  NAND2_X1 U4573 ( .A1(n4051), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4064) );
  AND2_X1 U4574 ( .A1(n4065), .A2(n4064), .ZN(n4066) );
  NAND2_X1 U4575 ( .A1(n4067), .A2(n4066), .ZN(n4776) );
  OAI21_X1 U4576 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n4068), .ZN(n7152) );
  AOI22_X1 U4577 ( .A1(n4582), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3628), 
        .B2(n7152), .ZN(n4070) );
  NAND2_X1 U4578 ( .A1(n4482), .A2(EAX_REG_2__SCAN_IN), .ZN(n4069) );
  OAI211_X1 U4579 ( .C1(n4098), .C2(n6248), .A(n4070), .B(n4069), .ZN(n4075)
         );
  NAND2_X1 U4580 ( .A1(n4783), .A2(n4075), .ZN(n4074) );
  INV_X1 U4581 ( .A(n4071), .ZN(n4072) );
  AOI21_X1 U4582 ( .B1(n4666), .B2(n4270), .A(n4582), .ZN(n4971) );
  NAND2_X1 U4583 ( .A1(n4074), .A2(n4971), .ZN(n4078) );
  INV_X1 U4584 ( .A(n4783), .ZN(n4077) );
  INV_X1 U4585 ( .A(n4075), .ZN(n4076) );
  NAND2_X1 U4586 ( .A1(n4078), .A2(n4969), .ZN(n4917) );
  NAND2_X1 U4587 ( .A1(n4080), .A2(n4079), .ZN(n4889) );
  AOI22_X1 U4588 ( .A1(n3678), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U4589 ( .A1(n3673), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4590 ( .A1(n3677), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U4591 ( .A1(n3935), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4081) );
  NAND4_X1 U4592 ( .A1(n4084), .A2(n4083), .A3(n4082), .A4(n4081), .ZN(n4090)
         );
  AOI22_X1 U4593 ( .A1(n3668), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4594 ( .A1(n4565), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4595 ( .A1(n4381), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U4596 ( .A1(n4497), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4085) );
  NAND4_X1 U4597 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4089)
         );
  NAND2_X1 U4598 ( .A1(n4632), .A2(n4689), .ZN(n4092) );
  NAND2_X1 U4599 ( .A1(n4622), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4091) );
  NAND2_X1 U4600 ( .A1(n4092), .A2(n4091), .ZN(n4102) );
  NOR2_X1 U4601 ( .A1(n4093), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4094)
         );
  NOR2_X1 U4602 ( .A1(n4118), .A2(n4094), .ZN(n7170) );
  INV_X1 U4603 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4097) );
  NAND2_X1 U4604 ( .A1(n7505), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4096)
         );
  NAND2_X1 U4605 ( .A1(n4482), .A2(EAX_REG_4__SCAN_IN), .ZN(n4095) );
  OAI211_X1 U4606 ( .C1(n4098), .C2(n4097), .A(n4096), .B(n4095), .ZN(n4099)
         );
  NAND2_X1 U4607 ( .A1(n4099), .A2(n4581), .ZN(n4100) );
  OAI21_X1 U4608 ( .B1(n7170), .B2(n4581), .A(n4100), .ZN(n4101) );
  INV_X1 U4609 ( .A(n4102), .ZN(n4115) );
  AOI22_X1 U4610 ( .A1(n3935), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U4611 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n4185), .B1(n3672), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U4612 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n4380), .B1(n3676), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U4613 ( .A1(n4540), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4103) );
  NAND4_X1 U4614 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4112)
         );
  AOI22_X1 U4615 ( .A1(n3668), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U4616 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n3678), .B1(n4451), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U4617 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n4564), .B1(n4497), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U4618 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n3666), .B1(n4559), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4107) );
  NAND4_X1 U4619 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4111)
         );
  AOI22_X1 U4620 ( .A1(n4632), .A2(n4692), .B1(INSTQUEUE_REG_0__5__SCAN_IN), 
        .B2(n4622), .ZN(n4114) );
  INV_X1 U4621 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n7181) );
  INV_X1 U4622 ( .A(n4582), .ZN(n4123) );
  INV_X1 U4623 ( .A(n4150), .ZN(n4121) );
  INV_X1 U4624 ( .A(n4118), .ZN(n4119) );
  NAND2_X1 U4625 ( .A1(n4119), .A2(n7181), .ZN(n4120) );
  NAND2_X1 U4626 ( .A1(n4121), .A2(n4120), .ZN(n7195) );
  NAND2_X1 U4627 ( .A1(n7195), .A2(n3628), .ZN(n4122) );
  OAI21_X1 U4628 ( .B1(n7181), .B2(n4123), .A(n4122), .ZN(n4124) );
  AOI21_X1 U4629 ( .B1(n4482), .B2(EAX_REG_5__SCAN_IN), .A(n4124), .ZN(n4125)
         );
  NAND2_X1 U4630 ( .A1(n4890), .A2(n4959), .ZN(n4958) );
  INV_X1 U4631 ( .A(n4958), .ZN(n4142) );
  AOI22_X1 U4632 ( .A1(n3678), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U4633 ( .A1(n3673), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U4634 ( .A1(n3676), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U4635 ( .A1(n3935), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4127) );
  NAND4_X1 U4636 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(n4136)
         );
  AOI22_X1 U4637 ( .A1(n4393), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U4638 ( .A1(n4185), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U4639 ( .A1(n4381), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U4640 ( .A1(n4497), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4131) );
  NAND4_X1 U4641 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4135)
         );
  AOI22_X1 U4642 ( .A1(n4632), .A2(n4709), .B1(n4622), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4144) );
  NAND2_X1 U4643 ( .A1(n4143), .A2(n4144), .ZN(n4699) );
  XNOR2_X1 U4644 ( .A(n4150), .B(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n7199) );
  INV_X1 U4645 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4138) );
  INV_X1 U4646 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4137) );
  OAI22_X1 U4647 ( .A1(n4579), .A2(n4138), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4137), .ZN(n4139) );
  MUX2_X1 U4648 ( .A(n7199), .B(n4139), .S(n4581), .Z(n4140) );
  INV_X1 U4649 ( .A(n4144), .ZN(n4145) );
  INV_X1 U4650 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n7683) );
  NAND2_X1 U4651 ( .A1(n4632), .A2(n4720), .ZN(n4147) );
  OAI21_X1 U4652 ( .B1(n4603), .B2(n7683), .A(n4147), .ZN(n4148) );
  INV_X1 U4653 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4155) );
  INV_X1 U4654 ( .A(n4171), .ZN(n4153) );
  NAND2_X1 U4655 ( .A1(n4150), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4151)
         );
  INV_X1 U4656 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n7208) );
  NAND2_X1 U4657 ( .A1(n4151), .A2(n7208), .ZN(n4152) );
  NAND2_X1 U4658 ( .A1(n4153), .A2(n4152), .ZN(n7216) );
  AOI22_X1 U4659 ( .A1(n7216), .A2(n3628), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4154) );
  OAI21_X1 U4660 ( .B1(n4579), .B2(n4155), .A(n4154), .ZN(n4156) );
  AOI22_X1 U4661 ( .A1(n3669), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U4662 ( .A1(n4558), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U4663 ( .A1(n4533), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U4664 ( .A1(n3678), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4157) );
  NAND4_X1 U4665 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4166)
         );
  AOI22_X1 U4666 ( .A1(n4380), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4667 ( .A1(n4565), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U4668 ( .A1(n3677), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U4669 ( .A1(n3666), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4161) );
  NAND4_X1 U4670 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), .ZN(n4165)
         );
  OAI21_X1 U4671 ( .B1(n4166), .B2(n4165), .A(n4270), .ZN(n4170) );
  NAND2_X1 U4672 ( .A1(n4482), .A2(EAX_REG_8__SCAN_IN), .ZN(n4169) );
  XNOR2_X1 U4673 ( .A(n4171), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U4674 ( .A1(n5367), .A2(n3628), .ZN(n4168) );
  NAND2_X1 U4675 ( .A1(n4582), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4167)
         );
  NAND4_X1 U4676 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n5352)
         );
  XOR2_X1 U4677 ( .A(n5443), .B(n4184), .Z(n5603) );
  AOI22_X1 U4678 ( .A1(n4482), .A2(EAX_REG_9__SCAN_IN), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U4679 ( .A1(n4380), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U4680 ( .A1(n4558), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U4681 ( .A1(n3678), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U4682 ( .A1(n3667), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4172) );
  NAND4_X1 U4683 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4181)
         );
  AOI22_X1 U4684 ( .A1(n4565), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U4685 ( .A1(n4564), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U4686 ( .A1(n3673), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U4687 ( .A1(n3668), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4176) );
  NAND4_X1 U4688 ( .A1(n4179), .A2(n4178), .A3(n4177), .A4(n4176), .ZN(n4180)
         );
  OAI21_X1 U4689 ( .B1(n4181), .B2(n4180), .A(n4270), .ZN(n4182) );
  OAI211_X1 U4690 ( .C1(n5603), .C2(n4581), .A(n4183), .B(n4182), .ZN(n5377)
         );
  XNOR2_X1 U4691 ( .A(n4201), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5644)
         );
  AOI22_X1 U4692 ( .A1(n4380), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4185), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U4693 ( .A1(n3672), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U4694 ( .A1(n3669), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U4695 ( .A1(n4558), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4186) );
  NAND4_X1 U4696 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4195)
         );
  AOI22_X1 U4697 ( .A1(n3678), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U4698 ( .A1(n3677), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U4699 ( .A1(n4564), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U4700 ( .A1(n4559), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4190) );
  NAND4_X1 U4701 ( .A1(n4193), .A2(n4192), .A3(n4191), .A4(n4190), .ZN(n4194)
         );
  OAI21_X1 U4702 ( .B1(n4195), .B2(n4194), .A(n4270), .ZN(n4198) );
  NAND2_X1 U4703 ( .A1(n4482), .A2(EAX_REG_10__SCAN_IN), .ZN(n4197) );
  NAND2_X1 U4704 ( .A1(n4582), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4196)
         );
  NAND3_X1 U4705 ( .A1(n4198), .A2(n4197), .A3(n4196), .ZN(n4199) );
  AOI21_X1 U4706 ( .B1(n5644), .B2(n3628), .A(n4199), .ZN(n5424) );
  XOR2_X1 U4707 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4215), .Z(n5665) );
  AOI22_X1 U4708 ( .A1(n4482), .A2(EAX_REG_11__SCAN_IN), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U4709 ( .A1(n4393), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U4710 ( .A1(n4565), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U4711 ( .A1(n4533), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U4712 ( .A1(n4564), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4202) );
  NAND4_X1 U4713 ( .A1(n4205), .A2(n4204), .A3(n4203), .A4(n4202), .ZN(n4211)
         );
  AOI22_X1 U4714 ( .A1(n3673), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U4715 ( .A1(n3678), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U4716 ( .A1(n4558), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U4717 ( .A1(n4381), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4206) );
  NAND4_X1 U4718 ( .A1(n4209), .A2(n4208), .A3(n4207), .A4(n4206), .ZN(n4210)
         );
  OAI21_X1 U4719 ( .B1(n4211), .B2(n4210), .A(n4270), .ZN(n4212) );
  OAI211_X1 U4720 ( .C1(n5665), .C2(n4581), .A(n4213), .B(n4212), .ZN(n5575)
         );
  INV_X1 U4721 ( .A(n5575), .ZN(n4214) );
  XNOR2_X1 U4722 ( .A(n4244), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n7228)
         );
  NAND2_X1 U4723 ( .A1(n7228), .A2(n3628), .ZN(n4220) );
  INV_X1 U4724 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4218) );
  INV_X1 U4725 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n7223) );
  AOI21_X1 U4726 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n7223), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4216) );
  INV_X1 U4727 ( .A(n4216), .ZN(n4217) );
  OAI21_X1 U4728 ( .B1(n4579), .B2(n4218), .A(n4217), .ZN(n4219) );
  NAND2_X1 U4729 ( .A1(n4220), .A2(n4219), .ZN(n4232) );
  AOI22_X1 U4730 ( .A1(n3669), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U4731 ( .A1(n4380), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4223) );
  AOI22_X1 U4732 ( .A1(n3672), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U4733 ( .A1(n4558), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4221) );
  NAND4_X1 U4734 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(n4230)
         );
  AOI22_X1 U4735 ( .A1(n4565), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U4736 ( .A1(n4533), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4227) );
  AOI22_X1 U4737 ( .A1(n3678), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4226) );
  AOI22_X1 U4738 ( .A1(n4564), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4225) );
  NAND4_X1 U4739 ( .A1(n4228), .A2(n4227), .A3(n4226), .A4(n4225), .ZN(n4229)
         );
  OAI21_X1 U4740 ( .B1(n4230), .B2(n4229), .A(n4270), .ZN(n4231) );
  NAND2_X1 U4741 ( .A1(n4232), .A2(n4231), .ZN(n5650) );
  AOI22_X1 U4742 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n4558), .B1(n3673), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U4743 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n4533), .B1(n3667), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U4744 ( .A1(n3666), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U4745 ( .A1(n3668), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4233) );
  NAND4_X1 U4746 ( .A1(n4236), .A2(n4235), .A3(n4234), .A4(n4233), .ZN(n4242)
         );
  AOI22_X1 U4747 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n4185), .B1(n4564), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U4748 ( .A1(n3678), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U4749 ( .A1(n4380), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U4750 ( .A1(n3675), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4237) );
  NAND4_X1 U4751 ( .A1(n4240), .A2(n4239), .A3(n4238), .A4(n4237), .ZN(n4241)
         );
  OR2_X1 U4752 ( .A1(n4242), .A2(n4241), .ZN(n4243) );
  AND2_X1 U4753 ( .A1(n4270), .A2(n4243), .ZN(n4248) );
  NAND2_X1 U4754 ( .A1(n4063), .A2(EAX_REG_13__SCAN_IN), .ZN(n4247) );
  OAI21_X1 U4755 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4245), .A(n4261), 
        .ZN(n7236) );
  AOI22_X1 U4756 ( .A1(n3628), .A2(n7236), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4246) );
  NAND2_X1 U4757 ( .A1(n4247), .A2(n4246), .ZN(n5671) );
  INV_X1 U4758 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n7246) );
  XOR2_X1 U4759 ( .A(n7246), .B(n4261), .Z(n7248) );
  AOI22_X1 U4760 ( .A1(n4482), .A2(EAX_REG_14__SCAN_IN), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4260) );
  AOI22_X1 U4761 ( .A1(n3678), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U4762 ( .A1(n3677), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4763 ( .A1(n4564), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U4764 ( .A1(n3666), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4249) );
  NAND4_X1 U4765 ( .A1(n4252), .A2(n4251), .A3(n4250), .A4(n4249), .ZN(n4258)
         );
  AOI22_X1 U4766 ( .A1(n4393), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U4767 ( .A1(n3672), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U4768 ( .A1(n4565), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U4769 ( .A1(n4558), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4253) );
  NAND4_X1 U4770 ( .A1(n4256), .A2(n4255), .A3(n4254), .A4(n4253), .ZN(n4257)
         );
  OAI21_X1 U4771 ( .B1(n4258), .B2(n4257), .A(n4270), .ZN(n4259) );
  OAI211_X1 U4772 ( .C1(n7248), .C2(n4581), .A(n4260), .B(n4259), .ZN(n6450)
         );
  XNOR2_X1 U4773 ( .A(n4278), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6585)
         );
  AOI22_X1 U4774 ( .A1(n3673), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4265) );
  AOI22_X1 U4775 ( .A1(n3668), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4264) );
  AOI22_X1 U4776 ( .A1(n4558), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U4777 ( .A1(n4381), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4262) );
  NAND4_X1 U4778 ( .A1(n4265), .A2(n4264), .A3(n4263), .A4(n4262), .ZN(n4272)
         );
  AOI22_X1 U4779 ( .A1(n4565), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4269) );
  AOI22_X1 U4780 ( .A1(n3678), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U4781 ( .A1(n3676), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U4782 ( .A1(n4380), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4266) );
  NAND4_X1 U4783 ( .A1(n4269), .A2(n4268), .A3(n4267), .A4(n4266), .ZN(n4271)
         );
  OAI21_X1 U4784 ( .B1(n4272), .B2(n4271), .A(n4270), .ZN(n4275) );
  NAND2_X1 U4785 ( .A1(n4063), .A2(EAX_REG_15__SCAN_IN), .ZN(n4274) );
  NAND2_X1 U4786 ( .A1(n4582), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4273)
         );
  NAND3_X1 U4787 ( .A1(n4275), .A2(n4274), .A3(n4273), .ZN(n4276) );
  AOI21_X1 U4788 ( .B1(n6585), .B2(n3628), .A(n4276), .ZN(n6376) );
  INV_X1 U4789 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n7260) );
  NAND2_X1 U4790 ( .A1(n4278), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4293)
         );
  XOR2_X1 U4791 ( .A(n7260), .B(n4293), .Z(n7255) );
  INV_X1 U4792 ( .A(n7255), .ZN(n6579) );
  AOI22_X1 U4793 ( .A1(n4380), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4282) );
  AOI22_X1 U4794 ( .A1(n4558), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U4795 ( .A1(n4565), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4280) );
  AOI22_X1 U4796 ( .A1(n4393), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4279) );
  NAND4_X1 U4797 ( .A1(n4282), .A2(n4281), .A3(n4280), .A4(n4279), .ZN(n4288)
         );
  AOI22_X1 U4798 ( .A1(n3678), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4286) );
  AOI22_X1 U4799 ( .A1(n3666), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4285) );
  AOI22_X1 U4800 ( .A1(n3677), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U4801 ( .A1(n4533), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4283) );
  NAND4_X1 U4802 ( .A1(n4286), .A2(n4285), .A3(n4284), .A4(n4283), .ZN(n4287)
         );
  NOR2_X1 U4803 ( .A1(n4288), .A2(n4287), .ZN(n4290) );
  AOI22_X1 U4804 ( .A1(n4063), .A2(EAX_REG_16__SCAN_IN), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4289) );
  OAI21_X1 U4805 ( .B1(n4525), .B2(n4290), .A(n4289), .ZN(n4291) );
  AOI21_X1 U4806 ( .B1(n6579), .B2(n3628), .A(n4291), .ZN(n6442) );
  XNOR2_X1 U4807 ( .A(n4324), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7271)
         );
  NAND2_X1 U4808 ( .A1(n7271), .A2(n3628), .ZN(n4308) );
  AOI22_X1 U4809 ( .A1(n3678), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4297) );
  AOI22_X1 U4810 ( .A1(n4558), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3673), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4296) );
  AOI22_X1 U4811 ( .A1(n4393), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4381), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U4812 ( .A1(n4564), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4294) );
  NAND4_X1 U4813 ( .A1(n4297), .A2(n4296), .A3(n4295), .A4(n4294), .ZN(n4303)
         );
  AOI22_X1 U4814 ( .A1(n3676), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4301) );
  AOI22_X1 U4815 ( .A1(n4565), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4300) );
  AOI22_X1 U4816 ( .A1(n3675), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4299) );
  AOI22_X1 U4817 ( .A1(n4380), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4298) );
  NAND4_X1 U4818 ( .A1(n4301), .A2(n4300), .A3(n4299), .A4(n4298), .ZN(n4302)
         );
  NOR2_X1 U4819 ( .A1(n4303), .A2(n4302), .ZN(n4306) );
  INV_X1 U4820 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7269) );
  AOI21_X1 U4821 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n7269), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4304) );
  AOI21_X1 U4822 ( .B1(n4482), .B2(EAX_REG_17__SCAN_IN), .A(n4304), .ZN(n4305)
         );
  OAI21_X1 U4823 ( .B1(n4525), .B2(n4306), .A(n4305), .ZN(n4307) );
  NAND2_X1 U4824 ( .A1(n4308), .A2(n4307), .ZN(n6436) );
  AOI22_X1 U4825 ( .A1(n3668), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4313) );
  AOI22_X1 U4826 ( .A1(n4533), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U4827 ( .A1(n3678), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4311) );
  AOI22_X1 U4828 ( .A1(n3666), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4310) );
  NAND4_X1 U4829 ( .A1(n4313), .A2(n4312), .A3(n4311), .A4(n4310), .ZN(n4319)
         );
  AOI22_X1 U4830 ( .A1(n4565), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U4831 ( .A1(n4380), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4316) );
  AOI22_X1 U4832 ( .A1(n4564), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4315) );
  AOI22_X1 U4833 ( .A1(n4558), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4314) );
  NAND4_X1 U4834 ( .A1(n4317), .A2(n4316), .A3(n4315), .A4(n4314), .ZN(n4318)
         );
  NOR2_X1 U4835 ( .A1(n4319), .A2(n4318), .ZN(n4323) );
  NAND2_X1 U4836 ( .A1(n7505), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4320)
         );
  NAND2_X1 U4837 ( .A1(n4581), .A2(n4320), .ZN(n4321) );
  AOI21_X1 U4838 ( .B1(n4482), .B2(EAX_REG_18__SCAN_IN), .A(n4321), .ZN(n4322)
         );
  OAI21_X1 U4839 ( .B1(n4525), .B2(n4323), .A(n4322), .ZN(n4327) );
  OAI21_X1 U4840 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n4325), .A(n4357), 
        .ZN(n7288) );
  OR2_X1 U4841 ( .A1(n4581), .A2(n7288), .ZN(n4326) );
  NAND2_X1 U4842 ( .A1(n4327), .A2(n4326), .ZN(n6429) );
  AOI22_X1 U4843 ( .A1(n3672), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U4844 ( .A1(n3678), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4330) );
  AOI22_X1 U4845 ( .A1(n4380), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U4846 ( .A1(n4558), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4328) );
  NAND4_X1 U4847 ( .A1(n4331), .A2(n4330), .A3(n4329), .A4(n4328), .ZN(n4337)
         );
  AOI22_X1 U4848 ( .A1(n4565), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4335) );
  AOI22_X1 U4849 ( .A1(n4533), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4334) );
  AOI22_X1 U4850 ( .A1(n3668), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U4851 ( .A1(n4381), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4332) );
  NAND4_X1 U4852 ( .A1(n4335), .A2(n4334), .A3(n4333), .A4(n4332), .ZN(n4336)
         );
  NOR2_X1 U4853 ( .A1(n4337), .A2(n4336), .ZN(n4340) );
  INV_X1 U4854 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n7293) );
  AOI21_X1 U4855 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n7293), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4338) );
  AOI21_X1 U4856 ( .B1(n4482), .B2(EAX_REG_19__SCAN_IN), .A(n4338), .ZN(n4339)
         );
  OAI21_X1 U4857 ( .B1(n4525), .B2(n4340), .A(n4339), .ZN(n4342) );
  XNOR2_X1 U4858 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4357), .ZN(n7300)
         );
  NAND2_X1 U4859 ( .A1(n7300), .A2(n3628), .ZN(n4341) );
  AOI22_X1 U4860 ( .A1(n3669), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U4861 ( .A1(n3672), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4345) );
  AOI22_X1 U4862 ( .A1(n4451), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U4863 ( .A1(n4558), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4343) );
  NAND4_X1 U4864 ( .A1(n4346), .A2(n4345), .A3(n4344), .A4(n4343), .ZN(n4352)
         );
  AOI22_X1 U4865 ( .A1(n3678), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U4866 ( .A1(n4185), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3676), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U4867 ( .A1(n4564), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4868 ( .A1(n3666), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4347) );
  NAND4_X1 U4869 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(n4351)
         );
  NOR2_X1 U4870 ( .A1(n4352), .A2(n4351), .ZN(n4356) );
  NAND2_X1 U4871 ( .A1(n7505), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4353)
         );
  NAND2_X1 U4872 ( .A1(n4581), .A2(n4353), .ZN(n4354) );
  AOI21_X1 U4873 ( .B1(n4482), .B2(EAX_REG_20__SCAN_IN), .A(n4354), .ZN(n4355)
         );
  OAI21_X1 U4874 ( .B1(n4525), .B2(n4356), .A(n4355), .ZN(n4364) );
  INV_X1 U4875 ( .A(n4485), .ZN(n4362) );
  INV_X1 U4876 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4360) );
  INV_X1 U4877 ( .A(n4358), .ZN(n4359) );
  NAND2_X1 U4878 ( .A1(n4360), .A2(n4359), .ZN(n4361) );
  NAND2_X1 U4879 ( .A1(n4362), .A2(n4361), .ZN(n7307) );
  OR2_X1 U4880 ( .A1(n7307), .A2(n4581), .ZN(n4363) );
  AOI22_X1 U4881 ( .A1(n4380), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4368) );
  AOI22_X1 U4882 ( .A1(n4185), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U4883 ( .A1(n3675), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4366) );
  AOI22_X1 U4884 ( .A1(n4497), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4365) );
  NAND4_X1 U4885 ( .A1(n4368), .A2(n4367), .A3(n4366), .A4(n4365), .ZN(n4375)
         );
  AOI22_X1 U4886 ( .A1(n3672), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U4887 ( .A1(n3678), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4372) );
  AOI22_X1 U4888 ( .A1(n3669), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4371) );
  AOI22_X1 U4889 ( .A1(n3935), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4370) );
  NAND4_X1 U4890 ( .A1(n4373), .A2(n4372), .A3(n4371), .A4(n4370), .ZN(n4374)
         );
  NOR2_X1 U4891 ( .A1(n4375), .A2(n4374), .ZN(n4439) );
  AOI22_X1 U4892 ( .A1(n3678), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4379) );
  AOI22_X1 U4893 ( .A1(n3672), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U4894 ( .A1(n3677), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U4895 ( .A1(n3935), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4376) );
  NAND4_X1 U4896 ( .A1(n4379), .A2(n4378), .A3(n4377), .A4(n4376), .ZN(n4387)
         );
  AOI22_X1 U4897 ( .A1(n4393), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U4898 ( .A1(n4565), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4384) );
  AOI22_X1 U4899 ( .A1(n4381), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U4900 ( .A1(n4497), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4382) );
  NAND4_X1 U4901 ( .A1(n4385), .A2(n4384), .A3(n4383), .A4(n4382), .ZN(n4386)
         );
  OR2_X1 U4902 ( .A1(n4387), .A2(n4386), .ZN(n4445) );
  AOI22_X1 U4903 ( .A1(n3678), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U4904 ( .A1(n3672), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U4905 ( .A1(n3676), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U4906 ( .A1(n3935), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4389) );
  NAND4_X1 U4907 ( .A1(n4392), .A2(n4391), .A3(n4390), .A4(n4389), .ZN(n4399)
         );
  AOI22_X1 U4908 ( .A1(n3668), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4397) );
  AOI22_X1 U4909 ( .A1(n4185), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U4910 ( .A1(n4381), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4395) );
  AOI22_X1 U4911 ( .A1(n4497), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4394) );
  NAND4_X1 U4912 ( .A1(n4397), .A2(n4396), .A3(n4395), .A4(n4394), .ZN(n4398)
         );
  OR2_X1 U4913 ( .A1(n4399), .A2(n4398), .ZN(n4444) );
  NAND2_X1 U4914 ( .A1(n4445), .A2(n4444), .ZN(n4440) );
  NOR2_X1 U4915 ( .A1(n4439), .A2(n4440), .ZN(n4438) );
  AOI22_X1 U4916 ( .A1(n3678), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4403) );
  AOI22_X1 U4917 ( .A1(n3672), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4402) );
  AOI22_X1 U4918 ( .A1(n3676), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3667), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U4919 ( .A1(n4558), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4400) );
  NAND4_X1 U4920 ( .A1(n4403), .A2(n4402), .A3(n4401), .A4(n4400), .ZN(n4409)
         );
  AOI22_X1 U4921 ( .A1(n3669), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U4922 ( .A1(n4185), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U4923 ( .A1(n3666), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U4924 ( .A1(n4497), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4404) );
  NAND4_X1 U4925 ( .A1(n4407), .A2(n4406), .A3(n4405), .A4(n4404), .ZN(n4408)
         );
  OR2_X1 U4926 ( .A1(n4409), .A2(n4408), .ZN(n4430) );
  NAND2_X1 U4927 ( .A1(n4438), .A2(n4430), .ZN(n4491) );
  AOI22_X1 U4928 ( .A1(n3669), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U4929 ( .A1(n4533), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4412) );
  AOI22_X1 U4930 ( .A1(n4185), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U4931 ( .A1(n4558), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4410) );
  NAND4_X1 U4932 ( .A1(n4413), .A2(n4412), .A3(n4411), .A4(n4410), .ZN(n4419)
         );
  AOI22_X1 U4933 ( .A1(n3673), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4417) );
  AOI22_X1 U4934 ( .A1(n4380), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4416) );
  AOI22_X1 U4935 ( .A1(n3677), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U4936 ( .A1(n3666), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4414) );
  NAND4_X1 U4937 ( .A1(n4417), .A2(n4416), .A3(n4415), .A4(n4414), .ZN(n4418)
         );
  NOR2_X1 U4938 ( .A1(n4419), .A2(n4418), .ZN(n4492) );
  XNOR2_X1 U4939 ( .A(n4491), .B(n4492), .ZN(n4423) );
  NAND2_X1 U4940 ( .A1(n7505), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4420)
         );
  NAND2_X1 U4941 ( .A1(n4581), .A2(n4420), .ZN(n4421) );
  AOI21_X1 U4942 ( .B1(n4482), .B2(EAX_REG_26__SCAN_IN), .A(n4421), .ZN(n4422)
         );
  OAI21_X1 U4943 ( .B1(n4423), .B2(n4525), .A(n4422), .ZN(n4429) );
  INV_X1 U4944 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6552) );
  INV_X1 U4945 ( .A(n4425), .ZN(n4426) );
  INV_X1 U4946 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U4947 ( .A1(n4426), .A2(n6511), .ZN(n4427) );
  AND2_X1 U4948 ( .A1(n4527), .A2(n4427), .ZN(n6509) );
  NAND2_X1 U4949 ( .A1(n6509), .A2(n3628), .ZN(n4428) );
  NAND2_X1 U4950 ( .A1(n4429), .A2(n4428), .ZN(n6322) );
  INV_X1 U4951 ( .A(n6322), .ZN(n4489) );
  XNOR2_X1 U4952 ( .A(n4430), .B(n4438), .ZN(n4433) );
  INV_X1 U4953 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6517) );
  AOI21_X1 U4954 ( .B1(n6517), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4431) );
  AOI21_X1 U4955 ( .B1(n4482), .B2(EAX_REG_25__SCAN_IN), .A(n4431), .ZN(n4432)
         );
  OAI21_X1 U4956 ( .B1(n4525), .B2(n4433), .A(n4432), .ZN(n4436) );
  XNOR2_X1 U4957 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4434), .ZN(n6521)
         );
  NAND2_X1 U4958 ( .A1(n3628), .A2(n6521), .ZN(n4435) );
  AND2_X1 U4959 ( .A1(n4436), .A2(n4435), .ZN(n6336) );
  INV_X1 U4960 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6530) );
  XNOR2_X1 U4961 ( .A(n4437), .B(n6530), .ZN(n7340) );
  INV_X1 U4962 ( .A(n4525), .ZN(n4574) );
  AOI21_X1 U4963 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(n4441) );
  NAND2_X1 U4964 ( .A1(n4574), .A2(n4441), .ZN(n4443) );
  AOI22_X1 U4965 ( .A1(n4482), .A2(EAX_REG_24__SCAN_IN), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4442) );
  OAI211_X1 U4966 ( .C1(n7340), .C2(n4581), .A(n4443), .B(n4442), .ZN(n6532)
         );
  INV_X1 U4967 ( .A(n6532), .ZN(n4470) );
  XNOR2_X1 U4968 ( .A(n4445), .B(n4444), .ZN(n4448) );
  INV_X1 U4969 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6544) );
  OAI21_X1 U4970 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6544), .A(n4581), .ZN(
        n4446) );
  AOI21_X1 U4971 ( .B1(n4063), .B2(EAX_REG_23__SCAN_IN), .A(n4446), .ZN(n4447)
         );
  OAI21_X1 U4972 ( .B1(n4525), .B2(n4448), .A(n4447), .ZN(n4450) );
  XNOR2_X1 U4973 ( .A(n4467), .B(n6544), .ZN(n6542) );
  NAND2_X1 U4974 ( .A1(n6542), .A2(n3628), .ZN(n4449) );
  NAND2_X1 U4975 ( .A1(n4450), .A2(n4449), .ZN(n6352) );
  AOI22_X1 U4976 ( .A1(n4451), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4455) );
  AOI22_X1 U4977 ( .A1(n3673), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4454) );
  AOI22_X1 U4978 ( .A1(n3675), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3676), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4453) );
  AOI22_X1 U4979 ( .A1(n4381), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4452) );
  NAND4_X1 U4980 ( .A1(n4455), .A2(n4454), .A3(n4453), .A4(n4452), .ZN(n4461)
         );
  AOI22_X1 U4981 ( .A1(n4185), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4459) );
  AOI22_X1 U4982 ( .A1(n4380), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U4983 ( .A1(n4558), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4457) );
  AOI22_X1 U4984 ( .A1(n3668), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4456) );
  NAND4_X1 U4985 ( .A1(n4459), .A2(n4458), .A3(n4457), .A4(n4456), .ZN(n4460)
         );
  NOR2_X1 U4986 ( .A1(n4461), .A2(n4460), .ZN(n4464) );
  OAI21_X1 U4987 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6552), .A(n4581), .ZN(
        n4462) );
  AOI21_X1 U4988 ( .B1(n4482), .B2(EAX_REG_22__SCAN_IN), .A(n4462), .ZN(n4463)
         );
  OAI21_X1 U4989 ( .B1(n4525), .B2(n4464), .A(n4463), .ZN(n4469) );
  AND2_X1 U4990 ( .A1(n4465), .A2(n6552), .ZN(n4466) );
  NOR2_X1 U4991 ( .A1(n4467), .A2(n4466), .ZN(n7322) );
  NAND2_X1 U4992 ( .A1(n7322), .A2(n3628), .ZN(n4468) );
  NAND2_X1 U4993 ( .A1(n4469), .A2(n4468), .ZN(n6397) );
  OR2_X1 U4994 ( .A1(n6352), .A2(n6397), .ZN(n6350) );
  NOR2_X1 U4995 ( .A1(n4470), .A2(n6350), .ZN(n6333) );
  AND2_X1 U4996 ( .A1(n6336), .A2(n6333), .ZN(n4488) );
  AOI22_X1 U4997 ( .A1(n4393), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U4998 ( .A1(n3672), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U4999 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n3667), .B1(n4564), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5000 ( .A1(n4497), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4471) );
  NAND4_X1 U5001 ( .A1(n4474), .A2(n4473), .A3(n4472), .A4(n4471), .ZN(n4480)
         );
  AOI22_X1 U5002 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n4533), .B1(n3675), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4478) );
  AOI22_X1 U5003 ( .A1(n4185), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3676), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4477) );
  AOI22_X1 U5004 ( .A1(n4380), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4476) );
  AOI22_X1 U5005 ( .A1(n4558), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4475) );
  NAND4_X1 U5006 ( .A1(n4478), .A2(n4477), .A3(n4476), .A4(n4475), .ZN(n4479)
         );
  NOR2_X1 U5007 ( .A1(n4480), .A2(n4479), .ZN(n4484) );
  INV_X1 U5008 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6559) );
  OAI21_X1 U5009 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6559), .A(n4581), .ZN(
        n4481) );
  AOI21_X1 U5010 ( .B1(n4482), .B2(EAX_REG_21__SCAN_IN), .A(n4481), .ZN(n4483)
         );
  OAI21_X1 U5011 ( .B1(n4525), .B2(n4484), .A(n4483), .ZN(n4487) );
  XNOR2_X1 U5012 ( .A(n4485), .B(n6559), .ZN(n6561) );
  NAND2_X1 U5013 ( .A1(n6561), .A2(n3628), .ZN(n4486) );
  NOR2_X1 U5014 ( .A1(n4492), .A2(n4491), .ZN(n4510) );
  AOI22_X1 U5015 ( .A1(n3678), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3675), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4496) );
  AOI22_X1 U5016 ( .A1(n3673), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5017 ( .A1(n3677), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4494) );
  AOI22_X1 U5018 ( .A1(n4558), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4493) );
  NAND4_X1 U5019 ( .A1(n4496), .A2(n4495), .A3(n4494), .A4(n4493), .ZN(n4503)
         );
  AOI22_X1 U5020 ( .A1(n3669), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5021 ( .A1(n4185), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5022 ( .A1(n4381), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5023 ( .A1(n4497), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4559), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4498) );
  NAND4_X1 U5024 ( .A1(n4501), .A2(n4500), .A3(n4499), .A4(n4498), .ZN(n4502)
         );
  OR2_X1 U5025 ( .A1(n4503), .A2(n4502), .ZN(n4509) );
  XNOR2_X1 U5026 ( .A(n4510), .B(n4509), .ZN(n4506) );
  INV_X1 U5027 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6503) );
  OAI21_X1 U5028 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6503), .A(n4581), .ZN(
        n4504) );
  AOI21_X1 U5029 ( .B1(n4063), .B2(EAX_REG_27__SCAN_IN), .A(n4504), .ZN(n4505)
         );
  OAI21_X1 U5030 ( .B1(n4506), .B2(n4525), .A(n4505), .ZN(n4508) );
  XNOR2_X1 U5031 ( .A(n4527), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6506)
         );
  NAND2_X1 U5032 ( .A1(n6506), .A2(n3628), .ZN(n4507) );
  NAND2_X1 U5033 ( .A1(n4508), .A2(n4507), .ZN(n6305) );
  NAND2_X1 U5034 ( .A1(n4510), .A2(n4509), .ZN(n4547) );
  AOI22_X1 U5035 ( .A1(n3669), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U5036 ( .A1(n4185), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4451), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4513) );
  AOI22_X1 U5037 ( .A1(n4497), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4535), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4512) );
  AOI22_X1 U5038 ( .A1(n3673), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4511) );
  NAND4_X1 U5039 ( .A1(n4514), .A2(n4513), .A3(n4512), .A4(n4511), .ZN(n4521)
         );
  AOI22_X1 U5040 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n3678), .B1(n3675), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4519) );
  AOI22_X1 U5041 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n4533), .B1(n4558), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4518) );
  AOI22_X1 U5042 ( .A1(n3676), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4517) );
  AOI22_X1 U5043 ( .A1(n3666), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4516) );
  NAND4_X1 U5044 ( .A1(n4519), .A2(n4518), .A3(n4517), .A4(n4516), .ZN(n4520)
         );
  NOR2_X1 U5045 ( .A1(n4521), .A2(n4520), .ZN(n4548) );
  XNOR2_X1 U5046 ( .A(n4547), .B(n4548), .ZN(n4526) );
  NAND2_X1 U5047 ( .A1(n7505), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4522)
         );
  NAND2_X1 U5048 ( .A1(n4581), .A2(n4522), .ZN(n4523) );
  AOI21_X1 U5049 ( .B1(n4063), .B2(EAX_REG_28__SCAN_IN), .A(n4523), .ZN(n4524)
         );
  OAI21_X1 U5050 ( .B1(n4526), .B2(n4525), .A(n4524), .ZN(n4532) );
  NAND2_X1 U5051 ( .A1(n4528), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4554)
         );
  INV_X1 U5052 ( .A(n4528), .ZN(n4529) );
  INV_X1 U5053 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U5054 ( .A1(n4529), .A2(n6297), .ZN(n4530) );
  NAND2_X1 U5055 ( .A1(n4554), .A2(n4530), .ZN(n6496) );
  AOI22_X1 U5056 ( .A1(n4185), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3678), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5057 ( .A1(n3673), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5058 ( .A1(n4381), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4537) );
  AOI22_X1 U5059 ( .A1(n4497), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4535), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4536) );
  NAND4_X1 U5060 ( .A1(n4539), .A2(n4538), .A3(n4537), .A4(n4536), .ZN(n4546)
         );
  AOI22_X1 U5061 ( .A1(n4393), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4380), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4544) );
  AOI22_X1 U5062 ( .A1(n3667), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3875), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U5063 ( .A1(n3675), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3676), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4542) );
  AOI22_X1 U5064 ( .A1(n4558), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4541) );
  NAND4_X1 U5065 ( .A1(n4544), .A2(n4543), .A3(n4542), .A4(n4541), .ZN(n4545)
         );
  NOR2_X1 U5066 ( .A1(n4546), .A2(n4545), .ZN(n4556) );
  OR2_X1 U5067 ( .A1(n4548), .A2(n4547), .ZN(n4557) );
  XOR2_X1 U5068 ( .A(n4556), .B(n4557), .Z(n4549) );
  NAND2_X1 U5069 ( .A1(n4549), .A2(n4574), .ZN(n4553) );
  INV_X1 U5070 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5822) );
  AOI21_X1 U5071 ( .B1(n5822), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4550) );
  AOI21_X1 U5072 ( .B1(n4063), .B2(EAX_REG_29__SCAN_IN), .A(n4550), .ZN(n4552)
         );
  XNOR2_X1 U5073 ( .A(n4554), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6283)
         );
  AND2_X1 U5074 ( .A1(n6283), .A2(n3628), .ZN(n4551) );
  AOI21_X1 U5075 ( .B1(n4553), .B2(n4552), .A(n4551), .ZN(n5824) );
  INV_X1 U5076 ( .A(n4554), .ZN(n4555) );
  XNOR2_X1 U5077 ( .A(n4646), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6488)
         );
  INV_X1 U5078 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4578) );
  NOR2_X1 U5079 ( .A1(n4557), .A2(n4556), .ZN(n4573) );
  AOI22_X1 U5080 ( .A1(n3678), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4533), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5081 ( .A1(n4558), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5082 ( .A1(n4559), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4534), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U5083 ( .A1(n4451), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4560) );
  NAND4_X1 U5084 ( .A1(n4563), .A2(n4562), .A3(n4561), .A4(n4560), .ZN(n4571)
         );
  AOI22_X1 U5085 ( .A1(n3668), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3666), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5086 ( .A1(n4380), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4564), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5087 ( .A1(n4565), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4567) );
  AOI22_X1 U5088 ( .A1(n3675), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4540), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4566) );
  NAND4_X1 U5089 ( .A1(n4569), .A2(n4568), .A3(n4567), .A4(n4566), .ZN(n4570)
         );
  NOR2_X1 U5090 ( .A1(n4571), .A2(n4570), .ZN(n4572) );
  XNOR2_X1 U5091 ( .A(n4573), .B(n4572), .ZN(n4575) );
  NAND2_X1 U5092 ( .A1(n4575), .A2(n4574), .ZN(n4577) );
  AOI21_X1 U5093 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n7505), .A(n3628), 
        .ZN(n4576) );
  OAI211_X1 U5094 ( .C1(n4579), .C2(n4578), .A(n4577), .B(n4576), .ZN(n4580)
         );
  OAI21_X1 U5095 ( .B1(n4581), .B2(n6488), .A(n4580), .ZN(n6273) );
  AOI22_X1 U5096 ( .A1(n4063), .A2(EAX_REG_31__SCAN_IN), .B1(n4582), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4583) );
  NOR2_X2 U5097 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7499) );
  NOR2_X1 U5098 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5266), .ZN(n5261) );
  NAND2_X1 U5099 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5261), .ZN(n6991) );
  INV_X1 U5100 ( .A(n6991), .ZN(n4584) );
  AND2_X2 U5101 ( .A1(n7499), .A2(n4584), .ZN(n6970) );
  XNOR2_X1 U5102 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4600) );
  NAND2_X1 U5103 ( .A1(n4599), .A2(n4600), .ZN(n4586) );
  NAND2_X1 U5104 ( .A1(n7496), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U5105 ( .A1(n4586), .A2(n4585), .ZN(n4590) );
  XNOR2_X1 U5106 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U5107 ( .A1(n4590), .A2(n4589), .ZN(n4588) );
  NAND2_X1 U5108 ( .A1(n7363), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4587) );
  NAND2_X1 U5109 ( .A1(n4588), .A2(n4587), .ZN(n4619) );
  XNOR2_X1 U5110 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4618) );
  XNOR2_X1 U5111 ( .A(n4619), .B(n4618), .ZN(n4754) );
  NAND2_X1 U5112 ( .A1(n4603), .A2(n4754), .ZN(n4617) );
  XNOR2_X1 U5113 ( .A(n4590), .B(n4589), .ZN(n4753) );
  NAND2_X1 U5114 ( .A1(n5139), .A2(n4653), .ZN(n4591) );
  NAND2_X1 U5115 ( .A1(n6261), .A2(n4591), .ZN(n4611) );
  AOI21_X1 U5116 ( .B1(n4622), .B2(n4753), .A(n4611), .ZN(n4615) );
  AND2_X1 U5117 ( .A1(n7354), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4592)
         );
  NOR2_X1 U5118 ( .A1(n4599), .A2(n4592), .ZN(n4595) );
  NAND2_X1 U5119 ( .A1(n4632), .A2(n4595), .ZN(n4593) );
  NAND2_X1 U5120 ( .A1(n4623), .A2(n4593), .ZN(n4598) );
  AOI21_X1 U5121 ( .B1(n4594), .B2(n4595), .A(n3947), .ZN(n4596) );
  NAND2_X1 U5122 ( .A1(n4598), .A2(n4597), .ZN(n4607) );
  XNOR2_X1 U5123 ( .A(n4600), .B(n4599), .ZN(n4752) );
  OR2_X1 U5124 ( .A1(n4752), .A2(n7400), .ZN(n4606) );
  INV_X1 U5125 ( .A(n4752), .ZN(n4602) );
  NAND2_X1 U5126 ( .A1(n4632), .A2(n3864), .ZN(n4601) );
  OAI211_X1 U5127 ( .C1(n4603), .C2(n4602), .A(n4601), .B(n4653), .ZN(n4604)
         );
  INV_X1 U5128 ( .A(n4604), .ZN(n4605) );
  OAI21_X1 U5129 ( .B1(n4607), .B2(n4606), .A(n4605), .ZN(n4609) );
  NAND3_X1 U5130 ( .A1(n4607), .A2(n4623), .A3(n4606), .ZN(n4608) );
  INV_X1 U5131 ( .A(n4612), .ZN(n4614) );
  INV_X1 U5132 ( .A(n4753), .ZN(n4610) );
  OAI211_X1 U5133 ( .C1(n4612), .C2(n4611), .A(n4610), .B(n4632), .ZN(n4613)
         );
  OAI21_X1 U5134 ( .B1(n4615), .B2(n4614), .A(n4613), .ZN(n4616) );
  AOI22_X1 U5135 ( .A1(n4617), .A2(n4616), .B1(n4635), .B2(n4754), .ZN(n4625)
         );
  NAND2_X1 U5136 ( .A1(n4619), .A2(n4618), .ZN(n4621) );
  NAND2_X1 U5137 ( .A1(n7364), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5138 ( .A1(n4621), .A2(n4620), .ZN(n4629) );
  INV_X1 U5139 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4628) );
  NOR2_X1 U5140 ( .A1(n4622), .A2(n4756), .ZN(n4624) );
  OAI22_X1 U5141 ( .A1(n4625), .A2(n4624), .B1(n4623), .B2(n4756), .ZN(n4626)
         );
  AOI21_X1 U5142 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7400), .A(n4626), 
        .ZN(n4634) );
  NAND2_X1 U5143 ( .A1(n4627), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U5144 ( .A1(n4629), .A2(n4628), .ZN(n4630) );
  NAND2_X1 U5145 ( .A1(n4631), .A2(n4630), .ZN(n4751) );
  NAND2_X1 U5146 ( .A1(n4632), .A2(n4751), .ZN(n4633) );
  NAND2_X1 U5147 ( .A1(n4634), .A2(n4633), .ZN(n4637) );
  NAND2_X1 U5148 ( .A1(n4635), .A2(n4751), .ZN(n4636) );
  NAND2_X1 U5149 ( .A1(n3904), .A2(n3947), .ZN(n4639) );
  NAND2_X1 U5150 ( .A1(n4640), .A2(n4639), .ZN(n4771) );
  OR2_X1 U5151 ( .A1(n4771), .A2(n4594), .ZN(n4864) );
  INV_X1 U5152 ( .A(n7499), .ZN(n7511) );
  NAND2_X1 U5153 ( .A1(n7511), .A2(n4641), .ZN(n6998) );
  NAND2_X1 U5154 ( .A1(n6998), .A2(n7400), .ZN(n4642) );
  NAND2_X1 U5155 ( .A1(n7400), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4644) );
  INV_X1 U5156 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7497) );
  NAND2_X1 U5157 ( .A1(n7497), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4643) );
  AND2_X1 U5158 ( .A1(n4644), .A2(n4643), .ZN(n4807) );
  INV_X1 U5159 ( .A(n4807), .ZN(n4645) );
  NAND2_X1 U5160 ( .A1(n4646), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4648)
         );
  INV_X1 U5161 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4647) );
  XNOR2_X1 U5162 ( .A(n4648), .B(n4647), .ZN(n5277) );
  AND2_X1 U5163 ( .A1(n7499), .A2(n5266), .ZN(n6982) );
  AND2_X2 U5164 ( .A1(n6982), .A2(n7400), .ZN(n7073) );
  INV_X1 U5165 ( .A(n7073), .ZN(n7136) );
  INV_X1 U5166 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6880) );
  NOR2_X1 U5167 ( .A1(n7136), .A2(n6880), .ZN(n5802) );
  AOI21_X1 U5168 ( .B1(n6969), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5802), 
        .ZN(n4649) );
  OAI21_X1 U5169 ( .B1(n6975), .B2(n5277), .A(n4649), .ZN(n4650) );
  AOI21_X1 U5170 ( .B1(n5775), .B2(n6970), .A(n4650), .ZN(n4750) );
  NAND2_X1 U5171 ( .A1(n3679), .A2(n4706), .ZN(n4658) );
  NAND2_X1 U5172 ( .A1(n4660), .A2(n4652), .ZN(n4671) );
  OAI21_X1 U5173 ( .B1(n4660), .B2(n4652), .A(n4671), .ZN(n4655) );
  INV_X1 U5174 ( .A(n4826), .ZN(n4654) );
  OAI211_X1 U5175 ( .C1(n4655), .C2(n5778), .A(n4654), .B(n4653), .ZN(n4656)
         );
  INV_X1 U5176 ( .A(n4656), .ZN(n4657) );
  INV_X1 U5177 ( .A(n4706), .ZN(n4772) );
  INV_X1 U5178 ( .A(n4659), .ZN(n4663) );
  OAI21_X1 U5179 ( .B1(n5778), .B2(n4660), .A(n4663), .ZN(n4661) );
  INV_X1 U5180 ( .A(n4661), .ZN(n4662) );
  OAI21_X1 U5181 ( .B1(n3662), .B2(n4772), .A(n4662), .ZN(n4806) );
  NAND2_X1 U5182 ( .A1(n4806), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6712)
         );
  NAND2_X1 U5183 ( .A1(n6710), .A2(n6712), .ZN(n4667) );
  NAND3_X1 U5184 ( .A1(n4667), .A2(n6711), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6932) );
  XNOR2_X1 U5185 ( .A(n4671), .B(n4669), .ZN(n4664) );
  OAI21_X1 U5186 ( .B1(n4664), .B2(n5778), .A(n4663), .ZN(n4665) );
  NAND2_X1 U5187 ( .A1(n4667), .A2(n3647), .ZN(n4668) );
  INV_X1 U5188 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4897) );
  INV_X1 U5189 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4676) );
  NAND2_X1 U5190 ( .A1(n5526), .A2(n4706), .ZN(n4675) );
  INV_X1 U5191 ( .A(n4669), .ZN(n4670) );
  NAND2_X1 U5192 ( .A1(n4671), .A2(n4670), .ZN(n4681) );
  INV_X1 U5193 ( .A(n4680), .ZN(n4672) );
  XNOR2_X1 U5194 ( .A(n4681), .B(n4672), .ZN(n4673) );
  NAND2_X1 U5195 ( .A1(n4673), .A2(n6995), .ZN(n4674) );
  AND2_X1 U5196 ( .A1(n4675), .A2(n4674), .ZN(n4914) );
  NAND2_X1 U5197 ( .A1(n4912), .A2(n4914), .ZN(n4678) );
  NAND2_X1 U5198 ( .A1(n4677), .A2(n4676), .ZN(n4913) );
  NAND2_X1 U5199 ( .A1(n4679), .A2(n4706), .ZN(n4684) );
  NAND2_X1 U5200 ( .A1(n4681), .A2(n4680), .ZN(n4691) );
  XNOR2_X1 U5201 ( .A(n4691), .B(n4689), .ZN(n4682) );
  NAND2_X1 U5202 ( .A1(n4682), .A2(n6995), .ZN(n4683) );
  INV_X1 U5203 ( .A(n4685), .ZN(n4686) );
  INV_X1 U5204 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n7021) );
  OAI22_X1 U5205 ( .A1(n4963), .A2(n4964), .B1(n4686), .B2(n7021), .ZN(n6939)
         );
  INV_X1 U5206 ( .A(n4687), .ZN(n4688) );
  NAND2_X1 U5207 ( .A1(n4688), .A2(n4706), .ZN(n4695) );
  INV_X1 U5208 ( .A(n4689), .ZN(n4690) );
  NOR2_X1 U5209 ( .A1(n4691), .A2(n4690), .ZN(n4693) );
  NAND2_X1 U5210 ( .A1(n4693), .A2(n4692), .ZN(n4708) );
  OAI211_X1 U5211 ( .C1(n4693), .C2(n4692), .A(n4708), .B(n6995), .ZN(n4694)
         );
  NAND2_X1 U5212 ( .A1(n4695), .A2(n4694), .ZN(n4696) );
  INV_X1 U5213 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U5214 ( .A1(n6939), .A2(n6940), .ZN(n4698) );
  NAND2_X1 U5215 ( .A1(n4696), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4697)
         );
  NAND2_X1 U5216 ( .A1(n4698), .A2(n4697), .ZN(n6945) );
  NAND3_X1 U5217 ( .A1(n4719), .A2(n4706), .A3(n4699), .ZN(n4702) );
  XNOR2_X1 U5218 ( .A(n4708), .B(n4709), .ZN(n4700) );
  NAND2_X1 U5219 ( .A1(n4700), .A2(n6995), .ZN(n4701) );
  AND2_X1 U5220 ( .A1(n4702), .A2(n4701), .ZN(n4703) );
  INV_X1 U5221 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U5222 ( .A1(n6945), .A2(n6947), .ZN(n4705) );
  INV_X1 U5223 ( .A(n4703), .ZN(n4704) );
  NAND2_X1 U5224 ( .A1(n4704), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6946)
         );
  NAND2_X1 U5225 ( .A1(n4705), .A2(n6946), .ZN(n6952) );
  NAND2_X1 U5226 ( .A1(n4707), .A2(n4706), .ZN(n4713) );
  INV_X1 U5227 ( .A(n4708), .ZN(n4710) );
  NAND2_X1 U5228 ( .A1(n4710), .A2(n4709), .ZN(n4722) );
  XNOR2_X1 U5229 ( .A(n4722), .B(n4720), .ZN(n4711) );
  NAND2_X1 U5230 ( .A1(n4711), .A2(n6995), .ZN(n4712) );
  NAND2_X1 U5231 ( .A1(n4713), .A2(n4712), .ZN(n4714) );
  INV_X1 U5232 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n7077) );
  XNOR2_X1 U5233 ( .A(n4714), .B(n7077), .ZN(n6954) );
  NAND2_X1 U5234 ( .A1(n4714), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4715)
         );
  NAND2_X1 U5235 ( .A1(n4720), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4716) );
  NOR2_X1 U5236 ( .A1(n4717), .A2(n4716), .ZN(n4718) );
  NAND2_X1 U5237 ( .A1(n6995), .A2(n4720), .ZN(n4721) );
  OR2_X1 U5238 ( .A1(n4722), .A2(n4721), .ZN(n4723) );
  NAND2_X1 U5239 ( .A1(n6549), .A2(n4723), .ZN(n4724) );
  INV_X1 U5240 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5348) );
  XNOR2_X1 U5241 ( .A(n6549), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5599)
         );
  INV_X1 U5242 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4725) );
  INV_X1 U5243 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4728) );
  NAND3_X1 U5244 ( .A1(n5703), .A2(n4728), .A3(n4727), .ZN(n4729) );
  INV_X1 U5245 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U5246 ( .A1(n6668), .A2(n5703), .ZN(n5702) );
  XNOR2_X1 U5247 ( .A(n6668), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6961)
         );
  INV_X1 U5248 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U5249 ( .A1(n6668), .A2(n7010), .ZN(n4730) );
  INV_X1 U5250 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U5251 ( .A1(n6668), .A2(n5697), .ZN(n4732) );
  INV_X1 U5252 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4733) );
  INV_X1 U5253 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U5254 ( .A1(n6668), .A2(n6707), .ZN(n6576) );
  NAND2_X1 U5255 ( .A1(n6575), .A2(n6576), .ZN(n6569) );
  INV_X1 U5256 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U5257 ( .A1(n6569), .A2(n3750), .ZN(n4735) );
  INV_X1 U5258 ( .A(n6569), .ZN(n4737) );
  NAND2_X1 U5259 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6674) );
  INV_X1 U5260 ( .A(n6674), .ZN(n4736) );
  AND2_X1 U5261 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6525) );
  AND2_X1 U5262 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U5263 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5808) );
  INV_X1 U5264 ( .A(n5808), .ZN(n4738) );
  NOR2_X1 U5265 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6676) );
  NOR2_X1 U5266 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6652) );
  INV_X1 U5267 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5748) );
  INV_X1 U5268 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6645) );
  INV_X1 U5269 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n7139) );
  NAND2_X1 U5270 ( .A1(n6515), .A2(n4739), .ZN(n4740) );
  AND2_X1 U5271 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5809) );
  NAND3_X1 U5272 ( .A1(n5809), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4743) );
  OAI21_X1 U5273 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6526), .ZN(n5815) );
  INV_X1 U5274 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6600) );
  NAND3_X1 U5275 ( .A1(n6526), .A2(n6483), .A3(n6600), .ZN(n4747) );
  INV_X1 U5276 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U5277 ( .A1(n6500), .A2(n3737), .ZN(n5816) );
  NAND4_X1 U5278 ( .A1(n6668), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A4(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n4746) );
  XNOR2_X1 U5279 ( .A(n4748), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5814)
         );
  NAND2_X1 U5280 ( .A1(n4750), .A2(n4749), .ZN(U2955) );
  INV_X1 U5281 ( .A(n4751), .ZN(n4758) );
  NOR3_X1 U5282 ( .A1(n4754), .A2(n4753), .A3(n4752), .ZN(n4755) );
  NAND2_X1 U5283 ( .A1(n4756), .A2(n4755), .ZN(n4757) );
  INV_X1 U5284 ( .A(n6258), .ZN(n4761) );
  INV_X1 U5285 ( .A(n7397), .ZN(n7377) );
  OR3_X1 U5286 ( .A1(n4761), .A2(n7377), .A3(n4760), .ZN(n5259) );
  INV_X1 U5287 ( .A(n5259), .ZN(n4762) );
  INV_X1 U5288 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7423) );
  INV_X1 U5289 ( .A(n6982), .ZN(n5368) );
  OAI211_X1 U5290 ( .C1(n4762), .C2(n7423), .A(n5260), .B(n5368), .ZN(U2788)
         );
  INV_X1 U5291 ( .A(n5772), .ZN(n4767) );
  INV_X1 U5292 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U5293 ( .A1(n5579), .A2(EBX_REG_0__SCAN_IN), .ZN(n4765) );
  INV_X1 U5294 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4778) );
  NAND2_X1 U5295 ( .A1(n5672), .A2(n4778), .ZN(n4764) );
  NAND2_X1 U5296 ( .A1(n4765), .A2(n4764), .ZN(n4789) );
  INV_X1 U5297 ( .A(n4789), .ZN(n4766) );
  AOI21_X1 U5298 ( .B1(n4767), .B2(n7062), .A(n4766), .ZN(n7143) );
  INV_X1 U5299 ( .A(n7143), .ZN(n4779) );
  NAND2_X1 U5300 ( .A1(n4768), .A2(n6995), .ZN(n4770) );
  NAND3_X1 U5301 ( .A1(n3885), .A2(n3891), .A3(n3904), .ZN(n4769) );
  NAND2_X1 U5302 ( .A1(n4770), .A2(n4769), .ZN(n4818) );
  NOR2_X1 U5303 ( .A1(n4771), .A2(n4818), .ZN(n4844) );
  OR2_X1 U5304 ( .A1(n5269), .A2(n3887), .ZN(n4825) );
  NOR2_X1 U5305 ( .A1(n3908), .A2(n4772), .ZN(n4836) );
  NAND2_X1 U5306 ( .A1(n4838), .A2(n4836), .ZN(n4988) );
  NAND3_X1 U5307 ( .A1(n5717), .A2(n5129), .A3(n3888), .ZN(n4951) );
  AND2_X4 U5308 ( .A1(n3891), .A2(n3864), .ZN(n6263) );
  OR3_X1 U5309 ( .A1(n4951), .A2(n4773), .A3(n4786), .ZN(n4774) );
  OAI21_X1 U5310 ( .B1(n6255), .B2(n4988), .A(n4774), .ZN(n4775) );
  XNOR2_X1 U5311 ( .A(n4777), .B(n4776), .ZN(n7149) );
  OAI222_X1 U5312 ( .A1(n4779), .A2(n6916), .B1(n4778), .B2(n6927), .C1(n6454), 
        .C2(n7149), .ZN(U2859) );
  NOR2_X1 U5313 ( .A1(n4781), .A2(n4780), .ZN(n4782) );
  NOR2_X1 U5314 ( .A1(n4783), .A2(n4782), .ZN(n6928) );
  INV_X1 U5315 ( .A(n6928), .ZN(n4957) );
  INV_X1 U5316 ( .A(n4763), .ZN(n4815) );
  OR2_X1 U5317 ( .A1(n5763), .A2(EBX_REG_1__SCAN_IN), .ZN(n4788) );
  NAND2_X1 U5318 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4784)
         );
  NAND2_X1 U5319 ( .A1(n5579), .A2(n4784), .ZN(n4785) );
  OAI21_X1 U5320 ( .B1(EBX_REG_1__SCAN_IN), .B2(n4786), .A(n4785), .ZN(n4787)
         );
  NAND2_X1 U5321 ( .A1(n4788), .A2(n4787), .ZN(n4893) );
  XNOR2_X1 U5322 ( .A(n4893), .B(n4789), .ZN(n4790) );
  NAND2_X1 U5323 ( .A1(n4790), .A2(n6263), .ZN(n4894) );
  OAI21_X1 U5324 ( .B1(n4790), .B2(n6263), .A(n4894), .ZN(n6715) );
  AOI22_X1 U5325 ( .A1(n6924), .A2(n6715), .B1(EBX_REG_1__SCAN_IN), .B2(n6426), 
        .ZN(n4791) );
  OAI21_X1 U5326 ( .B1(n6454), .B2(n4957), .A(n4791), .ZN(U2858) );
  INV_X1 U5327 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4797) );
  AND2_X1 U5328 ( .A1(n4793), .A2(n4792), .ZN(n4859) );
  NAND2_X1 U5329 ( .A1(n4859), .A2(n6995), .ZN(n7380) );
  NOR2_X1 U5330 ( .A1(n4760), .A2(n5139), .ZN(n5007) );
  INV_X1 U5331 ( .A(n5007), .ZN(n7353) );
  OR2_X1 U5332 ( .A1(n4861), .A2(n7353), .ZN(n4794) );
  NAND2_X1 U5333 ( .A1(n5046), .A2(n4794), .ZN(n4795) );
  INV_X1 U5334 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6832) );
  INV_X1 U5335 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7415) );
  OAI221_X1 U5336 ( .B1(n6988), .B2(n6832), .C1(STATE_REG_1__SCAN_IN), .C2(
        STATE_REG_2__SCAN_IN), .A(n7415), .ZN(n6989) );
  INV_X1 U5337 ( .A(n6989), .ZN(n6264) );
  NAND2_X1 U5338 ( .A1(n6799), .A2(n3891), .ZN(n4949) );
  NAND2_X1 U5339 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5261), .ZN(n7376) );
  NOR2_X4 U5340 ( .A1(n6828), .A2(n6799), .ZN(n6812) );
  AOI22_X1 U5341 ( .A1(n6828), .A2(UWORD_REG_5__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4796) );
  OAI21_X1 U5342 ( .B1(n4797), .B2(n4949), .A(n4796), .ZN(U2902) );
  INV_X1 U5343 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U5344 ( .A1(n6828), .A2(UWORD_REG_6__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4798) );
  OAI21_X1 U5345 ( .B1(n4799), .B2(n4949), .A(n4798), .ZN(U2901) );
  INV_X1 U5346 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4801) );
  AOI22_X1 U5347 ( .A1(n6828), .A2(UWORD_REG_8__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4800) );
  OAI21_X1 U5348 ( .B1(n4801), .B2(n4949), .A(n4800), .ZN(U2899) );
  INV_X1 U5349 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4803) );
  AOI22_X1 U5350 ( .A1(n6828), .A2(UWORD_REG_7__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4802) );
  OAI21_X1 U5351 ( .B1(n4803), .B2(n4949), .A(n4802), .ZN(U2900) );
  INV_X1 U5352 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4805) );
  AOI22_X1 U5353 ( .A1(n6828), .A2(UWORD_REG_9__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4804) );
  OAI21_X1 U5354 ( .B1(n4805), .B2(n4949), .A(n4804), .ZN(U2898) );
  OAI21_X1 U5355 ( .B1(n4806), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6712), 
        .ZN(n4883) );
  NAND2_X1 U5356 ( .A1(n4807), .A2(n6965), .ZN(n4810) );
  INV_X1 U5357 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4808) );
  NOR2_X1 U5358 ( .A1(n7136), .A2(n4808), .ZN(n4880) );
  NOR2_X1 U5359 ( .A1(n7149), .A2(n6962), .ZN(n4809) );
  AOI211_X1 U5360 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4810), .A(n4880), 
        .B(n4809), .ZN(n4811) );
  OAI21_X1 U5361 ( .B1(n7345), .B2(n4883), .A(n4811), .ZN(U2986) );
  NOR2_X1 U5362 ( .A1(n4812), .A2(n4813), .ZN(n4834) );
  AND2_X1 U5363 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  NOR2_X1 U5364 ( .A1(n4818), .A2(n4817), .ZN(n4819) );
  AND2_X1 U5365 ( .A1(n4820), .A2(n4819), .ZN(n4873) );
  INV_X1 U5366 ( .A(n4859), .ZN(n4824) );
  NAND3_X1 U5367 ( .A1(n4824), .A2(n4823), .A3(n3907), .ZN(n4830) );
  INV_X1 U5368 ( .A(n4825), .ZN(n4827) );
  OAI21_X1 U5369 ( .B1(n4827), .B2(n5772), .A(n4826), .ZN(n4829) );
  OAI21_X1 U5370 ( .B1(n3923), .B2(n3664), .A(n3887), .ZN(n4828) );
  NAND2_X1 U5371 ( .A1(n4829), .A2(n4828), .ZN(n4871) );
  NOR2_X1 U5372 ( .A1(n4830), .A2(n4871), .ZN(n4831) );
  AND2_X1 U5373 ( .A1(n4821), .A2(n4831), .ZN(n4832) );
  NAND2_X1 U5374 ( .A1(n4873), .A2(n4832), .ZN(n5015) );
  NAND2_X1 U5375 ( .A1(n4814), .A2(n5015), .ZN(n4833) );
  NAND2_X1 U5376 ( .A1(n5007), .A2(n3757), .ZN(n5008) );
  OAI211_X1 U5377 ( .C1(n4834), .C2(n3908), .A(n4833), .B(n5008), .ZN(n7355)
         );
  INV_X1 U5378 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5811) );
  AOI22_X1 U5379 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5811), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3653), .ZN(n6243) );
  NOR2_X1 U5380 ( .A1(n5266), .A2(n7062), .ZN(n6241) );
  INV_X1 U5381 ( .A(n4834), .ZN(n4835) );
  INV_X1 U5382 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7390) );
  AOI222_X1 U5383 ( .A1(n7355), .A2(n7383), .B1(n6243), .B2(n6241), .C1(n4835), 
        .C2(n6721), .ZN(n4849) );
  INV_X1 U5384 ( .A(n4836), .ZN(n4837) );
  OR2_X1 U5385 ( .A1(n6255), .A2(n4837), .ZN(n4856) );
  INV_X1 U5386 ( .A(n4838), .ZN(n4842) );
  OAI21_X1 U5387 ( .B1(n5007), .B2(n4859), .A(n6264), .ZN(n4840) );
  NAND2_X1 U5388 ( .A1(n4859), .A2(n6263), .ZN(n4868) );
  INV_X1 U5389 ( .A(READY_N), .ZN(n7414) );
  NAND2_X1 U5390 ( .A1(n6255), .A2(n7414), .ZN(n4839) );
  AOI21_X1 U5391 ( .B1(n4840), .B2(n4868), .A(n4839), .ZN(n4841) );
  NOR2_X1 U5392 ( .A1(n4842), .A2(n4841), .ZN(n4843) );
  NAND2_X1 U5393 ( .A1(n4856), .A2(n4843), .ZN(n4847) );
  AND2_X1 U5394 ( .A1(n4844), .A2(n3921), .ZN(n4986) );
  NAND2_X1 U5395 ( .A1(n6255), .A2(n4986), .ZN(n4846) );
  NAND2_X1 U5396 ( .A1(n6258), .A2(n7414), .ZN(n4850) );
  OR2_X1 U5397 ( .A1(n4821), .A2(n4850), .ZN(n4845) );
  NAND2_X1 U5398 ( .A1(n4846), .A2(n4845), .ZN(n4953) );
  NOR2_X1 U5399 ( .A1(n7505), .A2(n5266), .ZN(n5253) );
  INV_X1 U5400 ( .A(n5253), .ZN(n7388) );
  NOR2_X1 U5401 ( .A1(n7400), .A2(n7388), .ZN(n6993) );
  INV_X1 U5402 ( .A(n6993), .ZN(n7389) );
  INV_X1 U5403 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7373) );
  OAI22_X1 U5404 ( .A1(n5004), .A2(n7377), .B1(n7389), .B2(n7373), .ZN(n7349)
         );
  AOI21_X1 U5405 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7400), .A(n7349), .ZN(
        n6250) );
  NAND2_X1 U5406 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n6250), .ZN(n4848) );
  OAI21_X1 U5407 ( .B1(n4849), .B2(n6250), .A(n4848), .ZN(U3460) );
  NAND2_X1 U5408 ( .A1(n3864), .A2(n6989), .ZN(n4852) );
  INV_X1 U5409 ( .A(n4850), .ZN(n4851) );
  NAND3_X1 U5410 ( .A1(n4852), .A2(n3887), .A3(n4851), .ZN(n4853) );
  AND2_X1 U5411 ( .A1(n4854), .A2(n4853), .ZN(n4855) );
  AOI21_X1 U5412 ( .B1(n4856), .B2(n4855), .A(n7377), .ZN(n4863) );
  NOR2_X1 U5413 ( .A1(n3864), .A2(n6264), .ZN(n5273) );
  NOR2_X1 U5414 ( .A1(n5273), .A2(READY_N), .ZN(n4858) );
  AOI21_X1 U5415 ( .B1(n3923), .B2(n3891), .A(n3887), .ZN(n4857) );
  AOI21_X1 U5416 ( .B1(n4859), .B2(n4858), .A(n4857), .ZN(n4860) );
  NOR2_X1 U5417 ( .A1(n4861), .A2(n4860), .ZN(n4862) );
  INV_X1 U5418 ( .A(n4864), .ZN(n7370) );
  NOR2_X1 U5419 ( .A1(n4986), .A2(n7370), .ZN(n6252) );
  INV_X1 U5420 ( .A(n4865), .ZN(n4866) );
  NAND2_X1 U5421 ( .A1(n4866), .A2(n3889), .ZN(n4867) );
  NAND4_X1 U5422 ( .A1(n6252), .A2(n4868), .A3(n4821), .A4(n4867), .ZN(n4869)
         );
  INV_X1 U5423 ( .A(n4988), .ZN(n6254) );
  OAI21_X1 U5424 ( .B1(n3907), .B2(n3664), .A(n5012), .ZN(n4870) );
  NOR2_X1 U5425 ( .A1(n4871), .A2(n4870), .ZN(n4872) );
  NAND2_X1 U5426 ( .A1(n4873), .A2(n4872), .ZN(n4874) );
  NAND2_X1 U5427 ( .A1(n4879), .A2(n4874), .ZN(n5344) );
  NAND2_X1 U5428 ( .A1(n7063), .A2(n5344), .ZN(n5686) );
  NAND2_X1 U5429 ( .A1(n4879), .A2(n5007), .ZN(n5688) );
  INV_X1 U5430 ( .A(n5688), .ZN(n7013) );
  INV_X1 U5431 ( .A(n5344), .ZN(n5684) );
  NAND2_X1 U5432 ( .A1(n5684), .A2(n7062), .ZN(n4877) );
  INV_X1 U5433 ( .A(n4879), .ZN(n4875) );
  NAND2_X1 U5434 ( .A1(n4875), .A2(n7136), .ZN(n4876) );
  OAI21_X1 U5435 ( .B1(n7063), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n7088), 
        .ZN(n6709) );
  OAI22_X1 U5436 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5686), .B1(n7013), 
        .B2(n6709), .ZN(n4882) );
  OAI21_X1 U5437 ( .B1(n4865), .B2(n3889), .A(n7380), .ZN(n4878) );
  AOI21_X1 U5438 ( .B1(n7132), .B2(n7143), .A(n4880), .ZN(n4881) );
  OAI211_X1 U5439 ( .C1(n7055), .C2(n4883), .A(n4882), .B(n4881), .ZN(U3018)
         );
  INV_X1 U5440 ( .A(n4062), .ZN(n5452) );
  AOI22_X1 U5441 ( .A1(n5452), .A2(n5015), .B1(n4884), .B2(n7354), .ZN(n7352)
         );
  INV_X1 U5442 ( .A(n7383), .ZN(n6723) );
  AOI22_X1 U5443 ( .A1(n7354), .A2(n6721), .B1(n7062), .B2(
        STATE2_REG_1__SCAN_IN), .ZN(n4885) );
  OAI21_X1 U5444 ( .B1(n7352), .B2(n6723), .A(n4885), .ZN(n4887) );
  INV_X1 U5445 ( .A(n6250), .ZN(n7351) );
  OAI21_X1 U5446 ( .B1(n7353), .B2(n6723), .A(n7351), .ZN(n4886) );
  AOI22_X1 U5447 ( .A1(n4887), .A2(n7351), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4886), .ZN(n4888) );
  INV_X1 U5448 ( .A(n4888), .ZN(U3461) );
  AOI21_X1 U5449 ( .B1(n4891), .B2(n4918), .A(n4890), .ZN(n4892) );
  INV_X1 U5450 ( .A(n4892), .ZN(n7173) );
  NAND2_X1 U5451 ( .A1(n4894), .A2(n4893), .ZN(n4927) );
  MUX2_X1 U5452 ( .A(n5745), .B(n5672), .S(EBX_REG_3__SCAN_IN), .Z(n4896) );
  OR2_X1 U5453 ( .A1(n5772), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4895)
         );
  AND2_X1 U5454 ( .A1(n4896), .A2(n4895), .ZN(n4928) );
  OR2_X1 U5455 ( .A1(n5763), .A2(EBX_REG_2__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U5456 ( .A1(n5579), .A2(n4897), .ZN(n4899) );
  INV_X1 U5457 ( .A(EBX_REG_2__SCAN_IN), .ZN(n7164) );
  NAND2_X1 U5458 ( .A1(n6263), .A2(n7164), .ZN(n4898) );
  NAND3_X1 U5459 ( .A1(n4899), .A2(n5672), .A3(n4898), .ZN(n4900) );
  NAND2_X1 U5460 ( .A1(n4901), .A2(n4900), .ZN(n6912) );
  NAND2_X1 U5461 ( .A1(n4928), .A2(n6912), .ZN(n4902) );
  OR2_X1 U5462 ( .A1(n5763), .A2(EBX_REG_4__SCAN_IN), .ZN(n4907) );
  NAND2_X1 U5463 ( .A1(n5579), .A2(n7021), .ZN(n4905) );
  INV_X1 U5464 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U5465 ( .A1(n6263), .A2(n4903), .ZN(n4904) );
  NAND3_X1 U5466 ( .A1(n4905), .A2(n5672), .A3(n4904), .ZN(n4906) );
  NAND2_X1 U5467 ( .A1(n4907), .A2(n4906), .ZN(n4908) );
  NAND2_X1 U5468 ( .A1(n4930), .A2(n4908), .ZN(n5031) );
  OR2_X1 U5469 ( .A1(n4930), .A2(n4908), .ZN(n4909) );
  NAND2_X1 U5470 ( .A1(n5031), .A2(n4909), .ZN(n7169) );
  INV_X1 U5471 ( .A(n7169), .ZN(n4910) );
  AOI22_X1 U5472 ( .A1(n6924), .A2(n4910), .B1(EBX_REG_4__SCAN_IN), .B2(n6426), 
        .ZN(n4911) );
  OAI21_X1 U5473 ( .B1(n7173), .B2(n6454), .A(n4911), .ZN(U2855) );
  NAND2_X1 U5474 ( .A1(n4912), .A2(n4913), .ZN(n4916) );
  INV_X1 U5475 ( .A(n4914), .ZN(n4915) );
  XNOR2_X1 U5476 ( .A(n4916), .B(n4915), .ZN(n7032) );
  INV_X1 U5477 ( .A(n7032), .ZN(n4924) );
  INV_X1 U5478 ( .A(n4918), .ZN(n4919) );
  AOI21_X1 U5479 ( .B1(n4920), .B2(n4917), .A(n4919), .ZN(n5289) );
  AOI22_X1 U5480 ( .A1(n6969), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n7073), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4921) );
  OAI21_X1 U5481 ( .B1(n5290), .B2(n6975), .A(n4921), .ZN(n4922) );
  AOI21_X1 U5482 ( .B1(n5289), .B2(n6970), .A(n4922), .ZN(n4923) );
  OAI21_X1 U5483 ( .B1(n4924), .B2(n7345), .A(n4923), .ZN(U2983) );
  INV_X1 U5484 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4926) );
  AOI22_X1 U5485 ( .A1(n6828), .A2(UWORD_REG_2__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4925) );
  OAI21_X1 U5486 ( .B1(n4926), .B2(n4949), .A(n4925), .ZN(U2905) );
  INV_X1 U5487 ( .A(n5289), .ZN(n4962) );
  INV_X1 U5488 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4932) );
  INV_X1 U5489 ( .A(n4927), .ZN(n4929) );
  AOI21_X1 U5490 ( .B1(n4929), .B2(n6912), .A(n4928), .ZN(n4931) );
  OR2_X1 U5491 ( .A1(n4931), .A2(n4930), .ZN(n7030) );
  OAI222_X1 U5492 ( .A1(n4962), .A2(n6454), .B1(n4932), .B2(n6927), .C1(n6916), 
        .C2(n7030), .ZN(U2856) );
  INV_X1 U5493 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U5494 ( .A1(n6828), .A2(UWORD_REG_0__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4933) );
  OAI21_X1 U5495 ( .B1(n4934), .B2(n4949), .A(n4933), .ZN(U2907) );
  AOI22_X1 U5496 ( .A1(n6828), .A2(UWORD_REG_14__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4935) );
  OAI21_X1 U5497 ( .B1(n4578), .B2(n4949), .A(n4935), .ZN(U2893) );
  INV_X1 U5498 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U5499 ( .A1(n6828), .A2(UWORD_REG_1__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4936) );
  OAI21_X1 U5500 ( .B1(n4937), .B2(n4949), .A(n4936), .ZN(U2906) );
  INV_X1 U5501 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4939) );
  AOI22_X1 U5502 ( .A1(n6828), .A2(UWORD_REG_3__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4938) );
  OAI21_X1 U5503 ( .B1(n4939), .B2(n4949), .A(n4938), .ZN(U2904) );
  INV_X1 U5504 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U5505 ( .A1(n6828), .A2(UWORD_REG_4__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4940) );
  OAI21_X1 U5506 ( .B1(n4941), .B2(n4949), .A(n4940), .ZN(U2903) );
  INV_X1 U5507 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4943) );
  AOI22_X1 U5508 ( .A1(n6828), .A2(UWORD_REG_10__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4942) );
  OAI21_X1 U5509 ( .B1(n4943), .B2(n4949), .A(n4942), .ZN(U2897) );
  INV_X1 U5510 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U5511 ( .A1(n6828), .A2(UWORD_REG_11__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4944) );
  OAI21_X1 U5512 ( .B1(n4945), .B2(n4949), .A(n4944), .ZN(U2896) );
  INV_X1 U5513 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4947) );
  AOI22_X1 U5514 ( .A1(n6828), .A2(UWORD_REG_12__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4946) );
  OAI21_X1 U5515 ( .B1(n4947), .B2(n4949), .A(n4946), .ZN(U2895) );
  INV_X1 U5516 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4950) );
  AOI22_X1 U5517 ( .A1(n6828), .A2(UWORD_REG_13__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4948) );
  OAI21_X1 U5518 ( .B1(n4950), .B2(n4949), .A(n4948), .ZN(U2894) );
  NOR2_X1 U5519 ( .A1(n4823), .A2(n4951), .ZN(n4952) );
  OAI21_X1 U5520 ( .B1(n4953), .B2(n4952), .A(n7397), .ZN(n4954) );
  INV_X1 U5521 ( .A(n4955), .ZN(n4956) );
  INV_X1 U5522 ( .A(DATAI_1_), .ZN(n5077) );
  INV_X1 U5523 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6803) );
  OAI222_X1 U5524 ( .A1(n4957), .A2(n7581), .B1(n6481), .B2(n5077), .C1(n6479), 
        .C2(n6803), .ZN(U2890) );
  OR2_X1 U5525 ( .A1(n4890), .A2(n4959), .ZN(n4960) );
  AND2_X1 U5526 ( .A1(n4958), .A2(n4960), .ZN(n7191) );
  INV_X1 U5527 ( .A(n7191), .ZN(n4961) );
  INV_X1 U5528 ( .A(DATAI_5_), .ZN(n5059) );
  INV_X1 U5529 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6811) );
  OAI222_X1 U5530 ( .A1(n4961), .A2(n7581), .B1(n6481), .B2(n5059), .C1(n6479), 
        .C2(n6811), .ZN(U2886) );
  INV_X1 U5531 ( .A(DATAI_3_), .ZN(n5056) );
  INV_X1 U5532 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6807) );
  OAI222_X1 U5533 ( .A1(n4962), .A2(n7581), .B1(n6481), .B2(n5056), .C1(n6479), 
        .C2(n6807), .ZN(U2888) );
  XOR2_X1 U5534 ( .A(n4964), .B(n4963), .Z(n7024) );
  NAND2_X1 U5535 ( .A1(n7024), .A2(n6971), .ZN(n4968) );
  INV_X1 U5536 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U5537 ( .A1(n7073), .A2(REIP_REG_4__SCAN_IN), .ZN(n7020) );
  OAI21_X1 U5538 ( .B1(n6965), .B2(n4965), .A(n7020), .ZN(n4966) );
  AOI21_X1 U5539 ( .B1(n6941), .B2(n7170), .A(n4966), .ZN(n4967) );
  OAI211_X1 U5540 ( .C1(n7173), .C2(n6962), .A(n4968), .B(n4967), .ZN(U2982)
         );
  INV_X1 U5541 ( .A(DATAI_0_), .ZN(n7425) );
  INV_X1 U5542 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6801) );
  OAI222_X1 U5543 ( .A1(n6481), .A2(n7425), .B1(n6479), .B2(n6801), .C1(n7581), 
        .C2(n7149), .ZN(U2891) );
  INV_X1 U5544 ( .A(DATAI_2_), .ZN(n7434) );
  INV_X1 U5545 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6805) );
  INV_X1 U5546 ( .A(n4969), .ZN(n4970) );
  NAND2_X1 U5547 ( .A1(n4971), .A2(n4970), .ZN(n4972) );
  NAND2_X1 U5548 ( .A1(n4917), .A2(n4972), .ZN(n7156) );
  OAI222_X1 U5549 ( .A1(n6481), .A2(n7434), .B1(n6479), .B2(n6805), .C1(n7581), 
        .C2(n7156), .ZN(U2889) );
  INV_X1 U5550 ( .A(DATAI_4_), .ZN(n4973) );
  INV_X1 U5551 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6809) );
  OAI222_X1 U5552 ( .A1(n6481), .A2(n4973), .B1(n6479), .B2(n6809), .C1(n7581), 
        .C2(n7173), .ZN(U2887) );
  MUX2_X1 U5553 ( .A(n7373), .B(n5004), .S(n5266), .Z(n4974) );
  NAND2_X1 U5554 ( .A1(n4974), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U5555 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7373), .ZN(n4983) );
  INV_X1 U5556 ( .A(n4975), .ZN(n4982) );
  INV_X1 U5557 ( .A(n4976), .ZN(n4977) );
  NOR2_X1 U5558 ( .A1(n4978), .A2(n4977), .ZN(n4979) );
  XNOR2_X1 U5559 ( .A(n4979), .B(n4097), .ZN(n7347) );
  NOR2_X1 U5560 ( .A1(n4821), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U5561 ( .A1(n7347), .A2(n4980), .ZN(n4981) );
  OAI21_X1 U5562 ( .B1(n4983), .B2(n4982), .A(n4981), .ZN(n4984) );
  INV_X1 U5563 ( .A(n4984), .ZN(n4985) );
  AND2_X1 U5564 ( .A1(n5021), .A2(n4985), .ZN(n5019) );
  NAND2_X1 U5565 ( .A1(n7460), .A2(n5015), .ZN(n5003) );
  INV_X1 U5566 ( .A(n4986), .ZN(n4987) );
  NAND2_X1 U5567 ( .A1(n4988), .A2(n4987), .ZN(n5005) );
  MUX2_X1 U5568 ( .A(n4990), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4989), 
        .Z(n4991) );
  NOR2_X1 U5569 ( .A1(n4991), .A2(n4975), .ZN(n5001) );
  INV_X1 U5570 ( .A(n4992), .ZN(n4993) );
  OAI21_X1 U5571 ( .B1(n4989), .B2(n4994), .A(n4993), .ZN(n4995) );
  NOR2_X1 U5572 ( .A1(n4995), .A2(n3667), .ZN(n6722) );
  AND2_X1 U5573 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4997) );
  INV_X1 U5574 ( .A(n4997), .ZN(n4996) );
  MUX2_X1 U5575 ( .A(n4997), .B(n4996), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4998) );
  NAND2_X1 U5576 ( .A1(n5007), .A2(n4998), .ZN(n4999) );
  OAI21_X1 U5577 ( .B1(n6722), .B2(n5012), .A(n4999), .ZN(n5000) );
  AOI21_X1 U5578 ( .B1(n5005), .B2(n5001), .A(n5000), .ZN(n5002) );
  NAND2_X1 U5579 ( .A1(n5003), .A2(n5002), .ZN(n6720) );
  INV_X1 U5580 ( .A(n5004), .ZN(n7356) );
  MUX2_X1 U5581 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6720), .S(n7356), 
        .Z(n7365) );
  NAND2_X1 U5582 ( .A1(n5004), .A2(n6248), .ZN(n5017) );
  XNOR2_X1 U5583 ( .A(n4989), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5013)
         );
  NAND2_X1 U5584 ( .A1(n5005), .A2(n5013), .ZN(n5011) );
  NAND2_X1 U5585 ( .A1(n5007), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5009) );
  MUX2_X1 U5586 ( .A(n5009), .B(n5008), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n5010) );
  OAI211_X1 U5587 ( .C1(n5013), .C2(n5012), .A(n5011), .B(n5010), .ZN(n5014)
         );
  AOI21_X1 U5588 ( .B1(n5303), .B2(n5015), .A(n5014), .ZN(n6240) );
  NAND2_X1 U5589 ( .A1(n7356), .A2(n6240), .ZN(n5016) );
  AND2_X1 U5590 ( .A1(n5017), .A2(n5016), .ZN(n7360) );
  NAND3_X1 U5591 ( .A1(n7365), .A2(n7360), .A3(n5266), .ZN(n5018) );
  NAND2_X1 U5592 ( .A1(n5019), .A2(n5018), .ZN(n7369) );
  NAND2_X1 U5593 ( .A1(n5020), .A2(n5021), .ZN(n5022) );
  NAND2_X1 U5594 ( .A1(n7369), .A2(n5022), .ZN(n5254) );
  NAND2_X1 U5595 ( .A1(n5254), .A2(n7373), .ZN(n5023) );
  NAND2_X1 U5596 ( .A1(n5023), .A2(n6993), .ZN(n5024) );
  NAND2_X1 U5597 ( .A1(n7505), .A2(n5266), .ZN(n7393) );
  INV_X1 U5598 ( .A(n5388), .ZN(n5450) );
  AOI21_X1 U5599 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n7390), .A(n6796), .ZN(
        n5025) );
  INV_X1 U5600 ( .A(n5025), .ZN(n5255) );
  INV_X1 U5601 ( .A(n4814), .ZN(n5275) );
  NAND2_X1 U5602 ( .A1(n5045), .A2(n7499), .ZN(n5258) );
  XNOR2_X1 U5603 ( .A(n3679), .B(STATEBS16_REG_SCAN_IN), .ZN(n5026) );
  OAI222_X1 U5604 ( .A1(n5255), .A2(n5275), .B1(n5258), .B2(n5026), .C1(n7496), 
        .C2(n5045), .ZN(U3464) );
  INV_X1 U5605 ( .A(n5103), .ZN(n5027) );
  AOI21_X1 U5606 ( .B1(n5028), .B2(n4958), .A(n5027), .ZN(n6949) );
  INV_X1 U5607 ( .A(n6949), .ZN(n7200) );
  NAND2_X1 U5608 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5029)
         );
  OAI211_X1 U5609 ( .C1(n4786), .C2(EBX_REG_5__SCAN_IN), .A(n5579), .B(n5029), 
        .ZN(n5030) );
  OAI21_X1 U5610 ( .B1(n5745), .B2(EBX_REG_5__SCAN_IN), .A(n5030), .ZN(n6921)
         );
  INV_X1 U5611 ( .A(n5763), .ZN(n5651) );
  INV_X1 U5612 ( .A(EBX_REG_6__SCAN_IN), .ZN(n7197) );
  NAND2_X1 U5613 ( .A1(n5651), .A2(n7197), .ZN(n5035) );
  NAND2_X1 U5614 ( .A1(n5579), .A2(n7047), .ZN(n5033) );
  NAND2_X1 U5615 ( .A1(n6263), .A2(n7197), .ZN(n5032) );
  NAND3_X1 U5616 ( .A1(n5033), .A2(n5672), .A3(n5032), .ZN(n5034) );
  NAND2_X1 U5617 ( .A1(n6923), .A2(n5036), .ZN(n5037) );
  NAND2_X1 U5618 ( .A1(n5107), .A2(n5037), .ZN(n7196) );
  INV_X1 U5619 ( .A(n7196), .ZN(n5038) );
  AOI22_X1 U5620 ( .A1(n6924), .A2(n5038), .B1(EBX_REG_6__SCAN_IN), .B2(n6426), 
        .ZN(n5039) );
  OAI21_X1 U5621 ( .B1(n7200), .B2(n6454), .A(n5039), .ZN(U2853) );
  INV_X1 U5622 ( .A(n5303), .ZN(n7159) );
  INV_X1 U5623 ( .A(n3665), .ZN(n5041) );
  NAND2_X1 U5624 ( .A1(n3679), .A2(STATEBS16_REG_SCAN_IN), .ZN(n7482) );
  XNOR2_X1 U5625 ( .A(n5041), .B(n7482), .ZN(n5040) );
  OAI222_X1 U5626 ( .A1(n5045), .A2(n7363), .B1(n5255), .B2(n7159), .C1(n5258), 
        .C2(n5040), .ZN(U3463) );
  INV_X1 U5627 ( .A(n7460), .ZN(n5528) );
  NAND2_X1 U5628 ( .A1(n5526), .A2(n5041), .ZN(n7446) );
  OAI21_X1 U5629 ( .B1(n5112), .B2(STATEBS16_REG_SCAN_IN), .A(n7446), .ZN(
        n5043) );
  INV_X1 U5630 ( .A(n3679), .ZN(n5111) );
  NAND2_X1 U5631 ( .A1(n3665), .A2(n5111), .ZN(n5146) );
  NOR2_X1 U5632 ( .A1(n5503), .A2(n7497), .ZN(n5497) );
  NAND2_X1 U5633 ( .A1(n3665), .A2(n5042), .ZN(n5302) );
  NOR2_X1 U5634 ( .A1(n5302), .A2(n7482), .ZN(n7459) );
  NOR3_X1 U5635 ( .A1(n5043), .A2(n5497), .A3(n7459), .ZN(n5044) );
  OAI222_X1 U5636 ( .A1(n5045), .A2(n7364), .B1(n5255), .B2(n5528), .C1(n5258), 
        .C2(n5044), .ZN(U3462) );
  OAI222_X1 U5637 ( .A1(n7200), .A2(n7581), .B1(n6481), .B2(n7441), .C1(n6479), 
        .C2(n4138), .ZN(U2885) );
  NAND2_X1 U5638 ( .A1(n5065), .A2(DATAI_0_), .ZN(n5062) );
  INV_X2 U5639 ( .A(n5046), .ZN(n5092) );
  NOR2_X1 U5640 ( .A1(n5047), .A2(n5092), .ZN(n5057) );
  AOI22_X1 U5641 ( .A1(n5092), .A2(EAX_REG_16__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U5642 ( .A1(n5062), .A2(n5048), .ZN(U2924) );
  INV_X1 U5643 ( .A(DATAI_14_), .ZN(n6480) );
  OR2_X1 U5644 ( .A1(n5078), .A2(n6480), .ZN(n5098) );
  AOI22_X1 U5645 ( .A1(n5092), .A2(EAX_REG_14__SCAN_IN), .B1(n5057), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U5646 ( .A1(n5098), .A2(n5049), .ZN(U2953) );
  NAND2_X1 U5647 ( .A1(n5065), .A2(DATAI_10_), .ZN(n5087) );
  AOI22_X1 U5648 ( .A1(n5092), .A2(EAX_REG_10__SCAN_IN), .B1(n5057), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U5649 ( .A1(n5087), .A2(n5050), .ZN(U2949) );
  NAND2_X1 U5650 ( .A1(n5065), .A2(DATAI_12_), .ZN(n5074) );
  AOI22_X1 U5651 ( .A1(n5092), .A2(EAX_REG_12__SCAN_IN), .B1(n5057), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U5652 ( .A1(n5074), .A2(n5051), .ZN(U2951) );
  NAND2_X1 U5653 ( .A1(n5065), .A2(DATAI_13_), .ZN(n5101) );
  AOI22_X1 U5654 ( .A1(n5092), .A2(EAX_REG_13__SCAN_IN), .B1(n5057), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U5655 ( .A1(n5101), .A2(n5052), .ZN(U2952) );
  NAND2_X1 U5656 ( .A1(n5065), .A2(DATAI_11_), .ZN(n5096) );
  AOI22_X1 U5657 ( .A1(n5092), .A2(EAX_REG_11__SCAN_IN), .B1(n5057), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U5658 ( .A1(n5096), .A2(n5053), .ZN(U2950) );
  NAND2_X1 U5659 ( .A1(n5065), .A2(DATAI_9_), .ZN(n5091) );
  AOI22_X1 U5660 ( .A1(n5092), .A2(EAX_REG_9__SCAN_IN), .B1(n5057), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U5661 ( .A1(n5091), .A2(n5054), .ZN(U2948) );
  INV_X1 U5662 ( .A(DATAI_15_), .ZN(n6478) );
  AOI22_X1 U5663 ( .A1(n5092), .A2(EAX_REG_15__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n5055) );
  OAI21_X1 U5664 ( .B1(n5078), .B2(n6478), .A(n5055), .ZN(U2954) );
  OR2_X1 U5665 ( .A1(n5078), .A2(n5056), .ZN(n5076) );
  AOI22_X1 U5666 ( .A1(n5092), .A2(EAX_REG_3__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U5667 ( .A1(n5076), .A2(n5058), .ZN(U2942) );
  OR2_X1 U5668 ( .A1(n5078), .A2(n5059), .ZN(n5069) );
  AOI22_X1 U5669 ( .A1(n5092), .A2(EAX_REG_21__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U5670 ( .A1(n5069), .A2(n5060), .ZN(U2929) );
  AOI22_X1 U5671 ( .A1(n5092), .A2(EAX_REG_0__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U5672 ( .A1(n5062), .A2(n5061), .ZN(U2939) );
  NAND2_X1 U5673 ( .A1(n5065), .A2(DATAI_2_), .ZN(n5085) );
  AOI22_X1 U5674 ( .A1(n5092), .A2(EAX_REG_18__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U5675 ( .A1(n5085), .A2(n5063), .ZN(U2926) );
  NAND2_X1 U5676 ( .A1(n5065), .A2(DATAI_4_), .ZN(n5089) );
  AOI22_X1 U5677 ( .A1(n5092), .A2(EAX_REG_20__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U5678 ( .A1(n5089), .A2(n5064), .ZN(U2928) );
  NAND2_X1 U5679 ( .A1(n5065), .A2(DATAI_8_), .ZN(n5094) );
  AOI22_X1 U5680 ( .A1(n5092), .A2(EAX_REG_8__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U5681 ( .A1(n5094), .A2(n5066), .ZN(U2947) );
  OR2_X1 U5682 ( .A1(n5078), .A2(n7441), .ZN(n5071) );
  AOI22_X1 U5683 ( .A1(n5092), .A2(EAX_REG_22__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U5684 ( .A1(n5071), .A2(n5067), .ZN(U2930) );
  AOI22_X1 U5685 ( .A1(n5092), .A2(EAX_REG_5__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U5686 ( .A1(n5069), .A2(n5068), .ZN(U2944) );
  AOI22_X1 U5687 ( .A1(n5092), .A2(EAX_REG_6__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U5688 ( .A1(n5071), .A2(n5070), .ZN(U2945) );
  INV_X1 U5689 ( .A(DATAI_7_), .ZN(n5143) );
  OR2_X1 U5690 ( .A1(n5078), .A2(n5143), .ZN(n5081) );
  AOI22_X1 U5691 ( .A1(n5092), .A2(EAX_REG_7__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U5692 ( .A1(n5081), .A2(n5072), .ZN(U2946) );
  AOI22_X1 U5693 ( .A1(n5092), .A2(EAX_REG_28__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5073) );
  NAND2_X1 U5694 ( .A1(n5074), .A2(n5073), .ZN(U2936) );
  AOI22_X1 U5695 ( .A1(n5092), .A2(EAX_REG_19__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U5696 ( .A1(n5076), .A2(n5075), .ZN(U2927) );
  OR2_X1 U5697 ( .A1(n5078), .A2(n5077), .ZN(n5083) );
  AOI22_X1 U5698 ( .A1(n5092), .A2(EAX_REG_17__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U5699 ( .A1(n5083), .A2(n5079), .ZN(U2925) );
  AOI22_X1 U5700 ( .A1(n5092), .A2(EAX_REG_23__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5701 ( .A1(n5081), .A2(n5080), .ZN(U2931) );
  AOI22_X1 U5702 ( .A1(n5092), .A2(EAX_REG_1__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U5703 ( .A1(n5083), .A2(n5082), .ZN(U2940) );
  AOI22_X1 U5704 ( .A1(n5092), .A2(EAX_REG_2__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U5705 ( .A1(n5085), .A2(n5084), .ZN(U2941) );
  AOI22_X1 U5706 ( .A1(n5092), .A2(EAX_REG_26__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U5707 ( .A1(n5087), .A2(n5086), .ZN(U2934) );
  AOI22_X1 U5708 ( .A1(n5092), .A2(EAX_REG_4__SCAN_IN), .B1(n5099), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U5709 ( .A1(n5089), .A2(n5088), .ZN(U2943) );
  AOI22_X1 U5710 ( .A1(n5092), .A2(EAX_REG_25__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U5711 ( .A1(n5091), .A2(n5090), .ZN(U2933) );
  AOI22_X1 U5712 ( .A1(n5092), .A2(EAX_REG_24__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U5713 ( .A1(n5094), .A2(n5093), .ZN(U2932) );
  AOI22_X1 U5714 ( .A1(n5092), .A2(EAX_REG_27__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U5715 ( .A1(n5096), .A2(n5095), .ZN(U2935) );
  AOI22_X1 U5716 ( .A1(n5092), .A2(EAX_REG_30__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U5717 ( .A1(n5098), .A2(n5097), .ZN(U2938) );
  AOI22_X1 U5718 ( .A1(n5092), .A2(EAX_REG_29__SCAN_IN), .B1(n5099), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U5719 ( .A1(n5101), .A2(n5100), .ZN(U2937) );
  AND2_X1 U5720 ( .A1(n5103), .A2(n5102), .ZN(n5105) );
  OR2_X1 U5721 ( .A1(n5105), .A2(n3632), .ZN(n6956) );
  MUX2_X1 U5722 ( .A(n5745), .B(n5672), .S(EBX_REG_7__SCAN_IN), .Z(n5106) );
  OAI21_X1 U5723 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5772), .A(n5106), 
        .ZN(n5108) );
  AOI21_X1 U5724 ( .B1(n5108), .B2(n5107), .A(n5342), .ZN(n7206) );
  AOI22_X1 U5725 ( .A1(n6924), .A2(n7206), .B1(EBX_REG_7__SCAN_IN), .B2(n6426), 
        .ZN(n5109) );
  OAI21_X1 U5726 ( .B1(n6956), .B2(n6454), .A(n5109), .ZN(U2852) );
  NOR2_X1 U5727 ( .A1(n5387), .A2(n3947), .ZN(n7507) );
  NAND2_X1 U5728 ( .A1(n7364), .A2(n7363), .ZN(n7501) );
  INV_X1 U5729 ( .A(n7501), .ZN(n7495) );
  NAND2_X1 U5730 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7495), .ZN(n7489) );
  NOR2_X1 U5731 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7489), .ZN(n5115)
         );
  INV_X1 U5732 ( .A(n5115), .ZN(n5423) );
  NOR2_X1 U5733 ( .A1(n5526), .A2(n3665), .ZN(n7484) );
  NAND2_X1 U5734 ( .A1(n7484), .A2(n5111), .ZN(n7498) );
  OR2_X1 U5735 ( .A1(n7498), .A2(n3662), .ZN(n5418) );
  NAND2_X1 U5736 ( .A1(n3679), .A2(n3662), .ZN(n5301) );
  NOR2_X1 U5737 ( .A1(n3665), .A2(n5301), .ZN(n5525) );
  AND2_X1 U5738 ( .A1(n5112), .A2(n5525), .ZN(n7659) );
  NAND2_X1 U5739 ( .A1(n7499), .A2(n7497), .ZN(n5451) );
  OAI21_X1 U5740 ( .B1(n7667), .B2(n7659), .A(n5451), .ZN(n5114) );
  OR2_X1 U5741 ( .A1(n5303), .A2(n5275), .ZN(n7450) );
  INV_X1 U5742 ( .A(n7450), .ZN(n7486) );
  NAND2_X1 U5743 ( .A1(n5528), .A2(n7486), .ZN(n5113) );
  AOI21_X1 U5744 ( .B1(n5114), .B2(n5113), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5116) );
  NAND2_X1 U5745 ( .A1(n5529), .A2(n7364), .ZN(n5309) );
  NAND2_X1 U5746 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5309), .ZN(n5306) );
  NAND2_X1 U5747 ( .A1(n5117), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U5748 ( .A1(n5388), .A2(n6737), .ZN(n5533) );
  NAND2_X1 U5749 ( .A1(n5416), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U5750 ( .A1(DATAI_0_), .A2(n5388), .ZN(n7519) );
  NAND2_X1 U5751 ( .A1(n5528), .A2(n7499), .ZN(n5311) );
  INV_X1 U5752 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U5753 ( .A1(n5118), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5180) );
  OAI22_X1 U5754 ( .A1(n5311), .A2(n7450), .B1(n5309), .B2(n5180), .ZN(n5420)
         );
  AND2_X1 U5755 ( .A1(n6970), .A2(DATAI_24_), .ZN(n7516) );
  INV_X1 U5756 ( .A(n7516), .ZN(n5562) );
  AND2_X1 U5757 ( .A1(n6970), .A2(DATAI_16_), .ZN(n7508) );
  INV_X1 U5758 ( .A(n7508), .ZN(n5483) );
  OAI22_X1 U5759 ( .A1(n5418), .A2(n5562), .B1(n5417), .B2(n5483), .ZN(n5119)
         );
  AOI21_X1 U5760 ( .B1(n6740), .B2(n5420), .A(n5119), .ZN(n5120) );
  OAI211_X1 U5761 ( .C1(n5642), .C2(n5423), .A(n5121), .B(n5120), .ZN(U3036)
         );
  NOR2_X1 U5762 ( .A1(n5387), .A2(n3900), .ZN(n7554) );
  NAND2_X1 U5763 ( .A1(n5416), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U5764 ( .A1(DATAI_2_), .A2(n5388), .ZN(n7553) );
  AND2_X1 U5765 ( .A1(n6970), .A2(DATAI_26_), .ZN(n7556) );
  INV_X1 U5766 ( .A(n7556), .ZN(n5538) );
  AND2_X1 U5767 ( .A1(n6970), .A2(DATAI_18_), .ZN(n7557) );
  INV_X1 U5768 ( .A(n7557), .ZN(n5479) );
  OAI22_X1 U5769 ( .A1(n5418), .A2(n5538), .B1(n5417), .B2(n5479), .ZN(n5122)
         );
  AOI21_X1 U5770 ( .B1(n7555), .B2(n5420), .A(n5122), .ZN(n5123) );
  OAI211_X1 U5771 ( .C1(n5423), .C2(n5634), .A(n5124), .B(n5123), .ZN(U3038)
         );
  NAND2_X1 U5772 ( .A1(n5416), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U5773 ( .A1(DATAI_3_), .A2(n5388), .ZN(n7571) );
  AND2_X1 U5774 ( .A1(n6970), .A2(DATAI_27_), .ZN(n7574) );
  INV_X1 U5775 ( .A(n7574), .ZN(n5550) );
  AND2_X1 U5776 ( .A1(n6970), .A2(DATAI_19_), .ZN(n7575) );
  INV_X1 U5777 ( .A(n7575), .ZN(n5463) );
  OAI22_X1 U5778 ( .A1(n5418), .A2(n5550), .B1(n5417), .B2(n5463), .ZN(n5126)
         );
  AOI21_X1 U5779 ( .B1(n7573), .B2(n5420), .A(n5126), .ZN(n5127) );
  OAI211_X1 U5780 ( .C1(n5423), .C2(n5631), .A(n5128), .B(n5127), .ZN(U3039)
         );
  NAND2_X1 U5781 ( .A1(n5416), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U5782 ( .A1(DATAI_4_), .A2(n5388), .ZN(n7598) );
  AND2_X1 U5783 ( .A1(n6970), .A2(DATAI_28_), .ZN(n7601) );
  INV_X1 U5784 ( .A(n7601), .ZN(n5542) );
  AND2_X1 U5785 ( .A1(n6970), .A2(DATAI_20_), .ZN(n7602) );
  INV_X1 U5786 ( .A(n7602), .ZN(n5459) );
  OAI22_X1 U5787 ( .A1(n5418), .A2(n5542), .B1(n5417), .B2(n5459), .ZN(n5130)
         );
  AOI21_X1 U5788 ( .B1(n7600), .B2(n5420), .A(n5130), .ZN(n5131) );
  OAI211_X1 U5789 ( .C1(n5423), .C2(n5628), .A(n5132), .B(n5131), .ZN(U3040)
         );
  NOR2_X1 U5790 ( .A1(n5387), .A2(n3865), .ZN(n7632) );
  NAND2_X1 U5791 ( .A1(n5416), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U5792 ( .A1(DATAI_6_), .A2(n5388), .ZN(n7637) );
  AND2_X1 U5793 ( .A1(n6970), .A2(DATAI_30_), .ZN(n7634) );
  INV_X1 U5794 ( .A(n7634), .ZN(n5558) );
  AND2_X1 U5795 ( .A1(n6970), .A2(DATAI_22_), .ZN(n7633) );
  INV_X1 U5796 ( .A(n7633), .ZN(n5475) );
  OAI22_X1 U5797 ( .A1(n5418), .A2(n5558), .B1(n5417), .B2(n5475), .ZN(n5133)
         );
  AOI21_X1 U5798 ( .B1(n6765), .B2(n5420), .A(n5133), .ZN(n5134) );
  OAI211_X1 U5799 ( .C1(n5423), .C2(n5622), .A(n5135), .B(n5134), .ZN(U3042)
         );
  NAND2_X1 U5800 ( .A1(n5416), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U5801 ( .A1(DATAI_7_), .A2(n5388), .ZN(n7671) );
  AND2_X1 U5802 ( .A1(n6970), .A2(DATAI_31_), .ZN(n7678) );
  INV_X1 U5803 ( .A(n7678), .ZN(n5546) );
  AND2_X1 U5804 ( .A1(n6970), .A2(DATAI_23_), .ZN(n7679) );
  INV_X1 U5805 ( .A(n7679), .ZN(n5467) );
  OAI22_X1 U5806 ( .A1(n5418), .A2(n5546), .B1(n5417), .B2(n5467), .ZN(n5136)
         );
  AOI21_X1 U5807 ( .B1(n7676), .B2(n5420), .A(n5136), .ZN(n5137) );
  OAI211_X1 U5808 ( .C1(n5423), .C2(n5616), .A(n5138), .B(n5137), .ZN(U3043)
         );
  NAND2_X1 U5809 ( .A1(n5416), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U5810 ( .A1(DATAI_1_), .A2(n5388), .ZN(n7535) );
  AND2_X1 U5811 ( .A1(n6970), .A2(DATAI_25_), .ZN(n7538) );
  INV_X1 U5812 ( .A(n7538), .ZN(n5554) );
  AND2_X1 U5813 ( .A1(n6970), .A2(DATAI_17_), .ZN(n7539) );
  INV_X1 U5814 ( .A(n7539), .ZN(n5489) );
  OAI22_X1 U5815 ( .A1(n5418), .A2(n5554), .B1(n5417), .B2(n5489), .ZN(n5140)
         );
  AOI21_X1 U5816 ( .B1(n7537), .B2(n5420), .A(n5140), .ZN(n5141) );
  OAI211_X1 U5817 ( .C1(n5423), .C2(n5619), .A(n5142), .B(n5141), .ZN(U3037)
         );
  OAI222_X1 U5818 ( .A1(n6956), .A2(n7581), .B1(n6481), .B2(n5143), .C1(n6479), 
        .C2(n4155), .ZN(U2884) );
  NAND3_X1 U5819 ( .A1(n7364), .A2(n7496), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7476) );
  NOR2_X1 U5820 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7476), .ZN(n5151)
         );
  INV_X1 U5821 ( .A(n5151), .ZN(n5400) );
  AND2_X1 U5822 ( .A1(n7460), .A2(n7499), .ZN(n6735) );
  AND2_X1 U5823 ( .A1(n5303), .A2(n5275), .ZN(n7473) );
  NOR2_X1 U5824 ( .A1(n7473), .A2(n7511), .ZN(n5193) );
  INV_X1 U5825 ( .A(n7484), .ZN(n5144) );
  NAND2_X1 U5826 ( .A1(n3679), .A2(n5300), .ZN(n5223) );
  NOR2_X2 U5827 ( .A1(n5144), .A2(n5223), .ZN(n7661) );
  NOR2_X1 U5828 ( .A1(n5146), .A2(n5145), .ZN(n7471) );
  OAI21_X1 U5829 ( .B1(n7661), .B2(n7652), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5147) );
  OAI21_X1 U5830 ( .B1(n6735), .B2(n5193), .A(n5147), .ZN(n5150) );
  NAND2_X1 U5831 ( .A1(n5388), .A2(n5180), .ZN(n6727) );
  INV_X1 U5832 ( .A(n6727), .ZN(n5148) );
  OAI21_X1 U5833 ( .B1(n5529), .B2(n5195), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n5176) );
  AND2_X1 U5834 ( .A1(n5148), .A2(n5176), .ZN(n5149) );
  OAI211_X1 U5835 ( .C1(n5151), .C2(n7390), .A(n5150), .B(n5149), .ZN(n5398)
         );
  INV_X1 U5836 ( .A(n5311), .ZN(n6731) );
  NOR3_X1 U5837 ( .A1(n5195), .A2(n6737), .A3(n5529), .ZN(n5152) );
  AOI21_X1 U5838 ( .B1(n6731), .B2(n7473), .A(n5152), .ZN(n5396) );
  AOI22_X1 U5839 ( .A1(n7661), .A2(n7574), .B1(n7575), .B2(n7652), .ZN(n5153)
         );
  OAI21_X1 U5840 ( .B1(n7571), .B2(n5396), .A(n5153), .ZN(n5154) );
  AOI21_X1 U5841 ( .B1(INSTQUEUE_REG_4__3__SCAN_IN), .B2(n5398), .A(n5154), 
        .ZN(n5155) );
  OAI21_X1 U5842 ( .B1(n5631), .B2(n5400), .A(n5155), .ZN(U3055) );
  AOI22_X1 U5843 ( .A1(n7661), .A2(n7601), .B1(n7602), .B2(n7652), .ZN(n5156)
         );
  OAI21_X1 U5844 ( .B1(n7598), .B2(n5396), .A(n5156), .ZN(n5157) );
  AOI21_X1 U5845 ( .B1(INSTQUEUE_REG_4__4__SCAN_IN), .B2(n5398), .A(n5157), 
        .ZN(n5158) );
  OAI21_X1 U5846 ( .B1(n5628), .B2(n5400), .A(n5158), .ZN(U3056) );
  AOI22_X1 U5847 ( .A1(n7661), .A2(n7516), .B1(n7508), .B2(n7652), .ZN(n5159)
         );
  OAI21_X1 U5848 ( .B1(n7519), .B2(n5396), .A(n5159), .ZN(n5160) );
  AOI21_X1 U5849 ( .B1(INSTQUEUE_REG_4__0__SCAN_IN), .B2(n5398), .A(n5160), 
        .ZN(n5161) );
  OAI21_X1 U5850 ( .B1(n5642), .B2(n5400), .A(n5161), .ZN(U3052) );
  AOI22_X1 U5851 ( .A1(n7661), .A2(n7634), .B1(n7633), .B2(n7652), .ZN(n5162)
         );
  OAI21_X1 U5852 ( .B1(n7637), .B2(n5396), .A(n5162), .ZN(n5163) );
  AOI21_X1 U5853 ( .B1(INSTQUEUE_REG_4__6__SCAN_IN), .B2(n5398), .A(n5163), 
        .ZN(n5164) );
  OAI21_X1 U5854 ( .B1(n5622), .B2(n5400), .A(n5164), .ZN(U3058) );
  AOI22_X1 U5855 ( .A1(n7661), .A2(n7538), .B1(n7539), .B2(n7652), .ZN(n5165)
         );
  OAI21_X1 U5856 ( .B1(n7535), .B2(n5396), .A(n5165), .ZN(n5166) );
  AOI21_X1 U5857 ( .B1(INSTQUEUE_REG_4__1__SCAN_IN), .B2(n5398), .A(n5166), 
        .ZN(n5167) );
  OAI21_X1 U5858 ( .B1(n5619), .B2(n5400), .A(n5167), .ZN(U3053) );
  AOI22_X1 U5859 ( .A1(n7661), .A2(n7556), .B1(n7557), .B2(n7652), .ZN(n5168)
         );
  OAI21_X1 U5860 ( .B1(n7553), .B2(n5396), .A(n5168), .ZN(n5169) );
  AOI21_X1 U5861 ( .B1(INSTQUEUE_REG_4__2__SCAN_IN), .B2(n5398), .A(n5169), 
        .ZN(n5170) );
  OAI21_X1 U5862 ( .B1(n5634), .B2(n5400), .A(n5170), .ZN(U3054) );
  AOI22_X1 U5863 ( .A1(n7661), .A2(n7678), .B1(n7679), .B2(n7652), .ZN(n5171)
         );
  OAI21_X1 U5864 ( .B1(n7671), .B2(n5396), .A(n5171), .ZN(n5172) );
  AOI21_X1 U5865 ( .B1(INSTQUEUE_REG_4__7__SCAN_IN), .B2(n5398), .A(n5172), 
        .ZN(n5173) );
  OAI21_X1 U5866 ( .B1(n5616), .B2(n5400), .A(n5173), .ZN(U3059) );
  INV_X1 U5867 ( .A(n7498), .ZN(n5174) );
  AND2_X1 U5868 ( .A1(n3679), .A2(n5145), .ZN(n5175) );
  NAND2_X1 U5869 ( .A1(n5458), .A2(n5300), .ZN(n5488) );
  OAI21_X1 U5870 ( .B1(n7680), .B2(n7677), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5179) );
  OR2_X1 U5871 ( .A1(n5303), .A2(n4814), .ZN(n5182) );
  INV_X1 U5872 ( .A(n5182), .ZN(n7503) );
  NOR2_X1 U5873 ( .A1(n7503), .A2(n7511), .ZN(n5225) );
  OR2_X1 U5874 ( .A1(n5225), .A2(n6735), .ZN(n5178) );
  OAI211_X1 U5875 ( .C1(n7673), .C2(n7390), .A(n5227), .B(n5176), .ZN(n5177)
         );
  INV_X1 U5876 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5186) );
  INV_X1 U5877 ( .A(n5180), .ZN(n5530) );
  INV_X1 U5878 ( .A(n5529), .ZN(n5194) );
  NAND2_X1 U5879 ( .A1(n5530), .A2(n5194), .ZN(n5181) );
  OAI22_X1 U5880 ( .A1(n5311), .A2(n5182), .B1(n5195), .B2(n5181), .ZN(n7675)
         );
  INV_X1 U5881 ( .A(n7680), .ZN(n5187) );
  OAI22_X1 U5882 ( .A1(n5187), .A2(n5483), .B1(n5562), .B2(n5488), .ZN(n5183)
         );
  AOI21_X1 U5883 ( .B1(n6740), .B2(n7675), .A(n5183), .ZN(n5185) );
  NAND2_X1 U5884 ( .A1(n7507), .A2(n7673), .ZN(n5184) );
  OAI211_X1 U5885 ( .C1(n7684), .C2(n5186), .A(n5185), .B(n5184), .ZN(U3020)
         );
  INV_X1 U5886 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5191) );
  OAI22_X1 U5887 ( .A1(n5187), .A2(n5475), .B1(n5558), .B2(n5488), .ZN(n5188)
         );
  AOI21_X1 U5888 ( .B1(n6765), .B2(n7675), .A(n5188), .ZN(n5190) );
  NAND2_X1 U5889 ( .A1(n7632), .A2(n7673), .ZN(n5189) );
  OAI211_X1 U5890 ( .C1(n7684), .C2(n5191), .A(n5190), .B(n5189), .ZN(U3026)
         );
  NAND3_X1 U5891 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n7496), .ZN(n5500) );
  NOR2_X1 U5892 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5500), .ZN(n5199)
         );
  INV_X1 U5893 ( .A(n5199), .ZN(n5394) );
  NOR2_X2 U5894 ( .A1(n7446), .A2(n5223), .ZN(n7638) );
  NOR2_X2 U5895 ( .A1(n5503), .A2(n5300), .ZN(n5520) );
  OAI21_X1 U5896 ( .B1(n7638), .B2(n5520), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5192) );
  OAI21_X1 U5897 ( .B1(n6731), .B2(n5193), .A(n5192), .ZN(n5198) );
  NAND2_X1 U5898 ( .A1(n5195), .A2(n5194), .ZN(n5200) );
  NAND2_X1 U5899 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5200), .ZN(n5226) );
  INV_X1 U5900 ( .A(n5226), .ZN(n5196) );
  NOR2_X1 U5901 ( .A1(n5196), .A2(n6727), .ZN(n5197) );
  OAI211_X1 U5902 ( .C1(n7390), .C2(n5199), .A(n5198), .B(n5197), .ZN(n5392)
         );
  INV_X1 U5903 ( .A(n6737), .ZN(n5201) );
  INV_X1 U5904 ( .A(n5200), .ZN(n5231) );
  AOI22_X1 U5905 ( .A1(n6735), .A2(n7473), .B1(n5201), .B2(n5231), .ZN(n5390)
         );
  AOI22_X1 U5906 ( .A1(n7638), .A2(n7556), .B1(n5520), .B2(n7557), .ZN(n5202)
         );
  OAI21_X1 U5907 ( .B1(n7553), .B2(n5390), .A(n5202), .ZN(n5203) );
  AOI21_X1 U5908 ( .B1(INSTQUEUE_REG_12__2__SCAN_IN), .B2(n5392), .A(n5203), 
        .ZN(n5204) );
  OAI21_X1 U5909 ( .B1(n5634), .B2(n5394), .A(n5204), .ZN(U3118) );
  AOI22_X1 U5910 ( .A1(n7638), .A2(n7516), .B1(n5520), .B2(n7508), .ZN(n5205)
         );
  OAI21_X1 U5911 ( .B1(n7519), .B2(n5390), .A(n5205), .ZN(n5206) );
  AOI21_X1 U5912 ( .B1(INSTQUEUE_REG_12__0__SCAN_IN), .B2(n5392), .A(n5206), 
        .ZN(n5207) );
  OAI21_X1 U5913 ( .B1(n5642), .B2(n5394), .A(n5207), .ZN(U3116) );
  AOI22_X1 U5914 ( .A1(n7638), .A2(n7574), .B1(n5520), .B2(n7575), .ZN(n5208)
         );
  OAI21_X1 U5915 ( .B1(n7571), .B2(n5390), .A(n5208), .ZN(n5209) );
  AOI21_X1 U5916 ( .B1(INSTQUEUE_REG_12__3__SCAN_IN), .B2(n5392), .A(n5209), 
        .ZN(n5210) );
  OAI21_X1 U5917 ( .B1(n5631), .B2(n5394), .A(n5210), .ZN(U3119) );
  AOI22_X1 U5918 ( .A1(n7638), .A2(n7538), .B1(n5520), .B2(n7539), .ZN(n5211)
         );
  OAI21_X1 U5919 ( .B1(n7535), .B2(n5390), .A(n5211), .ZN(n5212) );
  AOI21_X1 U5920 ( .B1(INSTQUEUE_REG_12__1__SCAN_IN), .B2(n5392), .A(n5212), 
        .ZN(n5213) );
  OAI21_X1 U5921 ( .B1(n5619), .B2(n5394), .A(n5213), .ZN(U3117) );
  AOI22_X1 U5922 ( .A1(n7638), .A2(n7678), .B1(n5520), .B2(n7679), .ZN(n5214)
         );
  OAI21_X1 U5923 ( .B1(n7671), .B2(n5390), .A(n5214), .ZN(n5215) );
  AOI21_X1 U5924 ( .B1(INSTQUEUE_REG_12__7__SCAN_IN), .B2(n5392), .A(n5215), 
        .ZN(n5216) );
  OAI21_X1 U5925 ( .B1(n5616), .B2(n5394), .A(n5216), .ZN(U3123) );
  AOI22_X1 U5926 ( .A1(n7638), .A2(n7634), .B1(n5520), .B2(n7633), .ZN(n5217)
         );
  OAI21_X1 U5927 ( .B1(n7637), .B2(n5390), .A(n5217), .ZN(n5218) );
  AOI21_X1 U5928 ( .B1(INSTQUEUE_REG_12__6__SCAN_IN), .B2(n5392), .A(n5218), 
        .ZN(n5219) );
  OAI21_X1 U5929 ( .B1(n5622), .B2(n5394), .A(n5219), .ZN(U3122) );
  AOI22_X1 U5930 ( .A1(n7638), .A2(n7601), .B1(n5520), .B2(n7602), .ZN(n5220)
         );
  OAI21_X1 U5931 ( .B1(n7598), .B2(n5390), .A(n5220), .ZN(n5221) );
  AOI21_X1 U5932 ( .B1(INSTQUEUE_REG_12__4__SCAN_IN), .B2(n5392), .A(n5221), 
        .ZN(n5222) );
  OAI21_X1 U5933 ( .B1(n5628), .B2(n5394), .A(n5222), .ZN(U3120) );
  NOR3_X1 U5934 ( .A1(n7364), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5610) );
  INV_X1 U5935 ( .A(n5610), .ZN(n5611) );
  NOR2_X1 U5936 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5611), .ZN(n5230)
         );
  INV_X1 U5937 ( .A(n5230), .ZN(n5406) );
  NOR2_X2 U5938 ( .A1(n5605), .A2(n5300), .ZN(n5638) );
  NOR2_X2 U5939 ( .A1(n5302), .A2(n5223), .ZN(n7647) );
  OAI21_X1 U5940 ( .B1(n5638), .B2(n7647), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5224) );
  OAI21_X1 U5941 ( .B1(n6731), .B2(n5225), .A(n5224), .ZN(n5229) );
  AND2_X1 U5942 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  AOI22_X1 U5943 ( .A1(n6735), .A2(n7503), .B1(n5530), .B2(n5231), .ZN(n5402)
         );
  AOI22_X1 U5944 ( .A1(n5638), .A2(n7557), .B1(n7556), .B2(n7647), .ZN(n5232)
         );
  OAI21_X1 U5945 ( .B1(n7553), .B2(n5402), .A(n5232), .ZN(n5233) );
  AOI21_X1 U5946 ( .B1(INSTQUEUE_REG_8__2__SCAN_IN), .B2(n5404), .A(n5233), 
        .ZN(n5234) );
  OAI21_X1 U5947 ( .B1(n5634), .B2(n5406), .A(n5234), .ZN(U3086) );
  AOI22_X1 U5948 ( .A1(n5638), .A2(n7539), .B1(n7538), .B2(n7647), .ZN(n5235)
         );
  OAI21_X1 U5949 ( .B1(n7535), .B2(n5402), .A(n5235), .ZN(n5236) );
  AOI21_X1 U5950 ( .B1(INSTQUEUE_REG_8__1__SCAN_IN), .B2(n5404), .A(n5236), 
        .ZN(n5237) );
  OAI21_X1 U5951 ( .B1(n5619), .B2(n5406), .A(n5237), .ZN(U3085) );
  AOI22_X1 U5952 ( .A1(n5638), .A2(n7602), .B1(n7601), .B2(n7647), .ZN(n5238)
         );
  OAI21_X1 U5953 ( .B1(n7598), .B2(n5402), .A(n5238), .ZN(n5239) );
  AOI21_X1 U5954 ( .B1(INSTQUEUE_REG_8__4__SCAN_IN), .B2(n5404), .A(n5239), 
        .ZN(n5240) );
  OAI21_X1 U5955 ( .B1(n5628), .B2(n5406), .A(n5240), .ZN(U3088) );
  AOI22_X1 U5956 ( .A1(n5638), .A2(n7633), .B1(n7634), .B2(n7647), .ZN(n5241)
         );
  OAI21_X1 U5957 ( .B1(n7637), .B2(n5402), .A(n5241), .ZN(n5242) );
  AOI21_X1 U5958 ( .B1(INSTQUEUE_REG_8__6__SCAN_IN), .B2(n5404), .A(n5242), 
        .ZN(n5243) );
  OAI21_X1 U5959 ( .B1(n5622), .B2(n5406), .A(n5243), .ZN(U3090) );
  AOI22_X1 U5960 ( .A1(n5638), .A2(n7575), .B1(n7574), .B2(n7647), .ZN(n5244)
         );
  OAI21_X1 U5961 ( .B1(n7571), .B2(n5402), .A(n5244), .ZN(n5245) );
  AOI21_X1 U5962 ( .B1(INSTQUEUE_REG_8__3__SCAN_IN), .B2(n5404), .A(n5245), 
        .ZN(n5246) );
  OAI21_X1 U5963 ( .B1(n5631), .B2(n5406), .A(n5246), .ZN(U3087) );
  AOI22_X1 U5964 ( .A1(n5638), .A2(n7508), .B1(n7516), .B2(n7647), .ZN(n5247)
         );
  OAI21_X1 U5965 ( .B1(n7519), .B2(n5402), .A(n5247), .ZN(n5248) );
  AOI21_X1 U5966 ( .B1(INSTQUEUE_REG_8__0__SCAN_IN), .B2(n5404), .A(n5248), 
        .ZN(n5249) );
  OAI21_X1 U5967 ( .B1(n5642), .B2(n5406), .A(n5249), .ZN(U3084) );
  AOI22_X1 U5968 ( .A1(n5638), .A2(n7679), .B1(n7678), .B2(n7647), .ZN(n5250)
         );
  OAI21_X1 U5969 ( .B1(n7671), .B2(n5402), .A(n5250), .ZN(n5251) );
  AOI21_X1 U5970 ( .B1(INSTQUEUE_REG_8__7__SCAN_IN), .B2(n5404), .A(n5251), 
        .ZN(n5252) );
  OAI21_X1 U5971 ( .B1(n5616), .B2(n5406), .A(n5252), .ZN(U3091) );
  NAND2_X1 U5972 ( .A1(n5254), .A2(n5253), .ZN(n7399) );
  OAI22_X1 U5973 ( .A1(n6796), .A2(n7399), .B1(n4062), .B2(n5255), .ZN(n5256)
         );
  AOI21_X1 U5974 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6796), .A(n5256), 
        .ZN(n5257) );
  OAI21_X1 U5975 ( .B1(n3662), .B2(n5258), .A(n5257), .ZN(U3465) );
  INV_X1 U5976 ( .A(n4790), .ZN(n5288) );
  NOR3_X1 U5977 ( .A1(n7400), .A2(n7390), .A3(n7393), .ZN(n7395) );
  AND2_X1 U5978 ( .A1(n3628), .A2(n5261), .ZN(n7381) );
  OR3_X1 U5979 ( .A1(n7073), .A2(n7395), .A3(n7381), .ZN(n5263) );
  NAND2_X1 U5980 ( .A1(n7414), .A2(n7497), .ZN(n5279) );
  NAND2_X1 U5981 ( .A1(n5279), .A2(EBX_REG_31__SCAN_IN), .ZN(n5264) );
  NOR2_X1 U5982 ( .A1(n4786), .A2(n5264), .ZN(n5265) );
  NOR2_X1 U5983 ( .A1(n5277), .A2(n5266), .ZN(n5267) );
  NAND2_X1 U5984 ( .A1(n5776), .A2(n3921), .ZN(n5268) );
  INV_X1 U5985 ( .A(n7172), .ZN(n7190) );
  INV_X1 U5986 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U5987 ( .A1(n5776), .A2(n5270), .ZN(n7167) );
  INV_X1 U5988 ( .A(n5279), .ZN(n5271) );
  NAND2_X1 U5989 ( .A1(n3891), .A2(n5271), .ZN(n5272) );
  NOR2_X1 U5990 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  OAI22_X1 U5991 ( .A1(n5275), .A2(n7167), .B1(n7316), .B2(REIP_REG_1__SCAN_IN), .ZN(n5276) );
  AOI21_X1 U5992 ( .B1(n6928), .B2(n7190), .A(n5276), .ZN(n5287) );
  AND2_X1 U5993 ( .A1(n5277), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5278) );
  INV_X1 U5994 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5285) );
  NOR2_X1 U5995 ( .A1(n5279), .A2(n6989), .ZN(n5779) );
  INV_X1 U5996 ( .A(n5779), .ZN(n7379) );
  NAND2_X1 U5997 ( .A1(n6995), .A2(n7379), .ZN(n5281) );
  INV_X1 U5998 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5777) );
  NAND3_X1 U5999 ( .A1(n3664), .A2(n5777), .A3(n5279), .ZN(n5280) );
  NAND2_X1 U6000 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  AOI22_X1 U6001 ( .A1(EBX_REG_1__SCAN_IN), .A2(n7332), .B1(n7268), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5283) );
  OAI21_X1 U6002 ( .B1(n7294), .B2(n5285), .A(n5283), .ZN(n5284) );
  AOI21_X1 U6003 ( .B1(n7339), .B2(n5285), .A(n5284), .ZN(n5286) );
  OAI211_X1 U6004 ( .C1(n5288), .C2(n7329), .A(n5287), .B(n5286), .ZN(U2826)
         );
  NAND2_X1 U6005 ( .A1(n5289), .A2(n7190), .ZN(n5299) );
  INV_X1 U6006 ( .A(n5290), .ZN(n5295) );
  INV_X1 U6007 ( .A(REIP_REG_3__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U6008 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n7150) );
  NAND3_X1 U6009 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n7165) );
  NAND2_X1 U6010 ( .A1(n7316), .A2(n6366), .ZN(n7266) );
  OAI21_X1 U6011 ( .B1(n7268), .B2(n7165), .A(n7266), .ZN(n7178) );
  AOI221_X1 U6012 ( .B1(n7268), .B2(n7029), .C1(n7150), .C2(n7029), .A(n7178), 
        .ZN(n5291) );
  INV_X1 U6013 ( .A(n5291), .ZN(n5293) );
  AOI22_X1 U6014 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n7335), .B1(
        EBX_REG_3__SCAN_IN), .B2(n7332), .ZN(n5292) );
  NAND2_X1 U6015 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  AOI21_X1 U6016 ( .B1(n7339), .B2(n5295), .A(n5294), .ZN(n5296) );
  OAI21_X1 U6017 ( .B1(n7167), .B2(n5528), .A(n5296), .ZN(n5297) );
  INV_X1 U6018 ( .A(n5297), .ZN(n5298) );
  OAI211_X1 U6019 ( .C1(n7030), .C2(n7329), .A(n5299), .B(n5298), .ZN(U2824)
         );
  NOR3_X1 U6020 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n7363), .A3(n7496), 
        .ZN(n7464) );
  INV_X1 U6021 ( .A(n7464), .ZN(n7465) );
  NOR2_X1 U6022 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7465), .ZN(n5308)
         );
  INV_X1 U6023 ( .A(n5308), .ZN(n5415) );
  NAND2_X1 U6024 ( .A1(n7471), .A2(n5300), .ZN(n5410) );
  OAI21_X1 U6025 ( .B1(n7654), .B2(n7645), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5305) );
  NAND2_X1 U6026 ( .A1(n5303), .A2(n4814), .ZN(n5310) );
  INV_X1 U6027 ( .A(n5310), .ZN(n7462) );
  NOR2_X1 U6028 ( .A1(n7462), .A2(n7511), .ZN(n6730) );
  OR2_X1 U6029 ( .A1(n6730), .A2(n6735), .ZN(n5304) );
  AOI21_X1 U6030 ( .B1(n5305), .B2(n5304), .A(n6727), .ZN(n5307) );
  NAND2_X1 U6031 ( .A1(n5408), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5314) );
  OAI22_X1 U6032 ( .A1(n5311), .A2(n5310), .B1(n5309), .B2(n6737), .ZN(n5412)
         );
  OAI22_X1 U6033 ( .A1(n5410), .A2(n5546), .B1(n5467), .B2(n5409), .ZN(n5312)
         );
  AOI21_X1 U6034 ( .B1(n7676), .B2(n5412), .A(n5312), .ZN(n5313) );
  OAI211_X1 U6035 ( .C1(n5415), .C2(n5616), .A(n5314), .B(n5313), .ZN(U3075)
         );
  NAND2_X1 U6036 ( .A1(n5408), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5317) );
  OAI22_X1 U6037 ( .A1(n5410), .A2(n5562), .B1(n5483), .B2(n5409), .ZN(n5315)
         );
  AOI21_X1 U6038 ( .B1(n6740), .B2(n5412), .A(n5315), .ZN(n5316) );
  OAI211_X1 U6039 ( .C1(n5415), .C2(n5642), .A(n5317), .B(n5316), .ZN(U3068)
         );
  NAND2_X1 U6040 ( .A1(n5408), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5320) );
  OAI22_X1 U6041 ( .A1(n5410), .A2(n5542), .B1(n5459), .B2(n5409), .ZN(n5318)
         );
  AOI21_X1 U6042 ( .B1(n7600), .B2(n5412), .A(n5318), .ZN(n5319) );
  OAI211_X1 U6043 ( .C1(n5415), .C2(n5628), .A(n5320), .B(n5319), .ZN(U3072)
         );
  NAND2_X1 U6044 ( .A1(n5408), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5323) );
  OAI22_X1 U6045 ( .A1(n5410), .A2(n5554), .B1(n5489), .B2(n5409), .ZN(n5321)
         );
  AOI21_X1 U6046 ( .B1(n7537), .B2(n5412), .A(n5321), .ZN(n5322) );
  OAI211_X1 U6047 ( .C1(n5619), .C2(n5415), .A(n5323), .B(n5322), .ZN(U3069)
         );
  NAND2_X1 U6048 ( .A1(n5408), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5326) );
  OAI22_X1 U6049 ( .A1(n5410), .A2(n5558), .B1(n5475), .B2(n5409), .ZN(n5324)
         );
  AOI21_X1 U6050 ( .B1(n6765), .B2(n5412), .A(n5324), .ZN(n5325) );
  OAI211_X1 U6051 ( .C1(n5415), .C2(n5622), .A(n5326), .B(n5325), .ZN(U3074)
         );
  NAND2_X1 U6052 ( .A1(n5408), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5329) );
  OAI22_X1 U6053 ( .A1(n5410), .A2(n5538), .B1(n5479), .B2(n5409), .ZN(n5327)
         );
  AOI21_X1 U6054 ( .B1(n7555), .B2(n5412), .A(n5327), .ZN(n5328) );
  OAI211_X1 U6055 ( .C1(n5415), .C2(n5634), .A(n5329), .B(n5328), .ZN(U3070)
         );
  NAND2_X1 U6056 ( .A1(n5408), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5332) );
  OAI22_X1 U6057 ( .A1(n5410), .A2(n5550), .B1(n5463), .B2(n5409), .ZN(n5330)
         );
  AOI21_X1 U6058 ( .B1(n7573), .B2(n5412), .A(n5330), .ZN(n5331) );
  OAI211_X1 U6059 ( .C1(n5415), .C2(n5631), .A(n5332), .B(n5331), .ZN(U3071)
         );
  OAI21_X1 U6060 ( .B1(n5333), .B2(n5335), .A(n5334), .ZN(n5360) );
  OR2_X1 U6061 ( .A1(n5763), .A2(EBX_REG_8__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6062 ( .A1(n5579), .A2(n5348), .ZN(n5338) );
  INV_X1 U6063 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6064 ( .A1(n6263), .A2(n5336), .ZN(n5337) );
  NAND3_X1 U6065 ( .A1(n5338), .A2(n5672), .A3(n5337), .ZN(n5339) );
  NAND2_X1 U6066 ( .A1(n5340), .A2(n5339), .ZN(n5341) );
  NOR2_X1 U6067 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  OR2_X1 U6068 ( .A1(n5384), .A2(n5343), .ZN(n5370) );
  INV_X1 U6069 ( .A(n5370), .ZN(n5362) );
  AND2_X1 U6070 ( .A1(n7073), .A2(REIP_REG_8__SCAN_IN), .ZN(n5356) );
  NOR2_X1 U6071 ( .A1(n5348), .A2(n7077), .ZN(n7080) );
  NOR2_X1 U6072 ( .A1(n7021), .A2(n4676), .ZN(n7041) );
  OAI21_X1 U6073 ( .B1(n3653), .B2(n7062), .A(n4897), .ZN(n7027) );
  NAND2_X1 U6074 ( .A1(n7041), .A2(n7027), .ZN(n5345) );
  INV_X1 U6075 ( .A(n5345), .ZN(n7052) );
  NAND2_X1 U6076 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n7061) );
  NOR2_X1 U6077 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n7013), .ZN(n6708)
         );
  INV_X1 U6078 ( .A(n7068), .ZN(n7038) );
  AOI21_X1 U6079 ( .B1(n7061), .B2(n7063), .A(n5799), .ZN(n7028) );
  NAND3_X1 U6080 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n7052), .A3(n7028), 
        .ZN(n7048) );
  NOR2_X1 U6081 ( .A1(n7047), .A2(n7048), .ZN(n7079) );
  OAI21_X1 U6082 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n7079), .ZN(n5349) );
  INV_X1 U6083 ( .A(n7088), .ZN(n5347) );
  INV_X1 U6084 ( .A(n7061), .ZN(n7018) );
  NAND2_X1 U6085 ( .A1(n7018), .A2(n7041), .ZN(n7037) );
  NOR3_X1 U6086 ( .A1(n7047), .A2(n7051), .A3(n7037), .ZN(n5682) );
  NOR3_X1 U6087 ( .A1(n7047), .A2(n7051), .A3(n5345), .ZN(n5681) );
  OAI22_X1 U6088 ( .A1(n7019), .A2(n5682), .B1(n5681), .B2(n7063), .ZN(n5346)
         );
  NOR2_X1 U6089 ( .A1(n5347), .A2(n5346), .ZN(n7078) );
  OAI22_X1 U6090 ( .A1(n7080), .A2(n5349), .B1(n7078), .B2(n5348), .ZN(n5350)
         );
  AOI211_X1 U6091 ( .C1(n7132), .C2(n5362), .A(n5356), .B(n5350), .ZN(n5351)
         );
  OAI21_X1 U6092 ( .B1(n7055), .B2(n5360), .A(n5351), .ZN(U3010) );
  INV_X1 U6093 ( .A(n5352), .ZN(n5355) );
  INV_X1 U6094 ( .A(n3632), .ZN(n5354) );
  AOI21_X1 U6095 ( .B1(n5355), .B2(n5354), .A(n5353), .ZN(n5361) );
  AOI21_X1 U6096 ( .B1(n6969), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5356), 
        .ZN(n5357) );
  OAI21_X1 U6097 ( .B1(n5367), .B2(n6975), .A(n5357), .ZN(n5358) );
  AOI21_X1 U6098 ( .B1(n5361), .B2(n6970), .A(n5358), .ZN(n5359) );
  OAI21_X1 U6099 ( .B1(n5360), .B2(n7345), .A(n5359), .ZN(U2978) );
  INV_X1 U6100 ( .A(n5361), .ZN(n5375) );
  AOI22_X1 U6101 ( .A1(n6924), .A2(n5362), .B1(EBX_REG_8__SCAN_IN), .B2(n6426), 
        .ZN(n5363) );
  OAI21_X1 U6102 ( .B1(n5375), .B2(n6454), .A(n5363), .ZN(U2851) );
  NAND3_X1 U6104 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_8__SCAN_IN), .ZN(n5432) );
  INV_X1 U6105 ( .A(REIP_REG_4__SCAN_IN), .ZN(n7179) );
  NOR2_X1 U6106 ( .A1(n7165), .A2(n7179), .ZN(n7187) );
  NAND2_X1 U6107 ( .A1(n7187), .A2(REIP_REG_5__SCAN_IN), .ZN(n7184) );
  OR3_X1 U6108 ( .A1(n7268), .A2(n5432), .A3(n7184), .ZN(n6383) );
  NAND2_X1 U6109 ( .A1(n6383), .A2(n7266), .ZN(n5436) );
  INV_X1 U6110 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U6111 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n5364) );
  NAND3_X1 U6112 ( .A1(n7151), .A2(REIP_REG_5__SCAN_IN), .A3(n7187), .ZN(n7205) );
  OAI33_X1 U6113 ( .A1(1'b0), .A2(n5436), .A3(n6844), .B1(REIP_REG_8__SCAN_IN), 
        .B2(n5364), .B3(n7205), .ZN(n5366) );
  INV_X1 U6114 ( .A(n5366), .ZN(n5374) );
  INV_X1 U6115 ( .A(n5367), .ZN(n5372) );
  AOI22_X1 U6116 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n7335), .B1(
        EBX_REG_8__SCAN_IN), .B2(n7332), .ZN(n5369) );
  OAI211_X1 U6117 ( .C1(n7329), .C2(n5370), .A(n5369), .B(n7291), .ZN(n5371)
         );
  AOI21_X1 U6118 ( .B1(n7339), .B2(n5372), .A(n5371), .ZN(n5373) );
  OAI211_X1 U6119 ( .C1(n5375), .C2(n7325), .A(n5374), .B(n5373), .ZN(U2819)
         );
  INV_X1 U6120 ( .A(DATAI_8_), .ZN(n5888) );
  INV_X1 U6121 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6816) );
  OAI222_X1 U6122 ( .A1(n5375), .A2(n7581), .B1(n6481), .B2(n5888), .C1(n6479), 
        .C2(n6816), .ZN(U2883) );
  OR2_X1 U6123 ( .A1(n5353), .A2(n5377), .ZN(n5378) );
  NAND2_X1 U6124 ( .A1(n5376), .A2(n5378), .ZN(n5600) );
  INV_X1 U6125 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6126 ( .A1(n5759), .A2(n5379), .ZN(n5382) );
  NAND2_X1 U6127 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5380)
         );
  OAI211_X1 U6128 ( .C1(n4786), .C2(EBX_REG_9__SCAN_IN), .A(n5579), .B(n5380), 
        .ZN(n5381) );
  OR2_X1 U6129 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  AND2_X1 U6130 ( .A1(n5586), .A2(n5385), .ZN(n7096) );
  AOI22_X1 U6131 ( .A1(n6924), .A2(n7096), .B1(EBX_REG_9__SCAN_IN), .B2(n6426), 
        .ZN(n5386) );
  OAI21_X1 U6132 ( .B1(n5600), .B2(n6454), .A(n5386), .ZN(U2850) );
  NAND2_X1 U6133 ( .A1(DATAI_5_), .A2(n5388), .ZN(n7616) );
  AND2_X1 U6134 ( .A1(n6970), .A2(DATAI_29_), .ZN(n7619) );
  AND2_X1 U6135 ( .A1(n6970), .A2(DATAI_21_), .ZN(n7620) );
  AOI22_X1 U6136 ( .A1(n7638), .A2(n7619), .B1(n5520), .B2(n7620), .ZN(n5389)
         );
  OAI21_X1 U6137 ( .B1(n7616), .B2(n5390), .A(n5389), .ZN(n5391) );
  AOI21_X1 U6138 ( .B1(INSTQUEUE_REG_12__5__SCAN_IN), .B2(n5392), .A(n5391), 
        .ZN(n5393) );
  OAI21_X1 U6139 ( .B1(n5625), .B2(n5394), .A(n5393), .ZN(U3121) );
  AOI22_X1 U6140 ( .A1(n7661), .A2(n7619), .B1(n7620), .B2(n7652), .ZN(n5395)
         );
  OAI21_X1 U6141 ( .B1(n7616), .B2(n5396), .A(n5395), .ZN(n5397) );
  AOI21_X1 U6142 ( .B1(INSTQUEUE_REG_4__5__SCAN_IN), .B2(n5398), .A(n5397), 
        .ZN(n5399) );
  OAI21_X1 U6143 ( .B1(n5625), .B2(n5400), .A(n5399), .ZN(U3057) );
  AOI22_X1 U6144 ( .A1(n5638), .A2(n7620), .B1(n7619), .B2(n7647), .ZN(n5401)
         );
  OAI21_X1 U6145 ( .B1(n7616), .B2(n5402), .A(n5401), .ZN(n5403) );
  AOI21_X1 U6146 ( .B1(INSTQUEUE_REG_8__5__SCAN_IN), .B2(n5404), .A(n5403), 
        .ZN(n5405) );
  OAI21_X1 U6147 ( .B1(n5625), .B2(n5406), .A(n5405), .ZN(U3089) );
  INV_X1 U6148 ( .A(DATAI_9_), .ZN(n5407) );
  INV_X1 U6149 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6818) );
  OAI222_X1 U6150 ( .A1(n6481), .A2(n5407), .B1(n6479), .B2(n6818), .C1(n7581), 
        .C2(n5600), .ZN(U2882) );
  NAND2_X1 U6151 ( .A1(n5408), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5414) );
  INV_X1 U6152 ( .A(n7619), .ZN(n5567) );
  INV_X1 U6153 ( .A(n7620), .ZN(n5471) );
  OAI22_X1 U6154 ( .A1(n5410), .A2(n5567), .B1(n5471), .B2(n5409), .ZN(n5411)
         );
  AOI21_X1 U6155 ( .B1(n7618), .B2(n5412), .A(n5411), .ZN(n5413) );
  OAI211_X1 U6156 ( .C1(n5415), .C2(n5625), .A(n5414), .B(n5413), .ZN(U3073)
         );
  NAND2_X1 U6157 ( .A1(n5416), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5422) );
  OAI22_X1 U6158 ( .A1(n5418), .A2(n5567), .B1(n5417), .B2(n5471), .ZN(n5419)
         );
  AOI21_X1 U6159 ( .B1(n7618), .B2(n5420), .A(n5419), .ZN(n5421) );
  OAI211_X1 U6160 ( .C1(n5423), .C2(n5625), .A(n5422), .B(n5421), .ZN(U3041)
         );
  INV_X1 U6161 ( .A(n5376), .ZN(n5426) );
  OAI21_X1 U6162 ( .B1(n5426), .B2(n4200), .A(n5425), .ZN(n5648) );
  OR2_X1 U6163 ( .A1(n5763), .A2(EBX_REG_10__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6164 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6165 ( .A1(n5579), .A2(n5427), .ZN(n5428) );
  OAI21_X1 U6166 ( .B1(EBX_REG_10__SCAN_IN), .B2(n4786), .A(n5428), .ZN(n5429)
         );
  NAND2_X1 U6167 ( .A1(n5430), .A2(n5429), .ZN(n5584) );
  XNOR2_X1 U6168 ( .A(n5586), .B(n5584), .ZN(n7083) );
  AOI22_X1 U6169 ( .A1(n6924), .A2(n7083), .B1(EBX_REG_10__SCAN_IN), .B2(n6426), .ZN(n5431) );
  OAI21_X1 U6170 ( .B1(n5648), .B2(n6454), .A(n5431), .ZN(U2849) );
  INV_X1 U6171 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6846) );
  NOR2_X1 U6172 ( .A1(n5432), .A2(n7184), .ZN(n5781) );
  INV_X1 U6173 ( .A(n5781), .ZN(n5433) );
  INV_X1 U6174 ( .A(n7218), .ZN(n7230) );
  NOR3_X1 U6175 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6846), .A3(n7230), .ZN(n5440) );
  INV_X1 U6176 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5435) );
  AOI22_X1 U6177 ( .A1(EBX_REG_10__SCAN_IN), .A2(n7332), .B1(n7337), .B2(n7083), .ZN(n5434) );
  OAI211_X1 U6178 ( .C1(n7294), .C2(n5435), .A(n5434), .B(n7291), .ZN(n5439)
         );
  INV_X1 U6179 ( .A(n5436), .ZN(n5577) );
  NOR2_X1 U6180 ( .A1(REIP_REG_9__SCAN_IN), .A2(n7230), .ZN(n5444) );
  OAI21_X1 U6181 ( .B1(n5577), .B2(n5444), .A(REIP_REG_10__SCAN_IN), .ZN(n5437) );
  OAI21_X1 U6182 ( .B1(n7323), .B2(n5644), .A(n5437), .ZN(n5438) );
  NOR3_X1 U6183 ( .A1(n5440), .A2(n5439), .A3(n5438), .ZN(n5441) );
  OAI21_X1 U6184 ( .B1(n5648), .B2(n7325), .A(n5441), .ZN(U2817) );
  AOI22_X1 U6185 ( .A1(EBX_REG_9__SCAN_IN), .A2(n7332), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5577), .ZN(n5442) );
  OAI211_X1 U6186 ( .C1(n7294), .C2(n5443), .A(n5442), .B(n7291), .ZN(n5448)
         );
  AOI21_X1 U6187 ( .B1(n7339), .B2(n5603), .A(n5444), .ZN(n5446) );
  NAND2_X1 U6188 ( .A1(n7337), .A2(n7096), .ZN(n5445) );
  OAI211_X1 U6189 ( .C1(n5600), .C2(n7325), .A(n5446), .B(n5445), .ZN(n5447)
         );
  OR2_X1 U6190 ( .A1(n5448), .A2(n5447), .ZN(U2818) );
  INV_X1 U6191 ( .A(DATAI_10_), .ZN(n5890) );
  INV_X1 U6192 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6820) );
  OAI222_X1 U6193 ( .A1(n5648), .A2(n7581), .B1(n6481), .B2(n5890), .C1(n6479), 
        .C2(n6820), .ZN(U2881) );
  AND2_X1 U6194 ( .A1(n5449), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5453)
         );
  INV_X1 U6195 ( .A(n5453), .ZN(n5495) );
  NOR3_X1 U6196 ( .A1(n7364), .A2(n7363), .A3(n7496), .ZN(n6726) );
  OAI21_X1 U6197 ( .B1(n5458), .B2(n6962), .A(n5451), .ZN(n5454) );
  NAND2_X1 U6198 ( .A1(n7460), .A2(n5452), .ZN(n7451) );
  INV_X1 U6199 ( .A(n7451), .ZN(n5607) );
  AOI21_X1 U6200 ( .B1(n5607), .B2(n7462), .A(n5453), .ZN(n5457) );
  NAND2_X1 U6201 ( .A1(n5454), .A2(n5457), .ZN(n5455) );
  OAI211_X1 U6202 ( .C1(n7499), .C2(n6726), .A(n7513), .B(n5455), .ZN(n5487)
         );
  NAND2_X1 U6203 ( .A1(n5487), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5462)
         );
  INV_X1 U6204 ( .A(n6726), .ZN(n5456) );
  OAI22_X1 U6205 ( .A1(n5457), .A2(n7511), .B1(n5456), .B2(n7505), .ZN(n5492)
         );
  INV_X1 U6206 ( .A(n6771), .ZN(n5490) );
  OAI22_X1 U6207 ( .A1(n5490), .A2(n5542), .B1(n5459), .B2(n5488), .ZN(n5460)
         );
  AOI21_X1 U6208 ( .B1(n7600), .B2(n5492), .A(n5460), .ZN(n5461) );
  OAI211_X1 U6209 ( .C1(n5495), .C2(n5628), .A(n5462), .B(n5461), .ZN(U3144)
         );
  NAND2_X1 U6210 ( .A1(n5487), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5466)
         );
  OAI22_X1 U6211 ( .A1(n5490), .A2(n5550), .B1(n5463), .B2(n5488), .ZN(n5464)
         );
  AOI21_X1 U6212 ( .B1(n7573), .B2(n5492), .A(n5464), .ZN(n5465) );
  OAI211_X1 U6213 ( .C1(n5495), .C2(n5631), .A(n5466), .B(n5465), .ZN(U3143)
         );
  NAND2_X1 U6214 ( .A1(n5487), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5470)
         );
  OAI22_X1 U6215 ( .A1(n5490), .A2(n5546), .B1(n5467), .B2(n5488), .ZN(n5468)
         );
  AOI21_X1 U6216 ( .B1(n7676), .B2(n5492), .A(n5468), .ZN(n5469) );
  OAI211_X1 U6217 ( .C1(n5495), .C2(n5616), .A(n5470), .B(n5469), .ZN(U3147)
         );
  NAND2_X1 U6218 ( .A1(n5487), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5474)
         );
  OAI22_X1 U6219 ( .A1(n5490), .A2(n5567), .B1(n5471), .B2(n5488), .ZN(n5472)
         );
  AOI21_X1 U6220 ( .B1(n7618), .B2(n5492), .A(n5472), .ZN(n5473) );
  OAI211_X1 U6221 ( .C1(n5495), .C2(n5625), .A(n5474), .B(n5473), .ZN(U3145)
         );
  NAND2_X1 U6222 ( .A1(n5487), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5478)
         );
  OAI22_X1 U6223 ( .A1(n5490), .A2(n5558), .B1(n5475), .B2(n5488), .ZN(n5476)
         );
  AOI21_X1 U6224 ( .B1(n6765), .B2(n5492), .A(n5476), .ZN(n5477) );
  OAI211_X1 U6225 ( .C1(n5495), .C2(n5622), .A(n5478), .B(n5477), .ZN(U3146)
         );
  NAND2_X1 U6226 ( .A1(n5487), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5482)
         );
  OAI22_X1 U6227 ( .A1(n5490), .A2(n5538), .B1(n5479), .B2(n5488), .ZN(n5480)
         );
  AOI21_X1 U6228 ( .B1(n7555), .B2(n5492), .A(n5480), .ZN(n5481) );
  OAI211_X1 U6229 ( .C1(n5495), .C2(n5634), .A(n5482), .B(n5481), .ZN(U3142)
         );
  NAND2_X1 U6230 ( .A1(n5487), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5486)
         );
  OAI22_X1 U6231 ( .A1(n5490), .A2(n5562), .B1(n5483), .B2(n5488), .ZN(n5484)
         );
  AOI21_X1 U6232 ( .B1(n6740), .B2(n5492), .A(n5484), .ZN(n5485) );
  OAI211_X1 U6233 ( .C1(n5495), .C2(n5642), .A(n5486), .B(n5485), .ZN(U3140)
         );
  NAND2_X1 U6234 ( .A1(n5487), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5494)
         );
  OAI22_X1 U6235 ( .A1(n5490), .A2(n5554), .B1(n5489), .B2(n5488), .ZN(n5491)
         );
  AOI21_X1 U6236 ( .B1(n7537), .B2(n5492), .A(n5491), .ZN(n5493) );
  OAI211_X1 U6237 ( .C1(n5495), .C2(n5619), .A(n5494), .B(n5493), .ZN(U3141)
         );
  NOR2_X1 U6238 ( .A1(n7502), .A2(n5500), .ZN(n5496) );
  INV_X1 U6239 ( .A(n5496), .ZN(n5523) );
  AOI21_X1 U6240 ( .B1(n5607), .B2(n7473), .A(n5496), .ZN(n5502) );
  NOR2_X1 U6241 ( .A1(n5497), .A2(n7511), .ZN(n5499) );
  AOI22_X1 U6242 ( .A1(n5502), .A2(n5499), .B1(n7511), .B2(n5500), .ZN(n5498)
         );
  NAND2_X1 U6243 ( .A1(n7513), .A2(n5498), .ZN(n5519) );
  INV_X1 U6244 ( .A(n5499), .ZN(n5501) );
  OAI22_X1 U6245 ( .A1(n5502), .A2(n5501), .B1(n7505), .B2(n5500), .ZN(n5518)
         );
  AOI22_X1 U6246 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5519), .B1(n7555), 
        .B2(n5518), .ZN(n5505) );
  NOR2_X2 U6247 ( .A1(n5503), .A2(n3662), .ZN(n6772) );
  AOI22_X1 U6248 ( .A1(n5520), .A2(n7556), .B1(n6772), .B2(n7557), .ZN(n5504)
         );
  OAI211_X1 U6249 ( .C1(n5523), .C2(n5634), .A(n5505), .B(n5504), .ZN(U3126)
         );
  AOI22_X1 U6250 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5519), .B1(n7618), 
        .B2(n5518), .ZN(n5507) );
  AOI22_X1 U6251 ( .A1(n5520), .A2(n7619), .B1(n6772), .B2(n7620), .ZN(n5506)
         );
  OAI211_X1 U6252 ( .C1(n5523), .C2(n5625), .A(n5507), .B(n5506), .ZN(U3129)
         );
  AOI22_X1 U6253 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5519), .B1(n7600), 
        .B2(n5518), .ZN(n5509) );
  AOI22_X1 U6254 ( .A1(n5520), .A2(n7601), .B1(n6772), .B2(n7602), .ZN(n5508)
         );
  OAI211_X1 U6255 ( .C1(n5523), .C2(n5628), .A(n5509), .B(n5508), .ZN(U3128)
         );
  AOI22_X1 U6256 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5519), .B1(n6740), 
        .B2(n5518), .ZN(n5511) );
  AOI22_X1 U6257 ( .A1(n7516), .A2(n5520), .B1(n6772), .B2(n7508), .ZN(n5510)
         );
  OAI211_X1 U6258 ( .C1(n5523), .C2(n5642), .A(n5511), .B(n5510), .ZN(U3124)
         );
  AOI22_X1 U6259 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5519), .B1(n7573), 
        .B2(n5518), .ZN(n5513) );
  AOI22_X1 U6260 ( .A1(n5520), .A2(n7574), .B1(n6772), .B2(n7575), .ZN(n5512)
         );
  OAI211_X1 U6261 ( .C1(n5523), .C2(n5631), .A(n5513), .B(n5512), .ZN(U3127)
         );
  AOI22_X1 U6262 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5519), .B1(n7537), 
        .B2(n5518), .ZN(n5515) );
  AOI22_X1 U6263 ( .A1(n5520), .A2(n7538), .B1(n6772), .B2(n7539), .ZN(n5514)
         );
  OAI211_X1 U6264 ( .C1(n5523), .C2(n5619), .A(n5515), .B(n5514), .ZN(U3125)
         );
  AOI22_X1 U6265 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5519), .B1(n7676), 
        .B2(n5518), .ZN(n5517) );
  AOI22_X1 U6266 ( .A1(n5520), .A2(n7678), .B1(n6772), .B2(n7679), .ZN(n5516)
         );
  OAI211_X1 U6267 ( .C1(n5523), .C2(n5616), .A(n5517), .B(n5516), .ZN(U3131)
         );
  AOI22_X1 U6268 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5519), .B1(n6765), 
        .B2(n5518), .ZN(n5522) );
  AOI22_X1 U6269 ( .A1(n5520), .A2(n7634), .B1(n6772), .B2(n7633), .ZN(n5521)
         );
  OAI211_X1 U6270 ( .C1(n5523), .C2(n5622), .A(n5522), .B(n5521), .ZN(U3130)
         );
  NOR2_X1 U6271 ( .A1(n5605), .A2(n3662), .ZN(n5637) );
  AOI21_X1 U6272 ( .B1(n5527), .B2(STATEBS16_REG_SCAN_IN), .A(n7511), .ZN(
        n5535) );
  NOR2_X1 U6273 ( .A1(n5528), .A2(n7450), .ZN(n5531) );
  NAND2_X1 U6274 ( .A1(n5529), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6736) );
  INV_X1 U6275 ( .A(n6736), .ZN(n5532) );
  AOI22_X1 U6276 ( .A1(n5535), .A2(n5531), .B1(n5532), .B2(n5530), .ZN(n5572)
         );
  NOR3_X1 U6277 ( .A1(n7364), .A2(n7496), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n7453) );
  INV_X1 U6278 ( .A(n7453), .ZN(n7448) );
  NOR2_X1 U6279 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7448), .ZN(n5570)
         );
  INV_X1 U6280 ( .A(n5531), .ZN(n5534) );
  NOR2_X1 U6281 ( .A1(n5532), .A2(n7505), .ZN(n6728) );
  AOI211_X1 U6282 ( .C1(n5535), .C2(n5534), .A(n5533), .B(n6728), .ZN(n5536)
         );
  AOI22_X1 U6283 ( .A1(n7640), .A2(n7557), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5565), .ZN(n5537) );
  OAI21_X1 U6284 ( .B1(n5568), .B2(n5538), .A(n5537), .ZN(n5539) );
  AOI21_X1 U6285 ( .B1(n7554), .B2(n5570), .A(n5539), .ZN(n5540) );
  OAI21_X1 U6286 ( .B1(n5572), .B2(n7553), .A(n5540), .ZN(U3102) );
  AOI22_X1 U6287 ( .A1(n7640), .A2(n7602), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5565), .ZN(n5541) );
  OAI21_X1 U6288 ( .B1(n5568), .B2(n5542), .A(n5541), .ZN(n5543) );
  AOI21_X1 U6289 ( .B1(n7599), .B2(n5570), .A(n5543), .ZN(n5544) );
  OAI21_X1 U6290 ( .B1(n5572), .B2(n7598), .A(n5544), .ZN(U3104) );
  AOI22_X1 U6291 ( .A1(n7640), .A2(n7679), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5565), .ZN(n5545) );
  OAI21_X1 U6292 ( .B1(n5568), .B2(n5546), .A(n5545), .ZN(n5547) );
  AOI21_X1 U6293 ( .B1(n7674), .B2(n5570), .A(n5547), .ZN(n5548) );
  OAI21_X1 U6294 ( .B1(n5572), .B2(n7671), .A(n5548), .ZN(U3107) );
  AOI22_X1 U6295 ( .A1(n7640), .A2(n7575), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5565), .ZN(n5549) );
  OAI21_X1 U6296 ( .B1(n5568), .B2(n5550), .A(n5549), .ZN(n5551) );
  AOI21_X1 U6297 ( .B1(n7572), .B2(n5570), .A(n5551), .ZN(n5552) );
  OAI21_X1 U6298 ( .B1(n5572), .B2(n7571), .A(n5552), .ZN(U3103) );
  AOI22_X1 U6299 ( .A1(n7640), .A2(n7539), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5565), .ZN(n5553) );
  OAI21_X1 U6300 ( .B1(n5568), .B2(n5554), .A(n5553), .ZN(n5555) );
  AOI21_X1 U6301 ( .B1(n7536), .B2(n5570), .A(n5555), .ZN(n5556) );
  OAI21_X1 U6302 ( .B1(n5572), .B2(n7535), .A(n5556), .ZN(U3101) );
  AOI22_X1 U6303 ( .A1(n7640), .A2(n7633), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5565), .ZN(n5557) );
  OAI21_X1 U6304 ( .B1(n5568), .B2(n5558), .A(n5557), .ZN(n5559) );
  AOI21_X1 U6305 ( .B1(n7632), .B2(n5570), .A(n5559), .ZN(n5560) );
  OAI21_X1 U6306 ( .B1(n5572), .B2(n7637), .A(n5560), .ZN(U3106) );
  AOI22_X1 U6307 ( .A1(n7640), .A2(n7508), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5565), .ZN(n5561) );
  OAI21_X1 U6308 ( .B1(n5568), .B2(n5562), .A(n5561), .ZN(n5563) );
  AOI21_X1 U6309 ( .B1(n7507), .B2(n5570), .A(n5563), .ZN(n5564) );
  OAI21_X1 U6310 ( .B1(n5572), .B2(n7519), .A(n5564), .ZN(U3100) );
  AOI22_X1 U6311 ( .A1(n7640), .A2(n7620), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5565), .ZN(n5566) );
  OAI21_X1 U6312 ( .B1(n5568), .B2(n5567), .A(n5566), .ZN(n5569) );
  AOI21_X1 U6313 ( .B1(n7617), .B2(n5570), .A(n5569), .ZN(n5571) );
  OAI21_X1 U6314 ( .B1(n5572), .B2(n7616), .A(n5571), .ZN(U3105) );
  INV_X1 U6315 ( .A(n5425), .ZN(n5576) );
  INV_X1 U6316 ( .A(n5573), .ZN(n5574) );
  OAI21_X1 U6317 ( .B1(n5576), .B2(n5575), .A(n5574), .ZN(n5668) );
  NAND3_X1 U6318 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        n7218), .ZN(n5591) );
  INV_X1 U6319 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6850) );
  NAND3_X1 U6320 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_11__SCAN_IN), .ZN(n7232) );
  AOI21_X1 U6321 ( .B1(n7232), .B2(n7151), .A(n5577), .ZN(n7242) );
  INV_X1 U6322 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5588) );
  INV_X1 U6323 ( .A(n5584), .ZN(n5583) );
  NAND2_X1 U6324 ( .A1(n5759), .A2(n5588), .ZN(n5581) );
  NAND2_X1 U6325 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5578) );
  OAI211_X1 U6326 ( .C1(n4786), .C2(EBX_REG_11__SCAN_IN), .A(n5579), .B(n5578), 
        .ZN(n5580) );
  AND2_X1 U6327 ( .A1(n5581), .A2(n5580), .ZN(n5585) );
  INV_X1 U6328 ( .A(n5585), .ZN(n5582) );
  OAI21_X1 U6329 ( .B1(n5586), .B2(n5583), .A(n5582), .ZN(n5587) );
  NAND2_X1 U6330 ( .A1(n5587), .A2(n5657), .ZN(n5594) );
  OAI22_X1 U6331 ( .A1(n5588), .A2(n7312), .B1(n7329), .B2(n5594), .ZN(n5589)
         );
  AOI211_X1 U6332 ( .C1(n7335), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n7279), 
        .B(n5589), .ZN(n5590) );
  OAI221_X1 U6333 ( .B1(REIP_REG_11__SCAN_IN), .B2(n5591), .C1(n6850), .C2(
        n7242), .A(n5590), .ZN(n5592) );
  AOI21_X1 U6334 ( .B1(n5665), .B2(n7339), .A(n5592), .ZN(n5593) );
  OAI21_X1 U6335 ( .B1(n5668), .B2(n7325), .A(n5593), .ZN(U2816) );
  INV_X1 U6336 ( .A(n5594), .ZN(n7105) );
  AOI22_X1 U6337 ( .A1(n6924), .A2(n7105), .B1(EBX_REG_11__SCAN_IN), .B2(n6426), .ZN(n5595) );
  OAI21_X1 U6338 ( .B1(n5668), .B2(n6454), .A(n5595), .ZN(U2848) );
  OAI21_X1 U6339 ( .B1(n5596), .B2(n5599), .A(n5597), .ZN(n7097) );
  NAND2_X1 U6340 ( .A1(n7073), .A2(REIP_REG_9__SCAN_IN), .ZN(n7094) );
  OAI21_X1 U6341 ( .B1(n6965), .B2(n5443), .A(n7094), .ZN(n5602) );
  NOR2_X1 U6342 ( .A1(n5600), .A2(n6962), .ZN(n5601) );
  AOI211_X1 U6343 ( .C1(n6941), .C2(n5603), .A(n5602), .B(n5601), .ZN(n5604)
         );
  OAI21_X1 U6344 ( .B1(n7345), .B2(n7097), .A(n5604), .ZN(U2977) );
  NOR2_X1 U6345 ( .A1(n7502), .A2(n5611), .ZN(n5606) );
  INV_X1 U6346 ( .A(n5606), .ZN(n5641) );
  OAI21_X1 U6347 ( .B1(n5605), .B2(n7497), .A(n7499), .ZN(n5612) );
  INV_X1 U6348 ( .A(n5612), .ZN(n5608) );
  AOI21_X1 U6349 ( .B1(n5607), .B2(n7503), .A(n5606), .ZN(n5613) );
  NAND2_X1 U6350 ( .A1(n5608), .A2(n5613), .ZN(n5609) );
  OAI211_X1 U6351 ( .C1(n7499), .C2(n5610), .A(n7513), .B(n5609), .ZN(n5636)
         );
  OAI22_X1 U6352 ( .A1(n5613), .A2(n5612), .B1(n7505), .B2(n5611), .ZN(n5635)
         );
  AOI22_X1 U6353 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5636), .B1(n7676), 
        .B2(n5635), .ZN(n5615) );
  AOI22_X1 U6354 ( .A1(n7678), .A2(n5638), .B1(n5637), .B2(n7679), .ZN(n5614)
         );
  OAI211_X1 U6355 ( .C1(n5616), .C2(n5641), .A(n5615), .B(n5614), .ZN(U3099)
         );
  AOI22_X1 U6356 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5636), .B1(n7537), 
        .B2(n5635), .ZN(n5618) );
  AOI22_X1 U6357 ( .A1(n7538), .A2(n5638), .B1(n5637), .B2(n7539), .ZN(n5617)
         );
  OAI211_X1 U6358 ( .C1(n5619), .C2(n5641), .A(n5618), .B(n5617), .ZN(U3093)
         );
  AOI22_X1 U6359 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5636), .B1(n6765), 
        .B2(n5635), .ZN(n5621) );
  AOI22_X1 U6360 ( .A1(n7634), .A2(n5638), .B1(n5637), .B2(n7633), .ZN(n5620)
         );
  OAI211_X1 U6361 ( .C1(n5622), .C2(n5641), .A(n5621), .B(n5620), .ZN(U3098)
         );
  AOI22_X1 U6362 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5636), .B1(n7618), 
        .B2(n5635), .ZN(n5624) );
  AOI22_X1 U6363 ( .A1(n7619), .A2(n5638), .B1(n5637), .B2(n7620), .ZN(n5623)
         );
  OAI211_X1 U6364 ( .C1(n5625), .C2(n5641), .A(n5624), .B(n5623), .ZN(U3097)
         );
  AOI22_X1 U6365 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5636), .B1(n7600), 
        .B2(n5635), .ZN(n5627) );
  AOI22_X1 U6366 ( .A1(n7601), .A2(n5638), .B1(n5637), .B2(n7602), .ZN(n5626)
         );
  OAI211_X1 U6367 ( .C1(n5628), .C2(n5641), .A(n5627), .B(n5626), .ZN(U3096)
         );
  AOI22_X1 U6368 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5636), .B1(n7573), 
        .B2(n5635), .ZN(n5630) );
  AOI22_X1 U6369 ( .A1(n7574), .A2(n5638), .B1(n5637), .B2(n7575), .ZN(n5629)
         );
  OAI211_X1 U6370 ( .C1(n5631), .C2(n5641), .A(n5630), .B(n5629), .ZN(U3095)
         );
  AOI22_X1 U6371 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5636), .B1(n7555), 
        .B2(n5635), .ZN(n5633) );
  AOI22_X1 U6372 ( .A1(n7556), .A2(n5638), .B1(n5637), .B2(n7557), .ZN(n5632)
         );
  OAI211_X1 U6373 ( .C1(n5634), .C2(n5641), .A(n5633), .B(n5632), .ZN(U3094)
         );
  AOI22_X1 U6374 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5636), .B1(n6740), 
        .B2(n5635), .ZN(n5640) );
  AOI22_X1 U6375 ( .A1(n7516), .A2(n5638), .B1(n5637), .B2(n7508), .ZN(n5639)
         );
  OAI211_X1 U6376 ( .C1(n5642), .C2(n5641), .A(n5640), .B(n5639), .ZN(U3092)
         );
  INV_X1 U6377 ( .A(DATAI_11_), .ZN(n7579) );
  INV_X1 U6378 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6822) );
  OAI222_X1 U6379 ( .A1(n6481), .A2(n7579), .B1(n6479), .B2(n6822), .C1(n7581), 
        .C2(n5668), .ZN(U2880) );
  XNOR2_X1 U6380 ( .A(n6526), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5643)
         );
  NOR2_X1 U6381 ( .A1(n3687), .A2(n5643), .ZN(n5660) );
  AOI21_X1 U6382 ( .B1(n3687), .B2(n5643), .A(n5660), .ZN(n7090) );
  NAND2_X1 U6383 ( .A1(n7090), .A2(n6971), .ZN(n5647) );
  AND2_X1 U6384 ( .A1(n7073), .A2(REIP_REG_10__SCAN_IN), .ZN(n7082) );
  NOR2_X1 U6385 ( .A1(n6975), .A2(n5644), .ZN(n5645) );
  AOI211_X1 U6386 ( .C1(n6969), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n7082), 
        .B(n5645), .ZN(n5646) );
  OAI211_X1 U6387 ( .C1(n6962), .C2(n5648), .A(n5647), .B(n5646), .ZN(U2976)
         );
  OAI21_X1 U6388 ( .B1(n5573), .B2(n5650), .A(n5649), .ZN(n7226) );
  INV_X1 U6389 ( .A(EBX_REG_12__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U6390 ( .A1(n5651), .A2(n7220), .ZN(n5655) );
  NAND2_X1 U6391 ( .A1(n5579), .A2(n5703), .ZN(n5653) );
  NAND2_X1 U6392 ( .A1(n6263), .A2(n7220), .ZN(n5652) );
  NAND3_X1 U6393 ( .A1(n5653), .A2(n5672), .A3(n5652), .ZN(n5654) );
  AND2_X1 U6394 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  OR2_X1 U6395 ( .A1(n5658), .A2(n5675), .ZN(n7219) );
  INV_X1 U6396 ( .A(n7219), .ZN(n5709) );
  AOI22_X1 U6397 ( .A1(n6924), .A2(n5709), .B1(EBX_REG_12__SCAN_IN), .B2(n6426), .ZN(n5659) );
  OAI21_X1 U6398 ( .B1(n7226), .B2(n6454), .A(n5659), .ZN(U2847) );
  INV_X1 U6399 ( .A(DATAI_12_), .ZN(n5886) );
  OAI222_X1 U6400 ( .A1(n6481), .A2(n5886), .B1(n6479), .B2(n4218), .C1(n7581), 
        .C2(n7226), .ZN(U2879) );
  AOI21_X1 U6401 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6526), .A(n5660), 
        .ZN(n5662) );
  MUX2_X1 U6402 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .B(n4727), .S(n6668), 
        .Z(n5661) );
  NOR2_X1 U6403 ( .A1(n5662), .A2(n5661), .ZN(n5701) );
  AOI21_X1 U6404 ( .B1(n5662), .B2(n5661), .A(n5701), .ZN(n7107) );
  NAND2_X1 U6405 ( .A1(n7107), .A2(n6971), .ZN(n5667) );
  INV_X1 U6406 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6407 ( .A1(n7073), .A2(REIP_REG_11__SCAN_IN), .ZN(n7103) );
  OAI21_X1 U6408 ( .B1(n6965), .B2(n5663), .A(n7103), .ZN(n5664) );
  AOI21_X1 U6409 ( .B1(n6941), .B2(n5665), .A(n5664), .ZN(n5666) );
  OAI211_X1 U6410 ( .C1(n6962), .C2(n5668), .A(n5667), .B(n5666), .ZN(U2975)
         );
  OAI21_X1 U6411 ( .B1(n5669), .B2(n5671), .A(n5670), .ZN(n7237) );
  MUX2_X1 U6412 ( .A(n5745), .B(n5672), .S(EBX_REG_13__SCAN_IN), .Z(n5673) );
  OAI21_X1 U6413 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5772), .A(n5673), 
        .ZN(n5677) );
  INV_X1 U6414 ( .A(n5675), .ZN(n5676) );
  INV_X1 U6415 ( .A(n5677), .ZN(n5674) );
  AOI21_X1 U6416 ( .B1(n5677), .B2(n5676), .A(n5694), .ZN(n7233) );
  AOI22_X1 U6417 ( .A1(n6924), .A2(n7233), .B1(EBX_REG_13__SCAN_IN), .B2(n6426), .ZN(n5678) );
  OAI21_X1 U6418 ( .B1(n7237), .B2(n6454), .A(n5678), .ZN(U2846) );
  XNOR2_X1 U6419 ( .A(n6668), .B(n5697), .ZN(n5680) );
  XNOR2_X1 U6420 ( .A(n5679), .B(n5680), .ZN(n6594) );
  NAND2_X1 U6421 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5706) );
  NOR2_X1 U6422 ( .A1(n7010), .A2(n5706), .ZN(n5792) );
  NAND2_X1 U6423 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U6424 ( .A1(n7080), .A2(n5681), .ZN(n7086) );
  NOR2_X1 U6425 ( .A1(n7081), .A2(n7086), .ZN(n5793) );
  INV_X1 U6426 ( .A(n5793), .ZN(n5683) );
  NAND2_X1 U6427 ( .A1(n5682), .A2(n7080), .ZN(n7084) );
  NOR2_X1 U6428 ( .A1(n7084), .A2(n7081), .ZN(n7012) );
  OAI21_X1 U6429 ( .B1(n7019), .B2(n7012), .A(n7088), .ZN(n5795) );
  AOI21_X1 U6430 ( .B1(n7087), .B2(n5683), .A(n5795), .ZN(n7110) );
  NAND2_X1 U6431 ( .A1(n7087), .A2(n5793), .ZN(n5696) );
  NAND3_X1 U6432 ( .A1(n5684), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n7012), 
        .ZN(n5685) );
  AOI211_X1 U6433 ( .C1(n5696), .C2(n5685), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n5706), .ZN(n7009) );
  AOI21_X1 U6434 ( .B1(n5706), .B2(n5686), .A(n7009), .ZN(n5687) );
  OAI211_X1 U6435 ( .C1(n5792), .C2(n5688), .A(n7110), .B(n5687), .ZN(n7008)
         );
  OR2_X1 U6436 ( .A1(n5763), .A2(EBX_REG_14__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U6437 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U6438 ( .A1(n5579), .A2(n5689), .ZN(n5690) );
  OAI21_X1 U6439 ( .B1(EBX_REG_14__SCAN_IN), .B2(n4786), .A(n5690), .ZN(n5691)
         );
  NAND2_X1 U6440 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  NAND2_X1 U6441 ( .A1(n5694), .A2(n5693), .ZN(n5721) );
  OR2_X1 U6442 ( .A1(n5694), .A2(n5693), .ZN(n5695) );
  NAND2_X1 U6443 ( .A1(n5721), .A2(n5695), .ZN(n7245) );
  INV_X1 U6444 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6854) );
  OAI22_X1 U6445 ( .A1(n7042), .A2(n7245), .B1(n6854), .B2(n7136), .ZN(n5699)
         );
  NAND2_X1 U6446 ( .A1(n7068), .A2(n7012), .ZN(n6689) );
  AND3_X1 U6447 ( .A1(n5792), .A2(n5697), .A3(n7106), .ZN(n5698) );
  AOI211_X1 U6448 ( .C1(n7008), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5699), .B(n5698), .ZN(n5700) );
  OAI21_X1 U6449 ( .B1(n6594), .B2(n7055), .A(n5700), .ZN(U3004) );
  AOI21_X1 U6450 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6526), .A(n5701), 
        .ZN(n5705) );
  OAI21_X1 U6451 ( .B1(n5703), .B2(n6668), .A(n5702), .ZN(n5704) );
  XNOR2_X1 U6452 ( .A(n5705), .B(n5704), .ZN(n5716) );
  INV_X1 U6453 ( .A(n5706), .ZN(n7011) );
  OAI221_X1 U6454 ( .B1(n7011), .B2(n6689), .C1(n7011), .C2(n7063), .A(n7110), 
        .ZN(n5707) );
  OAI221_X1 U6455 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .C1(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .C2(n7106), .A(n5707), .ZN(n5711) );
  NAND2_X1 U6456 ( .A1(n7073), .A2(REIP_REG_12__SCAN_IN), .ZN(n5712) );
  INV_X1 U6457 ( .A(n5712), .ZN(n5708) );
  AOI21_X1 U6458 ( .B1(n7132), .B2(n5709), .A(n5708), .ZN(n5710) );
  OAI211_X1 U6459 ( .C1(n5716), .C2(n7055), .A(n5711), .B(n5710), .ZN(U3006)
         );
  INV_X1 U6460 ( .A(DATAI_13_), .ZN(n5882) );
  INV_X1 U6461 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6825) );
  OAI222_X1 U6462 ( .A1(n7237), .A2(n7581), .B1(n6481), .B2(n5882), .C1(n6479), 
        .C2(n6825), .ZN(U2878) );
  OAI21_X1 U6463 ( .B1(n6965), .B2(n7223), .A(n5712), .ZN(n5714) );
  NOR2_X1 U6464 ( .A1(n7226), .A2(n6962), .ZN(n5713) );
  AOI211_X1 U6465 ( .C1(n6941), .C2(n7228), .A(n5714), .B(n5713), .ZN(n5715)
         );
  OAI21_X1 U6466 ( .B1(n5716), .B2(n7345), .A(n5715), .ZN(U2974) );
  NAND3_X1 U6467 ( .A1(n5775), .A2(n5717), .A3(n6479), .ZN(n5719) );
  NOR2_X2 U6468 ( .A1(n7584), .A2(n3923), .ZN(n7585) );
  AOI22_X1 U6469 ( .A1(DATAI_31_), .A2(n7585), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7584), .ZN(n5718) );
  NAND2_X1 U6470 ( .A1(n5719), .A2(n5718), .ZN(U2860) );
  MUX2_X1 U6471 ( .A(n5745), .B(n5672), .S(EBX_REG_15__SCAN_IN), .Z(n5720) );
  OAI21_X1 U6472 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5772), .A(n5720), 
        .ZN(n6380) );
  OR2_X2 U6473 ( .A1(n5721), .A2(n6380), .ZN(n6445) );
  OR2_X1 U6474 ( .A1(n5763), .A2(EBX_REG_16__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U6475 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U6476 ( .A1(n5579), .A2(n5722), .ZN(n5723) );
  OAI21_X1 U6477 ( .B1(EBX_REG_16__SCAN_IN), .B2(n4786), .A(n5723), .ZN(n5724)
         );
  AND2_X1 U6478 ( .A1(n5725), .A2(n5724), .ZN(n6444) );
  OR2_X2 U6479 ( .A1(n6445), .A2(n6444), .ZN(n6447) );
  NAND2_X1 U6480 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5726) );
  OAI211_X1 U6481 ( .C1(n4786), .C2(EBX_REG_17__SCAN_IN), .A(n5579), .B(n5726), 
        .ZN(n5727) );
  OAI21_X1 U6482 ( .B1(n5745), .B2(EBX_REG_17__SCAN_IN), .A(n5727), .ZN(n6438)
         );
  NOR2_X4 U6483 ( .A1(n6447), .A2(n6438), .ZN(n6440) );
  OR2_X1 U6484 ( .A1(n5763), .A2(EBX_REG_18__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U6485 ( .A1(n5579), .A2(n6686), .ZN(n5729) );
  INV_X1 U6486 ( .A(EBX_REG_18__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U6487 ( .A1(n6263), .A2(n7277), .ZN(n5728) );
  NAND3_X1 U6488 ( .A1(n5729), .A2(n5672), .A3(n5728), .ZN(n5730) );
  NAND2_X1 U6489 ( .A1(n5731), .A2(n5730), .ZN(n6431) );
  MUX2_X1 U6490 ( .A(n5745), .B(n5672), .S(EBX_REG_19__SCAN_IN), .Z(n5732) );
  OAI21_X1 U6491 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5772), .A(n5732), 
        .ZN(n6425) );
  OR2_X1 U6492 ( .A1(n5763), .A2(EBX_REG_20__SCAN_IN), .ZN(n5736) );
  INV_X1 U6493 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U6494 ( .A1(n5579), .A2(n6667), .ZN(n5734) );
  INV_X1 U6495 ( .A(EBX_REG_20__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U6496 ( .A1(n6263), .A2(n7313), .ZN(n5733) );
  NAND3_X1 U6497 ( .A1(n5734), .A2(n5672), .A3(n5733), .ZN(n5735) );
  AND2_X1 U6498 ( .A1(n5736), .A2(n5735), .ZN(n6414) );
  INV_X1 U6499 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U6500 ( .A1(n5759), .A2(n6407), .ZN(n5739) );
  NAND2_X1 U6501 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U6502 ( .C1(n4786), .C2(EBX_REG_21__SCAN_IN), .A(n5579), .B(n5737), 
        .ZN(n5738) );
  AND2_X1 U6503 ( .A1(n5739), .A2(n5738), .ZN(n6367) );
  OR2_X1 U6504 ( .A1(n5763), .A2(EBX_REG_22__SCAN_IN), .ZN(n5743) );
  INV_X1 U6505 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U6506 ( .A1(n5579), .A2(n6548), .ZN(n5741) );
  INV_X1 U6507 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U6508 ( .A1(n6263), .A2(n6404), .ZN(n5740) );
  NAND3_X1 U6509 ( .A1(n5741), .A2(n5672), .A3(n5740), .ZN(n5742) );
  NAND2_X1 U6510 ( .A1(n5743), .A2(n5742), .ZN(n6401) );
  MUX2_X1 U6511 ( .A(n5745), .B(n5672), .S(EBX_REG_23__SCAN_IN), .Z(n5744) );
  OAI21_X1 U6512 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5772), .A(n5744), 
        .ZN(n6356) );
  MUX2_X1 U6513 ( .A(n5745), .B(n5672), .S(EBX_REG_25__SCAN_IN), .Z(n5747) );
  OR2_X1 U6514 ( .A1(n5772), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5746)
         );
  AND2_X1 U6515 ( .A1(n5747), .A2(n5746), .ZN(n6337) );
  OR2_X1 U6516 ( .A1(n5763), .A2(EBX_REG_24__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U6517 ( .A1(n5579), .A2(n5748), .ZN(n5750) );
  INV_X1 U6518 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U6519 ( .A1(n6263), .A2(n6915), .ZN(n5749) );
  NAND3_X1 U6520 ( .A1(n5750), .A2(n5672), .A3(n5749), .ZN(n5751) );
  NAND2_X1 U6521 ( .A1(n5752), .A2(n5751), .ZN(n6631) );
  NAND2_X1 U6522 ( .A1(n6337), .A2(n6631), .ZN(n5753) );
  OR2_X1 U6523 ( .A1(n5763), .A2(EBX_REG_26__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U6524 ( .A1(n5579), .A2(n6623), .ZN(n5756) );
  INV_X1 U6525 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U6526 ( .A1(n6263), .A2(n5754), .ZN(n5755) );
  NAND3_X1 U6527 ( .A1(n5756), .A2(n5672), .A3(n5755), .ZN(n5757) );
  INV_X1 U6528 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U6529 ( .A1(n5759), .A2(n6920), .ZN(n5762) );
  NAND2_X1 U6530 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5760) );
  OAI211_X1 U6531 ( .C1(n4786), .C2(EBX_REG_27__SCAN_IN), .A(n5579), .B(n5760), 
        .ZN(n5761) );
  AND2_X1 U6532 ( .A1(n5762), .A2(n5761), .ZN(n6307) );
  OR2_X1 U6533 ( .A1(n5763), .A2(EBX_REG_28__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U6534 ( .A1(n5672), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U6535 ( .A1(n5579), .A2(n5764), .ZN(n5765) );
  OAI21_X1 U6536 ( .B1(EBX_REG_28__SCAN_IN), .B2(n4786), .A(n5765), .ZN(n5766)
         );
  AND2_X1 U6537 ( .A1(n5767), .A2(n5766), .ZN(n6296) );
  INV_X1 U6538 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U6539 ( .A1(n6263), .A2(n6391), .ZN(n5769) );
  OR2_X1 U6540 ( .A1(n5772), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5768)
         );
  NAND2_X1 U6541 ( .A1(n5768), .A2(n5769), .ZN(n6267) );
  MUX2_X1 U6542 ( .A(n5769), .B(n6267), .S(n5672), .Z(n5817) );
  OAI22_X1 U6543 ( .A1(n5772), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n4786), .ZN(n6270) );
  NAND2_X1 U6544 ( .A1(n6268), .A2(n6270), .ZN(n5770) );
  OAI22_X1 U6545 ( .A1(n5772), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4786), .ZN(n5773) );
  OAI22_X1 U6546 ( .A1(n5803), .A2(n6916), .B1(n6927), .B2(n5777), .ZN(U2828)
         );
  INV_X1 U6547 ( .A(n5776), .ZN(n5780) );
  NOR4_X1 U6548 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n5789)
         );
  INV_X1 U6549 ( .A(REIP_REG_25__SCAN_IN), .ZN(n7135) );
  INV_X1 U6550 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6867) );
  INV_X1 U6551 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7320) );
  INV_X1 U6552 ( .A(REIP_REG_20__SCAN_IN), .ZN(n7304) );
  INV_X1 U6553 ( .A(REIP_REG_18__SCAN_IN), .ZN(n7280) );
  INV_X1 U6554 ( .A(REIP_REG_13__SCAN_IN), .ZN(n7243) );
  INV_X1 U6555 ( .A(REIP_REG_12__SCAN_IN), .ZN(n7231) );
  NOR4_X1 U6556 ( .A1(n7232), .A2(n7243), .A3(n6854), .A4(n7231), .ZN(n6382)
         );
  INV_X1 U6557 ( .A(REIP_REG_17__SCAN_IN), .ZN(n7123) );
  INV_X1 U6558 ( .A(REIP_REG_16__SCAN_IN), .ZN(n7258) );
  NOR2_X1 U6559 ( .A1(n7123), .A2(n7258), .ZN(n7282) );
  NAND4_X1 U6560 ( .A1(n5781), .A2(n6382), .A3(n7282), .A4(
        REIP_REG_15__SCAN_IN), .ZN(n7267) );
  NOR2_X1 U6561 ( .A1(n7280), .A2(n7267), .ZN(n7290) );
  NAND2_X1 U6562 ( .A1(REIP_REG_19__SCAN_IN), .A2(n7290), .ZN(n7305) );
  NOR2_X1 U6563 ( .A1(n7304), .A2(n7305), .ZN(n6370) );
  NAND2_X1 U6564 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6370), .ZN(n6359) );
  NOR3_X1 U6565 ( .A1(n6867), .A2(n7320), .A3(n6359), .ZN(n7334) );
  NAND2_X1 U6566 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7334), .ZN(n6343) );
  NOR2_X1 U6567 ( .A1(n7135), .A2(n6343), .ZN(n6325) );
  NAND2_X1 U6568 ( .A1(n6325), .A2(REIP_REG_26__SCAN_IN), .ZN(n5782) );
  NOR2_X1 U6569 ( .A1(n7316), .A2(n5782), .ZN(n6311) );
  AND2_X1 U6570 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n5784) );
  NAND2_X1 U6571 ( .A1(n6311), .A2(n5784), .ZN(n6282) );
  NAND2_X1 U6572 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .ZN(
        n5783) );
  NOR2_X1 U6573 ( .A1(n6282), .A2(n5783), .ZN(n5787) );
  INV_X1 U6574 ( .A(n5783), .ZN(n5786) );
  NAND2_X1 U6575 ( .A1(n6366), .A2(n6325), .ZN(n6324) );
  INV_X1 U6576 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6872) );
  NOR2_X1 U6577 ( .A1(n6324), .A2(n6872), .ZN(n6310) );
  NAND2_X1 U6578 ( .A1(n6310), .A2(n5784), .ZN(n5785) );
  NAND2_X1 U6579 ( .A1(n7266), .A2(n5785), .ZN(n6301) );
  OAI21_X1 U6580 ( .B1(n5786), .B2(n7316), .A(n6301), .ZN(n6278) );
  MUX2_X1 U6581 ( .A(n5787), .B(n6278), .S(REIP_REG_31__SCAN_IN), .Z(n5788) );
  AOI211_X1 U6582 ( .C1(PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n7335), .A(n5789), 
        .B(n5788), .ZN(n5790) );
  OAI211_X1 U6583 ( .C1(n5803), .C2(n7329), .A(n5791), .B(n5790), .ZN(U2796)
         );
  AND2_X1 U6584 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6626) );
  INV_X1 U6585 ( .A(n6651), .ZN(n5798) );
  INV_X1 U6586 ( .A(n7040), .ZN(n6698) );
  NAND2_X1 U6587 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5792), .ZN(n6697) );
  NAND2_X1 U6588 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6700) );
  NOR2_X1 U6589 ( .A1(n6697), .A2(n6700), .ZN(n5794) );
  NAND2_X1 U6590 ( .A1(n5793), .A2(n5794), .ZN(n6671) );
  INV_X1 U6591 ( .A(n6525), .ZN(n6677) );
  NOR3_X1 U6592 ( .A1(n6671), .A2(n6677), .A3(n6674), .ZN(n5797) );
  INV_X1 U6593 ( .A(n7019), .ZN(n7085) );
  INV_X1 U6594 ( .A(n5794), .ZN(n5796) );
  AOI21_X1 U6595 ( .B1(n7085), .B2(n5796), .A(n5795), .ZN(n6672) );
  OAI21_X1 U6596 ( .B1(n7040), .B2(n5797), .A(n6672), .ZN(n6661) );
  AOI21_X1 U6597 ( .B1(n5798), .B2(n6698), .A(n6661), .ZN(n6643) );
  OAI21_X1 U6598 ( .B1(n4738), .B2(n5799), .A(n6643), .ZN(n7138) );
  INV_X1 U6599 ( .A(n7138), .ZN(n6634) );
  OAI21_X1 U6600 ( .B1(n6626), .B2(n7040), .A(n6634), .ZN(n6618) );
  AOI21_X1 U6601 ( .B1(n5809), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n7040), 
        .ZN(n5800) );
  NOR2_X1 U6602 ( .A1(n6618), .A2(n5800), .ZN(n6597) );
  OAI21_X1 U6603 ( .B1(n7040), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n6597), 
        .ZN(n5801) );
  INV_X1 U6604 ( .A(n5801), .ZN(n5805) );
  INV_X1 U6605 ( .A(n5802), .ZN(n5804) );
  INV_X1 U6606 ( .A(n5806), .ZN(n5813) );
  INV_X1 U6607 ( .A(n6697), .ZN(n5807) );
  NAND2_X1 U6608 ( .A1(n7127), .A2(n4736), .ZN(n7006) );
  NAND2_X1 U6609 ( .A1(n6650), .A2(n6651), .ZN(n6633) );
  NAND2_X1 U6610 ( .A1(n7140), .A2(n6626), .ZN(n6610) );
  INV_X1 U6611 ( .A(n5809), .ZN(n5810) );
  NOR2_X1 U6612 ( .A1(n6610), .A2(n5810), .ZN(n6601) );
  NAND4_X1 U6613 ( .A1(n6601), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n5811), .ZN(n5812) );
  OAI211_X1 U6614 ( .C1(n5814), .C2(n7055), .A(n5813), .B(n5812), .ZN(U2987)
         );
  NAND2_X1 U6615 ( .A1(n5816), .A2(n5815), .ZN(n6492) );
  NOR2_X1 U6616 ( .A1(n6492), .A2(n6494), .ZN(n6493) );
  XNOR2_X1 U6617 ( .A(n6294), .B(n5817), .ZN(n6390) );
  NOR2_X1 U6618 ( .A1(n6390), .A2(n7042), .ZN(n5819) );
  NAND2_X1 U6619 ( .A1(n7073), .A2(REIP_REG_29__SCAN_IN), .ZN(n5821) );
  OAI21_X1 U6620 ( .B1(n6597), .B2(n6483), .A(n5821), .ZN(n5818) );
  AOI211_X1 U6621 ( .C1(n6601), .C2(n6483), .A(n5819), .B(n5818), .ZN(n5820)
         );
  INV_X1 U6622 ( .A(n6283), .ZN(n5827) );
  OAI21_X1 U6623 ( .B1(n6965), .B2(n5822), .A(n5821), .ZN(n5823) );
  INV_X1 U6624 ( .A(n5823), .ZN(n5826) );
  INV_X1 U6625 ( .A(n5828), .ZN(n5829) );
  OAI21_X1 U6626 ( .B1(n5830), .B2(n7345), .A(n5829), .ZN(U2957) );
  AOI22_X1 U6627 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput_252), .B1(
        DATAWIDTH_REG_19__SCAN_IN), .B2(keyinput_251), .ZN(n5831) );
  OAI221_X1 U6628 ( .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput_252), .C1(
        DATAWIDTH_REG_19__SCAN_IN), .C2(keyinput_251), .A(n5831), .ZN(n6054)
         );
  OAI22_X1 U6629 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(keyinput_250), .B1(
        DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput_249), .ZN(n5832) );
  AOI221_X1 U6630 ( .B1(DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput_250), .C1(
        keyinput_249), .C2(DATAWIDTH_REG_17__SCAN_IN), .A(n5832), .ZN(n6053)
         );
  INV_X1 U6631 ( .A(keyinput_224), .ZN(n6013) );
  INV_X1 U6632 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6839) );
  INV_X1 U6633 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6862) );
  AOI22_X1 U6634 ( .A1(keyinput_208), .A2(ADDRESS_REG_20__SCAN_IN), .B1(n6862), 
        .B2(keyinput_209), .ZN(n5833) );
  OAI221_X1 U6635 ( .B1(keyinput_208), .B2(ADDRESS_REG_20__SCAN_IN), .C1(n6862), .C2(keyinput_209), .A(n5833), .ZN(n5990) );
  INV_X1 U6636 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6873) );
  INV_X1 U6637 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6876) );
  INV_X1 U6638 ( .A(keyinput_182), .ZN(n5944) );
  INV_X1 U6639 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6901) );
  XOR2_X1 U6640 ( .A(n6901), .B(keyinput_177), .Z(n5942) );
  INV_X1 U6641 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7422) );
  AND2_X1 U6642 ( .A1(keyinput_168), .A2(n7422), .ZN(n5923) );
  AOI22_X1 U6643 ( .A1(BS16_N), .A2(keyinput_162), .B1(READY_N), .B2(
        keyinput_163), .ZN(n5834) );
  OAI221_X1 U6644 ( .B1(BS16_N), .B2(keyinput_162), .C1(READY_N), .C2(
        keyinput_163), .A(n5834), .ZN(n5908) );
  INV_X1 U6645 ( .A(keyinput_161), .ZN(n5906) );
  INV_X1 U6646 ( .A(NA_N), .ZN(n7412) );
  OAI22_X1 U6647 ( .A1(n7425), .A2(keyinput_159), .B1(DATAI_1_), .B2(
        keyinput_158), .ZN(n5835) );
  AOI221_X1 U6648 ( .B1(n7425), .B2(keyinput_159), .C1(keyinput_158), .C2(
        DATAI_1_), .A(n5835), .ZN(n5903) );
  INV_X1 U6649 ( .A(DATAI_16_), .ZN(n5876) );
  INV_X1 U6650 ( .A(DATAI_19_), .ZN(n5871) );
  INV_X1 U6651 ( .A(keyinput_140), .ZN(n5870) );
  INV_X1 U6652 ( .A(DATAI_20_), .ZN(n5868) );
  INV_X1 U6653 ( .A(keyinput_139), .ZN(n5867) );
  INV_X1 U6654 ( .A(DATAI_21_), .ZN(n5863) );
  INV_X1 U6655 ( .A(DATAI_23_), .ZN(n5838) );
  INV_X1 U6656 ( .A(DATAI_22_), .ZN(n5837) );
  AOI22_X1 U6657 ( .A1(n5838), .A2(keyinput_136), .B1(keyinput_137), .B2(n5837), .ZN(n5836) );
  OAI221_X1 U6658 ( .B1(n5838), .B2(keyinput_136), .C1(n5837), .C2(
        keyinput_137), .A(n5836), .ZN(n5862) );
  OAI22_X1 U6659 ( .A1(DATAI_30_), .A2(keyinput_129), .B1(DATAI_31_), .B2(
        keyinput_128), .ZN(n5839) );
  INV_X1 U6660 ( .A(n5839), .ZN(n5847) );
  INV_X1 U6661 ( .A(DATAI_29_), .ZN(n5841) );
  OAI22_X1 U6662 ( .A1(n5841), .A2(keyinput_130), .B1(n5840), .B2(DATAI_29_), 
        .ZN(n5842) );
  INV_X1 U6663 ( .A(n5842), .ZN(n5846) );
  NAND2_X1 U6664 ( .A1(DATAI_31_), .A2(keyinput_128), .ZN(n5844) );
  AND2_X1 U6665 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  NAND3_X1 U6666 ( .A1(n5847), .A2(n5846), .A3(n5845), .ZN(n5851) );
  INV_X1 U6667 ( .A(DATAI_28_), .ZN(n6464) );
  INV_X1 U6668 ( .A(keyinput_131), .ZN(n5848) );
  OAI22_X1 U6669 ( .A1(n6464), .A2(keyinput_131), .B1(n5848), .B2(DATAI_28_), 
        .ZN(n5849) );
  INV_X1 U6670 ( .A(n5849), .ZN(n5850) );
  NAND2_X1 U6671 ( .A1(n5851), .A2(n5850), .ZN(n5856) );
  INV_X1 U6672 ( .A(DATAI_27_), .ZN(n5853) );
  INV_X1 U6673 ( .A(keyinput_132), .ZN(n5852) );
  INV_X1 U6674 ( .A(n5854), .ZN(n5855) );
  NAND2_X1 U6675 ( .A1(n5856), .A2(n5855), .ZN(n5861) );
  OAI22_X1 U6676 ( .A1(DATAI_24_), .A2(keyinput_135), .B1(DATAI_25_), .B2(
        keyinput_134), .ZN(n5858) );
  AOI221_X1 U6677 ( .B1(DATAI_24_), .B2(keyinput_135), .C1(keyinput_134), .C2(
        DATAI_25_), .A(n5858), .ZN(n5859) );
  OAI22_X1 U6678 ( .A1(keyinput_138), .A2(n5863), .B1(n5862), .B2(n3740), .ZN(
        n5865) );
  AND2_X1 U6679 ( .A1(keyinput_138), .A2(n5863), .ZN(n5864) );
  NOR2_X1 U6680 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  AOI221_X1 U6681 ( .B1(DATAI_20_), .B2(keyinput_139), .C1(n5868), .C2(n5867), 
        .A(n5866), .ZN(n5869) );
  AOI221_X1 U6682 ( .B1(DATAI_19_), .B2(keyinput_140), .C1(n5871), .C2(n5870), 
        .A(n5869), .ZN(n5875) );
  INV_X1 U6683 ( .A(DATAI_17_), .ZN(n5873) );
  AOI22_X1 U6684 ( .A1(DATAI_18_), .A2(keyinput_141), .B1(n5873), .B2(
        keyinput_142), .ZN(n5872) );
  OAI221_X1 U6685 ( .B1(DATAI_18_), .B2(keyinput_141), .C1(n5873), .C2(
        keyinput_142), .A(n5872), .ZN(n5874) );
  OAI22_X1 U6686 ( .A1(keyinput_143), .A2(n5876), .B1(n5875), .B2(n5874), .ZN(
        n5877) );
  INV_X1 U6687 ( .A(n5877), .ZN(n5878) );
  AOI22_X1 U6688 ( .A1(DATAI_14_), .A2(keyinput_145), .B1(n6478), .B2(
        keyinput_144), .ZN(n5879) );
  OAI221_X1 U6689 ( .B1(DATAI_14_), .B2(keyinput_145), .C1(n6478), .C2(
        keyinput_144), .A(n5879), .ZN(n5880) );
  INV_X1 U6690 ( .A(n5880), .ZN(n5884) );
  XNOR2_X1 U6691 ( .A(n5886), .B(keyinput_147), .ZN(n5893) );
  AOI22_X1 U6692 ( .A1(n5888), .A2(keyinput_151), .B1(keyinput_148), .B2(n7579), .ZN(n5887) );
  OAI221_X1 U6693 ( .B1(n5888), .B2(keyinput_151), .C1(n7579), .C2(
        keyinput_148), .A(n5887), .ZN(n5892) );
  AOI22_X1 U6694 ( .A1(DATAI_9_), .A2(keyinput_150), .B1(n5890), .B2(
        keyinput_149), .ZN(n5889) );
  OAI221_X1 U6695 ( .B1(DATAI_9_), .B2(keyinput_150), .C1(n5890), .C2(
        keyinput_149), .A(n5889), .ZN(n5891) );
  AOI211_X1 U6696 ( .C1(n5894), .C2(n5893), .A(n5892), .B(n5891), .ZN(n5901)
         );
  AOI22_X1 U6697 ( .A1(DATAI_7_), .A2(keyinput_152), .B1(DATAI_6_), .B2(
        keyinput_153), .ZN(n5895) );
  OAI221_X1 U6698 ( .B1(DATAI_7_), .B2(keyinput_152), .C1(DATAI_6_), .C2(
        keyinput_153), .A(n5895), .ZN(n5900) );
  OAI22_X1 U6699 ( .A1(n7434), .A2(keyinput_157), .B1(DATAI_4_), .B2(
        keyinput_155), .ZN(n5896) );
  AOI221_X1 U6700 ( .B1(n7434), .B2(keyinput_157), .C1(keyinput_155), .C2(
        DATAI_4_), .A(n5896), .ZN(n5899) );
  OAI22_X1 U6701 ( .A1(DATAI_5_), .A2(keyinput_154), .B1(DATAI_3_), .B2(
        keyinput_156), .ZN(n5897) );
  AOI221_X1 U6702 ( .B1(DATAI_5_), .B2(keyinput_154), .C1(keyinput_156), .C2(
        DATAI_3_), .A(n5897), .ZN(n5898) );
  OAI211_X1 U6703 ( .C1(n5901), .C2(n5900), .A(n5899), .B(n5898), .ZN(n5902)
         );
  OAI211_X1 U6704 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_160), .A(n5903), 
        .B(n5902), .ZN(n5904) );
  AOI21_X1 U6705 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_160), .A(n5904), 
        .ZN(n5905) );
  AOI221_X1 U6706 ( .B1(NA_N), .B2(n5906), .C1(n7412), .C2(keyinput_161), .A(
        n5905), .ZN(n5907) );
  OAI22_X1 U6707 ( .A1(n5908), .A2(n5907), .B1(keyinput_164), .B2(HOLD), .ZN(
        n5909) );
  AOI21_X1 U6708 ( .B1(keyinput_164), .B2(HOLD), .A(n5909), .ZN(n5910) );
  INV_X1 U6709 ( .A(n5910), .ZN(n5914) );
  INV_X1 U6710 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6984) );
  INV_X1 U6711 ( .A(keyinput_165), .ZN(n5911) );
  NAND2_X1 U6712 ( .A1(n6984), .A2(n5911), .ZN(n5913) );
  INV_X1 U6713 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6977) );
  INV_X1 U6714 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6797) );
  AOI22_X1 U6715 ( .A1(n6977), .A2(keyinput_167), .B1(keyinput_166), .B2(n6797), .ZN(n5915) );
  OAI221_X1 U6716 ( .B1(n6977), .B2(keyinput_167), .C1(n6797), .C2(
        keyinput_166), .A(n5915), .ZN(n5916) );
  INV_X1 U6717 ( .A(n5916), .ZN(n5917) );
  NAND2_X1 U6718 ( .A1(n5918), .A2(n5917), .ZN(n5921) );
  NAND2_X1 U6719 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  NOR2_X1 U6720 ( .A1(n5923), .A2(n5922), .ZN(n5929) );
  INV_X1 U6721 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6987) );
  INV_X1 U6722 ( .A(D_C_N_REG_SCAN_IN), .ZN(n5925) );
  AOI22_X1 U6723 ( .A1(n6987), .A2(keyinput_170), .B1(keyinput_169), .B2(n5925), .ZN(n5924) );
  OAI221_X1 U6724 ( .B1(n6987), .B2(keyinput_170), .C1(n5925), .C2(
        keyinput_169), .A(n5924), .ZN(n5928) );
  INV_X1 U6725 ( .A(MORE_REG_SCAN_IN), .ZN(n7374) );
  OAI22_X1 U6726 ( .A1(n7374), .A2(keyinput_172), .B1(STATEBS16_REG_SCAN_IN), 
        .B2(keyinput_171), .ZN(n5926) );
  AOI221_X1 U6727 ( .B1(n7374), .B2(keyinput_172), .C1(keyinput_171), .C2(
        STATEBS16_REG_SCAN_IN), .A(n5926), .ZN(n5927) );
  OAI21_X1 U6728 ( .B1(n5929), .B2(n5928), .A(n5927), .ZN(n5933) );
  INV_X1 U6729 ( .A(keyinput_173), .ZN(n5930) );
  OAI22_X1 U6730 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_174), .B1(
        BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_175), .ZN(n5934) );
  AOI221_X1 U6731 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_174), .C1(
        keyinput_175), .C2(BYTEENABLE_REG_0__SCAN_IN), .A(n5934), .ZN(n5935)
         );
  INV_X1 U6732 ( .A(n5935), .ZN(n5936) );
  INV_X1 U6733 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6906) );
  INV_X1 U6734 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6877) );
  INV_X1 U6735 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6882) );
  AOI22_X1 U6736 ( .A1(n6877), .A2(keyinput_181), .B1(keyinput_180), .B2(n6882), .ZN(n5937) );
  OAI221_X1 U6737 ( .B1(n6877), .B2(keyinput_181), .C1(n6882), .C2(
        keyinput_180), .A(n5937), .ZN(n5940) );
  AOI22_X1 U6738 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_178), .B1(
        REIP_REG_31__SCAN_IN), .B2(keyinput_179), .ZN(n5938) );
  OAI221_X1 U6739 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_178), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput_179), .A(n5938), .ZN(n5939) );
  AOI211_X1 U6740 ( .C1(n5942), .C2(n5941), .A(n5940), .B(n5939), .ZN(n5943)
         );
  AOI221_X1 U6741 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_182), .C1(n6876), 
        .C2(n5944), .A(n5943), .ZN(n5955) );
  AOI22_X1 U6742 ( .A1(n7135), .A2(keyinput_185), .B1(keyinput_184), .B2(n6872), .ZN(n5945) );
  OAI221_X1 U6743 ( .B1(n7135), .B2(keyinput_185), .C1(n6872), .C2(
        keyinput_184), .A(n5945), .ZN(n5946) );
  INV_X1 U6744 ( .A(n5946), .ZN(n5950) );
  INV_X1 U6745 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6874) );
  OR2_X1 U6746 ( .A1(n6874), .A2(keyinput_183), .ZN(n5948) );
  AND2_X1 U6747 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  NAND2_X1 U6748 ( .A1(n5950), .A2(n5949), .ZN(n5954) );
  INV_X1 U6749 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6868) );
  INV_X1 U6750 ( .A(keyinput_186), .ZN(n5951) );
  INV_X1 U6751 ( .A(n5952), .ZN(n5953) );
  OAI21_X1 U6752 ( .B1(n5955), .B2(n5954), .A(n5953), .ZN(n5959) );
  INV_X1 U6753 ( .A(keyinput_187), .ZN(n5956) );
  INV_X1 U6754 ( .A(keyinput_188), .ZN(n5960) );
  OAI22_X1 U6755 ( .A1(n7320), .A2(keyinput_188), .B1(n5960), .B2(
        REIP_REG_22__SCAN_IN), .ZN(n5962) );
  INV_X1 U6756 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6864) );
  XNOR2_X1 U6757 ( .A(n6864), .B(keyinput_189), .ZN(n5961) );
  NAND2_X1 U6758 ( .A1(n5965), .A2(n5964), .ZN(n5972) );
  AOI22_X1 U6759 ( .A1(keyinput_190), .A2(REIP_REG_20__SCAN_IN), .B1(n7280), 
        .B2(keyinput_192), .ZN(n5966) );
  OAI221_X1 U6760 ( .B1(keyinput_190), .B2(REIP_REG_20__SCAN_IN), .C1(n7280), 
        .C2(keyinput_192), .A(n5966), .ZN(n5971) );
  INV_X1 U6761 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6884) );
  OAI22_X1 U6762 ( .A1(n7258), .A2(keyinput_194), .B1(n6884), .B2(keyinput_195), .ZN(n5967) );
  AOI221_X1 U6763 ( .B1(n7258), .B2(keyinput_194), .C1(keyinput_195), .C2(
        n6884), .A(n5967), .ZN(n5970) );
  OAI22_X1 U6764 ( .A1(n7123), .A2(keyinput_193), .B1(BE_N_REG_2__SCAN_IN), 
        .B2(keyinput_196), .ZN(n5968) );
  AOI221_X1 U6765 ( .B1(n7123), .B2(keyinput_193), .C1(keyinput_196), .C2(
        BE_N_REG_2__SCAN_IN), .A(n5968), .ZN(n5969) );
  OAI211_X1 U6766 ( .C1(n5972), .C2(n5971), .A(n5970), .B(n5969), .ZN(n5973)
         );
  INV_X1 U6767 ( .A(n5973), .ZN(n5978) );
  INV_X1 U6768 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n6903) );
  OAI22_X1 U6769 ( .A1(n6903), .A2(keyinput_197), .B1(BE_N_REG_0__SCAN_IN), 
        .B2(keyinput_198), .ZN(n5974) );
  AOI221_X1 U6770 ( .B1(n6903), .B2(keyinput_197), .C1(keyinput_198), .C2(
        BE_N_REG_0__SCAN_IN), .A(n5974), .ZN(n5975) );
  INV_X1 U6771 ( .A(n5975), .ZN(n5977) );
  INV_X1 U6772 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6878) );
  XNOR2_X1 U6773 ( .A(n6878), .B(keyinput_200), .ZN(n5979) );
  OAI22_X1 U6774 ( .A1(n5980), .A2(n5979), .B1(n6873), .B2(keyinput_202), .ZN(
        n5981) );
  AOI21_X1 U6775 ( .B1(n6873), .B2(keyinput_202), .A(n5981), .ZN(n5988) );
  OAI22_X1 U6776 ( .A1(ADDRESS_REG_27__SCAN_IN), .A2(keyinput_201), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(keyinput_203), .ZN(n5982) );
  AOI221_X1 U6777 ( .B1(ADDRESS_REG_27__SCAN_IN), .B2(keyinput_201), .C1(
        keyinput_203), .C2(ADDRESS_REG_25__SCAN_IN), .A(n5982), .ZN(n5987) );
  AOI22_X1 U6778 ( .A1(ADDRESS_REG_23__SCAN_IN), .A2(keyinput_205), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(keyinput_207), .ZN(n5983) );
  OAI221_X1 U6779 ( .B1(ADDRESS_REG_23__SCAN_IN), .B2(keyinput_205), .C1(
        ADDRESS_REG_21__SCAN_IN), .C2(keyinput_207), .A(n5983), .ZN(n5986) );
  AOI22_X1 U6780 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput_204), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(keyinput_206), .ZN(n5984) );
  OAI221_X1 U6781 ( .B1(ADDRESS_REG_24__SCAN_IN), .B2(keyinput_204), .C1(
        ADDRESS_REG_22__SCAN_IN), .C2(keyinput_206), .A(n5984), .ZN(n5985) );
  AOI211_X1 U6782 ( .C1(n5988), .C2(n5987), .A(n5986), .B(n5985), .ZN(n5989)
         );
  OAI22_X1 U6783 ( .A1(n5990), .A2(n5989), .B1(keyinput_210), .B2(
        ADDRESS_REG_18__SCAN_IN), .ZN(n5991) );
  AOI21_X1 U6784 ( .B1(keyinput_210), .B2(ADDRESS_REG_18__SCAN_IN), .A(n5991), 
        .ZN(n5997) );
  INV_X1 U6785 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6857) );
  INV_X1 U6786 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6858) );
  AOI22_X1 U6787 ( .A1(n6857), .A2(keyinput_212), .B1(keyinput_211), .B2(n6858), .ZN(n5992) );
  OAI221_X1 U6788 ( .B1(n6857), .B2(keyinput_212), .C1(n6858), .C2(
        keyinput_211), .A(n5992), .ZN(n5996) );
  OAI22_X1 U6789 ( .A1(ADDRESS_REG_13__SCAN_IN), .A2(keyinput_215), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(keyinput_213), .ZN(n5993) );
  AOI221_X1 U6790 ( .B1(ADDRESS_REG_13__SCAN_IN), .B2(keyinput_215), .C1(
        keyinput_213), .C2(ADDRESS_REG_15__SCAN_IN), .A(n5993), .ZN(n5995) );
  INV_X1 U6791 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6855) );
  XOR2_X1 U6792 ( .A(n6855), .B(keyinput_214), .Z(n5994) );
  OAI211_X1 U6793 ( .C1(n5997), .C2(n5996), .A(n5995), .B(n5994), .ZN(n5998)
         );
  INV_X1 U6794 ( .A(n5998), .ZN(n6004) );
  INV_X1 U6795 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6852) );
  INV_X1 U6796 ( .A(keyinput_216), .ZN(n5999) );
  OAI22_X1 U6797 ( .A1(n6852), .A2(keyinput_216), .B1(n5999), .B2(
        ADDRESS_REG_12__SCAN_IN), .ZN(n6003) );
  INV_X1 U6798 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6851) );
  INV_X1 U6799 ( .A(keyinput_217), .ZN(n6000) );
  OAI22_X1 U6800 ( .A1(n6851), .A2(keyinput_217), .B1(n6000), .B2(
        ADDRESS_REG_11__SCAN_IN), .ZN(n6001) );
  OAI21_X1 U6801 ( .B1(n6004), .B2(n6003), .A(n6002), .ZN(n6011) );
  INV_X1 U6802 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6841) );
  INV_X1 U6803 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6845) );
  OAI22_X1 U6804 ( .A1(n6841), .A2(keyinput_222), .B1(n6845), .B2(keyinput_220), .ZN(n6005) );
  AOI221_X1 U6805 ( .B1(n6841), .B2(keyinput_222), .C1(keyinput_220), .C2(
        n6845), .A(n6005), .ZN(n6010) );
  INV_X1 U6806 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6840) );
  OAI22_X1 U6807 ( .A1(n6840), .A2(keyinput_223), .B1(ADDRESS_REG_7__SCAN_IN), 
        .B2(keyinput_221), .ZN(n6006) );
  AOI221_X1 U6808 ( .B1(n6840), .B2(keyinput_223), .C1(keyinput_221), .C2(
        ADDRESS_REG_7__SCAN_IN), .A(n6006), .ZN(n6009) );
  OAI22_X1 U6809 ( .A1(ADDRESS_REG_9__SCAN_IN), .A2(keyinput_219), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(keyinput_218), .ZN(n6007) );
  AOI221_X1 U6810 ( .B1(ADDRESS_REG_9__SCAN_IN), .B2(keyinput_219), .C1(
        keyinput_218), .C2(ADDRESS_REG_10__SCAN_IN), .A(n6007), .ZN(n6008) );
  NAND2_X1 U6811 ( .A1(n6011), .A2(n3749), .ZN(n6012) );
  OAI221_X1 U6812 ( .B1(ADDRESS_REG_4__SCAN_IN), .B2(n6013), .C1(n6839), .C2(
        keyinput_224), .A(n6012), .ZN(n6018) );
  INV_X1 U6813 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6838) );
  XOR2_X1 U6814 ( .A(n6838), .B(keyinput_225), .Z(n6017) );
  AOI22_X1 U6815 ( .A1(ADDRESS_REG_0__SCAN_IN), .A2(keyinput_228), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(keyinput_227), .ZN(n6014) );
  OAI221_X1 U6816 ( .B1(ADDRESS_REG_0__SCAN_IN), .B2(keyinput_228), .C1(
        ADDRESS_REG_1__SCAN_IN), .C2(keyinput_227), .A(n6014), .ZN(n6016) );
  INV_X1 U6817 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6837) );
  XNOR2_X1 U6818 ( .A(n6837), .B(keyinput_226), .ZN(n6015) );
  AOI21_X1 U6819 ( .B1(n6018), .B2(n6017), .A(n3735), .ZN(n6024) );
  AOI22_X1 U6820 ( .A1(STATE_REG_1__SCAN_IN), .A2(keyinput_230), .B1(
        STATE_REG_2__SCAN_IN), .B2(keyinput_229), .ZN(n6019) );
  OAI221_X1 U6821 ( .B1(STATE_REG_1__SCAN_IN), .B2(keyinput_230), .C1(
        STATE_REG_2__SCAN_IN), .C2(keyinput_229), .A(n6019), .ZN(n6023) );
  INV_X1 U6822 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6899) );
  OAI22_X1 U6823 ( .A1(n6899), .A2(keyinput_232), .B1(STATE_REG_0__SCAN_IN), 
        .B2(keyinput_231), .ZN(n6020) );
  AOI221_X1 U6824 ( .B1(n6899), .B2(keyinput_232), .C1(keyinput_231), .C2(
        STATE_REG_0__SCAN_IN), .A(n6020), .ZN(n6022) );
  XNOR2_X1 U6825 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_233), .ZN(n6021)
         );
  OAI211_X1 U6826 ( .C1(n6024), .C2(n6023), .A(n6022), .B(n6021), .ZN(n6030)
         );
  OAI22_X1 U6827 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(keyinput_234), .B1(
        DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput_235), .ZN(n6025) );
  AOI221_X1 U6828 ( .B1(DATAWIDTH_REG_2__SCAN_IN), .B2(keyinput_234), .C1(
        keyinput_235), .C2(DATAWIDTH_REG_3__SCAN_IN), .A(n6025), .ZN(n6029) );
  INV_X1 U6829 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6027) );
  AOI22_X1 U6830 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(keyinput_237), .B1(n6027), .B2(keyinput_236), .ZN(n6026) );
  OAI221_X1 U6831 ( .B1(DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput_237), .C1(
        n6027), .C2(keyinput_236), .A(n6026), .ZN(n6028) );
  AOI21_X1 U6832 ( .B1(n6030), .B2(n6029), .A(n6028), .ZN(n6042) );
  INV_X1 U6833 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6781) );
  INV_X1 U6834 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6782) );
  OAI22_X1 U6835 ( .A1(n6781), .A2(keyinput_238), .B1(n6782), .B2(keyinput_239), .ZN(n6031) );
  AOI221_X1 U6836 ( .B1(n6781), .B2(keyinput_238), .C1(keyinput_239), .C2(
        n6782), .A(n6031), .ZN(n6032) );
  INV_X1 U6837 ( .A(n6032), .ZN(n6041) );
  INV_X1 U6838 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6783) );
  OAI22_X1 U6839 ( .A1(n6783), .A2(keyinput_240), .B1(
        DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput_243), .ZN(n6033) );
  AOI221_X1 U6840 ( .B1(n6783), .B2(keyinput_240), .C1(keyinput_243), .C2(
        DATAWIDTH_REG_11__SCAN_IN), .A(n6033), .ZN(n6036) );
  INV_X1 U6841 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6784) );
  OAI22_X1 U6842 ( .A1(n6784), .A2(keyinput_241), .B1(
        DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput_245), .ZN(n6034) );
  AOI221_X1 U6843 ( .B1(n6784), .B2(keyinput_241), .C1(keyinput_245), .C2(
        DATAWIDTH_REG_13__SCAN_IN), .A(n6034), .ZN(n6035) );
  INV_X1 U6844 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6785) );
  INV_X1 U6845 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6787) );
  OAI22_X1 U6846 ( .A1(n6785), .A2(keyinput_242), .B1(n6787), .B2(keyinput_244), .ZN(n6037) );
  AOI221_X1 U6847 ( .B1(n6785), .B2(keyinput_242), .C1(keyinput_244), .C2(
        n6787), .A(n6037), .ZN(n6038) );
  OAI21_X1 U6848 ( .B1(n6042), .B2(n6041), .A(n6040), .ZN(n6046) );
  INV_X1 U6849 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6789) );
  OAI22_X1 U6850 ( .A1(n6789), .A2(keyinput_247), .B1(
        DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput_246), .ZN(n6043) );
  AOI221_X1 U6851 ( .B1(n6789), .B2(keyinput_247), .C1(keyinput_246), .C2(
        DATAWIDTH_REG_14__SCAN_IN), .A(n6043), .ZN(n6045) );
  INV_X1 U6852 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6790) );
  AND2_X1 U6853 ( .A1(n6790), .A2(keyinput_248), .ZN(n6044) );
  AOI21_X1 U6854 ( .B1(n6046), .B2(n6045), .A(n6044), .ZN(n6049) );
  NAND2_X1 U6855 ( .A1(n6049), .A2(n6048), .ZN(n6052) );
  INV_X1 U6856 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6793) );
  OAI22_X1 U6857 ( .A1(n6793), .A2(keyinput_254), .B1(
        DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput_253), .ZN(n6050) );
  AOI221_X1 U6858 ( .B1(n6793), .B2(keyinput_254), .C1(keyinput_253), .C2(
        DATAWIDTH_REG_21__SCAN_IN), .A(n6050), .ZN(n6051) );
  OAI221_X1 U6859 ( .B1(n6054), .B2(n6053), .C1(n6052), .C2(n6054), .A(n6051), 
        .ZN(n6236) );
  XOR2_X1 U6860 ( .A(keyinput_127), .B(keyinput_255), .Z(n6235) );
  INV_X1 U6861 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6794) );
  XNOR2_X1 U6862 ( .A(n6794), .B(keyinput_127), .ZN(n6234) );
  XOR2_X1 U6863 ( .A(DATAI_30_), .B(keyinput_1), .Z(n6057) );
  XOR2_X1 U6864 ( .A(DATAI_31_), .B(keyinput_0), .Z(n6056) );
  XNOR2_X1 U6865 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n6055) );
  NAND3_X1 U6866 ( .A1(n6057), .A2(n6056), .A3(n6055), .ZN(n6060) );
  XNOR2_X1 U6867 ( .A(DATAI_28_), .B(keyinput_3), .ZN(n6059) );
  XNOR2_X1 U6868 ( .A(keyinput_4), .B(DATAI_27_), .ZN(n6058) );
  AOI21_X1 U6869 ( .B1(n6060), .B2(n6059), .A(n6058), .ZN(n6064) );
  XOR2_X1 U6870 ( .A(keyinput_5), .B(DATAI_26_), .Z(n6063) );
  XOR2_X1 U6871 ( .A(keyinput_6), .B(DATAI_25_), .Z(n6062) );
  XOR2_X1 U6872 ( .A(keyinput_7), .B(DATAI_24_), .Z(n6061) );
  NOR4_X1 U6873 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n6067)
         );
  XNOR2_X1 U6874 ( .A(keyinput_8), .B(DATAI_23_), .ZN(n6066) );
  XNOR2_X1 U6875 ( .A(keyinput_9), .B(DATAI_22_), .ZN(n6065) );
  NOR3_X1 U6876 ( .A1(n6067), .A2(n6066), .A3(n6065), .ZN(n6070) );
  XOR2_X1 U6877 ( .A(keyinput_10), .B(DATAI_21_), .Z(n6069) );
  XOR2_X1 U6878 ( .A(keyinput_11), .B(DATAI_20_), .Z(n6068) );
  OAI21_X1 U6879 ( .B1(n6070), .B2(n6069), .A(n6068), .ZN(n6074) );
  XOR2_X1 U6880 ( .A(keyinput_12), .B(DATAI_19_), .Z(n6073) );
  XOR2_X1 U6881 ( .A(keyinput_13), .B(DATAI_18_), .Z(n6072) );
  XNOR2_X1 U6882 ( .A(keyinput_14), .B(DATAI_17_), .ZN(n6071) );
  AOI211_X1 U6883 ( .C1(n6074), .C2(n6073), .A(n6072), .B(n6071), .ZN(n6080)
         );
  XNOR2_X1 U6884 ( .A(keyinput_15), .B(DATAI_16_), .ZN(n6079) );
  XOR2_X1 U6885 ( .A(keyinput_16), .B(DATAI_15_), .Z(n6077) );
  XNOR2_X1 U6886 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n6076) );
  XNOR2_X1 U6887 ( .A(DATAI_14_), .B(keyinput_17), .ZN(n6075) );
  NOR3_X1 U6888 ( .A1(n6077), .A2(n6076), .A3(n6075), .ZN(n6078) );
  OAI21_X1 U6889 ( .B1(n6080), .B2(n6079), .A(n6078), .ZN(n6087) );
  XNOR2_X1 U6890 ( .A(DATAI_12_), .B(keyinput_19), .ZN(n6086) );
  XOR2_X1 U6891 ( .A(keyinput_23), .B(DATAI_8_), .Z(n6084) );
  XOR2_X1 U6892 ( .A(keyinput_21), .B(DATAI_10_), .Z(n6083) );
  XNOR2_X1 U6893 ( .A(keyinput_20), .B(DATAI_11_), .ZN(n6082) );
  XNOR2_X1 U6894 ( .A(keyinput_22), .B(DATAI_9_), .ZN(n6081) );
  NAND4_X1 U6895 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), .ZN(n6085)
         );
  AOI21_X1 U6896 ( .B1(n6087), .B2(n6086), .A(n6085), .ZN(n6090) );
  XNOR2_X1 U6897 ( .A(keyinput_24), .B(DATAI_7_), .ZN(n6089) );
  XNOR2_X1 U6898 ( .A(keyinput_25), .B(DATAI_6_), .ZN(n6088) );
  NOR3_X1 U6899 ( .A1(n6090), .A2(n6089), .A3(n6088), .ZN(n6100) );
  XOR2_X1 U6900 ( .A(keyinput_26), .B(DATAI_5_), .Z(n6094) );
  XOR2_X1 U6901 ( .A(keyinput_28), .B(DATAI_3_), .Z(n6093) );
  XNOR2_X1 U6902 ( .A(keyinput_29), .B(DATAI_2_), .ZN(n6092) );
  XNOR2_X1 U6903 ( .A(keyinput_27), .B(DATAI_4_), .ZN(n6091) );
  NAND4_X1 U6904 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n6099)
         );
  XOR2_X1 U6905 ( .A(keyinput_32), .B(MEMORYFETCH_REG_SCAN_IN), .Z(n6097) );
  XOR2_X1 U6906 ( .A(keyinput_31), .B(DATAI_0_), .Z(n6096) );
  XNOR2_X1 U6907 ( .A(keyinput_30), .B(DATAI_1_), .ZN(n6095) );
  NOR3_X1 U6908 ( .A1(n6097), .A2(n6096), .A3(n6095), .ZN(n6098) );
  OAI21_X1 U6909 ( .B1(n6100), .B2(n6099), .A(n6098), .ZN(n6104) );
  XOR2_X1 U6910 ( .A(NA_N), .B(keyinput_33), .Z(n6103) );
  INV_X1 U6911 ( .A(BS16_N), .ZN(n6779) );
  XNOR2_X1 U6912 ( .A(n6779), .B(keyinput_34), .ZN(n6102) );
  XOR2_X1 U6913 ( .A(READY_N), .B(keyinput_35), .Z(n6101) );
  AOI211_X1 U6914 ( .C1(n6104), .C2(n6103), .A(n6102), .B(n6101), .ZN(n6107)
         );
  XNOR2_X1 U6915 ( .A(HOLD), .B(keyinput_36), .ZN(n6106) );
  XNOR2_X1 U6916 ( .A(keyinput_37), .B(READREQUEST_REG_SCAN_IN), .ZN(n6105) );
  OAI21_X1 U6917 ( .B1(n6107), .B2(n6106), .A(n6105), .ZN(n6110) );
  XOR2_X1 U6918 ( .A(ADS_N_REG_SCAN_IN), .B(keyinput_38), .Z(n6109) );
  XOR2_X1 U6919 ( .A(CODEFETCH_REG_SCAN_IN), .B(keyinput_39), .Z(n6108) );
  NAND3_X1 U6920 ( .A1(n6110), .A2(n6109), .A3(n6108), .ZN(n6114) );
  XNOR2_X1 U6921 ( .A(keyinput_40), .B(M_IO_N_REG_SCAN_IN), .ZN(n6113) );
  XOR2_X1 U6922 ( .A(keyinput_41), .B(D_C_N_REG_SCAN_IN), .Z(n6112) );
  XNOR2_X1 U6923 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(keyinput_42), .ZN(n6111)
         );
  AOI211_X1 U6924 ( .C1(n6114), .C2(n6113), .A(n6112), .B(n6111), .ZN(n6117)
         );
  XNOR2_X1 U6925 ( .A(STATEBS16_REG_SCAN_IN), .B(keyinput_43), .ZN(n6116) );
  XNOR2_X1 U6926 ( .A(keyinput_44), .B(MORE_REG_SCAN_IN), .ZN(n6115) );
  NOR3_X1 U6927 ( .A1(n6117), .A2(n6116), .A3(n6115), .ZN(n6121) );
  XOR2_X1 U6928 ( .A(keyinput_45), .B(FLUSH_REG_SCAN_IN), .Z(n6120) );
  XOR2_X1 U6929 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_47), .Z(n6119) );
  XNOR2_X1 U6930 ( .A(keyinput_46), .B(W_R_N_REG_SCAN_IN), .ZN(n6118) );
  OAI211_X1 U6931 ( .C1(n6121), .C2(n6120), .A(n6119), .B(n6118), .ZN(n6124)
         );
  XNOR2_X1 U6932 ( .A(keyinput_48), .B(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6123)
         );
  XOR2_X1 U6933 ( .A(keyinput_49), .B(BYTEENABLE_REG_2__SCAN_IN), .Z(n6122) );
  AOI21_X1 U6934 ( .B1(n6124), .B2(n6123), .A(n6122), .ZN(n6131) );
  XOR2_X1 U6935 ( .A(REIP_REG_30__SCAN_IN), .B(keyinput_52), .Z(n6128) );
  XOR2_X1 U6936 ( .A(REIP_REG_29__SCAN_IN), .B(keyinput_53), .Z(n6127) );
  XOR2_X1 U6937 ( .A(REIP_REG_31__SCAN_IN), .B(keyinput_51), .Z(n6126) );
  XNOR2_X1 U6938 ( .A(keyinput_50), .B(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6125)
         );
  NAND4_X1 U6939 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n6130)
         );
  XNOR2_X1 U6940 ( .A(REIP_REG_28__SCAN_IN), .B(keyinput_54), .ZN(n6129) );
  OAI21_X1 U6941 ( .B1(n6131), .B2(n6130), .A(n6129), .ZN(n6135) );
  XOR2_X1 U6942 ( .A(REIP_REG_27__SCAN_IN), .B(keyinput_55), .Z(n6134) );
  XOR2_X1 U6943 ( .A(keyinput_57), .B(REIP_REG_25__SCAN_IN), .Z(n6133) );
  XNOR2_X1 U6944 ( .A(REIP_REG_26__SCAN_IN), .B(keyinput_56), .ZN(n6132) );
  NAND4_X1 U6945 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n6138)
         );
  XNOR2_X1 U6946 ( .A(REIP_REG_24__SCAN_IN), .B(keyinput_58), .ZN(n6137) );
  XNOR2_X1 U6947 ( .A(keyinput_59), .B(REIP_REG_23__SCAN_IN), .ZN(n6136) );
  AOI21_X1 U6948 ( .B1(n6138), .B2(n6137), .A(n6136), .ZN(n6141) );
  XOR2_X1 U6949 ( .A(keyinput_60), .B(REIP_REG_22__SCAN_IN), .Z(n6140) );
  XOR2_X1 U6950 ( .A(keyinput_61), .B(REIP_REG_21__SCAN_IN), .Z(n6139) );
  OAI21_X1 U6951 ( .B1(n6141), .B2(n6140), .A(n6139), .ZN(n6145) );
  XNOR2_X1 U6952 ( .A(keyinput_63), .B(REIP_REG_19__SCAN_IN), .ZN(n6144) );
  XNOR2_X1 U6953 ( .A(keyinput_62), .B(REIP_REG_20__SCAN_IN), .ZN(n6143) );
  XNOR2_X1 U6954 ( .A(keyinput_64), .B(REIP_REG_18__SCAN_IN), .ZN(n6142) );
  NAND4_X1 U6955 ( .A1(n6145), .A2(n6144), .A3(n6143), .A4(n6142), .ZN(n6155)
         );
  XOR2_X1 U6956 ( .A(keyinput_65), .B(REIP_REG_17__SCAN_IN), .Z(n6149) );
  XNOR2_X1 U6957 ( .A(BE_N_REG_2__SCAN_IN), .B(keyinput_68), .ZN(n6148) );
  XNOR2_X1 U6958 ( .A(keyinput_66), .B(REIP_REG_16__SCAN_IN), .ZN(n6147) );
  XNOR2_X1 U6959 ( .A(BE_N_REG_3__SCAN_IN), .B(keyinput_67), .ZN(n6146) );
  NOR4_X1 U6960 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n6154)
         );
  XOR2_X1 U6961 ( .A(BE_N_REG_0__SCAN_IN), .B(keyinput_70), .Z(n6152) );
  XOR2_X1 U6962 ( .A(BE_N_REG_1__SCAN_IN), .B(keyinput_69), .Z(n6151) );
  XOR2_X1 U6963 ( .A(ADDRESS_REG_29__SCAN_IN), .B(keyinput_71), .Z(n6150) );
  NAND3_X1 U6964 ( .A1(n6152), .A2(n6151), .A3(n6150), .ZN(n6153) );
  AOI21_X1 U6965 ( .B1(n6155), .B2(n6154), .A(n6153), .ZN(n6161) );
  XOR2_X1 U6966 ( .A(keyinput_72), .B(ADDRESS_REG_28__SCAN_IN), .Z(n6160) );
  INV_X1 U6967 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6875) );
  XNOR2_X1 U6968 ( .A(n6875), .B(keyinput_73), .ZN(n6158) );
  INV_X1 U6969 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6871) );
  XNOR2_X1 U6970 ( .A(n6871), .B(keyinput_75), .ZN(n6157) );
  XNOR2_X1 U6971 ( .A(ADDRESS_REG_26__SCAN_IN), .B(keyinput_74), .ZN(n6156) );
  NOR3_X1 U6972 ( .A1(n6158), .A2(n6157), .A3(n6156), .ZN(n6159) );
  OAI21_X1 U6973 ( .B1(n6161), .B2(n6160), .A(n6159), .ZN(n6169) );
  INV_X1 U6974 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6865) );
  XNOR2_X1 U6975 ( .A(n6865), .B(keyinput_79), .ZN(n6165) );
  INV_X1 U6976 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6869) );
  XNOR2_X1 U6977 ( .A(n6869), .B(keyinput_77), .ZN(n6164) );
  XNOR2_X1 U6978 ( .A(ADDRESS_REG_24__SCAN_IN), .B(keyinput_76), .ZN(n6163) );
  XNOR2_X1 U6979 ( .A(ADDRESS_REG_22__SCAN_IN), .B(keyinput_78), .ZN(n6162) );
  NOR4_X1 U6980 ( .A1(n6165), .A2(n6164), .A3(n6163), .A4(n6162), .ZN(n6168)
         );
  XOR2_X1 U6981 ( .A(keyinput_81), .B(ADDRESS_REG_19__SCAN_IN), .Z(n6167) );
  XNOR2_X1 U6982 ( .A(ADDRESS_REG_20__SCAN_IN), .B(keyinput_80), .ZN(n6166) );
  AOI211_X1 U6983 ( .C1(n6169), .C2(n6168), .A(n6167), .B(n6166), .ZN(n6173)
         );
  INV_X1 U6984 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6861) );
  XNOR2_X1 U6985 ( .A(n6861), .B(keyinput_82), .ZN(n6172) );
  XOR2_X1 U6986 ( .A(ADDRESS_REG_16__SCAN_IN), .B(keyinput_84), .Z(n6171) );
  XNOR2_X1 U6987 ( .A(keyinput_83), .B(ADDRESS_REG_17__SCAN_IN), .ZN(n6170) );
  OAI211_X1 U6988 ( .C1(n6173), .C2(n6172), .A(n6171), .B(n6170), .ZN(n6177)
         );
  XOR2_X1 U6989 ( .A(ADDRESS_REG_13__SCAN_IN), .B(keyinput_87), .Z(n6176) );
  XNOR2_X1 U6990 ( .A(keyinput_85), .B(ADDRESS_REG_15__SCAN_IN), .ZN(n6175) );
  XNOR2_X1 U6991 ( .A(keyinput_86), .B(ADDRESS_REG_14__SCAN_IN), .ZN(n6174) );
  NAND4_X1 U6992 ( .A1(n6177), .A2(n6176), .A3(n6175), .A4(n6174), .ZN(n6180)
         );
  XNOR2_X1 U6993 ( .A(keyinput_88), .B(ADDRESS_REG_12__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U6994 ( .A(keyinput_89), .B(ADDRESS_REG_11__SCAN_IN), .ZN(n6178) );
  AOI21_X1 U6995 ( .B1(n6180), .B2(n6179), .A(n6178), .ZN(n6188) );
  XNOR2_X1 U6996 ( .A(ADDRESS_REG_10__SCAN_IN), .B(keyinput_90), .ZN(n6187) );
  XNOR2_X1 U6997 ( .A(ADDRESS_REG_7__SCAN_IN), .B(keyinput_93), .ZN(n6186) );
  XOR2_X1 U6998 ( .A(ADDRESS_REG_5__SCAN_IN), .B(keyinput_95), .Z(n6184) );
  XOR2_X1 U6999 ( .A(ADDRESS_REG_6__SCAN_IN), .B(keyinput_94), .Z(n6183) );
  XOR2_X1 U7000 ( .A(ADDRESS_REG_8__SCAN_IN), .B(keyinput_92), .Z(n6182) );
  XNOR2_X1 U7001 ( .A(keyinput_91), .B(ADDRESS_REG_9__SCAN_IN), .ZN(n6181) );
  NAND4_X1 U7002 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n6185)
         );
  NOR4_X1 U7003 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .ZN(n6191)
         );
  XNOR2_X1 U7004 ( .A(keyinput_96), .B(ADDRESS_REG_4__SCAN_IN), .ZN(n6190) );
  XOR2_X1 U7005 ( .A(keyinput_97), .B(ADDRESS_REG_3__SCAN_IN), .Z(n6189) );
  OAI21_X1 U7006 ( .B1(n6191), .B2(n6190), .A(n6189), .ZN(n6195) );
  XNOR2_X1 U7007 ( .A(keyinput_100), .B(ADDRESS_REG_0__SCAN_IN), .ZN(n6194) );
  XNOR2_X1 U7008 ( .A(keyinput_98), .B(ADDRESS_REG_2__SCAN_IN), .ZN(n6193) );
  XNOR2_X1 U7009 ( .A(keyinput_99), .B(ADDRESS_REG_1__SCAN_IN), .ZN(n6192) );
  NAND4_X1 U7010 ( .A1(n6195), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n6198)
         );
  XOR2_X1 U7011 ( .A(STATE_REG_1__SCAN_IN), .B(keyinput_102), .Z(n6197) );
  XOR2_X1 U7012 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput_101), .Z(n6196) );
  NAND3_X1 U7013 ( .A1(n6198), .A2(n6197), .A3(n6196), .ZN(n6202) );
  XOR2_X1 U7014 ( .A(DATAWIDTH_REG_1__SCAN_IN), .B(keyinput_105), .Z(n6201) );
  XNOR2_X1 U7015 ( .A(keyinput_103), .B(STATE_REG_0__SCAN_IN), .ZN(n6200) );
  XNOR2_X1 U7016 ( .A(keyinput_104), .B(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6199)
         );
  NAND4_X1 U7017 ( .A1(n6202), .A2(n6201), .A3(n6200), .A4(n6199), .ZN(n6205)
         );
  XOR2_X1 U7018 ( .A(DATAWIDTH_REG_3__SCAN_IN), .B(keyinput_107), .Z(n6204) );
  XNOR2_X1 U7019 ( .A(keyinput_106), .B(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6203)
         );
  NAND3_X1 U7020 ( .A1(n6205), .A2(n6204), .A3(n6203), .ZN(n6208) );
  XOR2_X1 U7021 ( .A(DATAWIDTH_REG_5__SCAN_IN), .B(keyinput_109), .Z(n6207) );
  XNOR2_X1 U7022 ( .A(keyinput_108), .B(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6206)
         );
  NAND3_X1 U7023 ( .A1(n6208), .A2(n6207), .A3(n6206), .ZN(n6211) );
  XOR2_X1 U7024 ( .A(DATAWIDTH_REG_6__SCAN_IN), .B(keyinput_110), .Z(n6210) );
  XNOR2_X1 U7025 ( .A(keyinput_111), .B(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6209)
         );
  NAND3_X1 U7026 ( .A1(n6211), .A2(n6210), .A3(n6209), .ZN(n6219) );
  XOR2_X1 U7027 ( .A(DATAWIDTH_REG_10__SCAN_IN), .B(keyinput_114), .Z(n6218)
         );
  XOR2_X1 U7028 ( .A(DATAWIDTH_REG_8__SCAN_IN), .B(keyinput_112), .Z(n6217) );
  XOR2_X1 U7029 ( .A(keyinput_116), .B(DATAWIDTH_REG_12__SCAN_IN), .Z(n6215)
         );
  XOR2_X1 U7030 ( .A(keyinput_113), .B(DATAWIDTH_REG_9__SCAN_IN), .Z(n6214) );
  INV_X1 U7031 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6788) );
  XNOR2_X1 U7032 ( .A(n6788), .B(keyinput_117), .ZN(n6213) );
  INV_X1 U7033 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6786) );
  XNOR2_X1 U7034 ( .A(n6786), .B(keyinput_115), .ZN(n6212) );
  NOR4_X1 U7035 ( .A1(n6215), .A2(n6214), .A3(n6213), .A4(n6212), .ZN(n6216)
         );
  NAND4_X1 U7036 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n6222)
         );
  XOR2_X1 U7037 ( .A(DATAWIDTH_REG_14__SCAN_IN), .B(keyinput_118), .Z(n6221)
         );
  XNOR2_X1 U7038 ( .A(keyinput_119), .B(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6220)
         );
  NAND3_X1 U7039 ( .A1(n6222), .A2(n6221), .A3(n6220), .ZN(n6226) );
  XNOR2_X1 U7040 ( .A(keyinput_120), .B(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6225)
         );
  INV_X1 U7041 ( .A(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6791) );
  XNOR2_X1 U7042 ( .A(n6791), .B(keyinput_122), .ZN(n6224) );
  XNOR2_X1 U7043 ( .A(DATAWIDTH_REG_17__SCAN_IN), .B(keyinput_121), .ZN(n6223)
         );
  AOI211_X1 U7044 ( .C1(n6226), .C2(n6225), .A(n6224), .B(n6223), .ZN(n6229)
         );
  INV_X1 U7045 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6792) );
  XNOR2_X1 U7046 ( .A(n6792), .B(keyinput_123), .ZN(n6228) );
  XNOR2_X1 U7047 ( .A(DATAWIDTH_REG_20__SCAN_IN), .B(keyinput_124), .ZN(n6227)
         );
  NOR3_X1 U7048 ( .A1(n6229), .A2(n6228), .A3(n6227), .ZN(n6232) );
  XOR2_X1 U7049 ( .A(keyinput_126), .B(DATAWIDTH_REG_22__SCAN_IN), .Z(n6231)
         );
  XNOR2_X1 U7050 ( .A(DATAWIDTH_REG_21__SCAN_IN), .B(keyinput_125), .ZN(n6230)
         );
  NOR3_X1 U7051 ( .A1(n6232), .A2(n6231), .A3(n6230), .ZN(n6233) );
  OR2_X1 U7052 ( .A1(n6988), .A2(STATE_REG_0__SCAN_IN), .ZN(n7421) );
  AOI21_X1 U7053 ( .B1(n6832), .B2(STATE_REG_1__SCAN_IN), .A(n7415), .ZN(n6798) );
  INV_X1 U7054 ( .A(n6798), .ZN(n6237) );
  NAND2_X1 U7055 ( .A1(n7421), .A2(n6237), .ZN(n7404) );
  NAND2_X1 U7056 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n7404), .ZN(n6238) );
  XNOR2_X1 U7057 ( .A(n6239), .B(n6238), .ZN(U3178) );
  INV_X1 U7058 ( .A(n6240), .ZN(n6246) );
  INV_X1 U7059 ( .A(n6241), .ZN(n6244) );
  NAND3_X1 U7060 ( .A1(n4989), .A2(n6721), .A3(n6248), .ZN(n6242) );
  OAI21_X1 U7061 ( .B1(n6244), .B2(n6243), .A(n6242), .ZN(n6245) );
  AOI21_X1 U7062 ( .B1(n6246), .B2(n7383), .A(n6245), .ZN(n6251) );
  INV_X1 U7063 ( .A(n4989), .ZN(n6247) );
  AOI21_X1 U7064 ( .B1(n6247), .B2(n6721), .A(n6250), .ZN(n6249) );
  OAI22_X1 U7065 ( .A1(n6251), .A2(n6250), .B1(n6249), .B2(n6248), .ZN(U3459)
         );
  AND2_X1 U7066 ( .A1(n6252), .A2(n6260), .ZN(n6253) );
  OR2_X1 U7067 ( .A1(n6255), .A2(n6253), .ZN(n6257) );
  NAND2_X1 U7068 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  OAI211_X1 U7069 ( .C1(n6258), .C2(n4760), .A(n6257), .B(n6256), .ZN(n7368)
         );
  NAND2_X1 U7070 ( .A1(n3920), .A2(n6258), .ZN(n6259) );
  AOI22_X1 U7071 ( .A1(n6262), .A2(n6261), .B1(n6260), .B2(n6259), .ZN(n6976)
         );
  NOR2_X1 U7072 ( .A1(n3921), .A2(n6263), .ZN(n6985) );
  INV_X1 U7073 ( .A(n6985), .ZN(n6265) );
  OAI21_X1 U7074 ( .B1(n6265), .B2(n6264), .A(n7414), .ZN(n6994) );
  NAND2_X1 U7075 ( .A1(n6976), .A2(n6994), .ZN(n7375) );
  INV_X1 U7076 ( .A(n7375), .ZN(n6266) );
  NOR2_X1 U7077 ( .A1(n6266), .A2(n7377), .ZN(n7346) );
  MUX2_X1 U7078 ( .A(MORE_REG_SCAN_IN), .B(n7368), .S(n7346), .Z(U3471) );
  OAI22_X1 U7079 ( .A1(n6268), .A2(n5672), .B1(n6267), .B2(n6294), .ZN(n6269)
         );
  XOR2_X1 U7080 ( .A(n6270), .B(n6269), .Z(n6595) );
  NAND2_X1 U7081 ( .A1(n6490), .A2(n7338), .ZN(n6280) );
  INV_X1 U7082 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6389) );
  INV_X1 U7083 ( .A(n6488), .ZN(n6274) );
  AOI22_X1 U7084 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n7335), .B1(n7339), 
        .B2(n6274), .ZN(n6275) );
  OAI21_X1 U7085 ( .B1(n7312), .B2(n6389), .A(n6275), .ZN(n6277) );
  NOR3_X1 U7086 ( .A1(n6282), .A2(REIP_REG_30__SCAN_IN), .A3(n6877), .ZN(n6276) );
  AOI211_X1 U7087 ( .C1(REIP_REG_30__SCAN_IN), .C2(n6278), .A(n6277), .B(n6276), .ZN(n6279) );
  OAI211_X1 U7088 ( .C1(n6595), .C2(n7329), .A(n6280), .B(n6279), .ZN(U2797)
         );
  INV_X1 U7089 ( .A(n6390), .ZN(n6287) );
  MUX2_X1 U7090 ( .A(n6282), .B(n6301), .S(REIP_REG_29__SCAN_IN), .Z(n6285) );
  AOI22_X1 U7091 ( .A1(n6283), .A2(n7339), .B1(n7335), .B2(
        PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6284) );
  OAI211_X1 U7092 ( .C1(n6391), .C2(n7312), .A(n6285), .B(n6284), .ZN(n6286)
         );
  AOI21_X1 U7093 ( .B1(n6287), .B2(n7337), .A(n6286), .ZN(n6288) );
  OAI21_X1 U7094 ( .B1(n6281), .B2(n7325), .A(n6288), .ZN(U2798) );
  INV_X1 U7095 ( .A(n6289), .ZN(n6293) );
  INV_X1 U7096 ( .A(n6290), .ZN(n6292) );
  AOI21_X1 U7097 ( .B1(n6293), .B2(n6292), .A(n3657), .ZN(n6498) );
  INV_X1 U7098 ( .A(n6498), .ZN(n6393) );
  INV_X1 U7099 ( .A(n6294), .ZN(n6295) );
  AOI21_X1 U7100 ( .B1(n6296), .B2(n6309), .A(n6295), .ZN(n6609) );
  OAI22_X1 U7101 ( .A1(n6297), .A2(n7294), .B1(n7323), .B2(n6496), .ZN(n6298)
         );
  AOI21_X1 U7102 ( .B1(n7332), .B2(EBX_REG_28__SCAN_IN), .A(n6298), .ZN(n6300)
         );
  NAND3_X1 U7103 ( .A1(n6311), .A2(REIP_REG_27__SCAN_IN), .A3(n6876), .ZN(
        n6299) );
  OAI211_X1 U7104 ( .C1(n6301), .C2(n6876), .A(n6300), .B(n6299), .ZN(n6302)
         );
  AOI21_X1 U7105 ( .B1(n6609), .B2(n7337), .A(n6302), .ZN(n6303) );
  OAI21_X1 U7106 ( .B1(n6393), .B2(n7325), .A(n6303), .ZN(U2799) );
  AND2_X1 U7107 ( .A1(n6304), .A2(n6305), .ZN(n6306) );
  OR2_X1 U7108 ( .A1(n6330), .A2(n6307), .ZN(n6308) );
  NAND2_X1 U7109 ( .A1(n6309), .A2(n6308), .ZN(n6917) );
  INV_X1 U7110 ( .A(n6917), .ZN(n6317) );
  INV_X1 U7111 ( .A(n7266), .ZN(n7186) );
  NOR3_X1 U7112 ( .A1(n7186), .A2(n6310), .A3(n6874), .ZN(n6316) );
  INV_X1 U7113 ( .A(n6311), .ZN(n6314) );
  OAI22_X1 U7114 ( .A1(n6503), .A2(n7294), .B1(n6920), .B2(n7312), .ZN(n6312)
         );
  AOI21_X1 U7115 ( .B1(n7339), .B2(n6506), .A(n6312), .ZN(n6313) );
  OAI21_X1 U7116 ( .B1(n6314), .B2(REIP_REG_27__SCAN_IN), .A(n6313), .ZN(n6315) );
  AOI211_X1 U7117 ( .C1(n6317), .C2(n7337), .A(n6316), .B(n6315), .ZN(n6318)
         );
  OAI21_X1 U7118 ( .B1(n7582), .B2(n7325), .A(n6318), .ZN(U2800) );
  NAND2_X1 U7119 ( .A1(n6319), .A2(n6320), .ZN(n6335) );
  INV_X1 U7120 ( .A(n6304), .ZN(n6321) );
  AOI21_X1 U7121 ( .B1(n6322), .B2(n6335), .A(n6321), .ZN(n6513) );
  INV_X1 U7122 ( .A(n6513), .ZN(n6468) );
  INV_X1 U7123 ( .A(n6509), .ZN(n6323) );
  OAI22_X1 U7124 ( .A1(n6511), .A2(n7294), .B1(n7323), .B2(n6323), .ZN(n6329)
         );
  INV_X1 U7125 ( .A(n6324), .ZN(n6327) );
  AOI21_X1 U7126 ( .B1(n7151), .B2(n6325), .A(REIP_REG_26__SCAN_IN), .ZN(n6326) );
  AOI211_X1 U7127 ( .C1(REIP_REG_26__SCAN_IN), .C2(n6327), .A(n7186), .B(n6326), .ZN(n6328) );
  AOI211_X1 U7128 ( .C1(n7332), .C2(EBX_REG_26__SCAN_IN), .A(n6329), .B(n6328), 
        .ZN(n6332) );
  AOI21_X1 U7129 ( .B1(n3690), .B2(n3696), .A(n6330), .ZN(n6625) );
  NAND2_X1 U7130 ( .A1(n6625), .A2(n7337), .ZN(n6331) );
  OAI211_X1 U7131 ( .C1(n6468), .C2(n7325), .A(n6332), .B(n6331), .ZN(U2801)
         );
  AND2_X1 U7132 ( .A1(n6319), .A2(n6365), .ZN(n6334) );
  INV_X1 U7133 ( .A(n6632), .ZN(n6355) );
  AOI21_X1 U7134 ( .B1(n6355), .B2(n6631), .A(n6337), .ZN(n6339) );
  NOR2_X1 U7135 ( .A1(n6339), .A2(n6338), .ZN(n7131) );
  INV_X1 U7136 ( .A(n7334), .ZN(n6340) );
  NAND2_X1 U7137 ( .A1(n7151), .A2(n6340), .ZN(n6341) );
  AND2_X1 U7138 ( .A1(n6341), .A2(n6366), .ZN(n6361) );
  INV_X1 U7139 ( .A(n6361), .ZN(n7331) );
  NOR2_X1 U7140 ( .A1(n7316), .A2(REIP_REG_24__SCAN_IN), .ZN(n7333) );
  NOR2_X1 U7141 ( .A1(n7331), .A2(n7333), .ZN(n6342) );
  OAI22_X1 U7142 ( .A1(n6342), .A2(n7135), .B1(n6517), .B2(n7294), .ZN(n6348)
         );
  INV_X1 U7143 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6346) );
  NOR3_X1 U7144 ( .A1(n7316), .A2(REIP_REG_25__SCAN_IN), .A3(n6343), .ZN(n6344) );
  AOI21_X1 U7145 ( .B1(n7339), .B2(n6521), .A(n6344), .ZN(n6345) );
  OAI21_X1 U7146 ( .B1(n7312), .B2(n6346), .A(n6345), .ZN(n6347) );
  AOI211_X1 U7147 ( .C1(n7131), .C2(n7337), .A(n6348), .B(n6347), .ZN(n6349)
         );
  OAI21_X1 U7148 ( .B1(n6518), .B2(n7325), .A(n6349), .ZN(U2802) );
  AOI21_X1 U7149 ( .B1(n6356), .B2(n6354), .A(n6355), .ZN(n6640) );
  INV_X1 U7150 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6358) );
  INV_X1 U7151 ( .A(n6542), .ZN(n6357) );
  OAI22_X1 U7152 ( .A1(n7312), .A2(n6358), .B1(n6357), .B2(n7323), .ZN(n6363)
         );
  NOR2_X1 U7153 ( .A1(n7316), .A2(n6359), .ZN(n7321) );
  AOI21_X1 U7154 ( .B1(REIP_REG_22__SCAN_IN), .B2(n7321), .A(
        REIP_REG_23__SCAN_IN), .ZN(n6360) );
  OAI22_X1 U7155 ( .A1(n6361), .A2(n6360), .B1(n6544), .B2(n7294), .ZN(n6362)
         );
  AOI211_X1 U7156 ( .C1(n6640), .C2(n7337), .A(n6363), .B(n6362), .ZN(n6364)
         );
  OAI21_X1 U7157 ( .B1(n6473), .B2(n7325), .A(n6364), .ZN(U2804) );
  OAI21_X1 U7158 ( .B1(n6319), .B2(n6365), .A(n6398), .ZN(n6564) );
  OAI21_X1 U7159 ( .B1(n7316), .B2(n6370), .A(n6366), .ZN(n7314) );
  NOR2_X1 U7160 ( .A1(n3629), .A2(n6367), .ZN(n6368) );
  OR2_X1 U7161 ( .A1(n6402), .A2(n6368), .ZN(n6659) );
  OAI22_X1 U7162 ( .A1(n6559), .A2(n7294), .B1(n6407), .B2(n7312), .ZN(n6369)
         );
  AOI21_X1 U7163 ( .B1(n7339), .B2(n6561), .A(n6369), .ZN(n6372) );
  NAND3_X1 U7164 ( .A1(n7151), .A2(n6370), .A3(n6864), .ZN(n6371) );
  OAI211_X1 U7165 ( .C1(n6659), .C2(n7329), .A(n6372), .B(n6371), .ZN(n6373)
         );
  AOI21_X1 U7166 ( .B1(REIP_REG_21__SCAN_IN), .B2(n7314), .A(n6373), .ZN(n6374) );
  OAI21_X1 U7167 ( .B1(n6564), .B2(n7325), .A(n6374), .ZN(U2806) );
  OAI21_X1 U7168 ( .B1(n6378), .B2(n4277), .A(n6377), .ZN(n6589) );
  INV_X1 U7169 ( .A(n6585), .ZN(n6387) );
  NAND2_X1 U7170 ( .A1(n6382), .A2(n7218), .ZN(n7256) );
  AOI22_X1 U7171 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n7335), .B1(
        EBX_REG_15__SCAN_IN), .B2(n7332), .ZN(n6379) );
  OAI211_X1 U7172 ( .C1(REIP_REG_15__SCAN_IN), .C2(n7256), .A(n6379), .B(n7291), .ZN(n6386) );
  NAND2_X1 U7173 ( .A1(n5721), .A2(n6380), .ZN(n6381) );
  NAND2_X1 U7174 ( .A1(n6445), .A2(n6381), .ZN(n7111) );
  INV_X1 U7175 ( .A(REIP_REG_15__SCAN_IN), .ZN(n7257) );
  INV_X1 U7176 ( .A(n6382), .ZN(n6384) );
  OAI21_X1 U7177 ( .B1(n6384), .B2(n6383), .A(n7266), .ZN(n7253) );
  OAI22_X1 U7178 ( .A1(n7329), .A2(n7111), .B1(n7257), .B2(n7253), .ZN(n6385)
         );
  AOI211_X1 U7179 ( .C1(n7339), .C2(n6387), .A(n6386), .B(n6385), .ZN(n6388)
         );
  OAI21_X1 U7180 ( .B1(n6589), .B2(n7325), .A(n6388), .ZN(U2812) );
  INV_X1 U7181 ( .A(n6490), .ZN(n6459) );
  OAI222_X1 U7182 ( .A1(n6459), .A2(n6454), .B1(n6389), .B2(n6927), .C1(n6916), 
        .C2(n6595), .ZN(U2829) );
  AOI22_X1 U7183 ( .A1(n6609), .A2(n6924), .B1(EBX_REG_28__SCAN_IN), .B2(n6426), .ZN(n6392) );
  OAI21_X1 U7184 ( .B1(n6393), .B2(n6454), .A(n6392), .ZN(U2831) );
  AOI22_X1 U7185 ( .A1(n6625), .A2(n6924), .B1(EBX_REG_26__SCAN_IN), .B2(n6426), .ZN(n6394) );
  OAI21_X1 U7186 ( .B1(n6468), .B2(n6454), .A(n6394), .ZN(U2833) );
  AOI22_X1 U7187 ( .A1(n7131), .A2(n6924), .B1(EBX_REG_25__SCAN_IN), .B2(n6426), .ZN(n6395) );
  OAI21_X1 U7188 ( .B1(n6518), .B2(n6454), .A(n6395), .ZN(U2834) );
  AOI22_X1 U7189 ( .A1(n6640), .A2(n6924), .B1(EBX_REG_23__SCAN_IN), .B2(n6426), .ZN(n6396) );
  OAI21_X1 U7190 ( .B1(n6473), .B2(n6454), .A(n6396), .ZN(U2836) );
  NAND2_X1 U7191 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  OR2_X1 U7192 ( .A1(n6402), .A2(n6401), .ZN(n6403) );
  NAND2_X1 U7193 ( .A1(n6354), .A2(n6403), .ZN(n7330) );
  OAI22_X1 U7194 ( .A1(n7330), .A2(n6916), .B1(n6404), .B2(n6927), .ZN(n6405)
         );
  INV_X1 U7195 ( .A(n6405), .ZN(n6406) );
  OAI21_X1 U7196 ( .B1(n7442), .B2(n6454), .A(n6406), .ZN(U2837) );
  OAI22_X1 U7197 ( .A1(n6659), .A2(n6916), .B1(n6407), .B2(n6927), .ZN(n6408)
         );
  INV_X1 U7198 ( .A(n6408), .ZN(n6409) );
  OAI21_X1 U7199 ( .B1(n6564), .B2(n6454), .A(n6409), .ZN(U2838) );
  NOR2_X1 U7200 ( .A1(n6410), .A2(n6411), .ZN(n6412) );
  INV_X1 U7201 ( .A(n6454), .ZN(n6925) );
  AND2_X1 U7202 ( .A1(n6423), .A2(n6414), .ZN(n6416) );
  OR2_X1 U7203 ( .A1(n6416), .A2(n3629), .ZN(n7308) );
  OAI22_X1 U7204 ( .A1(n7308), .A2(n6916), .B1(n7313), .B2(n6927), .ZN(n6417)
         );
  AOI21_X1 U7205 ( .B1(n6413), .B2(n6925), .A(n6417), .ZN(n6418) );
  INV_X1 U7206 ( .A(n6418), .ZN(U2839) );
  INV_X1 U7207 ( .A(n6410), .ZN(n6420) );
  OAI21_X1 U7208 ( .B1(n6421), .B2(n6419), .A(n6420), .ZN(n7297) );
  INV_X1 U7209 ( .A(n6423), .ZN(n6424) );
  AOI21_X1 U7210 ( .B1(n6425), .B2(n6422), .A(n6424), .ZN(n7295) );
  AOI22_X1 U7211 ( .A1(n7295), .A2(n6924), .B1(EBX_REG_19__SCAN_IN), .B2(n6426), .ZN(n6427) );
  OAI21_X1 U7212 ( .B1(n7297), .B2(n6454), .A(n6427), .ZN(U2840) );
  AND2_X1 U7213 ( .A1(n6428), .A2(n6429), .ZN(n6430) );
  OR2_X1 U7214 ( .A1(n6430), .A2(n6419), .ZN(n7435) );
  OR2_X1 U7215 ( .A1(n6440), .A2(n6431), .ZN(n6432) );
  NAND2_X1 U7216 ( .A1(n6422), .A2(n6432), .ZN(n7284) );
  OAI22_X1 U7217 ( .A1(n7284), .A2(n6916), .B1(n7277), .B2(n6927), .ZN(n6433)
         );
  AOI21_X1 U7218 ( .B1(n7286), .B2(n6925), .A(n6433), .ZN(n6434) );
  INV_X1 U7219 ( .A(n6434), .ZN(U2841) );
  NAND2_X1 U7220 ( .A1(n6435), .A2(n6436), .ZN(n6437) );
  NAND2_X1 U7221 ( .A1(n6428), .A2(n6437), .ZN(n7430) );
  INV_X1 U7222 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6441) );
  AND2_X1 U7223 ( .A1(n6447), .A2(n6438), .ZN(n6439) );
  NOR2_X1 U7224 ( .A1(n6440), .A2(n6439), .ZN(n7121) );
  INV_X1 U7225 ( .A(n7121), .ZN(n7272) );
  OAI222_X1 U7226 ( .A1(n7430), .A2(n6454), .B1(n6441), .B2(n6927), .C1(n7272), 
        .C2(n6916), .ZN(U2842) );
  NAND2_X1 U7227 ( .A1(n6377), .A2(n6442), .ZN(n6443) );
  NAND2_X1 U7228 ( .A1(n6435), .A2(n6443), .ZN(n7426) );
  INV_X1 U7229 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U7230 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  NAND2_X1 U7231 ( .A1(n6447), .A2(n6446), .ZN(n7265) );
  OAI222_X1 U7232 ( .A1(n7426), .A2(n6454), .B1(n6448), .B2(n6927), .C1(n6916), 
        .C2(n7265), .ZN(U2843) );
  INV_X1 U7233 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6449) );
  OAI222_X1 U7234 ( .A1(n6589), .A2(n6454), .B1(n6449), .B2(n6927), .C1(n6916), 
        .C2(n7111), .ZN(U2844) );
  OR2_X1 U7235 ( .A1(n6451), .A2(n6450), .ZN(n6452) );
  AND2_X1 U7236 ( .A1(n6375), .A2(n6452), .ZN(n7249) );
  INV_X1 U7237 ( .A(n7249), .ZN(n6482) );
  INV_X1 U7238 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6453) );
  OAI222_X1 U7239 ( .A1(n6482), .A2(n6454), .B1(n6453), .B2(n6927), .C1(n6916), 
        .C2(n7245), .ZN(U2845) );
  AOI22_X1 U7240 ( .A1(n7520), .A2(DATAI_14_), .B1(n7584), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U7241 ( .A1(n7585), .A2(DATAI_30_), .ZN(n6457) );
  OAI211_X1 U7242 ( .C1(n6459), .C2(n7581), .A(n6458), .B(n6457), .ZN(U2861)
         );
  AOI22_X1 U7243 ( .A1(n7520), .A2(DATAI_13_), .B1(n7584), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U7244 ( .A1(n7585), .A2(DATAI_29_), .ZN(n6460) );
  OAI211_X1 U7245 ( .C1(n6281), .C2(n7581), .A(n6461), .B(n6460), .ZN(U2862)
         );
  INV_X1 U7246 ( .A(n7585), .ZN(n6465) );
  NAND2_X1 U7247 ( .A1(n6498), .A2(n7521), .ZN(n6463) );
  AOI22_X1 U7248 ( .A1(n7520), .A2(DATAI_12_), .B1(n7584), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6462) );
  OAI211_X1 U7249 ( .C1(n6465), .C2(n6464), .A(n6463), .B(n6462), .ZN(U2863)
         );
  AOI22_X1 U7250 ( .A1(n7520), .A2(DATAI_10_), .B1(n7584), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7251 ( .A1(n7585), .A2(DATAI_26_), .ZN(n6466) );
  OAI211_X1 U7252 ( .C1(n6468), .C2(n7581), .A(n6467), .B(n6466), .ZN(U2865)
         );
  AOI22_X1 U7253 ( .A1(n7520), .A2(DATAI_9_), .B1(n7584), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U7254 ( .A1(n7585), .A2(DATAI_25_), .ZN(n6469) );
  OAI211_X1 U7255 ( .C1(n6518), .C2(n7581), .A(n6470), .B(n6469), .ZN(U2866)
         );
  AOI22_X1 U7256 ( .A1(n7520), .A2(DATAI_7_), .B1(n7584), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U7257 ( .A1(n7585), .A2(DATAI_23_), .ZN(n6471) );
  OAI211_X1 U7258 ( .C1(n6473), .C2(n7581), .A(n6472), .B(n6471), .ZN(U2868)
         );
  AOI22_X1 U7259 ( .A1(n7520), .A2(DATAI_5_), .B1(n7584), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7260 ( .A1(n7585), .A2(DATAI_21_), .ZN(n6474) );
  OAI211_X1 U7261 ( .C1(n6564), .C2(n7581), .A(n6475), .B(n6474), .ZN(U2870)
         );
  AOI22_X1 U7262 ( .A1(n7520), .A2(DATAI_3_), .B1(n7584), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U7263 ( .A1(n7585), .A2(DATAI_19_), .ZN(n6476) );
  OAI211_X1 U7264 ( .C1(n7297), .C2(n7581), .A(n6477), .B(n6476), .ZN(U2872)
         );
  INV_X1 U7265 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6831) );
  OAI222_X1 U7266 ( .A1(n6478), .A2(n6481), .B1(n6479), .B2(n6831), .C1(n7581), 
        .C2(n6589), .ZN(U2876) );
  INV_X1 U7267 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6827) );
  OAI222_X1 U7268 ( .A1(n6482), .A2(n7581), .B1(n6481), .B2(n6480), .C1(n6479), 
        .C2(n6827), .ZN(U2877) );
  NAND2_X1 U7269 ( .A1(n6485), .A2(n6526), .ZN(n6484) );
  NAND2_X1 U7270 ( .A1(n7073), .A2(REIP_REG_30__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U7271 ( .A1(n6969), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6487)
         );
  OAI211_X1 U7272 ( .C1(n6975), .C2(n6488), .A(n6596), .B(n6487), .ZN(n6489)
         );
  AOI21_X1 U7273 ( .B1(n6490), .B2(n6970), .A(n6489), .ZN(n6491) );
  OAI21_X1 U7274 ( .B1(n6604), .B2(n7345), .A(n6491), .ZN(U2956) );
  AOI21_X1 U7275 ( .B1(n6494), .B2(n6492), .A(n6493), .ZN(n6614) );
  NAND2_X1 U7276 ( .A1(n7073), .A2(REIP_REG_28__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U7277 ( .A1(n6969), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6495)
         );
  OAI211_X1 U7278 ( .C1(n6975), .C2(n6496), .A(n6605), .B(n6495), .ZN(n6497)
         );
  AOI21_X1 U7279 ( .B1(n6498), .B2(n6970), .A(n6497), .ZN(n6499) );
  OAI21_X1 U7280 ( .B1(n6614), .B2(n7345), .A(n6499), .ZN(U2958) );
  NOR2_X1 U7281 ( .A1(n6668), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6501)
         );
  MUX2_X1 U7282 ( .A(n6501), .B(n6668), .S(n6500), .Z(n6502) );
  XNOR2_X1 U7283 ( .A(n6502), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6621)
         );
  NAND2_X1 U7284 ( .A1(n7073), .A2(REIP_REG_27__SCAN_IN), .ZN(n6615) );
  OAI21_X1 U7285 ( .B1(n6965), .B2(n6503), .A(n6615), .ZN(n6505) );
  NOR2_X1 U7286 ( .A1(n7582), .A2(n6962), .ZN(n6504) );
  AOI211_X1 U7287 ( .C1(n6941), .C2(n6506), .A(n6505), .B(n6504), .ZN(n6507)
         );
  OAI21_X1 U7288 ( .B1(n7345), .B2(n6621), .A(n6507), .ZN(U2959) );
  XNOR2_X1 U7289 ( .A(n6549), .B(n6623), .ZN(n6508) );
  XNOR2_X1 U7290 ( .A(n4745), .B(n6508), .ZN(n6630) );
  NAND2_X1 U7291 ( .A1(n6941), .A2(n6509), .ZN(n6510) );
  NAND2_X1 U7292 ( .A1(n7073), .A2(REIP_REG_26__SCAN_IN), .ZN(n6622) );
  OAI211_X1 U7293 ( .C1(n6965), .C2(n6511), .A(n6510), .B(n6622), .ZN(n6512)
         );
  AOI21_X1 U7294 ( .B1(n6513), .B2(n6970), .A(n6512), .ZN(n6514) );
  OAI21_X1 U7295 ( .B1(n7345), .B2(n6630), .A(n6514), .ZN(U2960) );
  XNOR2_X1 U7296 ( .A(n6526), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6516)
         );
  XNOR2_X1 U7297 ( .A(n6515), .B(n6516), .ZN(n7130) );
  OAI22_X1 U7298 ( .A1(n6965), .A2(n6517), .B1(n7135), .B2(n7136), .ZN(n6520)
         );
  NOR2_X1 U7299 ( .A1(n6518), .A2(n6962), .ZN(n6519) );
  AOI211_X1 U7300 ( .C1(n6941), .C2(n6521), .A(n6520), .B(n6519), .ZN(n6522)
         );
  OAI21_X1 U7301 ( .B1(n7345), .B2(n7130), .A(n6522), .ZN(U2961) );
  XNOR2_X1 U7302 ( .A(n6526), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6565)
         );
  OAI21_X1 U7303 ( .B1(n6668), .B2(n6667), .A(n6665), .ZN(n6524) );
  XNOR2_X1 U7304 ( .A(n6526), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6557)
         );
  NOR2_X1 U7305 ( .A1(n6558), .A2(n6557), .ZN(n6556) );
  NAND3_X1 U7306 ( .A1(n6668), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6527) );
  NAND4_X1 U7307 ( .A1(n6665), .A2(n6526), .A3(n6652), .A4(n6667), .ZN(n6538)
         );
  OAI22_X1 U7308 ( .A1(n6551), .A2(n6527), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6538), .ZN(n6528) );
  XNOR2_X1 U7309 ( .A(n6528), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6639)
         );
  AND2_X1 U7310 ( .A1(n7073), .A2(REIP_REG_24__SCAN_IN), .ZN(n6637) );
  INV_X1 U7311 ( .A(n6637), .ZN(n6529) );
  OAI21_X1 U7312 ( .B1(n6965), .B2(n6530), .A(n6529), .ZN(n6531) );
  AOI21_X1 U7313 ( .B1(n6941), .B2(n7340), .A(n6531), .ZN(n6537) );
  NOR2_X1 U7314 ( .A1(n6533), .A2(n6532), .ZN(n6534) );
  NOR2_X2 U7315 ( .A1(n6535), .A2(n6534), .ZN(n7522) );
  NAND2_X1 U7316 ( .A1(n7522), .A2(n6970), .ZN(n6536) );
  OAI211_X1 U7317 ( .C1(n6639), .C2(n7345), .A(n6537), .B(n6536), .ZN(U2962)
         );
  NAND2_X1 U7318 ( .A1(n6668), .A2(n3693), .ZN(n6539) );
  OAI21_X1 U7319 ( .B1(n6540), .B2(n6539), .A(n6538), .ZN(n6541) );
  XNOR2_X1 U7320 ( .A(n6541), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6648)
         );
  NAND2_X1 U7321 ( .A1(n6941), .A2(n6542), .ZN(n6543) );
  NAND2_X1 U7322 ( .A1(n7073), .A2(REIP_REG_23__SCAN_IN), .ZN(n6641) );
  OAI211_X1 U7323 ( .C1(n6965), .C2(n6544), .A(n6543), .B(n6641), .ZN(n6545)
         );
  AOI21_X1 U7324 ( .B1(n6546), .B2(n6970), .A(n6545), .ZN(n6547) );
  OAI21_X1 U7325 ( .B1(n6648), .B2(n7345), .A(n6547), .ZN(U2963) );
  XNOR2_X1 U7326 ( .A(n6549), .B(n6548), .ZN(n6550) );
  XNOR2_X1 U7327 ( .A(n6551), .B(n6550), .ZN(n6656) );
  NAND2_X1 U7328 ( .A1(n7073), .A2(REIP_REG_22__SCAN_IN), .ZN(n6649) );
  OAI21_X1 U7329 ( .B1(n6965), .B2(n6552), .A(n6649), .ZN(n6554) );
  NOR2_X1 U7330 ( .A1(n7442), .A2(n6962), .ZN(n6553) );
  NAND2_X1 U7331 ( .A1(n6558), .A2(n6557), .ZN(n6657) );
  NAND3_X1 U7332 ( .A1(n3655), .A2(n6971), .A3(n6657), .ZN(n6563) );
  NAND2_X1 U7333 ( .A1(n7073), .A2(REIP_REG_21__SCAN_IN), .ZN(n6658) );
  OAI21_X1 U7334 ( .B1(n6965), .B2(n6559), .A(n6658), .ZN(n6560) );
  AOI21_X1 U7335 ( .B1(n6941), .B2(n6561), .A(n6560), .ZN(n6562) );
  OAI211_X1 U7336 ( .C1(n6962), .C2(n6564), .A(n6563), .B(n6562), .ZN(U2965)
         );
  AOI21_X1 U7337 ( .B1(n6523), .B2(n6565), .A(n6665), .ZN(n7002) );
  OAI22_X1 U7338 ( .A1(n6965), .A2(n7293), .B1(n7136), .B2(n5963), .ZN(n6567)
         );
  NOR2_X1 U7339 ( .A1(n7297), .A2(n6962), .ZN(n6566) );
  AOI211_X1 U7340 ( .C1(n6941), .C2(n7300), .A(n6567), .B(n6566), .ZN(n6568)
         );
  OAI21_X1 U7341 ( .B1(n7002), .B2(n7345), .A(n6568), .ZN(U2967) );
  OR2_X1 U7343 ( .A1(n6668), .A2(n6707), .ZN(n6578) );
  NAND2_X1 U7344 ( .A1(n6570), .A2(n6578), .ZN(n6683) );
  INV_X1 U7345 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n7126) );
  MUX2_X1 U7346 ( .A(n7126), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .S(n6668), 
        .Z(n6571) );
  XNOR2_X1 U7347 ( .A(n6683), .B(n6571), .ZN(n7120) );
  OAI22_X1 U7348 ( .A1(n6965), .A2(n7269), .B1(n7136), .B2(n7123), .ZN(n6573)
         );
  NOR2_X1 U7349 ( .A1(n7430), .A2(n6962), .ZN(n6572) );
  AOI211_X1 U7350 ( .C1(n6941), .C2(n7271), .A(n6573), .B(n6572), .ZN(n6574)
         );
  OAI21_X1 U7351 ( .B1(n7120), .B2(n7345), .A(n6574), .ZN(U2969) );
  AOI21_X1 U7352 ( .B1(n6576), .B2(n6578), .A(n6575), .ZN(n6577) );
  AOI21_X1 U7353 ( .B1(n4737), .B2(n6578), .A(n6577), .ZN(n6699) );
  NAND2_X1 U7354 ( .A1(n6699), .A2(n6971), .ZN(n6582) );
  AND2_X1 U7355 ( .A1(n7073), .A2(REIP_REG_16__SCAN_IN), .ZN(n6703) );
  NOR2_X1 U7356 ( .A1(n6975), .A2(n6579), .ZN(n6580) );
  AOI211_X1 U7357 ( .C1(n6969), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6703), 
        .B(n6580), .ZN(n6581) );
  OAI211_X1 U7358 ( .C1(n6962), .C2(n7426), .A(n6582), .B(n6581), .ZN(U2970)
         );
  XNOR2_X1 U7359 ( .A(n6668), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6584)
         );
  XNOR2_X1 U7360 ( .A(n6583), .B(n6584), .ZN(n7116) );
  NAND2_X1 U7361 ( .A1(n7116), .A2(n6971), .ZN(n6588) );
  AND2_X1 U7362 ( .A1(n7073), .A2(REIP_REG_15__SCAN_IN), .ZN(n7112) );
  NOR2_X1 U7363 ( .A1(n6975), .A2(n6585), .ZN(n6586) );
  AOI211_X1 U7364 ( .C1(n6969), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n7112), 
        .B(n6586), .ZN(n6587) );
  OAI211_X1 U7365 ( .C1(n6962), .C2(n6589), .A(n6588), .B(n6587), .ZN(U2971)
         );
  INV_X1 U7366 ( .A(n7248), .ZN(n6591) );
  AOI22_X1 U7367 ( .A1(n6969), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n7073), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n6590) );
  OAI21_X1 U7368 ( .B1(n6975), .B2(n6591), .A(n6590), .ZN(n6592) );
  AOI21_X1 U7369 ( .B1(n7249), .B2(n6970), .A(n6592), .ZN(n6593) );
  OAI21_X1 U7370 ( .B1(n6594), .B2(n7345), .A(n6593), .ZN(U2972) );
  INV_X1 U7371 ( .A(n6595), .ZN(n6599) );
  OAI21_X1 U7372 ( .B1(n6597), .B2(n6600), .A(n6596), .ZN(n6598) );
  AOI21_X1 U7373 ( .B1(n6599), .B2(n7132), .A(n6598), .ZN(n6603) );
  NAND3_X1 U7374 ( .A1(n6601), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n6600), .ZN(n6602) );
  OAI211_X1 U7375 ( .C1(n6604), .C2(n7055), .A(n6603), .B(n6602), .ZN(U2988)
         );
  INV_X1 U7376 ( .A(n6605), .ZN(n6608) );
  INV_X1 U7377 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6606) );
  NOR3_X1 U7378 ( .A1(n6610), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n6606), 
        .ZN(n6607) );
  AOI211_X1 U7379 ( .C1(n7132), .C2(n6609), .A(n6608), .B(n6607), .ZN(n6613)
         );
  OR2_X1 U7380 ( .A1(n6610), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6619)
         );
  INV_X1 U7381 ( .A(n6619), .ZN(n6611) );
  OAI21_X1 U7382 ( .B1(n6611), .B2(n6618), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n6612) );
  OAI211_X1 U7383 ( .C1(n6614), .C2(n7055), .A(n6613), .B(n6612), .ZN(U2990)
         );
  INV_X1 U7384 ( .A(n6615), .ZN(n6617) );
  NOR2_X1 U7385 ( .A1(n6917), .A2(n7042), .ZN(n6616) );
  AOI211_X1 U7386 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n6618), .A(n6617), .B(n6616), .ZN(n6620) );
  OAI211_X1 U7387 ( .C1(n6621), .C2(n7055), .A(n6620), .B(n6619), .ZN(U2991)
         );
  OAI21_X1 U7388 ( .B1(n6634), .B2(n6623), .A(n6622), .ZN(n6624) );
  AOI21_X1 U7389 ( .B1(n6625), .B2(n7132), .A(n6624), .ZN(n6629) );
  INV_X1 U7390 ( .A(n6626), .ZN(n6627) );
  OAI211_X1 U7391 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n7140), .B(n6627), .ZN(n6628) );
  OAI211_X1 U7392 ( .C1(n6630), .C2(n7055), .A(n6629), .B(n6628), .ZN(U2992)
         );
  XNOR2_X1 U7393 ( .A(n6632), .B(n6631), .ZN(n7336) );
  INV_X1 U7394 ( .A(n6633), .ZN(n6646) );
  AOI21_X1 U7395 ( .B1(n6646), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U7396 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  AOI211_X1 U7397 ( .C1(n7132), .C2(n7336), .A(n6637), .B(n6636), .ZN(n6638)
         );
  OAI21_X1 U7398 ( .B1(n6639), .B2(n7055), .A(n6638), .ZN(U2994) );
  NAND2_X1 U7399 ( .A1(n6640), .A2(n7132), .ZN(n6642) );
  OAI211_X1 U7400 ( .C1(n6643), .C2(n6645), .A(n6642), .B(n6641), .ZN(n6644)
         );
  AOI21_X1 U7401 ( .B1(n6646), .B2(n6645), .A(n6644), .ZN(n6647) );
  OAI21_X1 U7402 ( .B1(n6648), .B2(n7055), .A(n6647), .ZN(U2995) );
  OAI21_X1 U7403 ( .B1(n7330), .B2(n7042), .A(n6649), .ZN(n6654) );
  INV_X1 U7404 ( .A(n6650), .ZN(n6664) );
  NOR3_X1 U7405 ( .A1(n6664), .A2(n6652), .A3(n6651), .ZN(n6653) );
  AOI211_X1 U7406 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n6661), .A(n6654), .B(n6653), .ZN(n6655) );
  OAI21_X1 U7407 ( .B1(n6656), .B2(n7055), .A(n6655), .ZN(U2996) );
  NAND3_X1 U7408 ( .A1(n3655), .A2(n7133), .A3(n6657), .ZN(n6663) );
  OAI21_X1 U7409 ( .B1(n6659), .B2(n7042), .A(n6658), .ZN(n6660) );
  AOI21_X1 U7410 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n6661), .A(n6660), 
        .ZN(n6662) );
  OAI211_X1 U7411 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n6664), .A(n6663), .B(n6662), .ZN(U2997) );
  INV_X1 U7412 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6666) );
  AOI21_X1 U7413 ( .B1(n6668), .B2(n6666), .A(n6665), .ZN(n6670) );
  XNOR2_X1 U7414 ( .A(n6668), .B(n6667), .ZN(n6669) );
  XNOR2_X1 U7415 ( .A(n6670), .B(n6669), .ZN(n6972) );
  INV_X1 U7416 ( .A(n6972), .ZN(n6682) );
  NOR2_X1 U7417 ( .A1(n6671), .A2(n7126), .ZN(n6673) );
  OAI21_X1 U7418 ( .B1(n6673), .B2(n7063), .A(n6672), .ZN(n7125) );
  AOI21_X1 U7419 ( .B1(n6674), .B2(n7085), .A(n7125), .ZN(n6675) );
  OAI21_X1 U7420 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n7063), .A(n6675), 
        .ZN(n7001) );
  NOR2_X1 U7421 ( .A1(n6676), .A2(n7006), .ZN(n6678) );
  AOI22_X1 U7422 ( .A1(n7073), .A2(REIP_REG_20__SCAN_IN), .B1(n6678), .B2(
        n6677), .ZN(n6679) );
  OAI21_X1 U7423 ( .B1(n7308), .B2(n7042), .A(n6679), .ZN(n6680) );
  AOI21_X1 U7424 ( .B1(n7001), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n6680), 
        .ZN(n6681) );
  OAI21_X1 U7425 ( .B1(n6682), .B2(n7055), .A(n6681), .ZN(U2998) );
  NOR2_X1 U7426 ( .A1(n6570), .A2(n7126), .ZN(n6685) );
  NOR2_X1 U7427 ( .A1(n6683), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6684)
         );
  MUX2_X1 U7428 ( .A(n6685), .B(n6684), .S(n6526), .Z(n6687) );
  XNOR2_X1 U7429 ( .A(n6687), .B(n6686), .ZN(n6966) );
  INV_X1 U7430 ( .A(n6966), .ZN(n6695) );
  INV_X1 U7431 ( .A(n7125), .ZN(n6688) );
  OAI21_X1 U7432 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6689), .A(n6688), 
        .ZN(n6691) );
  OAI22_X1 U7433 ( .A1(n7284), .A2(n7042), .B1(n7136), .B2(n7280), .ZN(n6690)
         );
  AOI21_X1 U7434 ( .B1(n6691), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n6690), 
        .ZN(n6694) );
  NOR2_X1 U7435 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n7126), .ZN(n6692)
         );
  NAND2_X1 U7436 ( .A1(n7127), .A2(n6692), .ZN(n6693) );
  OAI211_X1 U7437 ( .C1(n6695), .C2(n7055), .A(n6694), .B(n6693), .ZN(U3000)
         );
  INV_X1 U7438 ( .A(n7110), .ZN(n6696) );
  AOI21_X1 U7439 ( .B1(n6698), .B2(n6697), .A(n6696), .ZN(n7114) );
  NAND2_X1 U7440 ( .A1(n6699), .A2(n7133), .ZN(n6706) );
  INV_X1 U7441 ( .A(n7265), .ZN(n6704) );
  OAI21_X1 U7442 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6700), .ZN(n6701) );
  NOR2_X1 U7443 ( .A1(n7119), .A2(n6701), .ZN(n6702) );
  AOI211_X1 U7444 ( .C1(n7132), .C2(n6704), .A(n6703), .B(n6702), .ZN(n6705)
         );
  OAI211_X1 U7445 ( .C1(n7114), .C2(n6707), .A(n6706), .B(n6705), .ZN(U3002)
         );
  OR3_X1 U7446 ( .A1(n7040), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6708), 
        .ZN(n6719) );
  AOI22_X1 U7447 ( .A1(n7073), .A2(REIP_REG_1__SCAN_IN), .B1(n6709), .B2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6718) );
  NAND2_X1 U7448 ( .A1(n3647), .A2(n6710), .ZN(n6714) );
  INV_X1 U7449 ( .A(n6712), .ZN(n6713) );
  XNOR2_X1 U7450 ( .A(n6714), .B(n6713), .ZN(n6929) );
  NAND2_X1 U7451 ( .A1(n6929), .A2(n7133), .ZN(n6717) );
  NAND2_X1 U7452 ( .A1(n7132), .A2(n6715), .ZN(n6716) );
  NAND4_X1 U7453 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(U3017)
         );
  INV_X1 U7454 ( .A(n6720), .ZN(n6724) );
  INV_X1 U7455 ( .A(n6721), .ZN(n7392) );
  OAI22_X1 U7456 ( .A1(n6724), .A2(n6723), .B1(n6722), .B2(n7392), .ZN(n6725)
         );
  MUX2_X1 U7457 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6725), .S(n7351), 
        .Z(U3456) );
  NAND2_X1 U7458 ( .A1(n7502), .A2(n6726), .ZN(n6734) );
  AOI211_X1 U7459 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6734), .A(n6728), .B(
        n6727), .ZN(n6733) );
  OAI21_X1 U7460 ( .B1(n6772), .B2(n6771), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6729) );
  OAI21_X1 U7461 ( .B1(n6731), .B2(n6730), .A(n6729), .ZN(n6732) );
  NAND2_X1 U7462 ( .A1(n6733), .A2(n6732), .ZN(n6770) );
  NAND2_X1 U7463 ( .A1(n6770), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6744)
         );
  AOI22_X1 U7464 ( .A1(n6772), .A2(n7516), .B1(n7508), .B2(n6771), .ZN(n6743)
         );
  INV_X1 U7465 ( .A(n6734), .ZN(n6773) );
  NAND2_X1 U7466 ( .A1(n7507), .A2(n6773), .ZN(n6742) );
  NAND2_X1 U7467 ( .A1(n6735), .A2(n7462), .ZN(n6739) );
  OR2_X1 U7468 ( .A1(n6737), .A2(n6736), .ZN(n6738) );
  NAND2_X1 U7469 ( .A1(n6739), .A2(n6738), .ZN(n6774) );
  NAND2_X1 U7470 ( .A1(n6740), .A2(n6774), .ZN(n6741) );
  NAND4_X1 U7471 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(U3132)
         );
  NAND2_X1 U7472 ( .A1(n6770), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6748)
         );
  AOI22_X1 U7473 ( .A1(n6772), .A2(n7538), .B1(n7539), .B2(n6771), .ZN(n6747)
         );
  NAND2_X1 U7474 ( .A1(n7536), .A2(n6773), .ZN(n6746) );
  NAND2_X1 U7475 ( .A1(n7537), .A2(n6774), .ZN(n6745) );
  NAND4_X1 U7476 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(U3133)
         );
  NAND2_X1 U7477 ( .A1(n6770), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6752)
         );
  AOI22_X1 U7478 ( .A1(n6772), .A2(n7556), .B1(n7557), .B2(n6771), .ZN(n6751)
         );
  NAND2_X1 U7479 ( .A1(n7554), .A2(n6773), .ZN(n6750) );
  NAND2_X1 U7480 ( .A1(n7555), .A2(n6774), .ZN(n6749) );
  NAND4_X1 U7481 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(U3134)
         );
  NAND2_X1 U7482 ( .A1(n6770), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6756)
         );
  AOI22_X1 U7483 ( .A1(n6772), .A2(n7574), .B1(n7575), .B2(n6771), .ZN(n6755)
         );
  NAND2_X1 U7484 ( .A1(n7572), .A2(n6773), .ZN(n6754) );
  NAND2_X1 U7485 ( .A1(n7573), .A2(n6774), .ZN(n6753) );
  NAND4_X1 U7486 ( .A1(n6756), .A2(n6755), .A3(n6754), .A4(n6753), .ZN(U3135)
         );
  NAND2_X1 U7487 ( .A1(n6770), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6760)
         );
  AOI22_X1 U7488 ( .A1(n6772), .A2(n7601), .B1(n7602), .B2(n6771), .ZN(n6759)
         );
  NAND2_X1 U7489 ( .A1(n7599), .A2(n6773), .ZN(n6758) );
  NAND2_X1 U7490 ( .A1(n7600), .A2(n6774), .ZN(n6757) );
  NAND4_X1 U7491 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(U3136)
         );
  NAND2_X1 U7492 ( .A1(n6770), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6764)
         );
  AOI22_X1 U7493 ( .A1(n6772), .A2(n7619), .B1(n7620), .B2(n6771), .ZN(n6763)
         );
  NAND2_X1 U7494 ( .A1(n7617), .A2(n6773), .ZN(n6762) );
  NAND2_X1 U7495 ( .A1(n7618), .A2(n6774), .ZN(n6761) );
  NAND4_X1 U7496 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(U3137)
         );
  NAND2_X1 U7497 ( .A1(n6770), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6769)
         );
  AOI22_X1 U7498 ( .A1(n6772), .A2(n7634), .B1(n7633), .B2(n6771), .ZN(n6768)
         );
  NAND2_X1 U7499 ( .A1(n7632), .A2(n6773), .ZN(n6767) );
  NAND2_X1 U7500 ( .A1(n6765), .A2(n6774), .ZN(n6766) );
  NAND4_X1 U7501 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(U3138)
         );
  NAND2_X1 U7502 ( .A1(n6770), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6778)
         );
  AOI22_X1 U7503 ( .A1(n6772), .A2(n7678), .B1(n7679), .B2(n6771), .ZN(n6777)
         );
  NAND2_X1 U7504 ( .A1(n7674), .A2(n6773), .ZN(n6776) );
  NAND2_X1 U7505 ( .A1(n7676), .A2(n6774), .ZN(n6775) );
  NAND4_X1 U7506 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(U3139)
         );
  NAND2_X1 U7507 ( .A1(n6832), .A2(n7415), .ZN(n6981) );
  AOI21_X1 U7508 ( .B1(n6779), .B2(n6981), .A(n7404), .ZN(n7403) );
  AOI21_X1 U7509 ( .B1(n7404), .B2(n6899), .A(n7403), .ZN(U3451) );
  INV_X1 U7510 ( .A(n7404), .ZN(n6795) );
  INV_X1 U7511 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6780) );
  NOR2_X1 U7512 ( .A1(n6795), .A2(n6780), .ZN(U3180) );
  AND2_X1 U7513 ( .A1(n7404), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7514 ( .A1(n7404), .A2(DATAWIDTH_REG_5__SCAN_IN), .ZN(U3177) );
  NOR2_X1 U7515 ( .A1(n6795), .A2(n6781), .ZN(U3176) );
  NOR2_X1 U7516 ( .A1(n6795), .A2(n6782), .ZN(U3175) );
  NOR2_X1 U7517 ( .A1(n6795), .A2(n6783), .ZN(U3174) );
  NOR2_X1 U7518 ( .A1(n6795), .A2(n6784), .ZN(U3173) );
  NOR2_X1 U7519 ( .A1(n6795), .A2(n6785), .ZN(U3172) );
  NOR2_X1 U7520 ( .A1(n6795), .A2(n6786), .ZN(U3171) );
  NOR2_X1 U7521 ( .A1(n6795), .A2(n6787), .ZN(U3170) );
  NOR2_X1 U7522 ( .A1(n6795), .A2(n6788), .ZN(U3169) );
  AND2_X1 U7523 ( .A1(n7404), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  NOR2_X1 U7524 ( .A1(n6795), .A2(n6789), .ZN(U3167) );
  NOR2_X1 U7525 ( .A1(n6795), .A2(n6790), .ZN(U3166) );
  AND2_X1 U7526 ( .A1(n7404), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  NOR2_X1 U7527 ( .A1(n6795), .A2(n6791), .ZN(U3164) );
  NOR2_X1 U7528 ( .A1(n6795), .A2(n6792), .ZN(U3163) );
  AND2_X1 U7529 ( .A1(n7404), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U7530 ( .A1(n7404), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  NOR2_X1 U7531 ( .A1(n6795), .A2(n6793), .ZN(U3160) );
  NOR2_X1 U7532 ( .A1(n6795), .A2(n6794), .ZN(U3159) );
  AND2_X1 U7533 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7404), .ZN(U3158) );
  AND2_X1 U7534 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n7404), .ZN(U3157) );
  AND2_X1 U7535 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7404), .ZN(U3156) );
  AND2_X1 U7536 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7404), .ZN(U3155) );
  AND2_X1 U7537 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7404), .ZN(U3154) );
  AND2_X1 U7538 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7404), .ZN(U3153) );
  AND2_X1 U7539 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7404), .ZN(U3152) );
  AND2_X1 U7540 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7404), .ZN(U3151) );
  AND2_X1 U7541 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6796), .ZN(U3019)
         );
  AND2_X1 U7542 ( .A1(n6812), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7543 ( .A(n7421), .ZN(n7411) );
  AOI21_X1 U7544 ( .B1(n6798), .B2(n6797), .A(n7411), .ZN(U2789) );
  AOI22_X1 U7545 ( .A1(n6828), .A2(LWORD_REG_0__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6800) );
  OAI21_X1 U7546 ( .B1(n6801), .B2(n6830), .A(n6800), .ZN(U2923) );
  AOI22_X1 U7547 ( .A1(n6828), .A2(LWORD_REG_1__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6802) );
  OAI21_X1 U7548 ( .B1(n6803), .B2(n6830), .A(n6802), .ZN(U2922) );
  AOI22_X1 U7549 ( .A1(n6828), .A2(LWORD_REG_2__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6804) );
  OAI21_X1 U7550 ( .B1(n6805), .B2(n6830), .A(n6804), .ZN(U2921) );
  AOI22_X1 U7551 ( .A1(n6828), .A2(LWORD_REG_3__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6806) );
  OAI21_X1 U7552 ( .B1(n6807), .B2(n6830), .A(n6806), .ZN(U2920) );
  AOI22_X1 U7553 ( .A1(n6828), .A2(LWORD_REG_4__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6808) );
  OAI21_X1 U7554 ( .B1(n6809), .B2(n6830), .A(n6808), .ZN(U2919) );
  AOI22_X1 U7555 ( .A1(n6828), .A2(LWORD_REG_5__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6810) );
  OAI21_X1 U7556 ( .B1(n6811), .B2(n6830), .A(n6810), .ZN(U2918) );
  AOI22_X1 U7557 ( .A1(n6828), .A2(LWORD_REG_6__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6813) );
  OAI21_X1 U7558 ( .B1(n4138), .B2(n6830), .A(n6813), .ZN(U2917) );
  AOI22_X1 U7559 ( .A1(n6828), .A2(LWORD_REG_7__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6814) );
  OAI21_X1 U7560 ( .B1(n4155), .B2(n6830), .A(n6814), .ZN(U2916) );
  AOI22_X1 U7561 ( .A1(n6828), .A2(LWORD_REG_8__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6815) );
  OAI21_X1 U7562 ( .B1(n6816), .B2(n6830), .A(n6815), .ZN(U2915) );
  AOI22_X1 U7563 ( .A1(n6828), .A2(LWORD_REG_9__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6817) );
  OAI21_X1 U7564 ( .B1(n6818), .B2(n6830), .A(n6817), .ZN(U2914) );
  AOI22_X1 U7565 ( .A1(n6828), .A2(LWORD_REG_10__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6819) );
  OAI21_X1 U7566 ( .B1(n6820), .B2(n6830), .A(n6819), .ZN(U2913) );
  AOI22_X1 U7567 ( .A1(n6828), .A2(LWORD_REG_11__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6821) );
  OAI21_X1 U7568 ( .B1(n6822), .B2(n6830), .A(n6821), .ZN(U2912) );
  AOI22_X1 U7569 ( .A1(n6828), .A2(LWORD_REG_12__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6823) );
  OAI21_X1 U7570 ( .B1(n4218), .B2(n6830), .A(n6823), .ZN(U2911) );
  AOI22_X1 U7571 ( .A1(n6828), .A2(LWORD_REG_13__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6824) );
  OAI21_X1 U7572 ( .B1(n6825), .B2(n6830), .A(n6824), .ZN(U2910) );
  AOI22_X1 U7573 ( .A1(n6828), .A2(LWORD_REG_14__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6826) );
  OAI21_X1 U7574 ( .B1(n6827), .B2(n6830), .A(n6826), .ZN(U2909) );
  AOI22_X1 U7575 ( .A1(n6828), .A2(LWORD_REG_15__SCAN_IN), .B1(n6812), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6829) );
  OAI21_X1 U7576 ( .B1(n6831), .B2(n6830), .A(n6829), .ZN(U2908) );
  NAND2_X1 U7577 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7411), .ZN(n6859) );
  CLKBUF_X1 U7578 ( .A(n6859), .Z(n6883) );
  INV_X1 U7579 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6834) );
  INV_X1 U7580 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U7581 ( .A1(n7411), .A2(n6832), .ZN(n6860) );
  INV_X1 U7582 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6836) );
  OAI222_X1 U7583 ( .A1(n6883), .A2(n6834), .B1(n6833), .B2(n7411), .C1(n6860), 
        .C2(n6836), .ZN(U3184) );
  INV_X1 U7584 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6835) );
  INV_X1 U7585 ( .A(n7421), .ZN(n7424) );
  CLKBUF_X1 U7586 ( .A(n6860), .Z(n6879) );
  OAI222_X1 U7587 ( .A1(n6859), .A2(n6836), .B1(n6835), .B2(n7424), .C1(n6879), 
        .C2(n7029), .ZN(U3185) );
  OAI222_X1 U7588 ( .A1(n6859), .A2(n7029), .B1(n6837), .B2(n7411), .C1(n6879), 
        .C2(n7179), .ZN(U3186) );
  INV_X1 U7589 ( .A(REIP_REG_5__SCAN_IN), .ZN(n7188) );
  OAI222_X1 U7590 ( .A1(n6859), .A2(n7179), .B1(n6838), .B2(n7424), .C1(n6860), 
        .C2(n7188), .ZN(U3187) );
  INV_X1 U7591 ( .A(REIP_REG_6__SCAN_IN), .ZN(n7204) );
  OAI222_X1 U7592 ( .A1(n6859), .A2(n7188), .B1(n6839), .B2(n7411), .C1(n6860), 
        .C2(n7204), .ZN(U3188) );
  INV_X1 U7593 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6842) );
  OAI222_X1 U7594 ( .A1(n6859), .A2(n7204), .B1(n6840), .B2(n7424), .C1(n6860), 
        .C2(n6842), .ZN(U3189) );
  OAI222_X1 U7595 ( .A1(n6859), .A2(n6842), .B1(n6841), .B2(n7424), .C1(n6860), 
        .C2(n6844), .ZN(U3190) );
  INV_X1 U7596 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6843) );
  OAI222_X1 U7597 ( .A1(n6883), .A2(n6844), .B1(n6843), .B2(n7424), .C1(n6860), 
        .C2(n6846), .ZN(U3191) );
  INV_X1 U7598 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6848) );
  OAI222_X1 U7599 ( .A1(n6883), .A2(n6846), .B1(n6845), .B2(n7424), .C1(n6860), 
        .C2(n6848), .ZN(U3192) );
  INV_X1 U7600 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6847) );
  OAI222_X1 U7601 ( .A1(n6883), .A2(n6848), .B1(n6847), .B2(n7424), .C1(n6860), 
        .C2(n6850), .ZN(U3193) );
  INV_X1 U7602 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6849) );
  OAI222_X1 U7603 ( .A1(n6883), .A2(n6850), .B1(n6849), .B2(n7424), .C1(n6860), 
        .C2(n7231), .ZN(U3194) );
  OAI222_X1 U7604 ( .A1(n6883), .A2(n7231), .B1(n6851), .B2(n7424), .C1(n6860), 
        .C2(n7243), .ZN(U3195) );
  OAI222_X1 U7605 ( .A1(n6883), .A2(n7243), .B1(n6852), .B2(n7424), .C1(n6879), 
        .C2(n6854), .ZN(U3196) );
  INV_X1 U7606 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6853) );
  OAI222_X1 U7607 ( .A1(n6883), .A2(n6854), .B1(n6853), .B2(n7424), .C1(n6860), 
        .C2(n7257), .ZN(U3197) );
  OAI222_X1 U7608 ( .A1(n6883), .A2(n7257), .B1(n6855), .B2(n7424), .C1(n6879), 
        .C2(n7258), .ZN(U3198) );
  INV_X1 U7609 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6856) );
  OAI222_X1 U7610 ( .A1(n6859), .A2(n7258), .B1(n6856), .B2(n7424), .C1(n6879), 
        .C2(n7123), .ZN(U3199) );
  OAI222_X1 U7611 ( .A1(n6859), .A2(n7123), .B1(n6857), .B2(n7424), .C1(n6879), 
        .C2(n7280), .ZN(U3200) );
  OAI222_X1 U7612 ( .A1(n6859), .A2(n7280), .B1(n6858), .B2(n7424), .C1(n6879), 
        .C2(n5963), .ZN(U3201) );
  OAI222_X1 U7613 ( .A1(n6883), .A2(n5963), .B1(n6861), .B2(n7424), .C1(n6860), 
        .C2(n7304), .ZN(U3202) );
  OAI222_X1 U7614 ( .A1(n6883), .A2(n7304), .B1(n6862), .B2(n7424), .C1(n6879), 
        .C2(n6864), .ZN(U3203) );
  INV_X1 U7615 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n6863) );
  OAI222_X1 U7616 ( .A1(n6883), .A2(n6864), .B1(n6863), .B2(n7411), .C1(n6879), 
        .C2(n7320), .ZN(U3204) );
  OAI222_X1 U7617 ( .A1(n6883), .A2(n7320), .B1(n6865), .B2(n7424), .C1(n6879), 
        .C2(n6867), .ZN(U3205) );
  INV_X1 U7618 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6866) );
  OAI222_X1 U7619 ( .A1(n6883), .A2(n6867), .B1(n6866), .B2(n7411), .C1(n6868), 
        .C2(n6879), .ZN(U3206) );
  OAI222_X1 U7620 ( .A1(n7135), .A2(n6879), .B1(n6869), .B2(n7411), .C1(n6868), 
        .C2(n6883), .ZN(U3207) );
  INV_X1 U7621 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6870) );
  OAI222_X1 U7622 ( .A1(n6883), .A2(n7135), .B1(n6870), .B2(n7424), .C1(n6879), 
        .C2(n6872), .ZN(U3208) );
  OAI222_X1 U7623 ( .A1(n6883), .A2(n6872), .B1(n6871), .B2(n7411), .C1(n6874), 
        .C2(n6879), .ZN(U3209) );
  OAI222_X1 U7624 ( .A1(n6883), .A2(n6874), .B1(n6873), .B2(n7424), .C1(n6876), 
        .C2(n6879), .ZN(U3210) );
  OAI222_X1 U7625 ( .A1(n6883), .A2(n6876), .B1(n6875), .B2(n7411), .C1(n6877), 
        .C2(n6879), .ZN(U3211) );
  OAI222_X1 U7626 ( .A1(n6879), .A2(n6882), .B1(n6878), .B2(n7411), .C1(n6877), 
        .C2(n6883), .ZN(U3212) );
  INV_X1 U7627 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6881) );
  OAI222_X1 U7628 ( .A1(n6883), .A2(n6882), .B1(n6881), .B2(n7411), .C1(n6880), 
        .C2(n6879), .ZN(U3213) );
  INV_X1 U7629 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U7630 ( .A1(n7411), .A2(n6896), .B1(n6884), .B2(n7421), .ZN(U3445)
         );
  NOR4_X1 U7631 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6888) );
  NOR4_X1 U7632 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_31__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n6887) );
  NOR4_X1 U7633 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(DATAWIDTH_REG_17__SCAN_IN), .ZN(
        n6886) );
  NOR4_X1 U7634 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n6885) );
  NAND4_X1 U7635 ( .A1(n6888), .A2(n6887), .A3(n6886), .A4(n6885), .ZN(n6894)
         );
  NOR4_X1 U7636 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_15__SCAN_IN), .ZN(
        n6892) );
  AOI211_X1 U7637 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_16__SCAN_IN), .B(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6891) );
  NOR4_X1 U7638 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6890)
         );
  NOR4_X1 U7639 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_18__SCAN_IN), .ZN(
        n6889) );
  NAND4_X1 U7640 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), .ZN(n6893)
         );
  NOR2_X1 U7641 ( .A1(n6894), .A2(n6893), .ZN(n6911) );
  NOR3_X1 U7642 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n6904) );
  NOR2_X1 U7643 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), 
        .ZN(n6900) );
  OAI21_X1 U7644 ( .B1(n6904), .B2(n6900), .A(n6911), .ZN(n6895) );
  OAI21_X1 U7645 ( .B1(n6911), .B2(n6896), .A(n6895), .ZN(U2795) );
  OAI22_X1 U7646 ( .A1(n7421), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(
        BE_N_REG_2__SCAN_IN), .B2(n7424), .ZN(n6897) );
  INV_X1 U7647 ( .A(n6897), .ZN(U3446) );
  NOR3_X1 U7648 ( .A1(n6899), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_0__SCAN_IN), .ZN(n6898) );
  AOI221_X1 U7649 ( .B1(n6900), .B2(n6899), .C1(REIP_REG_0__SCAN_IN), .C2(
        REIP_REG_1__SCAN_IN), .A(n6898), .ZN(n6902) );
  INV_X1 U7650 ( .A(n6911), .ZN(n6908) );
  AOI22_X1 U7651 ( .A1(n6911), .A2(n6902), .B1(n6901), .B2(n6908), .ZN(U3468)
         );
  AOI22_X1 U7652 ( .A1(n7424), .A2(n6906), .B1(n6903), .B2(n7421), .ZN(U3447)
         );
  OAI21_X1 U7653 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6904), .A(n6911), .ZN(n6905)
         );
  OAI21_X1 U7654 ( .B1(n6911), .B2(n6906), .A(n6905), .ZN(U2794) );
  OAI22_X1 U7655 ( .A1(n7421), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(n7424), .ZN(n6907) );
  INV_X1 U7656 ( .A(n6907), .ZN(U3448) );
  NOR2_X1 U7657 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6910) );
  INV_X1 U7658 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U7659 ( .A1(n6911), .A2(n6910), .B1(n6909), .B2(n6908), .ZN(U3469)
         );
  INV_X1 U7660 ( .A(n7156), .ZN(n6936) );
  XNOR2_X1 U7661 ( .A(n3631), .B(n6912), .ZN(n7157) );
  AOI22_X1 U7662 ( .A1(n6936), .A2(n6925), .B1(n6924), .B2(n7157), .ZN(n6913)
         );
  OAI21_X1 U7663 ( .B1(n6927), .B2(n7164), .A(n6913), .ZN(U2857) );
  AOI22_X1 U7664 ( .A1(n7522), .A2(n6925), .B1(n6924), .B2(n7336), .ZN(n6914)
         );
  OAI21_X1 U7665 ( .B1(n6927), .B2(n6915), .A(n6914), .ZN(U2835) );
  OAI22_X1 U7666 ( .A1(n7582), .A2(n6454), .B1(n6917), .B2(n6916), .ZN(n6918)
         );
  INV_X1 U7667 ( .A(n6918), .ZN(n6919) );
  OAI21_X1 U7668 ( .B1(n6927), .B2(n6920), .A(n6919), .ZN(U2832) );
  INV_X1 U7669 ( .A(EBX_REG_5__SCAN_IN), .ZN(n7180) );
  NAND2_X1 U7670 ( .A1(n5031), .A2(n6921), .ZN(n6922) );
  AND2_X1 U7671 ( .A1(n6923), .A2(n6922), .ZN(n7183) );
  AOI22_X1 U7672 ( .A1(n7191), .A2(n6925), .B1(n6924), .B2(n7183), .ZN(n6926)
         );
  OAI21_X1 U7673 ( .B1(n6927), .B2(n7180), .A(n6926), .ZN(U2854) );
  AOI22_X1 U7674 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6969), .B1(n7073), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6931) );
  AOI22_X1 U7675 ( .A1(n6971), .A2(n6929), .B1(n6928), .B2(n6970), .ZN(n6930)
         );
  OAI211_X1 U7676 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6975), .A(n6931), 
        .B(n6930), .ZN(U2985) );
  AOI22_X1 U7677 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6969), .B1(n7073), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6938) );
  NAND2_X1 U7678 ( .A1(n6932), .A2(n6933), .ZN(n6934) );
  XOR2_X1 U7679 ( .A(n6935), .B(n6934), .Z(n7066) );
  AOI22_X1 U7680 ( .A1(n7066), .A2(n6971), .B1(n6970), .B2(n6936), .ZN(n6937)
         );
  OAI211_X1 U7681 ( .C1(n6975), .C2(n7152), .A(n6938), .B(n6937), .ZN(U2984)
         );
  XNOR2_X1 U7682 ( .A(n6940), .B(n6939), .ZN(n7056) );
  INV_X1 U7683 ( .A(n7056), .ZN(n6943) );
  INV_X1 U7684 ( .A(n7195), .ZN(n6942) );
  AOI222_X1 U7685 ( .A1(n6943), .A2(n6971), .B1(n6970), .B2(n7191), .C1(n6942), 
        .C2(n6941), .ZN(n6944) );
  NAND2_X1 U7686 ( .A1(n7073), .A2(REIP_REG_5__SCAN_IN), .ZN(n7049) );
  OAI211_X1 U7687 ( .C1(n6965), .C2(n7181), .A(n6944), .B(n7049), .ZN(U2981)
         );
  AOI22_X1 U7688 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6969), .B1(n7073), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U7689 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  XNOR2_X1 U7690 ( .A(n6945), .B(n6948), .ZN(n7044) );
  AOI22_X1 U7691 ( .A1(n6971), .A2(n7044), .B1(n6949), .B2(n6970), .ZN(n6950)
         );
  OAI211_X1 U7692 ( .C1(n6975), .C2(n7199), .A(n6951), .B(n6950), .ZN(U2980)
         );
  AOI22_X1 U7693 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6969), .B1(n7073), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6958) );
  OAI21_X1 U7694 ( .B1(n6952), .B2(n6954), .A(n6953), .ZN(n6955) );
  INV_X1 U7695 ( .A(n6955), .ZN(n7074) );
  INV_X1 U7696 ( .A(n6956), .ZN(n7211) );
  AOI22_X1 U7697 ( .A1(n7074), .A2(n6971), .B1(n6970), .B2(n7211), .ZN(n6957)
         );
  OAI211_X1 U7698 ( .C1(n6975), .C2(n7216), .A(n6958), .B(n6957), .ZN(U2979)
         );
  INV_X1 U7699 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n7235) );
  OAI21_X1 U7700 ( .B1(n6959), .B2(n6961), .A(n3648), .ZN(n7007) );
  OAI22_X1 U7701 ( .A1(n7237), .A2(n6962), .B1(n7236), .B2(n6975), .ZN(n6963)
         );
  AOI21_X1 U7702 ( .B1(n6971), .B2(n7007), .A(n6963), .ZN(n6964) );
  NAND2_X1 U7703 ( .A1(n7073), .A2(REIP_REG_13__SCAN_IN), .ZN(n7016) );
  OAI211_X1 U7704 ( .C1(n6965), .C2(n7235), .A(n6964), .B(n7016), .ZN(U2973)
         );
  AOI22_X1 U7705 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6969), .B1(n7073), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n6968) );
  AOI22_X1 U7706 ( .A1(n6966), .A2(n6971), .B1(n6970), .B2(n7286), .ZN(n6967)
         );
  OAI211_X1 U7707 ( .C1(n6975), .C2(n7288), .A(n6968), .B(n6967), .ZN(U2968)
         );
  AOI22_X1 U7708 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6969), .B1(n7073), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n6974) );
  AOI22_X1 U7709 ( .A1(n6972), .A2(n6971), .B1(n6970), .B2(n6413), .ZN(n6973)
         );
  OAI211_X1 U7710 ( .C1(n6975), .C2(n7307), .A(n6974), .B(n6973), .ZN(U2966)
         );
  AND2_X1 U7711 ( .A1(n6976), .A2(n7397), .ZN(n6978) );
  OAI22_X1 U7712 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6979), .B1(n6978), .B2(
        n6977), .ZN(U2790) );
  NOR2_X1 U7713 ( .A1(n7411), .A2(D_C_N_REG_SCAN_IN), .ZN(n6980) );
  AOI22_X1 U7714 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7411), .B1(n6981), .B2(
        n6980), .ZN(U2791) );
  NOR2_X1 U7715 ( .A1(n6997), .A2(n6982), .ZN(n6983) );
  AOI22_X1 U7716 ( .A1(n6985), .A2(n6997), .B1(n6984), .B2(n6983), .ZN(U3474)
         );
  INV_X1 U7717 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6986) );
  AOI22_X1 U7718 ( .A1(n7411), .A2(READREQUEST_REG_SCAN_IN), .B1(n6986), .B2(
        n7421), .ZN(U3470) );
  AND2_X1 U7719 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n7408) );
  NOR2_X1 U7720 ( .A1(n7415), .A2(n6987), .ZN(n7413) );
  AOI21_X1 U7721 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7413), .ZN(n6990)
         );
  NOR2_X1 U7722 ( .A1(n6988), .A2(n7414), .ZN(n7406) );
  INV_X1 U7723 ( .A(n7406), .ZN(n7419) );
  OAI211_X1 U7724 ( .C1(n7408), .C2(n6990), .A(n6989), .B(n7419), .ZN(U3182)
         );
  NOR2_X1 U7725 ( .A1(n7400), .A2(READY_N), .ZN(n7382) );
  AOI21_X1 U7726 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n7382), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6992) );
  OAI21_X1 U7727 ( .B1(n6993), .B2(n6992), .A(n6991), .ZN(U3150) );
  AOI211_X1 U7728 ( .C1(n6995), .C2(n7497), .A(n7505), .B(n6994), .ZN(n6996)
         );
  OAI21_X1 U7729 ( .B1(n6996), .B2(n7400), .A(n7393), .ZN(n7000) );
  AOI211_X1 U7730 ( .C1(n6828), .C2(n7414), .A(n6998), .B(n6997), .ZN(n6999)
         );
  MUX2_X1 U7731 ( .A(n7000), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6999), .Z(
        U3472) );
  AOI22_X1 U7732 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n7001), .B1(n7073), .B2(REIP_REG_19__SCAN_IN), .ZN(n7005) );
  INV_X1 U7733 ( .A(n7002), .ZN(n7003) );
  AOI22_X1 U7734 ( .A1(n7003), .A2(n7133), .B1(n7132), .B2(n7295), .ZN(n7004)
         );
  OAI211_X1 U7735 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n7006), .A(n7005), .B(n7004), .ZN(U2999) );
  AOI22_X1 U7736 ( .A1(n7007), .A2(n7133), .B1(n7132), .B2(n7233), .ZN(n7017)
         );
  OAI21_X1 U7737 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n7009), .A(n7008), 
        .ZN(n7015) );
  NAND4_X1 U7738 ( .A1(n7013), .A2(n7012), .A3(n7011), .A4(n7010), .ZN(n7014)
         );
  NAND4_X1 U7739 ( .A1(n7017), .A2(n7016), .A3(n7015), .A4(n7014), .ZN(U3005)
         );
  OAI211_X1 U7740 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n7028), .B(n7027), .ZN(n7026) );
  NOR2_X1 U7741 ( .A1(n7042), .A2(n7169), .ZN(n7023) );
  NOR2_X1 U7742 ( .A1(n7063), .A2(n7027), .ZN(n7064) );
  OAI21_X1 U7743 ( .B1(n7019), .B2(n7018), .A(n7088), .ZN(n7067) );
  NOR2_X1 U7744 ( .A1(n7064), .A2(n7067), .ZN(n7039) );
  OAI21_X1 U7745 ( .B1(n7039), .B2(n7021), .A(n7020), .ZN(n7022) );
  AOI211_X1 U7746 ( .C1(n7024), .C2(n7133), .A(n7023), .B(n7022), .ZN(n7025)
         );
  OAI21_X1 U7747 ( .B1(n7041), .B2(n7026), .A(n7025), .ZN(U3014) );
  NAND2_X1 U7748 ( .A1(n7028), .A2(n7027), .ZN(n7034) );
  OAI22_X1 U7749 ( .A1(n7042), .A2(n7030), .B1(n7029), .B2(n7136), .ZN(n7031)
         );
  AOI21_X1 U7750 ( .B1(n7032), .B2(n7133), .A(n7031), .ZN(n7033) );
  OAI21_X1 U7751 ( .B1(n7034), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n7033), 
        .ZN(n7035) );
  INV_X1 U7752 ( .A(n7035), .ZN(n7036) );
  OAI21_X1 U7753 ( .B1(n7039), .B2(n4676), .A(n7036), .ZN(U3015) );
  NOR3_X1 U7754 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n7038), .A3(n7037), 
        .ZN(n7058) );
  OAI21_X1 U7755 ( .B1(n7041), .B2(n7040), .A(n7039), .ZN(n7059) );
  AOI211_X1 U7756 ( .C1(n7087), .C2(n7051), .A(n7058), .B(n7059), .ZN(n7046)
         );
  OAI22_X1 U7757 ( .A1(n7042), .A2(n7196), .B1(n7204), .B2(n7136), .ZN(n7043)
         );
  AOI21_X1 U7758 ( .B1(n7044), .B2(n7133), .A(n7043), .ZN(n7045) );
  OAI221_X1 U7759 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n7048), .C1(n7047), .C2(n7046), .A(n7045), .ZN(U3012) );
  INV_X1 U7760 ( .A(n7049), .ZN(n7050) );
  AOI21_X1 U7761 ( .B1(n7132), .B2(n7183), .A(n7050), .ZN(n7054) );
  NAND3_X1 U7762 ( .A1(n7087), .A2(n7052), .A3(n7051), .ZN(n7053) );
  OAI211_X1 U7763 ( .C1(n7056), .C2(n7055), .A(n7054), .B(n7053), .ZN(n7057)
         );
  AOI211_X1 U7764 ( .C1(INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n7059), .A(n7058), 
        .B(n7057), .ZN(n7060) );
  INV_X1 U7765 ( .A(n7060), .ZN(U3013) );
  NOR3_X1 U7766 ( .A1(n7063), .A2(n7062), .A3(n7061), .ZN(n7065) );
  AOI211_X1 U7767 ( .C1(n7132), .C2(n7157), .A(n7065), .B(n7064), .ZN(n7072)
         );
  AOI22_X1 U7768 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n7067), .B1(n7066), 
        .B2(n7133), .ZN(n7071) );
  NAND2_X1 U7769 ( .A1(n7073), .A2(REIP_REG_2__SCAN_IN), .ZN(n7070) );
  NAND3_X1 U7770 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n7068), .A3(n4897), 
        .ZN(n7069) );
  NAND4_X1 U7771 ( .A1(n7072), .A2(n7071), .A3(n7070), .A4(n7069), .ZN(U3016)
         );
  AOI22_X1 U7772 ( .A1(n7132), .A2(n7206), .B1(n7073), .B2(REIP_REG_7__SCAN_IN), .ZN(n7076) );
  AOI22_X1 U7773 ( .A1(n7079), .A2(n7077), .B1(n7133), .B2(n7074), .ZN(n7075)
         );
  OAI211_X1 U7774 ( .C1(n7078), .C2(n7077), .A(n7076), .B(n7075), .ZN(U3011)
         );
  NAND2_X1 U7775 ( .A1(n7080), .A2(n7079), .ZN(n7102) );
  OAI21_X1 U7776 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n7081), .ZN(n7093) );
  AOI21_X1 U7777 ( .B1(n7132), .B2(n7083), .A(n7082), .ZN(n7092) );
  AOI22_X1 U7778 ( .A1(n7087), .A2(n7086), .B1(n7085), .B2(n7084), .ZN(n7089)
         );
  NAND2_X1 U7779 ( .A1(n7089), .A2(n7088), .ZN(n7098) );
  AOI22_X1 U7780 ( .A1(n7090), .A2(n7133), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n7098), .ZN(n7091) );
  OAI211_X1 U7781 ( .C1(n7102), .C2(n7093), .A(n7092), .B(n7091), .ZN(U3008)
         );
  INV_X1 U7782 ( .A(n7094), .ZN(n7095) );
  AOI21_X1 U7783 ( .B1(n7132), .B2(n7096), .A(n7095), .ZN(n7101) );
  INV_X1 U7784 ( .A(n7097), .ZN(n7099) );
  AOI22_X1 U7785 ( .A1(n7099), .A2(n7133), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n7098), .ZN(n7100) );
  OAI211_X1 U7786 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n7102), .A(n7101), 
        .B(n7100), .ZN(U3009) );
  INV_X1 U7787 ( .A(n7103), .ZN(n7104) );
  AOI21_X1 U7788 ( .B1(n7132), .B2(n7105), .A(n7104), .ZN(n7109) );
  AOI22_X1 U7789 ( .A1(n7107), .A2(n7133), .B1(n4727), .B2(n7106), .ZN(n7108)
         );
  OAI211_X1 U7790 ( .C1(n7110), .C2(n4727), .A(n7109), .B(n7108), .ZN(U3007)
         );
  INV_X1 U7791 ( .A(n7111), .ZN(n7113) );
  AOI21_X1 U7792 ( .B1(n7132), .B2(n7113), .A(n7112), .ZN(n7118) );
  INV_X1 U7793 ( .A(n7114), .ZN(n7115) );
  AOI22_X1 U7794 ( .A1(n7116), .A2(n7133), .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n7115), .ZN(n7117) );
  OAI211_X1 U7795 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n7119), .A(n7118), .B(n7117), .ZN(U3003) );
  INV_X1 U7796 ( .A(n7120), .ZN(n7122) );
  AOI22_X1 U7797 ( .A1(n7122), .A2(n7133), .B1(n7132), .B2(n7121), .ZN(n7129)
         );
  NOR2_X1 U7798 ( .A1(n7136), .A2(n7123), .ZN(n7124) );
  AOI221_X1 U7799 ( .B1(n7127), .B2(n7126), .C1(n7125), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n7124), .ZN(n7128) );
  NAND2_X1 U7800 ( .A1(n7129), .A2(n7128), .ZN(U3001) );
  INV_X1 U7801 ( .A(n7130), .ZN(n7134) );
  AOI22_X1 U7802 ( .A1(n7134), .A2(n7133), .B1(n7132), .B2(n7131), .ZN(n7142)
         );
  NOR2_X1 U7803 ( .A1(n7136), .A2(n7135), .ZN(n7137) );
  AOI221_X1 U7804 ( .B1(n7140), .B2(n7139), .C1(n7138), .C2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n7137), .ZN(n7141) );
  NAND2_X1 U7805 ( .A1(n7142), .A2(n7141), .ZN(U2993) );
  AOI22_X1 U7806 ( .A1(n7337), .A2(n7143), .B1(REIP_REG_0__SCAN_IN), .B2(n7266), .ZN(n7148) );
  NAND2_X1 U7807 ( .A1(n7332), .A2(EBX_REG_0__SCAN_IN), .ZN(n7145) );
  OAI21_X1 U7808 ( .B1(n7335), .B2(n7339), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n7144) );
  OAI211_X1 U7809 ( .C1(n7167), .C2(n4062), .A(n7145), .B(n7144), .ZN(n7146)
         );
  INV_X1 U7810 ( .A(n7146), .ZN(n7147) );
  OAI211_X1 U7811 ( .C1(n7172), .C2(n7149), .A(n7148), .B(n7147), .ZN(U2827)
         );
  AOI22_X1 U7812 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n7335), .B1(n7268), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n7163) );
  OAI211_X1 U7813 ( .C1(REIP_REG_2__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        n7151), .B(n7150), .ZN(n7155) );
  INV_X1 U7814 ( .A(n7152), .ZN(n7153) );
  NAND2_X1 U7815 ( .A1(n7339), .A2(n7153), .ZN(n7154) );
  OAI211_X1 U7816 ( .C1(n7172), .C2(n7156), .A(n7155), .B(n7154), .ZN(n7161)
         );
  NAND2_X1 U7817 ( .A1(n7337), .A2(n7157), .ZN(n7158) );
  OAI21_X1 U7818 ( .B1(n7159), .B2(n7167), .A(n7158), .ZN(n7160) );
  NOR2_X1 U7819 ( .A1(n7161), .A2(n7160), .ZN(n7162) );
  OAI211_X1 U7820 ( .C1(n7164), .C2(n7312), .A(n7163), .B(n7162), .ZN(U2825)
         );
  NOR3_X1 U7821 ( .A1(n7316), .A2(n7165), .A3(REIP_REG_4__SCAN_IN), .ZN(n7166)
         );
  AOI211_X1 U7822 ( .C1(n7335), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n7279), 
        .B(n7166), .ZN(n7177) );
  INV_X1 U7823 ( .A(n7347), .ZN(n7168) );
  OAI22_X1 U7824 ( .A1(n7329), .A2(n7169), .B1(n7168), .B2(n7167), .ZN(n7175)
         );
  INV_X1 U7825 ( .A(n7170), .ZN(n7171) );
  OAI22_X1 U7826 ( .A1(n7173), .A2(n7172), .B1(n7171), .B2(n7323), .ZN(n7174)
         );
  AOI211_X1 U7827 ( .C1(EBX_REG_4__SCAN_IN), .C2(n7332), .A(n7175), .B(n7174), 
        .ZN(n7176) );
  OAI211_X1 U7828 ( .C1(n7179), .C2(n7178), .A(n7177), .B(n7176), .ZN(U2823)
         );
  OAI22_X1 U7829 ( .A1(n7181), .A2(n7294), .B1(n7180), .B2(n7312), .ZN(n7182)
         );
  AOI211_X1 U7830 ( .C1(n7337), .C2(n7183), .A(n7279), .B(n7182), .ZN(n7194)
         );
  NOR2_X1 U7831 ( .A1(n7268), .A2(n7184), .ZN(n7185) );
  NOR2_X1 U7832 ( .A1(n7186), .A2(n7185), .ZN(n7212) );
  INV_X1 U7833 ( .A(n7187), .ZN(n7189) );
  OAI21_X1 U7834 ( .B1(n7316), .B2(n7189), .A(n7188), .ZN(n7192) );
  AOI22_X1 U7835 ( .A1(n7212), .A2(n7192), .B1(n7191), .B2(n7190), .ZN(n7193)
         );
  OAI211_X1 U7836 ( .C1(n7195), .C2(n7323), .A(n7194), .B(n7193), .ZN(U2822)
         );
  OAI22_X1 U7837 ( .A1(n7197), .A2(n7312), .B1(n7329), .B2(n7196), .ZN(n7198)
         );
  AOI211_X1 U7838 ( .C1(n7335), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n7279), 
        .B(n7198), .ZN(n7203) );
  NOR2_X1 U7839 ( .A1(REIP_REG_6__SCAN_IN), .A2(n7205), .ZN(n7213) );
  OAI22_X1 U7840 ( .A1(n7200), .A2(n7325), .B1(n7199), .B2(n7323), .ZN(n7201)
         );
  AOI211_X1 U7841 ( .C1(REIP_REG_6__SCAN_IN), .C2(n7212), .A(n7213), .B(n7201), 
        .ZN(n7202) );
  NAND2_X1 U7842 ( .A1(n7203), .A2(n7202), .ZN(U2821) );
  NOR3_X1 U7843 ( .A1(n7205), .A2(n7204), .A3(REIP_REG_7__SCAN_IN), .ZN(n7210)
         );
  AOI22_X1 U7844 ( .A1(EBX_REG_7__SCAN_IN), .A2(n7332), .B1(n7337), .B2(n7206), 
        .ZN(n7207) );
  OAI211_X1 U7845 ( .C1(n7294), .C2(n7208), .A(n7207), .B(n7291), .ZN(n7209)
         );
  AOI211_X1 U7846 ( .C1(n7211), .C2(n7338), .A(n7210), .B(n7209), .ZN(n7215)
         );
  OAI21_X1 U7847 ( .B1(n7213), .B2(n7212), .A(REIP_REG_7__SCAN_IN), .ZN(n7214)
         );
  OAI211_X1 U7848 ( .C1(n7323), .C2(n7216), .A(n7215), .B(n7214), .ZN(U2820)
         );
  NOR2_X1 U7849 ( .A1(REIP_REG_12__SCAN_IN), .A2(n7232), .ZN(n7217) );
  NAND2_X1 U7850 ( .A1(n7218), .A2(n7217), .ZN(n7241) );
  OAI22_X1 U7851 ( .A1(n7220), .A2(n7312), .B1(n7329), .B2(n7219), .ZN(n7221)
         );
  NOR2_X1 U7852 ( .A1(n7279), .A2(n7221), .ZN(n7222) );
  OAI211_X1 U7853 ( .C1(n7223), .C2(n7294), .A(n7241), .B(n7222), .ZN(n7224)
         );
  INV_X1 U7854 ( .A(n7224), .ZN(n7225) );
  OAI21_X1 U7855 ( .B1(n7226), .B2(n7325), .A(n7225), .ZN(n7227) );
  AOI21_X1 U7856 ( .B1(n7228), .B2(n7339), .A(n7227), .ZN(n7229) );
  OAI21_X1 U7857 ( .B1(n7242), .B2(n7231), .A(n7229), .ZN(U2815) );
  NOR3_X1 U7858 ( .A1(n7232), .A2(n7231), .A3(n7230), .ZN(n7244) );
  AOI22_X1 U7859 ( .A1(n7337), .A2(n7233), .B1(n7244), .B2(n7243), .ZN(n7234)
         );
  OAI211_X1 U7860 ( .C1(n7294), .C2(n7235), .A(n7234), .B(n7291), .ZN(n7239)
         );
  OAI22_X1 U7861 ( .A1(n7237), .A2(n7325), .B1(n7236), .B2(n7323), .ZN(n7238)
         );
  AOI211_X1 U7862 ( .C1(EBX_REG_13__SCAN_IN), .C2(n7332), .A(n7239), .B(n7238), 
        .ZN(n7240) );
  OAI221_X1 U7863 ( .B1(n7243), .B2(n7242), .C1(n7243), .C2(n7241), .A(n7240), 
        .ZN(U2814) );
  AOI21_X1 U7864 ( .B1(REIP_REG_13__SCAN_IN), .B2(n7244), .A(
        REIP_REG_14__SCAN_IN), .ZN(n7252) );
  OAI22_X1 U7865 ( .A1(n7246), .A2(n7294), .B1(n7329), .B2(n7245), .ZN(n7247)
         );
  AOI211_X1 U7866 ( .C1(n7332), .C2(EBX_REG_14__SCAN_IN), .A(n7279), .B(n7247), 
        .ZN(n7251) );
  AOI22_X1 U7867 ( .A1(n7249), .A2(n7338), .B1(n7339), .B2(n7248), .ZN(n7250)
         );
  OAI211_X1 U7868 ( .C1(n7252), .C2(n7253), .A(n7251), .B(n7250), .ZN(U2813)
         );
  OAI21_X1 U7869 ( .B1(REIP_REG_15__SCAN_IN), .B2(n7256), .A(n7253), .ZN(n7254) );
  AOI22_X1 U7870 ( .A1(n7255), .A2(n7339), .B1(REIP_REG_16__SCAN_IN), .B2(
        n7254), .ZN(n7264) );
  INV_X1 U7871 ( .A(n7426), .ZN(n7262) );
  NOR2_X1 U7872 ( .A1(n7257), .A2(n7256), .ZN(n7281) );
  AOI22_X1 U7873 ( .A1(EBX_REG_16__SCAN_IN), .A2(n7332), .B1(n7281), .B2(n7258), .ZN(n7259) );
  OAI211_X1 U7874 ( .C1(n7260), .C2(n7294), .A(n7259), .B(n7291), .ZN(n7261)
         );
  AOI21_X1 U7875 ( .B1(n7262), .B2(n7338), .A(n7261), .ZN(n7263) );
  OAI211_X1 U7876 ( .C1(n7329), .C2(n7265), .A(n7264), .B(n7263), .ZN(U2811)
         );
  AOI21_X1 U7877 ( .B1(REIP_REG_16__SCAN_IN), .B2(n7281), .A(
        REIP_REG_17__SCAN_IN), .ZN(n7276) );
  OAI21_X1 U7878 ( .B1(n7268), .B2(n7267), .A(n7266), .ZN(n7302) );
  OAI22_X1 U7879 ( .A1(n7269), .A2(n7294), .B1(n6441), .B2(n7312), .ZN(n7270)
         );
  AOI211_X1 U7880 ( .C1(n7339), .C2(n7271), .A(n7279), .B(n7270), .ZN(n7275)
         );
  OAI22_X1 U7881 ( .A1(n7430), .A2(n7325), .B1(n7329), .B2(n7272), .ZN(n7273)
         );
  INV_X1 U7882 ( .A(n7273), .ZN(n7274) );
  OAI211_X1 U7883 ( .C1(n7276), .C2(n7302), .A(n7275), .B(n7274), .ZN(U2810)
         );
  OAI22_X1 U7884 ( .A1(n7277), .A2(n7312), .B1(n7280), .B2(n7302), .ZN(n7278)
         );
  AOI211_X1 U7885 ( .C1(n7335), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n7279), 
        .B(n7278), .ZN(n7283) );
  NAND3_X1 U7886 ( .A1(n7282), .A2(n7281), .A3(n7280), .ZN(n7303) );
  OAI211_X1 U7887 ( .C1(n7329), .C2(n7284), .A(n7283), .B(n7303), .ZN(n7285)
         );
  AOI21_X1 U7888 ( .B1(n7286), .B2(n7338), .A(n7285), .ZN(n7287) );
  OAI21_X1 U7889 ( .B1(n7288), .B2(n7323), .A(n7287), .ZN(U2809) );
  NOR2_X1 U7890 ( .A1(n7316), .A2(REIP_REG_19__SCAN_IN), .ZN(n7289) );
  AOI22_X1 U7891 ( .A1(EBX_REG_19__SCAN_IN), .A2(n7332), .B1(n7290), .B2(n7289), .ZN(n7292) );
  OAI211_X1 U7892 ( .C1(n7294), .C2(n7293), .A(n7292), .B(n7291), .ZN(n7299)
         );
  INV_X1 U7893 ( .A(n7295), .ZN(n7296) );
  OAI22_X1 U7894 ( .A1(n7297), .A2(n7325), .B1(n7329), .B2(n7296), .ZN(n7298)
         );
  AOI211_X1 U7895 ( .C1(n7300), .C2(n7339), .A(n7299), .B(n7298), .ZN(n7301)
         );
  OAI221_X1 U7896 ( .B1(n5963), .B2(n7303), .C1(n5963), .C2(n7302), .A(n7301), 
        .ZN(U2808) );
  OAI21_X1 U7897 ( .B1(n7316), .B2(n7305), .A(n7304), .ZN(n7306) );
  AOI22_X1 U7898 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n7335), .B1(n7314), 
        .B2(n7306), .ZN(n7311) );
  OAI22_X1 U7899 ( .A1(n7308), .A2(n7329), .B1(n7307), .B2(n7323), .ZN(n7309)
         );
  AOI21_X1 U7900 ( .B1(n6413), .B2(n7338), .A(n7309), .ZN(n7310) );
  OAI211_X1 U7901 ( .C1(n7313), .C2(n7312), .A(n7311), .B(n7310), .ZN(U2807)
         );
  INV_X1 U7902 ( .A(n7314), .ZN(n7315) );
  OAI21_X1 U7903 ( .B1(REIP_REG_21__SCAN_IN), .B2(n7316), .A(n7315), .ZN(n7319) );
  AOI22_X1 U7904 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n7335), .B1(
        EBX_REG_22__SCAN_IN), .B2(n7332), .ZN(n7317) );
  INV_X1 U7905 ( .A(n7317), .ZN(n7318) );
  AOI221_X1 U7906 ( .B1(n7321), .B2(n7320), .C1(n7319), .C2(
        REIP_REG_22__SCAN_IN), .A(n7318), .ZN(n7328) );
  INV_X1 U7907 ( .A(n7322), .ZN(n7324) );
  OAI22_X1 U7908 ( .A1(n7442), .A2(n7325), .B1(n7324), .B2(n7323), .ZN(n7326)
         );
  INV_X1 U7909 ( .A(n7326), .ZN(n7327) );
  OAI211_X1 U7910 ( .C1(n7330), .C2(n7329), .A(n7328), .B(n7327), .ZN(U2805)
         );
  AOI22_X1 U7911 ( .A1(EBX_REG_24__SCAN_IN), .A2(n7332), .B1(
        REIP_REG_24__SCAN_IN), .B2(n7331), .ZN(n7344) );
  AOI22_X1 U7912 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n7335), .B1(n7334), 
        .B2(n7333), .ZN(n7343) );
  AOI22_X1 U7913 ( .A1(n7522), .A2(n7338), .B1(n7337), .B2(n7336), .ZN(n7342)
         );
  NAND2_X1 U7914 ( .A1(n7340), .A2(n7339), .ZN(n7341) );
  NAND4_X1 U7915 ( .A1(n7344), .A2(n7343), .A3(n7342), .A4(n7341), .ZN(U2803)
         );
  OAI21_X1 U7916 ( .B1(n7346), .B2(n7373), .A(n7345), .ZN(U2793) );
  INV_X1 U7917 ( .A(n4821), .ZN(n7348) );
  NAND4_X1 U7918 ( .A1(n7349), .A2(n7383), .A3(n7348), .A4(n7347), .ZN(n7350)
         );
  OAI21_X1 U7919 ( .B1(n7351), .B2(n4097), .A(n7350), .ZN(U3455) );
  OAI211_X1 U7920 ( .C1(n7354), .C2(n7353), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n7352), .ZN(n7357) );
  OAI211_X1 U7921 ( .C1(n7496), .C2(n7357), .A(n7356), .B(n7355), .ZN(n7359)
         );
  NAND2_X1 U7922 ( .A1(n7496), .A2(n7357), .ZN(n7358) );
  NAND2_X1 U7923 ( .A1(n7359), .A2(n7358), .ZN(n7362) );
  AND2_X1 U7924 ( .A1(n7363), .A2(n7362), .ZN(n7361) );
  OAI222_X1 U7925 ( .A1(n7364), .A2(n7365), .B1(n7363), .B2(n7362), .C1(n7361), 
        .C2(n7360), .ZN(n7367) );
  NAND2_X1 U7926 ( .A1(n7365), .A2(n7364), .ZN(n7366) );
  AOI21_X1 U7927 ( .B1(n7367), .B2(n7366), .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .ZN(n7371) );
  NOR4_X1 U7928 ( .A1(n7371), .A2(n7370), .A3(n7369), .A4(n7368), .ZN(n7372)
         );
  OAI221_X1 U7929 ( .B1(n7375), .B2(n7374), .C1(n7375), .C2(n7373), .A(n7372), 
        .ZN(n7396) );
  OAI22_X1 U7930 ( .A1(n7396), .A2(n7377), .B1(n7376), .B2(n7414), .ZN(n7378)
         );
  AOI221_X1 U7931 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7391), .C1(n7414), .C2(
        n7391), .A(n7400), .ZN(n7394) );
  AOI21_X1 U7932 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n7394), .A(n7381), .ZN(
        n7387) );
  AOI21_X1 U7933 ( .B1(n7383), .B2(n7382), .A(n7397), .ZN(n7384) );
  INV_X1 U7934 ( .A(n7384), .ZN(n7385) );
  NAND2_X1 U7935 ( .A1(n7391), .A2(n7385), .ZN(n7386) );
  OAI211_X1 U7936 ( .C1(n7388), .C2(n7391), .A(n7387), .B(n7386), .ZN(U3149)
         );
  OAI221_X1 U7937 ( .B1(n7390), .B2(STATE2_REG_0__SCAN_IN), .C1(n7390), .C2(
        n7391), .A(n7389), .ZN(U3453) );
  OAI21_X1 U7938 ( .B1(n7393), .B2(n7392), .A(n7391), .ZN(n7401) );
  AOI211_X1 U7939 ( .C1(n7397), .C2(n7396), .A(n7395), .B(n7394), .ZN(n7398)
         );
  OAI221_X1 U7940 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n7401), .C1(n7400), .C2(
        n7399), .A(n7398), .ZN(U3148) );
  AOI21_X1 U7941 ( .B1(n7404), .B2(STATEBS16_REG_SCAN_IN), .A(n7403), .ZN(
        n7402) );
  INV_X1 U7942 ( .A(n7402), .ZN(U2792) );
  AOI21_X1 U7943 ( .B1(n7404), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(n7403), .ZN(
        n7405) );
  INV_X1 U7944 ( .A(n7405), .ZN(U3452) );
  NAND2_X1 U7945 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n7410) );
  NAND2_X1 U7946 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n7407) );
  AOI221_X1 U7947 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7412), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7418) );
  AOI221_X1 U7948 ( .B1(n7408), .B2(n7407), .C1(n7406), .C2(n7407), .A(n7418), 
        .ZN(n7409) );
  OAI221_X1 U7949 ( .B1(n7411), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7411), 
        .C2(n7410), .A(n7409), .ZN(U3181) );
  AOI21_X1 U7950 ( .B1(n7413), .B2(n7412), .A(STATE_REG_2__SCAN_IN), .ZN(n7420) );
  AOI221_X1 U7951 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7414), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7416) );
  AOI221_X1 U7952 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7416), .C2(HOLD), .A(n7415), .ZN(n7417) );
  OAI22_X1 U7953 ( .A1(n7420), .A2(n7419), .B1(n7418), .B2(n7417), .ZN(U3183)
         );
  AOI22_X1 U7954 ( .A1(n7424), .A2(n7423), .B1(n7422), .B2(n7421), .ZN(U3473)
         );
  INV_X1 U7955 ( .A(n7520), .ZN(n7580) );
  OAI22_X1 U7956 ( .A1(n7426), .A2(n7581), .B1(n7580), .B2(n7425), .ZN(n7427)
         );
  INV_X1 U7957 ( .A(n7427), .ZN(n7429) );
  AOI22_X1 U7958 ( .A1(n7585), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n7584), .ZN(n7428) );
  NAND2_X1 U7959 ( .A1(n7429), .A2(n7428), .ZN(U2875) );
  OAI22_X1 U7960 ( .A1(n7430), .A2(n7581), .B1(n5077), .B2(n7580), .ZN(n7431)
         );
  INV_X1 U7961 ( .A(n7431), .ZN(n7433) );
  AOI22_X1 U7962 ( .A1(n7585), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n7584), .ZN(n7432) );
  NAND2_X1 U7963 ( .A1(n7433), .A2(n7432), .ZN(U2874) );
  OAI22_X1 U7964 ( .A1(n7435), .A2(n7581), .B1(n7580), .B2(n7434), .ZN(n7436)
         );
  INV_X1 U7965 ( .A(n7436), .ZN(n7438) );
  AOI22_X1 U7966 ( .A1(n7585), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n7584), .ZN(n7437) );
  NAND2_X1 U7967 ( .A1(n7438), .A2(n7437), .ZN(U2873) );
  AOI22_X1 U7968 ( .A1(n6413), .A2(n7521), .B1(n7520), .B2(DATAI_4_), .ZN(
        n7440) );
  AOI22_X1 U7969 ( .A1(n7585), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n7584), .ZN(n7439) );
  NAND2_X1 U7970 ( .A1(n7440), .A2(n7439), .ZN(U2871) );
  INV_X1 U7971 ( .A(DATAI_6_), .ZN(n7441) );
  OAI22_X1 U7972 ( .A1(n7442), .A2(n7581), .B1(n7441), .B2(n7580), .ZN(n7443)
         );
  INV_X1 U7973 ( .A(n7443), .ZN(n7445) );
  AOI22_X1 U7974 ( .A1(n7585), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n7584), .ZN(n7444) );
  NAND2_X1 U7975 ( .A1(n7445), .A2(n7444), .ZN(U2869) );
  OR2_X1 U7976 ( .A1(n7446), .A2(n7482), .ZN(n7447) );
  NAND2_X1 U7977 ( .A1(n7447), .A2(n7499), .ZN(n7455) );
  INV_X1 U7978 ( .A(n7455), .ZN(n7452) );
  NOR2_X1 U7979 ( .A1(n7502), .A2(n7448), .ZN(n7639) );
  INV_X1 U7980 ( .A(n7639), .ZN(n7449) );
  OAI21_X1 U7981 ( .B1(n7451), .B2(n7450), .A(n7449), .ZN(n7456) );
  AOI22_X1 U7982 ( .A1(n7452), .A2(n7456), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7453), .ZN(n7644) );
  AOI22_X1 U7983 ( .A1(n7507), .A2(n7639), .B1(n7516), .B2(n7640), .ZN(n7458)
         );
  OR2_X1 U7984 ( .A1(n7499), .A2(n7453), .ZN(n7454) );
  OAI211_X1 U7985 ( .C1(n7456), .C2(n7455), .A(n7513), .B(n7454), .ZN(n7641)
         );
  AOI22_X1 U7986 ( .A1(n7641), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n7508), 
        .B2(n7638), .ZN(n7457) );
  OAI211_X1 U7987 ( .C1(n7644), .C2(n7519), .A(n7458), .B(n7457), .ZN(U3108)
         );
  NOR2_X1 U7988 ( .A1(n7459), .A2(n7511), .ZN(n7467) );
  NOR2_X1 U7989 ( .A1(n7460), .A2(n4062), .ZN(n7504) );
  INV_X1 U7990 ( .A(n7461), .ZN(n7646) );
  AOI21_X1 U7991 ( .B1(n7504), .B2(n7462), .A(n7646), .ZN(n7466) );
  INV_X1 U7992 ( .A(n7466), .ZN(n7463) );
  AOI22_X1 U7993 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7464), .B1(n7467), .B2(
        n7463), .ZN(n7651) );
  AOI22_X1 U7994 ( .A1(n7507), .A2(n7646), .B1(n7508), .B2(n7647), .ZN(n7470)
         );
  AOI22_X1 U7995 ( .A1(n7467), .A2(n7466), .B1(n7511), .B2(n7465), .ZN(n7468)
         );
  NAND2_X1 U7996 ( .A1(n7513), .A2(n7468), .ZN(n7648) );
  AOI22_X1 U7997 ( .A1(n7648), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n7516), 
        .B2(n7645), .ZN(n7469) );
  OAI211_X1 U7998 ( .C1(n7651), .C2(n7519), .A(n7470), .B(n7469), .ZN(U3076)
         );
  NAND2_X1 U7999 ( .A1(n7471), .A2(STATEBS16_REG_SCAN_IN), .ZN(n7472) );
  NAND2_X1 U8000 ( .A1(n7472), .A2(n7499), .ZN(n7478) );
  NOR2_X1 U8001 ( .A1(n7502), .A2(n7476), .ZN(n7653) );
  AOI21_X1 U8002 ( .B1(n7504), .B2(n7473), .A(n7653), .ZN(n7475) );
  OAI22_X1 U8003 ( .A1(n7505), .A2(n7476), .B1(n7478), .B2(n7475), .ZN(n7474)
         );
  AOI22_X1 U8004 ( .A1(n7507), .A2(n7653), .B1(n7508), .B2(n7654), .ZN(n7481)
         );
  INV_X1 U8005 ( .A(n7475), .ZN(n7479) );
  NAND2_X1 U8006 ( .A1(n7511), .A2(n7476), .ZN(n7477) );
  OAI211_X1 U8007 ( .C1(n7479), .C2(n7478), .A(n7513), .B(n7477), .ZN(n7655)
         );
  AOI22_X1 U8008 ( .A1(n7655), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n7516), 
        .B2(n7652), .ZN(n7480) );
  OAI211_X1 U8009 ( .C1(n7658), .C2(n7519), .A(n7481), .B(n7480), .ZN(U3060)
         );
  INV_X1 U8010 ( .A(n7482), .ZN(n7483) );
  AOI21_X1 U8011 ( .B1(n7484), .B2(n7483), .A(n7511), .ZN(n7491) );
  AND2_X1 U8012 ( .A1(n7495), .A2(n7485), .ZN(n7660) );
  AOI21_X1 U8013 ( .B1(n7504), .B2(n7486), .A(n7660), .ZN(n7490) );
  INV_X1 U8014 ( .A(n7490), .ZN(n7488) );
  INV_X1 U8015 ( .A(n7489), .ZN(n7487) );
  AOI22_X1 U8016 ( .A1(n7491), .A2(n7488), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7487), .ZN(n7665) );
  AOI22_X1 U8017 ( .A1(n7507), .A2(n7660), .B1(n7516), .B2(n7659), .ZN(n7494)
         );
  AOI22_X1 U8018 ( .A1(n7491), .A2(n7490), .B1(n7489), .B2(n7511), .ZN(n7492)
         );
  NAND2_X1 U8019 ( .A1(n7513), .A2(n7492), .ZN(n7662) );
  AOI22_X1 U8020 ( .A1(n7662), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n7508), 
        .B2(n7661), .ZN(n7493) );
  OAI211_X1 U8021 ( .C1(n7665), .C2(n7519), .A(n7494), .B(n7493), .ZN(U3044)
         );
  NAND2_X1 U8022 ( .A1(n7496), .A2(n7495), .ZN(n7510) );
  OR2_X1 U8023 ( .A1(n7498), .A2(n7497), .ZN(n7500) );
  NAND2_X1 U8024 ( .A1(n7500), .A2(n7499), .ZN(n7514) );
  AOI21_X1 U8025 ( .B1(n7504), .B2(n7503), .A(n7666), .ZN(n7509) );
  OAI22_X1 U8026 ( .A1(n7505), .A2(n7510), .B1(n7514), .B2(n7509), .ZN(n7506)
         );
  AOI22_X1 U8027 ( .A1(n7667), .A2(n7508), .B1(n7507), .B2(n7666), .ZN(n7518)
         );
  INV_X1 U8028 ( .A(n7509), .ZN(n7515) );
  NAND2_X1 U8029 ( .A1(n7511), .A2(n7510), .ZN(n7512) );
  OAI211_X1 U8030 ( .C1(n7515), .C2(n7514), .A(n7513), .B(n7512), .ZN(n7668)
         );
  AOI22_X1 U8031 ( .A1(n7668), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n7516), 
        .B2(n7680), .ZN(n7517) );
  OAI211_X1 U8032 ( .C1(n7672), .C2(n7519), .A(n7518), .B(n7517), .ZN(U3028)
         );
  AOI22_X1 U8033 ( .A1(n7522), .A2(n7521), .B1(DATAI_8_), .B2(n7520), .ZN(
        n7524) );
  AOI22_X1 U8034 ( .A1(n7585), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n7584), .ZN(n7523) );
  NAND2_X1 U8035 ( .A1(n7524), .A2(n7523), .ZN(U2867) );
  AOI22_X1 U8036 ( .A1(n7536), .A2(n7639), .B1(n7538), .B2(n7640), .ZN(n7526)
         );
  AOI22_X1 U8037 ( .A1(n7641), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n7539), 
        .B2(n7638), .ZN(n7525) );
  OAI211_X1 U8038 ( .C1(n7644), .C2(n7535), .A(n7526), .B(n7525), .ZN(U3109)
         );
  AOI22_X1 U8039 ( .A1(n7536), .A2(n7646), .B1(n7539), .B2(n7647), .ZN(n7528)
         );
  AOI22_X1 U8040 ( .A1(n7648), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n7538), 
        .B2(n7645), .ZN(n7527) );
  OAI211_X1 U8041 ( .C1(n7651), .C2(n7535), .A(n7528), .B(n7527), .ZN(U3077)
         );
  AOI22_X1 U8042 ( .A1(n7536), .A2(n7653), .B1(n7539), .B2(n7654), .ZN(n7530)
         );
  AOI22_X1 U8043 ( .A1(n7655), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n7538), 
        .B2(n7652), .ZN(n7529) );
  OAI211_X1 U8044 ( .C1(n7658), .C2(n7535), .A(n7530), .B(n7529), .ZN(U3061)
         );
  AOI22_X1 U8045 ( .A1(n7536), .A2(n7660), .B1(n7539), .B2(n7661), .ZN(n7532)
         );
  AOI22_X1 U8046 ( .A1(n7662), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n7538), 
        .B2(n7659), .ZN(n7531) );
  OAI211_X1 U8047 ( .C1(n7665), .C2(n7535), .A(n7532), .B(n7531), .ZN(U3045)
         );
  AOI22_X1 U8048 ( .A1(n7680), .A2(n7538), .B1(n7536), .B2(n7666), .ZN(n7534)
         );
  AOI22_X1 U8049 ( .A1(n7668), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n7539), 
        .B2(n7667), .ZN(n7533) );
  OAI211_X1 U8050 ( .C1(n7672), .C2(n7535), .A(n7534), .B(n7533), .ZN(U3029)
         );
  INV_X1 U8051 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n7542) );
  AOI22_X1 U8052 ( .A1(n7537), .A2(n7675), .B1(n7536), .B2(n7673), .ZN(n7541)
         );
  AOI22_X1 U8053 ( .A1(n7680), .A2(n7539), .B1(n7538), .B2(n7677), .ZN(n7540)
         );
  OAI211_X1 U8054 ( .C1(n7684), .C2(n7542), .A(n7541), .B(n7540), .ZN(U3021)
         );
  AOI22_X1 U8055 ( .A1(n7554), .A2(n7639), .B1(n7557), .B2(n7638), .ZN(n7544)
         );
  AOI22_X1 U8056 ( .A1(n7641), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n7556), 
        .B2(n7640), .ZN(n7543) );
  OAI211_X1 U8057 ( .C1(n7644), .C2(n7553), .A(n7544), .B(n7543), .ZN(U3110)
         );
  AOI22_X1 U8058 ( .A1(n7554), .A2(n7646), .B1(n7556), .B2(n7645), .ZN(n7546)
         );
  AOI22_X1 U8059 ( .A1(n7648), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n7557), 
        .B2(n7647), .ZN(n7545) );
  OAI211_X1 U8060 ( .C1(n7651), .C2(n7553), .A(n7546), .B(n7545), .ZN(U3078)
         );
  AOI22_X1 U8061 ( .A1(n7554), .A2(n7653), .B1(n7557), .B2(n7654), .ZN(n7548)
         );
  AOI22_X1 U8062 ( .A1(n7655), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n7556), 
        .B2(n7652), .ZN(n7547) );
  OAI211_X1 U8063 ( .C1(n7658), .C2(n7553), .A(n7548), .B(n7547), .ZN(U3062)
         );
  AOI22_X1 U8064 ( .A1(n7554), .A2(n7660), .B1(n7557), .B2(n7661), .ZN(n7550)
         );
  AOI22_X1 U8065 ( .A1(n7662), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n7556), 
        .B2(n7659), .ZN(n7549) );
  OAI211_X1 U8066 ( .C1(n7665), .C2(n7553), .A(n7550), .B(n7549), .ZN(U3046)
         );
  AOI22_X1 U8067 ( .A1(n7667), .A2(n7557), .B1(n7554), .B2(n7666), .ZN(n7552)
         );
  AOI22_X1 U8068 ( .A1(n7668), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n7556), 
        .B2(n7680), .ZN(n7551) );
  OAI211_X1 U8069 ( .C1(n7672), .C2(n7553), .A(n7552), .B(n7551), .ZN(U3030)
         );
  AOI22_X1 U8070 ( .A1(n7555), .A2(n7675), .B1(n7554), .B2(n7673), .ZN(n7559)
         );
  AOI22_X1 U8071 ( .A1(n7680), .A2(n7557), .B1(n7556), .B2(n7677), .ZN(n7558)
         );
  OAI211_X1 U8072 ( .C1(n7684), .C2(n7560), .A(n7559), .B(n7558), .ZN(U3022)
         );
  AOI22_X1 U8073 ( .A1(n7572), .A2(n7639), .B1(n7574), .B2(n7640), .ZN(n7562)
         );
  AOI22_X1 U8074 ( .A1(n7641), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n7575), 
        .B2(n7638), .ZN(n7561) );
  OAI211_X1 U8075 ( .C1(n7644), .C2(n7571), .A(n7562), .B(n7561), .ZN(U3111)
         );
  AOI22_X1 U8076 ( .A1(n7572), .A2(n7646), .B1(n7574), .B2(n7645), .ZN(n7564)
         );
  AOI22_X1 U8077 ( .A1(n7648), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n7575), 
        .B2(n7647), .ZN(n7563) );
  OAI211_X1 U8078 ( .C1(n7651), .C2(n7571), .A(n7564), .B(n7563), .ZN(U3079)
         );
  AOI22_X1 U8079 ( .A1(n7572), .A2(n7653), .B1(n7574), .B2(n7652), .ZN(n7566)
         );
  AOI22_X1 U8080 ( .A1(n7655), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n7575), 
        .B2(n7654), .ZN(n7565) );
  OAI211_X1 U8081 ( .C1(n7658), .C2(n7571), .A(n7566), .B(n7565), .ZN(U3063)
         );
  AOI22_X1 U8082 ( .A1(n7572), .A2(n7660), .B1(n7575), .B2(n7661), .ZN(n7568)
         );
  AOI22_X1 U8083 ( .A1(n7662), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n7574), 
        .B2(n7659), .ZN(n7567) );
  OAI211_X1 U8084 ( .C1(n7665), .C2(n7571), .A(n7568), .B(n7567), .ZN(U3047)
         );
  AOI22_X1 U8085 ( .A1(n7667), .A2(n7575), .B1(n7572), .B2(n7666), .ZN(n7570)
         );
  AOI22_X1 U8086 ( .A1(n7668), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n7574), 
        .B2(n7680), .ZN(n7569) );
  OAI211_X1 U8087 ( .C1(n7672), .C2(n7571), .A(n7570), .B(n7569), .ZN(U3031)
         );
  AOI22_X1 U8088 ( .A1(n7573), .A2(n7675), .B1(n7572), .B2(n7673), .ZN(n7577)
         );
  AOI22_X1 U8089 ( .A1(n7680), .A2(n7575), .B1(n7574), .B2(n7677), .ZN(n7576)
         );
  OAI211_X1 U8090 ( .C1(n7684), .C2(n7578), .A(n7577), .B(n7576), .ZN(U3023)
         );
  OAI22_X1 U8091 ( .A1(n7582), .A2(n7581), .B1(n7580), .B2(n7579), .ZN(n7583)
         );
  INV_X1 U8092 ( .A(n7583), .ZN(n7587) );
  AOI22_X1 U8093 ( .A1(n7585), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n7584), .ZN(n7586) );
  NAND2_X1 U8094 ( .A1(n7587), .A2(n7586), .ZN(U2864) );
  AOI22_X1 U8095 ( .A1(n7599), .A2(n7639), .B1(n7602), .B2(n7638), .ZN(n7589)
         );
  AOI22_X1 U8096 ( .A1(n7641), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n7601), 
        .B2(n7640), .ZN(n7588) );
  OAI211_X1 U8097 ( .C1(n7644), .C2(n7598), .A(n7589), .B(n7588), .ZN(U3112)
         );
  AOI22_X1 U8098 ( .A1(n7599), .A2(n7646), .B1(n7602), .B2(n7647), .ZN(n7591)
         );
  AOI22_X1 U8099 ( .A1(n7648), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n7601), 
        .B2(n7645), .ZN(n7590) );
  OAI211_X1 U8100 ( .C1(n7651), .C2(n7598), .A(n7591), .B(n7590), .ZN(U3080)
         );
  AOI22_X1 U8101 ( .A1(n7599), .A2(n7653), .B1(n7601), .B2(n7652), .ZN(n7593)
         );
  AOI22_X1 U8102 ( .A1(n7655), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n7602), 
        .B2(n7654), .ZN(n7592) );
  OAI211_X1 U8103 ( .C1(n7658), .C2(n7598), .A(n7593), .B(n7592), .ZN(U3064)
         );
  AOI22_X1 U8104 ( .A1(n7599), .A2(n7660), .B1(n7601), .B2(n7659), .ZN(n7595)
         );
  AOI22_X1 U8105 ( .A1(n7662), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n7602), 
        .B2(n7661), .ZN(n7594) );
  OAI211_X1 U8106 ( .C1(n7665), .C2(n7598), .A(n7595), .B(n7594), .ZN(U3048)
         );
  AOI22_X1 U8107 ( .A1(n7667), .A2(n7602), .B1(n7599), .B2(n7666), .ZN(n7597)
         );
  AOI22_X1 U8108 ( .A1(n7668), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n7601), 
        .B2(n7680), .ZN(n7596) );
  OAI211_X1 U8109 ( .C1(n7672), .C2(n7598), .A(n7597), .B(n7596), .ZN(U3032)
         );
  INV_X1 U8110 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n7605) );
  AOI22_X1 U8111 ( .A1(n7600), .A2(n7675), .B1(n7599), .B2(n7673), .ZN(n7604)
         );
  AOI22_X1 U8112 ( .A1(n7680), .A2(n7602), .B1(n7601), .B2(n7677), .ZN(n7603)
         );
  OAI211_X1 U8113 ( .C1(n7684), .C2(n7605), .A(n7604), .B(n7603), .ZN(U3024)
         );
  AOI22_X1 U8114 ( .A1(n7617), .A2(n7639), .B1(n7620), .B2(n7638), .ZN(n7607)
         );
  AOI22_X1 U8115 ( .A1(n7641), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n7619), 
        .B2(n7640), .ZN(n7606) );
  OAI211_X1 U8116 ( .C1(n7644), .C2(n7616), .A(n7607), .B(n7606), .ZN(U3113)
         );
  AOI22_X1 U8117 ( .A1(n7617), .A2(n7646), .B1(n7620), .B2(n7647), .ZN(n7609)
         );
  AOI22_X1 U8118 ( .A1(n7648), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n7619), 
        .B2(n7645), .ZN(n7608) );
  OAI211_X1 U8119 ( .C1(n7651), .C2(n7616), .A(n7609), .B(n7608), .ZN(U3081)
         );
  AOI22_X1 U8120 ( .A1(n7617), .A2(n7653), .B1(n7619), .B2(n7652), .ZN(n7611)
         );
  AOI22_X1 U8121 ( .A1(n7655), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n7620), 
        .B2(n7654), .ZN(n7610) );
  OAI211_X1 U8122 ( .C1(n7658), .C2(n7616), .A(n7611), .B(n7610), .ZN(U3065)
         );
  AOI22_X1 U8123 ( .A1(n7617), .A2(n7660), .B1(n7620), .B2(n7661), .ZN(n7613)
         );
  AOI22_X1 U8124 ( .A1(n7662), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n7619), 
        .B2(n7659), .ZN(n7612) );
  OAI211_X1 U8125 ( .C1(n7665), .C2(n7616), .A(n7613), .B(n7612), .ZN(U3049)
         );
  AOI22_X1 U8126 ( .A1(n7667), .A2(n7620), .B1(n7617), .B2(n7666), .ZN(n7615)
         );
  AOI22_X1 U8127 ( .A1(n7668), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n7619), 
        .B2(n7680), .ZN(n7614) );
  OAI211_X1 U8128 ( .C1(n7672), .C2(n7616), .A(n7615), .B(n7614), .ZN(U3033)
         );
  INV_X1 U8129 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n7623) );
  AOI22_X1 U8130 ( .A1(n7618), .A2(n7675), .B1(n7617), .B2(n7673), .ZN(n7622)
         );
  AOI22_X1 U8131 ( .A1(n7680), .A2(n7620), .B1(n7619), .B2(n7677), .ZN(n7621)
         );
  OAI211_X1 U8132 ( .C1(n7684), .C2(n7623), .A(n7622), .B(n7621), .ZN(U3025)
         );
  AOI22_X1 U8133 ( .A1(n7632), .A2(n7639), .B1(n7633), .B2(n7638), .ZN(n7625)
         );
  AOI22_X1 U8134 ( .A1(n7641), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n7634), 
        .B2(n7640), .ZN(n7624) );
  OAI211_X1 U8135 ( .C1(n7644), .C2(n7637), .A(n7625), .B(n7624), .ZN(U3114)
         );
  AOI22_X1 U8136 ( .A1(n7632), .A2(n7646), .B1(n7633), .B2(n7647), .ZN(n7627)
         );
  AOI22_X1 U8137 ( .A1(n7648), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n7634), 
        .B2(n7645), .ZN(n7626) );
  OAI211_X1 U8138 ( .C1(n7651), .C2(n7637), .A(n7627), .B(n7626), .ZN(U3082)
         );
  AOI22_X1 U8139 ( .A1(n7632), .A2(n7653), .B1(n7634), .B2(n7652), .ZN(n7629)
         );
  AOI22_X1 U8140 ( .A1(n7655), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n7633), 
        .B2(n7654), .ZN(n7628) );
  OAI211_X1 U8141 ( .C1(n7658), .C2(n7637), .A(n7629), .B(n7628), .ZN(U3066)
         );
  AOI22_X1 U8142 ( .A1(n7632), .A2(n7660), .B1(n7633), .B2(n7661), .ZN(n7631)
         );
  AOI22_X1 U8143 ( .A1(n7662), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n7634), 
        .B2(n7659), .ZN(n7630) );
  OAI211_X1 U8144 ( .C1(n7665), .C2(n7637), .A(n7631), .B(n7630), .ZN(U3050)
         );
  AOI22_X1 U8145 ( .A1(n7667), .A2(n7633), .B1(n7632), .B2(n7666), .ZN(n7636)
         );
  AOI22_X1 U8146 ( .A1(n7668), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n7634), 
        .B2(n7680), .ZN(n7635) );
  OAI211_X1 U8147 ( .C1(n7672), .C2(n7637), .A(n7636), .B(n7635), .ZN(U3034)
         );
  AOI22_X1 U8148 ( .A1(n7674), .A2(n7639), .B1(n7679), .B2(n7638), .ZN(n7643)
         );
  AOI22_X1 U8149 ( .A1(n7641), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n7678), 
        .B2(n7640), .ZN(n7642) );
  OAI211_X1 U8150 ( .C1(n7644), .C2(n7671), .A(n7643), .B(n7642), .ZN(U3115)
         );
  AOI22_X1 U8151 ( .A1(n7674), .A2(n7646), .B1(n7678), .B2(n7645), .ZN(n7650)
         );
  AOI22_X1 U8152 ( .A1(n7648), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n7679), 
        .B2(n7647), .ZN(n7649) );
  OAI211_X1 U8153 ( .C1(n7651), .C2(n7671), .A(n7650), .B(n7649), .ZN(U3083)
         );
  AOI22_X1 U8154 ( .A1(n7674), .A2(n7653), .B1(n7678), .B2(n7652), .ZN(n7657)
         );
  AOI22_X1 U8155 ( .A1(n7655), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n7679), 
        .B2(n7654), .ZN(n7656) );
  OAI211_X1 U8156 ( .C1(n7658), .C2(n7671), .A(n7657), .B(n7656), .ZN(U3067)
         );
  AOI22_X1 U8157 ( .A1(n7674), .A2(n7660), .B1(n7678), .B2(n7659), .ZN(n7664)
         );
  AOI22_X1 U8158 ( .A1(n7662), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n7679), 
        .B2(n7661), .ZN(n7663) );
  OAI211_X1 U8159 ( .C1(n7665), .C2(n7671), .A(n7664), .B(n7663), .ZN(U3051)
         );
  AOI22_X1 U8160 ( .A1(n7667), .A2(n7679), .B1(n7674), .B2(n7666), .ZN(n7670)
         );
  AOI22_X1 U8161 ( .A1(n7668), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n7678), 
        .B2(n7680), .ZN(n7669) );
  OAI211_X1 U8162 ( .C1(n7672), .C2(n7671), .A(n7670), .B(n7669), .ZN(U3035)
         );
  AOI22_X1 U8163 ( .A1(n7676), .A2(n7675), .B1(n7674), .B2(n7673), .ZN(n7682)
         );
  AOI22_X1 U8164 ( .A1(n7680), .A2(n7679), .B1(n7678), .B2(n7677), .ZN(n7681)
         );
  OAI211_X1 U8165 ( .C1(n7684), .C2(n7683), .A(n7682), .B(n7681), .ZN(U3027)
         );
  INV_X1 U3863 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3757) );
  CLKBUF_X2 U3699 ( .A(n4651), .Z(n3679) );
  CLKBUF_X1 U3704 ( .A(n4369), .Z(n3671) );
  CLKBUF_X1 U3727 ( .A(n3993), .Z(n3994) );
  CLKBUF_X1 U3731 ( .A(n6569), .Z(n6570) );
  NAND2_X1 U3734 ( .A1(n4719), .A2(n4718), .ZN(n6549) );
  CLKBUF_X1 U3736 ( .A(n6960), .Z(n3648) );
  CLKBUF_X1 U3737 ( .A(n5057), .Z(n5099) );
  XNOR2_X1 U3775 ( .A(n4724), .B(n5348), .ZN(n5335) );
  OR2_X1 U3834 ( .A1(n5814), .A2(n7345), .ZN(n4749) );
  CLKBUF_X1 U3837 ( .A(n5524), .Z(n3662) );
endmodule

