

module b20_C_gen_AntiSAT_k_128_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4349, n4350, n4351, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282;

  OR2_X1 U4855 ( .A1(n9269), .A2(n4487), .ZN(n4486) );
  INV_X2 U4856 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X2 U4857 ( .A(n5038), .ZN(n5188) );
  INV_X1 U4858 ( .A(n5994), .ZN(n6189) );
  INV_X1 U4859 ( .A(n5086), .ZN(n5774) );
  NAND2_X1 U4860 ( .A1(n5904), .A2(n7856), .ZN(n5052) );
  INV_X1 U4861 ( .A(n6263), .ZN(n6096) );
  INV_X1 U4862 ( .A(n5993), .ZN(n8544) );
  OAI21_X1 U4863 ( .B1(n6185), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6187) );
  INV_X1 U4864 ( .A(n5627), .ZN(n8035) );
  NAND2_X2 U4865 ( .A1(n4651), .A2(n4650), .ZN(n5716) );
  OAI21_X1 U4866 ( .B1(n8504), .B2(n8420), .A(n8505), .ZN(n8346) );
  AOI21_X1 U4867 ( .B1(n7838), .B2(n6419), .A(n4945), .ZN(n7895) );
  AOI22_X1 U4868 ( .A1(n7226), .A2(n7227), .B1(n6411), .B2(n7192), .ZN(n7273)
         );
  OAI21_X1 U4869 ( .B1(n7999), .B2(n8678), .A(n7997), .ZN(n9016) );
  AND4_X1 U4870 ( .A1(n5076), .A2(n5075), .A3(n5074), .A4(n5073), .ZN(n6750)
         );
  AOI21_X2 U4871 ( .B1(n8761), .B2(n8760), .A(n8759), .ZN(n8763) );
  XNOR2_X2 U4872 ( .A(n5025), .B(n5024), .ZN(n5028) );
  OAI21_X2 U4873 ( .B1(n4583), .B2(n4374), .A(n4580), .ZN(n7999) );
  NAND2_X4 U4874 ( .A1(n6400), .A2(n6399), .ZN(n6404) );
  NAND2_X1 U4875 ( .A1(n4651), .A2(n4650), .ZN(n4349) );
  NAND2_X1 U4876 ( .A1(n4651), .A2(n4650), .ZN(n4350) );
  INV_X1 U4877 ( .A(n5716), .ZN(n5206) );
  NOR2_X2 U4878 ( .A1(n6200), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6209) );
  NAND2_X2 U4879 ( .A1(n8806), .A2(n6334), .ZN(n5994) );
  OR2_X1 U4880 ( .A1(n9520), .A2(n9519), .ZN(n9522) );
  INV_X1 U4881 ( .A(n6300), .ZN(n10130) );
  NOR2_X1 U4882 ( .A1(n9302), .A2(n7252), .ZN(n6710) );
  INV_X1 U4883 ( .A(n10156), .ZN(n6406) );
  INV_X4 U4884 ( .A(n4354), .ZN(n8747) );
  OAI21_X1 U4885 ( .B1(n5289), .B2(n4961), .A(n5288), .ZN(n5313) );
  INV_X1 U4886 ( .A(n6012), .ZN(n6167) );
  INV_X8 U4887 ( .A(n5061), .ZN(n4351) );
  NAND2_X2 U4888 ( .A1(n5052), .A2(n4349), .ZN(n5110) );
  CLKBUF_X3 U4889 ( .A(n5097), .Z(n5907) );
  NAND3_X2 U4890 ( .A1(n5779), .A2(n5781), .A3(n7552), .ZN(n5036) );
  NOR2_X1 U4891 ( .A1(n6148), .A2(n6147), .ZN(n6159) );
  XNOR2_X1 U4892 ( .A(n4982), .B(n4983), .ZN(n5818) );
  INV_X1 U4893 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9166) );
  INV_X4 U4894 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AOI21_X1 U4895 ( .B1(n6522), .B2(n4963), .A(n6521), .ZN(n6523) );
  AND2_X1 U4896 ( .A1(n8347), .A2(n8348), .ZN(n6491) );
  MUX2_X1 U4897 ( .A(n8757), .B(n8756), .S(n8755), .Z(n8760) );
  OAI21_X1 U4898 ( .B1(n8554), .B2(n8549), .A(n8553), .ZN(n8761) );
  NAND2_X1 U4899 ( .A1(n4637), .A2(n4634), .ZN(n8751) );
  AND2_X1 U4900 ( .A1(n4877), .A2(n4876), .ZN(n9242) );
  NAND2_X1 U4901 ( .A1(n4473), .A2(n4472), .ZN(n4471) );
  AOI21_X1 U4902 ( .B1(n4484), .B2(n4384), .A(n4476), .ZN(n5576) );
  XNOR2_X1 U4903 ( .A(n8019), .B(SI_29_), .ZN(n8014) );
  OR2_X1 U4904 ( .A1(n8729), .A2(n8730), .ZN(n8881) );
  OR2_X1 U4905 ( .A1(n9095), .A2(n8509), .ZN(n8555) );
  OR2_X1 U4906 ( .A1(n7861), .A2(n5516), .ZN(n4484) );
  NAND2_X1 U4907 ( .A1(n5745), .A2(n5744), .ZN(n9486) );
  XNOR2_X1 U4908 ( .A(n8021), .B(n8020), .ZN(n8019) );
  AND2_X1 U4909 ( .A1(n5770), .A2(n5769), .ZN(n9496) );
  AOI21_X1 U4910 ( .B1(n9160), .B2(n9009), .A(n6319), .ZN(n9006) );
  NAND2_X1 U4911 ( .A1(n6727), .A2(n5137), .ZN(n6720) );
  INV_X1 U4912 ( .A(n8895), .ZN(n8420) );
  NAND2_X1 U4913 ( .A1(n7186), .A2(n6409), .ZN(n7226) );
  NAND2_X1 U4914 ( .A1(n6268), .A2(n6267), .ZN(n8883) );
  NAND3_X1 U4915 ( .A1(n4696), .A2(n7187), .A3(n4355), .ZN(n7186) );
  AND3_X1 U4916 ( .A1(n6248), .A2(n6247), .A3(n6246), .ZN(n8773) );
  AND2_X1 U4917 ( .A1(n6960), .A2(n9976), .ZN(n6959) );
  NAND2_X1 U4918 ( .A1(n5367), .A2(n5366), .ZN(n7380) );
  AOI21_X1 U4919 ( .B1(n7214), .B2(n4771), .A(n4770), .ZN(n4769) );
  AND2_X1 U4920 ( .A1(n6251), .A2(n8510), .ZN(n6261) );
  NAND2_X2 U4921 ( .A1(n7692), .A2(n6817), .ZN(n9629) );
  NAND2_X1 U4922 ( .A1(n4826), .A2(n4828), .ZN(n5467) );
  AND4_X1 U4923 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n8975)
         );
  NOR2_X2 U4924 ( .A1(n6913), .A2(n6786), .ZN(n6939) );
  NAND2_X1 U4925 ( .A1(n5240), .A2(n5239), .ZN(n9968) );
  INV_X1 U4926 ( .A(n6902), .ZN(n6904) );
  NAND2_X1 U4927 ( .A1(n6333), .A2(n8550), .ZN(n10134) );
  NAND2_X1 U4928 ( .A1(n4673), .A2(n4672), .ZN(n5348) );
  NAND2_X1 U4929 ( .A1(n8822), .A2(n8755), .ZN(n6399) );
  AND2_X2 U4930 ( .A1(n7355), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3893) );
  AND4_X1 U4932 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n6300)
         );
  INV_X1 U4933 ( .A(n6754), .ZN(n6837) );
  OAI211_X1 U4934 ( .C1(n6563), .C2(n7348), .A(n6010), .B(n6009), .ZN(n10156)
         );
  NAND4_X1 U4935 ( .A1(n5984), .A2(n5983), .A3(n5982), .A4(n5981), .ZN(n8783)
         );
  NAND3_X2 U4936 ( .A1(n5880), .A2(n5036), .A3(n5034), .ZN(n5038) );
  NAND4_X1 U4937 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n8782)
         );
  AND4_X1 U4938 ( .A1(n5263), .A2(n5262), .A3(n5261), .A4(n5260), .ZN(n6881)
         );
  NAND2_X1 U4939 ( .A1(n8767), .A2(n8592), .ZN(n4354) );
  OR2_X1 U4940 ( .A1(n5230), .A2(n5229), .ZN(n5289) );
  AND3_X1 U4941 ( .A1(n5085), .A2(n5084), .A3(n4951), .ZN(n6735) );
  NAND2_X1 U4942 ( .A1(n5555), .A2(n8326), .ZN(n5880) );
  AND3_X2 U4943 ( .A1(n5014), .A2(n5013), .A3(n5012), .ZN(n5835) );
  AND2_X2 U4944 ( .A1(n8358), .A2(n5975), .ZN(n6012) );
  AND2_X2 U4945 ( .A1(n9176), .A2(n8358), .ZN(n4958) );
  AND2_X2 U4946 ( .A1(n5974), .A2(n5975), .ZN(n6263) );
  NAND2_X1 U4947 ( .A1(n6163), .A2(n6162), .ZN(n6185) );
  AND2_X1 U4948 ( .A1(n6350), .A2(n6349), .ZN(n6351) );
  INV_X1 U4949 ( .A(n8539), .ZN(n6281) );
  AND2_X1 U4950 ( .A1(n6294), .A2(n4370), .ZN(n8592) );
  AND2_X1 U4951 ( .A1(n6159), .A2(n6158), .ZN(n6163) );
  NAND2_X2 U4952 ( .A1(n5052), .A2(n4840), .ZN(n8173) );
  XNOR2_X1 U4953 ( .A(n6290), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8767) );
  AND2_X2 U4954 ( .A1(n9176), .A2(n5974), .ZN(n8539) );
  XNOR2_X1 U4955 ( .A(n5973), .B(n5968), .ZN(n9176) );
  AND2_X1 U4956 ( .A1(n4993), .A2(n4992), .ZN(n5781) );
  NAND2_X1 U4957 ( .A1(n5966), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5967) );
  XNOR2_X1 U4958 ( .A(n5962), .B(n5963), .ZN(n8806) );
  NAND2_X1 U4959 ( .A1(n5023), .A2(n9778), .ZN(n8344) );
  OR2_X1 U4960 ( .A1(n6291), .A2(n9166), .ZN(n4713) );
  XNOR2_X1 U4961 ( .A(n5016), .B(n5005), .ZN(n7856) );
  INV_X2 U4962 ( .A(n9780), .ZN(n8017) );
  AND2_X1 U4963 ( .A1(n6288), .A2(n6286), .ZN(n6291) );
  OAI21_X1 U4964 ( .B1(n5025), .B2(n5019), .A(n5018), .ZN(n5023) );
  AND2_X1 U4965 ( .A1(n6028), .A2(n4564), .ZN(n6101) );
  XNOR2_X1 U4966 ( .A(n4985), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8264) );
  XNOR2_X1 U4967 ( .A(n5217), .B(SI_7_), .ZN(n5264) );
  NAND2_X1 U4968 ( .A1(n4840), .A2(P1_U3086), .ZN(n9775) );
  NOR2_X1 U4969 ( .A1(n4725), .A2(n4723), .ZN(n4564) );
  AND2_X1 U4970 ( .A1(n4368), .A2(n5004), .ZN(n4900) );
  AND4_X1 U4971 ( .A1(n5317), .A2(n4871), .A3(n4965), .A4(n4976), .ZN(n4358)
         );
  NAND3_X1 U4972 ( .A1(n4490), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4650) );
  INV_X1 U4973 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4965) );
  INV_X1 U4974 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4871) );
  INV_X1 U4975 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4492) );
  NOR2_X2 U4976 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6035) );
  AND2_X1 U4977 ( .A1(n6491), .A2(n8346), .ZN(n8354) );
  XNOR2_X1 U4979 ( .A(n6187), .B(n6186), .ZN(n8822) );
  XNOR2_X2 U4980 ( .A(n4999), .B(n5001), .ZN(n5904) );
  NAND2_X2 U4981 ( .A1(n6257), .A2(n6256), .ZN(n8895) );
  OR2_X1 U4982 ( .A1(n8689), .A2(n4644), .ZN(n8695) );
  NAND2_X1 U4983 ( .A1(n4919), .A2(n4388), .ZN(n4644) );
  NAND2_X1 U4984 ( .A1(n8737), .A2(n8738), .ZN(n4637) );
  NAND2_X1 U4985 ( .A1(n10111), .A2(n4531), .ZN(n8808) );
  NAND2_X1 U4986 ( .A1(n8805), .A2(n10108), .ZN(n4531) );
  OR2_X1 U4987 ( .A1(n6536), .A2(n8772), .ZN(n8746) );
  INV_X1 U4988 ( .A(n4883), .ZN(n4882) );
  OAI21_X1 U4989 ( .B1(n4885), .B2(n4884), .A(n5867), .ZN(n4883) );
  NAND2_X1 U4990 ( .A1(n4676), .A2(n4675), .ZN(n5554) );
  INV_X1 U4991 ( .A(n5525), .ZN(n4675) );
  INV_X1 U4992 ( .A(n5526), .ZN(n4676) );
  OAI21_X1 U4993 ( .B1(n9503), .B2(n4896), .A(n4894), .ZN(n5932) );
  NAND2_X1 U4994 ( .A1(n4376), .A2(n4895), .ZN(n4894) );
  NAND2_X1 U4995 ( .A1(n4376), .A2(n4897), .ZN(n4896) );
  NAND2_X1 U4996 ( .A1(n4796), .A2(n5869), .ZN(n4895) );
  NAND2_X1 U4997 ( .A1(n4467), .A2(n5859), .ZN(n9588) );
  NOR2_X1 U4998 ( .A1(n5858), .A2(n4469), .ZN(n4468) );
  AND2_X1 U4999 ( .A1(n4900), .A2(n4899), .ZN(n4898) );
  INV_X1 U5000 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4899) );
  OAI21_X1 U5001 ( .B1(n8695), .B2(n8694), .A(n8693), .ZN(n4643) );
  NOR2_X1 U5002 ( .A1(n4504), .A2(n4509), .ZN(n4503) );
  NAND2_X1 U5003 ( .A1(n8284), .A2(n8116), .ZN(n4509) );
  NOR2_X1 U5004 ( .A1(n4505), .A2(n4508), .ZN(n4504) );
  NOR2_X1 U5005 ( .A1(n4366), .A2(n4771), .ZN(n4508) );
  AND2_X1 U5006 ( .A1(n8138), .A2(n9545), .ZN(n4520) );
  OR2_X1 U5007 ( .A1(n5440), .A2(SI_13_), .ZN(n5441) );
  NAND2_X1 U5008 ( .A1(n8397), .A2(n8399), .ZN(n6451) );
  NAND2_X1 U5009 ( .A1(n8402), .A2(n6455), .ZN(n4707) );
  INV_X1 U5010 ( .A(n8113), .ZN(n4798) );
  INV_X1 U5011 ( .A(n5435), .ZN(n5444) );
  OR2_X1 U5012 ( .A1(n5226), .A2(n5264), .ZN(n5225) );
  OR2_X1 U5013 ( .A1(n6451), .A2(n8395), .ZN(n6460) );
  NAND2_X1 U5014 ( .A1(n6469), .A2(n6468), .ZN(n4654) );
  AND2_X1 U5015 ( .A1(n4704), .A2(n4706), .ZN(n6469) );
  NOR2_X1 U5016 ( .A1(n7506), .A2(n4720), .ZN(n4719) );
  INV_X1 U5017 ( .A(n4962), .ZN(n4720) );
  INV_X1 U5018 ( .A(n9176), .ZN(n5975) );
  INV_X1 U5019 ( .A(n8811), .ZN(n8799) );
  OR2_X1 U5020 ( .A1(n10067), .A2(n4732), .ZN(n4731) );
  NOR2_X1 U5021 ( .A1(n10058), .A2(n8009), .ZN(n4732) );
  OR2_X1 U5022 ( .A1(n8779), .A2(n10187), .ZN(n8641) );
  OR2_X1 U5023 ( .A1(n7961), .A2(n10201), .ZN(n8655) );
  AOI21_X1 U5024 ( .B1(n8725), .B2(n6327), .A(n4403), .ZN(n4932) );
  NOR2_X1 U5025 ( .A1(n4905), .A2(n4391), .ZN(n4904) );
  NOR2_X1 U5026 ( .A1(n4906), .A2(n8931), .ZN(n4905) );
  AND4_X1 U5027 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n6344), .ZN(n5964)
         );
  NAND3_X1 U5028 ( .A1(n4493), .A2(n4492), .A3(n4491), .ZN(n4651) );
  INV_X1 U5029 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4491) );
  NAND2_X1 U5030 ( .A1(n4724), .A2(n6029), .ZN(n4723) );
  INV_X1 U5031 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4724) );
  AND2_X1 U5032 ( .A1(n4359), .A2(n4562), .ZN(n4941) );
  AND2_X1 U5033 ( .A1(n5957), .A2(n5958), .ZN(n4562) );
  INV_X1 U5034 ( .A(n9197), .ZN(n4472) );
  INV_X1 U5035 ( .A(n9196), .ZN(n4473) );
  NOR2_X1 U5036 ( .A1(n5883), .A2(n8151), .ZN(n4751) );
  NAND2_X1 U5037 ( .A1(n4838), .A2(n4836), .ZN(n8167) );
  AND2_X1 U5038 ( .A1(n4837), .A2(n5878), .ZN(n4836) );
  AOI21_X1 U5039 ( .B1(n4793), .B2(n4796), .A(n8206), .ZN(n4792) );
  INV_X1 U5040 ( .A(n5853), .ZN(n4680) );
  NAND2_X1 U5041 ( .A1(n4808), .A2(n5692), .ZN(n5710) );
  NAND2_X1 U5042 ( .A1(n5689), .A2(n5688), .ZN(n4808) );
  INV_X1 U5043 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4901) );
  AOI21_X1 U5044 ( .B1(n4668), .B2(n4670), .A(n4434), .ZN(n4667) );
  INV_X1 U5045 ( .A(n5447), .ZN(n4668) );
  INV_X1 U5046 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4870) );
  INV_X1 U5047 ( .A(n4958), .ZN(n6280) );
  AOI22_X1 U5048 ( .A1(n8753), .A2(n8754), .B1(n4636), .B2(n4633), .ZN(n8756)
         );
  NAND2_X1 U5049 ( .A1(n8751), .A2(n8752), .ZN(n4633) );
  NOR2_X1 U5050 ( .A1(n8749), .A2(n8750), .ZN(n4636) );
  NAND2_X1 U5051 ( .A1(n4729), .A2(n4728), .ZN(n7791) );
  NAND2_X1 U5052 ( .A1(n10033), .A2(n4390), .ZN(n4728) );
  INV_X1 U5053 ( .A(n8808), .ZN(n8810) );
  INV_X1 U5054 ( .A(n9000), .ZN(n8973) );
  NAND2_X1 U5055 ( .A1(n6082), .A2(n6081), .ZN(n7696) );
  NAND2_X1 U5056 ( .A1(n5994), .A2(n4840), .ZN(n5993) );
  OAI21_X1 U5057 ( .B1(n8872), .B2(n6329), .A(n6328), .ZN(n8859) );
  NAND2_X1 U5058 ( .A1(n4909), .A2(n4907), .ZN(n8961) );
  OAI21_X1 U5059 ( .B1(n4912), .B2(n4398), .A(n4908), .ZN(n4907) );
  INV_X1 U5060 ( .A(n6008), .ZN(n6188) );
  XNOR2_X1 U5061 ( .A(n8663), .B(n8662), .ZN(n8660) );
  AND2_X1 U5062 ( .A1(n6018), .A2(n5951), .ZN(n4565) );
  NAND2_X1 U5063 ( .A1(n5196), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5256) );
  INV_X1 U5064 ( .A(n5198), .ZN(n5196) );
  AND2_X1 U5065 ( .A1(n5141), .A2(n4850), .ZN(n4847) );
  AND2_X1 U5066 ( .A1(n5059), .A2(n4959), .ZN(n5060) );
  AND2_X1 U5067 ( .A1(n4420), .A2(n4861), .ZN(n4858) );
  INV_X1 U5068 ( .A(n5094), .ZN(n5627) );
  NOR2_X1 U5069 ( .A1(n4886), .A2(n5866), .ZN(n4885) );
  INV_X1 U5070 ( .A(n5863), .ZN(n4886) );
  AOI21_X1 U5071 ( .B1(n9591), .B2(n4777), .A(n4776), .ZN(n4775) );
  INV_X1 U5072 ( .A(n8058), .ZN(n4777) );
  INV_X1 U5073 ( .A(n8131), .ZN(n4776) );
  INV_X1 U5074 ( .A(n9591), .ZN(n4778) );
  NOR2_X1 U5075 ( .A1(n5857), .A2(n4893), .ZN(n4892) );
  INV_X1 U5076 ( .A(n5856), .ZN(n4893) );
  NAND2_X1 U5077 ( .A1(n4768), .A2(n4393), .ZN(n7280) );
  NAND2_X1 U5078 ( .A1(n6950), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U5079 ( .A1(n4769), .A2(n8230), .ZN(n4767) );
  INV_X1 U5080 ( .A(n8173), .ZN(n5557) );
  INV_X1 U5081 ( .A(n6611), .ZN(n5556) );
  NAND2_X1 U5083 ( .A1(n4821), .A2(n4820), .ZN(n5873) );
  AOI21_X1 U5084 ( .B1(n4364), .B2(n4825), .A(n4446), .ZN(n4820) );
  NAND2_X1 U5085 ( .A1(n5740), .A2(n4364), .ZN(n4821) );
  NOR3_X1 U5086 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_IR_REG_18__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U5087 ( .A1(n4674), .A2(n5582), .ZN(n5598) );
  NAND2_X1 U5088 ( .A1(n5554), .A2(n4839), .ZN(n4674) );
  XNOR2_X1 U5089 ( .A(n4975), .B(n4974), .ZN(n5555) );
  NAND2_X1 U5090 ( .A1(n5531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U5091 ( .A1(n5224), .A2(n4783), .ZN(n4782) );
  INV_X1 U5092 ( .A(n5224), .ZN(n4784) );
  XNOR2_X1 U5093 ( .A(n5152), .B(n5129), .ZN(n5151) );
  CLKBUF_X1 U5094 ( .A(n5206), .Z(n4840) );
  OAI21_X1 U5095 ( .B1(n6525), .B2(n7622), .A(n6343), .ZN(n6527) );
  INV_X1 U5096 ( .A(n4486), .ZN(n6553) );
  AOI211_X1 U5097 ( .C1(n9461), .C2(n9286), .A(n8183), .B(n8177), .ZN(n8182)
         );
  OR2_X1 U5098 ( .A1(n5933), .A2(n5932), .ZN(n8343) );
  NAND2_X1 U5099 ( .A1(n5052), .A2(n4878), .ZN(n5014) );
  OAI21_X1 U5100 ( .B1(n8672), .B2(n4937), .A(n8671), .ZN(n8673) );
  OAI21_X1 U5101 ( .B1(n8085), .B2(n4489), .A(n8176), .ZN(n4488) );
  INV_X1 U5102 ( .A(n4506), .ZN(n4505) );
  AOI21_X1 U5103 ( .B1(n8115), .B2(n4507), .A(n8103), .ZN(n4506) );
  INV_X1 U5104 ( .A(n8102), .ZN(n4507) );
  INV_X1 U5105 ( .A(n8119), .ZN(n4502) );
  NAND2_X1 U5106 ( .A1(n8696), .A2(n4354), .ZN(n4645) );
  NAND2_X1 U5107 ( .A1(n4642), .A2(n8747), .ZN(n4641) );
  INV_X1 U5108 ( .A(n4799), .ZN(n8229) );
  AOI21_X1 U5109 ( .B1(n4520), .B2(n8139), .A(n4518), .ZN(n4517) );
  INV_X1 U5110 ( .A(n8140), .ZN(n4518) );
  NOR2_X1 U5111 ( .A1(n4519), .A2(n4774), .ZN(n4516) );
  INV_X1 U5112 ( .A(n4520), .ZN(n4519) );
  NOR2_X1 U5113 ( .A1(n6311), .A2(n6310), .ZN(n6314) );
  AND2_X1 U5114 ( .A1(n7543), .A2(n4856), .ZN(n4855) );
  OR2_X1 U5115 ( .A1(n7375), .A2(n4857), .ZN(n4856) );
  INV_X1 U5116 ( .A(n5383), .ZN(n4857) );
  AND2_X1 U5117 ( .A1(n4766), .A2(n4765), .ZN(n4764) );
  AOI21_X1 U5118 ( .B1(n4667), .B2(n4669), .A(n4665), .ZN(n4664) );
  INV_X1 U5119 ( .A(n5517), .ZN(n4665) );
  INV_X1 U5120 ( .A(n5495), .ZN(n5496) );
  INV_X1 U5121 ( .A(n5441), .ZN(n4831) );
  AND2_X1 U5122 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  NOR2_X1 U5123 ( .A1(n5441), .A2(n5403), .ZN(n4832) );
  AND2_X1 U5124 ( .A1(n5437), .A2(n4834), .ZN(n4833) );
  INV_X1 U5125 ( .A(n5403), .ZN(n4830) );
  NAND2_X1 U5126 ( .A1(n5353), .A2(SI_12_), .ZN(n5437) );
  INV_X1 U5127 ( .A(SI_8_), .ZN(n7028) );
  INV_X1 U5128 ( .A(n6424), .ZN(n4701) );
  NAND2_X1 U5129 ( .A1(n4409), .A2(n8400), .ZN(n6456) );
  INV_X1 U5130 ( .A(n4662), .ZN(n4661) );
  AOI21_X1 U5131 ( .B1(n6199), .B2(n6198), .A(n6405), .ZN(n4662) );
  NAND2_X1 U5132 ( .A1(n6199), .A2(n4659), .ZN(n4658) );
  NOR2_X1 U5133 ( .A1(n6404), .A2(n4660), .ZN(n4659) );
  INV_X1 U5134 ( .A(n6198), .ZN(n4660) );
  NOR2_X1 U5135 ( .A1(n4705), .A2(n4943), .ZN(n4704) );
  NOR2_X1 U5136 ( .A1(n8438), .A2(n4707), .ZN(n4705) );
  NAND2_X1 U5137 ( .A1(n8738), .A2(n4635), .ZN(n4634) );
  INV_X1 U5138 ( .A(n8740), .ZN(n4635) );
  OR2_X1 U5139 ( .A1(n7426), .A2(n10015), .ZN(n7427) );
  INV_X1 U5140 ( .A(n10037), .ZN(n4556) );
  NAND2_X1 U5141 ( .A1(n4539), .A2(n4538), .ZN(n4537) );
  INV_X1 U5142 ( .A(n4449), .ZN(n4538) );
  INV_X1 U5143 ( .A(n4541), .ZN(n4539) );
  OAI21_X1 U5144 ( .B1(n10090), .B2(n9071), .A(n10091), .ZN(n8837) );
  AOI21_X1 U5145 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8824), .A(n10099), .ZN(
        n8792) );
  AND2_X1 U5146 ( .A1(n4938), .A2(n4937), .ZN(n4936) );
  OR2_X1 U5147 ( .A1(n4939), .A2(n4357), .ZN(n4938) );
  OR2_X1 U5148 ( .A1(n8635), .A2(n6314), .ZN(n7698) );
  OR2_X1 U5149 ( .A1(n8779), .A2(n7904), .ZN(n7701) );
  XNOR2_X1 U5150 ( .A(n9089), .B(n8591), .ZN(n8585) );
  AND2_X1 U5151 ( .A1(n9095), .A2(n8509), .ZN(n8733) );
  NOR2_X1 U5152 ( .A1(n9101), .A2(n8420), .ZN(n8729) );
  INV_X1 U5153 ( .A(n4594), .ZN(n4590) );
  OR2_X1 U5154 ( .A1(n9107), .A2(n8773), .ZN(n8727) );
  OR2_X1 U5155 ( .A1(n8926), .A2(n8488), .ZN(n8719) );
  OR2_X1 U5156 ( .A1(n9126), .A2(n6443), .ZN(n8711) );
  INV_X1 U5157 ( .A(n4576), .ZN(n4569) );
  NAND2_X1 U5158 ( .A1(n8559), .A2(n4578), .ZN(n4576) );
  INV_X1 U5159 ( .A(n8688), .ZN(n4579) );
  OAI21_X1 U5160 ( .B1(n8683), .B2(n4579), .A(n6320), .ZN(n4577) );
  AND2_X1 U5161 ( .A1(n8660), .A2(n4377), .ZN(n4939) );
  NAND2_X1 U5162 ( .A1(n7716), .A2(n6317), .ZN(n4940) );
  AND2_X1 U5163 ( .A1(n6289), .A2(n6344), .ZN(n4714) );
  INV_X1 U5164 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4490) );
  NAND2_X1 U5165 ( .A1(n4726), .A2(n4394), .ZN(n4725) );
  INV_X1 U5166 ( .A(n4924), .ZN(n4726) );
  NAND2_X1 U5167 ( .A1(n5952), .A2(n6043), .ZN(n4924) );
  INV_X1 U5168 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5952) );
  INV_X1 U5169 ( .A(n9203), .ZN(n4865) );
  NAND2_X1 U5170 ( .A1(n5796), .A2(n6805), .ZN(n4987) );
  NAND2_X1 U5171 ( .A1(n4485), .A2(n8254), .ZN(n8176) );
  NAND2_X1 U5172 ( .A1(n5555), .A2(n5818), .ZN(n5796) );
  OR2_X1 U5173 ( .A1(n9486), .A2(n9280), .ZN(n8303) );
  NOR2_X1 U5174 ( .A1(n9529), .A2(n9676), .ZN(n4757) );
  NOR2_X1 U5175 ( .A1(n9709), .A2(n7866), .ZN(n4762) );
  AND2_X1 U5176 ( .A1(n4804), .A2(n8105), .ZN(n4803) );
  AND2_X1 U5177 ( .A1(n6904), .A2(n9964), .ZN(n4766) );
  INV_X1 U5178 ( .A(n5841), .ZN(n4465) );
  NAND2_X1 U5179 ( .A1(n9299), .A2(n6735), .ZN(n8266) );
  OR2_X1 U5180 ( .A1(n6605), .A2(n5110), .ZN(n4807) );
  NAND2_X1 U5181 ( .A1(n5715), .A2(n5714), .ZN(n5740) );
  NAND2_X1 U5182 ( .A1(n5710), .A2(n5709), .ZN(n5715) );
  NAND2_X1 U5183 ( .A1(n5665), .A2(n5664), .ZN(n5689) );
  AOI21_X1 U5184 ( .B1(n5598), .B2(n4812), .A(n4810), .ZN(n4809) );
  NAND2_X1 U5185 ( .A1(n4811), .A2(n5618), .ZN(n4810) );
  NAND2_X1 U5186 ( .A1(n5439), .A2(n5437), .ZN(n5404) );
  AOI21_X1 U5187 ( .B1(n5352), .B2(n4954), .A(n4949), .ZN(n5357) );
  INV_X1 U5188 ( .A(n5348), .ZN(n5352) );
  NAND2_X1 U5189 ( .A1(n5232), .A2(SI_9_), .ZN(n5288) );
  AND2_X1 U5190 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  INV_X1 U5191 ( .A(n5226), .ZN(n5227) );
  NAND2_X1 U5192 ( .A1(n4703), .A2(n8438), .ZN(n8383) );
  NAND2_X1 U5193 ( .A1(n8425), .A2(n8437), .ZN(n4703) );
  INV_X1 U5194 ( .A(n7201), .ZN(n4695) );
  INV_X1 U5195 ( .A(n7629), .ZN(n4718) );
  XNOR2_X1 U5196 ( .A(n6404), .B(n4927), .ZN(n6401) );
  NOR2_X1 U5197 ( .A1(n8532), .A2(n8531), .ZN(n8554) );
  AND4_X1 U5198 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n8431)
         );
  AND4_X1 U5199 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n8774)
         );
  AND4_X1 U5200 ( .A1(n6132), .A2(n6131), .A3(n6130), .A4(n6129), .ZN(n6433)
         );
  NAND2_X1 U5201 ( .A1(n6012), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U5202 ( .A(n7338), .B(n4734), .ZN(n9989) );
  OR2_X1 U5203 ( .A1(n4598), .A2(n7348), .ZN(n4733) );
  NAND2_X1 U5204 ( .A1(n7496), .A2(n7347), .ZN(n4598) );
  OR2_X1 U5205 ( .A1(n7327), .A2(n7328), .ZN(n4561) );
  AND2_X1 U5206 ( .A1(n4561), .A2(n4560), .ZN(n10005) );
  NAND2_X1 U5207 ( .A1(n7407), .A2(n7413), .ZN(n4560) );
  OR2_X1 U5208 ( .A1(n10005), .A2(n10006), .ZN(n4559) );
  NAND2_X1 U5209 ( .A1(n10021), .A2(n7748), .ZN(n7750) );
  AOI21_X1 U5210 ( .B1(n4553), .B2(n4555), .A(n4551), .ZN(n4550) );
  INV_X1 U5211 ( .A(n7802), .ZN(n4551) );
  NAND2_X1 U5212 ( .A1(n7752), .A2(n7753), .ZN(n7874) );
  INV_X1 U5213 ( .A(n4609), .ZN(n4608) );
  OAI21_X1 U5214 ( .B1(n10028), .B2(n4610), .A(n7749), .ZN(n4609) );
  INV_X1 U5215 ( .A(n7724), .ZN(n4610) );
  OR2_X1 U5216 ( .A1(n7881), .A2(n7882), .ZN(n4606) );
  NOR2_X1 U5217 ( .A1(n4535), .A2(n8800), .ZN(n4534) );
  INV_X1 U5218 ( .A(n10047), .ZN(n4535) );
  OR2_X1 U5219 ( .A1(n7973), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U5220 ( .A1(n4615), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U5221 ( .A1(n8787), .A2(n4615), .ZN(n4611) );
  INV_X1 U5222 ( .A(n10068), .ZN(n4615) );
  OR2_X1 U5223 ( .A1(n10052), .A2(n10051), .ZN(n4614) );
  NAND2_X1 U5224 ( .A1(n10062), .A2(n8802), .ZN(n10078) );
  NAND2_X1 U5225 ( .A1(n10078), .A2(n10079), .ZN(n10077) );
  XNOR2_X1 U5226 ( .A(n8792), .B(n10108), .ZN(n10120) );
  OAI21_X1 U5227 ( .B1(n10120), .B2(n4744), .A(n4743), .ZN(n9794) );
  NAND2_X1 U5228 ( .A1(n4745), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U5229 ( .A1(n8793), .A2(n4745), .ZN(n4743) );
  OR2_X1 U5230 ( .A1(n10120), .A2(n10119), .ZN(n4617) );
  INV_X1 U5231 ( .A(n8931), .ZN(n8939) );
  XNOR2_X1 U5232 ( .A(n8938), .B(n8921), .ZN(n8931) );
  AND2_X1 U5233 ( .A1(n6321), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U5234 ( .A1(n4412), .A2(n4920), .ZN(n4912) );
  NAND2_X1 U5235 ( .A1(n8503), .A2(n8973), .ZN(n4920) );
  INV_X1 U5236 ( .A(n6321), .ZN(n4914) );
  NAND2_X1 U5237 ( .A1(n4928), .A2(n4927), .ZN(n8595) );
  AOI21_X1 U5238 ( .B1(n7696), .B2(n8643), .A(n6093), .ZN(n7719) );
  NAND2_X1 U5239 ( .A1(n8655), .A2(n8656), .ZN(n8575) );
  NOR2_X1 U5240 ( .A1(n8660), .A2(n8657), .ZN(n4584) );
  NAND2_X1 U5241 ( .A1(n6279), .A2(n6278), .ZN(n6536) );
  NAND2_X1 U5242 ( .A1(n8860), .A2(n10131), .ZN(n8862) );
  INV_X1 U5243 ( .A(n8585), .ZN(n8858) );
  AOI21_X1 U5244 ( .B1(n4932), .B2(n4930), .A(n4407), .ZN(n4929) );
  INV_X1 U5245 ( .A(n4932), .ZN(n4931) );
  INV_X1 U5246 ( .A(n6327), .ZN(n4930) );
  OAI21_X1 U5247 ( .B1(n8880), .B2(n8729), .A(n8556), .ZN(n8870) );
  AND2_X1 U5248 ( .A1(n4595), .A2(n8724), .ZN(n4594) );
  NAND2_X1 U5249 ( .A1(n4593), .A2(n8724), .ZN(n4592) );
  INV_X1 U5250 ( .A(n8721), .ZN(n4593) );
  AND2_X1 U5251 ( .A1(n8719), .A2(n8702), .ZN(n4595) );
  NAND2_X1 U5252 ( .A1(n4903), .A2(n4902), .ZN(n8905) );
  AOI21_X1 U5253 ( .B1(n4904), .B2(n4906), .A(n4404), .ZN(n4902) );
  NAND2_X1 U5254 ( .A1(n8930), .A2(n8931), .ZN(n8929) );
  AOI21_X1 U5255 ( .B1(n8968), .B2(n8970), .A(n8698), .ZN(n8958) );
  AND2_X1 U5256 ( .A1(n8697), .A2(n8707), .ZN(n8970) );
  NOR2_X1 U5257 ( .A1(n4415), .A2(n4922), .ZN(n4916) );
  OR2_X1 U5258 ( .A1(n4918), .A2(n4415), .ZN(n4917) );
  AOI21_X1 U5259 ( .B1(n9007), .B2(n4921), .A(n4919), .ZN(n4918) );
  NAND2_X1 U5260 ( .A1(n4577), .A2(n8559), .ZN(n4575) );
  OR2_X1 U5261 ( .A1(n9148), .A2(n8431), .ZN(n8983) );
  NOR2_X1 U5262 ( .A1(n8681), .A2(n4579), .ZN(n4578) );
  INV_X1 U5263 ( .A(n4577), .ZN(n4573) );
  AND2_X1 U5264 ( .A1(n9160), .A2(n8366), .ZN(n8681) );
  INV_X1 U5265 ( .A(n4581), .ZN(n4580) );
  OAI21_X1 U5266 ( .B1(n4582), .B2(n4374), .A(n4586), .ZN(n4581) );
  OR2_X1 U5267 ( .A1(n8479), .A2(n8670), .ZN(n4586) );
  AND2_X1 U5268 ( .A1(n4940), .A2(n4939), .ZN(n7812) );
  INV_X1 U5269 ( .A(n8976), .ZN(n10131) );
  NAND2_X1 U5270 ( .A1(n6104), .A2(n6103), .ZN(n10201) );
  INV_X1 U5271 ( .A(n6080), .ZN(n4638) );
  INV_X1 U5272 ( .A(n6515), .ZN(n6532) );
  AND2_X1 U5273 ( .A1(n6566), .A2(n6764), .ZN(n6686) );
  XNOR2_X1 U5274 ( .A(n5969), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U5275 ( .A1(n9167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U5276 ( .A1(n6346), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6350) );
  INV_X1 U5277 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5951) );
  AND2_X2 U5278 ( .A1(n5986), .A2(n4566), .ZN(n5995) );
  INV_X1 U5279 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4566) );
  OR2_X1 U5280 ( .A1(n5086), .A2(n7252), .ZN(n5064) );
  NAND2_X1 U5281 ( .A1(n6720), .A2(n5141), .ZN(n4851) );
  NAND2_X1 U5282 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5144) );
  NAND2_X1 U5283 ( .A1(n6799), .A2(n6794), .ZN(n7579) );
  INV_X1 U5284 ( .A(n9189), .ZN(n4477) );
  NAND2_X1 U5285 ( .A1(n4482), .A2(n5551), .ZN(n4480) );
  NAND2_X1 U5286 ( .A1(n9189), .A2(n5515), .ZN(n4478) );
  NOR2_X1 U5287 ( .A1(n4482), .A2(n5551), .ZN(n4481) );
  INV_X1 U5288 ( .A(n9243), .ZN(n4876) );
  NAND2_X1 U5289 ( .A1(n4471), .A2(n5615), .ZN(n4470) );
  NAND2_X1 U5290 ( .A1(n5068), .A2(n5067), .ZN(n6692) );
  INV_X1 U5291 ( .A(n5168), .ZN(n5166) );
  NAND2_X1 U5292 ( .A1(n4848), .A2(n4850), .ZN(n4845) );
  INV_X1 U5293 ( .A(n4849), .ZN(n4848) );
  NAND2_X1 U5294 ( .A1(n6766), .A2(n6768), .ZN(n6767) );
  NAND2_X1 U5295 ( .A1(n5419), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5478) );
  INV_X1 U5296 ( .A(n5421), .ZN(n5419) );
  AND2_X1 U5297 ( .A1(n9458), .A2(n8038), .ZN(n8212) );
  AND4_X1 U5298 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n7605)
         );
  NAND2_X1 U5299 ( .A1(n5627), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4466) );
  NAND2_X1 U5300 ( .A1(n5626), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4691) );
  NOR2_X1 U5301 ( .A1(n4787), .A2(n8250), .ZN(n4786) );
  INV_X1 U5302 ( .A(n4793), .ZN(n4787) );
  NAND2_X1 U5303 ( .A1(n4790), .A2(n4789), .ZN(n4788) );
  OR2_X1 U5304 ( .A1(n4792), .A2(n4797), .ZN(n4789) );
  NAND2_X1 U5305 ( .A1(n4792), .A2(n4386), .ZN(n4790) );
  NAND2_X1 U5306 ( .A1(n4792), .A2(n8250), .ZN(n4791) );
  OR2_X1 U5307 ( .A1(n5746), .A2(n6554), .ZN(n9475) );
  AND2_X1 U5308 ( .A1(n4684), .A2(n5869), .ZN(n4683) );
  OR2_X1 U5309 ( .A1(n4378), .A2(n4685), .ZN(n4684) );
  OAI21_X1 U5310 ( .B1(n4455), .B2(n4454), .A(n5868), .ZN(n9503) );
  INV_X1 U5311 ( .A(n4378), .ZN(n4454) );
  AOI21_X1 U5312 ( .B1(n4882), .B2(n4884), .A(n4389), .ZN(n4879) );
  NOR2_X1 U5313 ( .A1(n4944), .A2(n9676), .ZN(n9537) );
  OR2_X1 U5314 ( .A1(n9588), .A2(n4436), .ZN(n5864) );
  AOI21_X1 U5315 ( .B1(n4775), .B2(n4778), .A(n4774), .ZN(n4773) );
  AND2_X1 U5316 ( .A1(n4889), .A2(n4888), .ZN(n4887) );
  OR2_X1 U5317 ( .A1(n9628), .A2(n9610), .ZN(n4888) );
  OR2_X1 U5318 ( .A1(n5857), .A2(n4890), .ZN(n4889) );
  NAND2_X1 U5319 ( .A1(n4375), .A2(n5856), .ZN(n4890) );
  AOI21_X1 U5320 ( .B1(n4459), .B2(n4461), .A(n4411), .ZN(n4456) );
  NOR2_X1 U5321 ( .A1(n7824), .A2(n7866), .ZN(n7930) );
  AND4_X1 U5322 ( .A1(n5395), .A2(n5394), .A3(n5393), .A4(n5392), .ZN(n7559)
         );
  INV_X1 U5323 ( .A(n8116), .ZN(n4770) );
  AND4_X1 U5324 ( .A1(n5305), .A2(n5304), .A3(n5303), .A4(n5302), .ZN(n6952)
         );
  AND2_X1 U5325 ( .A1(n8280), .A2(n8228), .ZN(n5894) );
  OR2_X1 U5326 ( .A1(n5256), .A2(n5255), .ZN(n5258) );
  NOR2_X1 U5327 ( .A1(n4443), .A2(n4950), .ZN(n6781) );
  AND4_X1 U5328 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n6932)
         );
  AND2_X1 U5329 ( .A1(n5902), .A2(n5901), .ZN(n9546) );
  NAND2_X1 U5330 ( .A1(n5645), .A2(n5644), .ZN(n9562) );
  NAND2_X1 U5331 ( .A1(n5415), .A2(n5414), .ZN(n9725) );
  INV_X1 U5332 ( .A(n9546), .ZN(n9640) );
  NAND2_X1 U5333 ( .A1(n8023), .A2(n8022), .ZN(n8171) );
  OR2_X1 U5334 ( .A1(n8021), .A2(n8020), .ZN(n8022) );
  OR2_X1 U5335 ( .A1(n8019), .A2(n8018), .ZN(n8023) );
  INV_X1 U5336 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5017) );
  AND2_X1 U5337 ( .A1(n4679), .A2(n4678), .ZN(n5025) );
  NAND2_X1 U5338 ( .A1(n5236), .A2(n5015), .ZN(n4678) );
  AND2_X1 U5339 ( .A1(n4368), .A2(n5015), .ZN(n4453) );
  XNOR2_X1 U5340 ( .A(n8171), .B(n8170), .ZN(n8533) );
  XNOR2_X1 U5341 ( .A(n5758), .B(n5757), .ZN(n7778) );
  NAND2_X1 U5342 ( .A1(n4822), .A2(n5743), .ZN(n5758) );
  NAND2_X1 U5343 ( .A1(n5740), .A2(n5739), .ZN(n4822) );
  INV_X1 U5344 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4988) );
  XNOR2_X1 U5345 ( .A(n5740), .B(n5739), .ZN(n7762) );
  XNOR2_X1 U5346 ( .A(n5689), .B(n5688), .ZN(n7553) );
  OAI21_X1 U5347 ( .B1(n5598), .B2(n4814), .A(n4813), .ZN(n5619) );
  NAND2_X1 U5348 ( .A1(n5554), .A2(n5553), .ZN(n5577) );
  AND2_X1 U5349 ( .A1(n4379), .A2(n4970), .ZN(n4867) );
  INV_X1 U5350 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U5351 ( .A1(n4663), .A2(n4667), .ZN(n5518) );
  OR2_X1 U5352 ( .A1(n5467), .A2(n4669), .ZN(n4663) );
  NAND2_X1 U5353 ( .A1(n4671), .A2(n5448), .ZN(n5497) );
  NAND2_X1 U5354 ( .A1(n5467), .A2(n5447), .ZN(n4671) );
  INV_X1 U5355 ( .A(n5264), .ZN(n4780) );
  XNOR2_X1 U5356 ( .A(n5205), .B(n5186), .ZN(n5224) );
  NAND2_X1 U5357 ( .A1(n5154), .A2(n5153), .ZN(n5182) );
  XNOR2_X1 U5358 ( .A(n5183), .B(n5155), .ZN(n5181) );
  XNOR2_X1 U5359 ( .A(n5122), .B(n5108), .ZN(n5126) );
  XNOR2_X1 U5360 ( .A(n5107), .B(n5082), .ZN(n5105) );
  XNOR2_X1 U5361 ( .A(n5079), .B(n5007), .ZN(n5078) );
  AND4_X1 U5362 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n7511)
         );
  INV_X1 U5363 ( .A(n8618), .ZN(n7594) );
  XNOR2_X1 U5364 ( .A(n6401), .B(n8783), .ZN(n7206) );
  INV_X1 U5365 ( .A(n8777), .ZN(n7961) );
  INV_X1 U5366 ( .A(n9113), .ZN(n8456) );
  AND4_X1 U5367 ( .A1(n6197), .A2(n6196), .A3(n6195), .A4(n6194), .ZN(n8498)
         );
  NAND2_X1 U5368 ( .A1(n7956), .A2(n6424), .ZN(n8474) );
  INV_X1 U5369 ( .A(n9142), .ZN(n8503) );
  NAND2_X1 U5370 ( .A1(n6359), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5962) );
  INV_X1 U5371 ( .A(n8366), .ZN(n9009) );
  INV_X1 U5372 ( .A(n6433), .ZN(n9019) );
  INV_X1 U5373 ( .A(n8662), .ZN(n8776) );
  INV_X1 U5374 ( .A(n4525), .ZN(n4524) );
  NAND2_X1 U5375 ( .A1(n10010), .A2(n4450), .ZN(n4528) );
  OR2_X1 U5376 ( .A1(n8813), .A2(n8817), .ZN(n4530) );
  AND2_X1 U5377 ( .A1(n8547), .A2(n8546), .ZN(n8852) );
  INV_X1 U5378 ( .A(n9119), .ZN(n8926) );
  OAI211_X1 U5379 ( .C1(n6563), .C2(n7413), .A(n6022), .B(n6021), .ZN(n10139)
         );
  INV_X1 U5380 ( .A(n9086), .ZN(n9029) );
  NAND2_X1 U5381 ( .A1(n6108), .A2(n6107), .ZN(n8663) );
  NOR2_X1 U5382 ( .A1(n6527), .A2(n6526), .ZN(n6548) );
  OR2_X1 U5383 ( .A1(n6549), .A2(n6550), .ZN(n4487) );
  INV_X1 U5384 ( .A(n6625), .ZN(n6785) );
  OAI211_X1 U5385 ( .C1(n4844), .C2(n5434), .A(n4841), .B(n5494), .ZN(n7861)
         );
  NAND2_X1 U5386 ( .A1(n5585), .A2(n5584), .ZN(n9615) );
  AND4_X1 U5387 ( .A1(n5375), .A2(n5374), .A3(n5373), .A4(n5372), .ZN(n7546)
         );
  INV_X1 U5388 ( .A(n9298), .ZN(n6910) );
  AND2_X1 U5389 ( .A1(n5805), .A2(n5803), .ZN(n9274) );
  NAND2_X1 U5390 ( .A1(n5475), .A2(n5474), .ZN(n7947) );
  AND2_X1 U5391 ( .A1(n8256), .A2(n4452), .ZN(n4498) );
  NOR2_X1 U5392 ( .A1(n4361), .A2(n8329), .ZN(n4495) );
  INV_X1 U5393 ( .A(n8258), .ZN(n4818) );
  AND2_X1 U5394 ( .A1(n8212), .A2(n4485), .ZN(n4496) );
  AOI21_X1 U5395 ( .B1(n4817), .B2(n8324), .A(n8323), .ZN(n4816) );
  INV_X1 U5396 ( .A(n9496), .ZN(n6874) );
  OR2_X1 U5397 ( .A1(n5057), .A2(n5056), .ZN(n9302) );
  NAND2_X1 U5398 ( .A1(n5762), .A2(n5761), .ZN(n8151) );
  INV_X1 U5399 ( .A(n6981), .ZN(n6786) );
  INV_X1 U5400 ( .A(n6735), .ZN(n6818) );
  AND2_X1 U5401 ( .A1(n8033), .A2(n8032), .ZN(n9734) );
  OAI21_X1 U5402 ( .B1(n8343), .B2(n9728), .A(n5943), .ZN(n5948) );
  NAND2_X1 U5403 ( .A1(n4998), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4999) );
  OAI211_X1 U5404 ( .C1(n8747), .C2(n4632), .A(n4629), .B(n8661), .ZN(n4628)
         );
  INV_X1 U5405 ( .A(n5893), .ZN(n8096) );
  AOI21_X1 U5406 ( .B1(n4503), .B2(n4505), .A(n4502), .ZN(n4501) );
  AND2_X1 U5407 ( .A1(n8721), .A2(n4418), .ZN(n4624) );
  INV_X1 U5408 ( .A(n4623), .ZN(n4622) );
  OAI21_X1 U5409 ( .B1(n8723), .B2(n8724), .A(n8725), .ZN(n4623) );
  AND2_X1 U5410 ( .A1(n8879), .A2(n8728), .ZN(n4625) );
  NAND2_X1 U5411 ( .A1(n4621), .A2(n4619), .ZN(n8736) );
  AND2_X1 U5412 ( .A1(n4625), .A2(n4620), .ZN(n4619) );
  NAND2_X1 U5413 ( .A1(n4626), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U5414 ( .A1(n4622), .A2(n8723), .ZN(n4620) );
  NOR2_X1 U5415 ( .A1(n5444), .A2(n5443), .ZN(n5440) );
  INV_X1 U5416 ( .A(n6451), .ZN(n6452) );
  AND2_X1 U5417 ( .A1(n8570), .A2(n7616), .ZN(n7615) );
  NAND2_X1 U5418 ( .A1(n10130), .A2(n6406), .ZN(n8612) );
  AND2_X1 U5419 ( .A1(n9062), .A2(n8991), .ZN(n6322) );
  INV_X1 U5420 ( .A(n4516), .ZN(n4512) );
  OR2_X1 U5421 ( .A1(n8136), .A2(n4514), .ZN(n4510) );
  NAND2_X1 U5422 ( .A1(n4515), .A2(n4517), .ZN(n8154) );
  NAND2_X1 U5423 ( .A1(n5893), .A2(n4387), .ZN(n4799) );
  AND2_X1 U5424 ( .A1(n4813), .A2(n4438), .ZN(n4812) );
  NAND2_X1 U5425 ( .A1(n4812), .A2(n4814), .ZN(n4811) );
  AND2_X1 U5426 ( .A1(n5448), .A2(n4437), .ZN(n4670) );
  NOR2_X1 U5427 ( .A1(n4707), .A2(n4708), .ZN(n4702) );
  OR2_X1 U5428 ( .A1(n9029), .A2(n8589), .ZN(n8748) );
  NAND2_X1 U5429 ( .A1(n7415), .A2(n7414), .ZN(n7417) );
  NAND2_X1 U5430 ( .A1(n4742), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U5431 ( .A1(n8833), .A2(n10059), .ZN(n8834) );
  OR2_X1 U5432 ( .A1(n6314), .A2(n6313), .ZN(n7700) );
  NAND2_X1 U5433 ( .A1(n8617), .A2(n8612), .ZN(n8562) );
  OR2_X1 U5434 ( .A1(n6363), .A2(n6377), .ZN(n6486) );
  AND2_X1 U5435 ( .A1(n8557), .A2(n8912), .ZN(n8721) );
  INV_X1 U5436 ( .A(n6325), .ZN(n4906) );
  OR2_X1 U5437 ( .A1(n9132), .A2(n8975), .ZN(n8710) );
  NOR2_X1 U5438 ( .A1(n6322), .A2(n4911), .ZN(n4910) );
  INV_X1 U5439 ( .A(n4915), .ZN(n4911) );
  INV_X1 U5440 ( .A(n6322), .ZN(n4908) );
  AOI21_X1 U5441 ( .B1(n4855), .B2(n4857), .A(n4397), .ZN(n4852) );
  NAND2_X1 U5442 ( .A1(n4484), .A2(n5515), .ZN(n4483) );
  OAI21_X1 U5443 ( .B1(n5141), .B2(n4850), .A(n6569), .ZN(n4849) );
  INV_X1 U5444 ( .A(n8212), .ZN(n8312) );
  AOI21_X1 U5445 ( .B1(n9493), .B2(n4795), .A(n4794), .ZN(n4793) );
  INV_X1 U5446 ( .A(n8205), .ZN(n4794) );
  AND2_X1 U5447 ( .A1(n8143), .A2(n8158), .ZN(n8248) );
  INV_X1 U5448 ( .A(n5870), .ZN(n4897) );
  NAND2_X1 U5449 ( .A1(n9492), .A2(n9493), .ZN(n9491) );
  NAND2_X1 U5450 ( .A1(n4757), .A2(n9508), .ZN(n4756) );
  INV_X1 U5451 ( .A(n5865), .ZN(n4884) );
  INV_X1 U5452 ( .A(n4887), .ZN(n4469) );
  NAND2_X1 U5453 ( .A1(n9765), .A2(n4762), .ZN(n4761) );
  NOR2_X1 U5454 ( .A1(n7218), .A2(n7380), .ZN(n4753) );
  NAND2_X1 U5455 ( .A1(n4799), .A2(n5892), .ZN(n8280) );
  NAND2_X1 U5456 ( .A1(n6848), .A2(n8082), .ZN(n8085) );
  AND2_X1 U5457 ( .A1(n6939), .A2(n4363), .ZN(n6960) );
  NAND2_X1 U5458 ( .A1(n6939), .A2(n4764), .ZN(n6970) );
  OR2_X1 U5459 ( .A1(n8176), .A2(n8324), .ZN(n5882) );
  NAND2_X1 U5460 ( .A1(n5877), .A2(n5876), .ZN(n8021) );
  NAND2_X1 U5461 ( .A1(n4824), .A2(n5743), .ZN(n4823) );
  INV_X1 U5462 ( .A(n5739), .ZN(n4824) );
  INV_X1 U5463 ( .A(n5743), .ZN(n4825) );
  OR2_X1 U5464 ( .A1(n4815), .A2(n5596), .ZN(n4813) );
  AND2_X1 U5465 ( .A1(n4815), .A2(n5596), .ZN(n4814) );
  AND2_X1 U5466 ( .A1(n5579), .A2(n5553), .ZN(n4839) );
  NAND2_X1 U5467 ( .A1(n4666), .A2(n4664), .ZN(n5523) );
  INV_X1 U5468 ( .A(n4670), .ZN(n4669) );
  NOR2_X1 U5469 ( .A1(n5446), .A2(n4955), .ZN(n5447) );
  INV_X1 U5470 ( .A(n5466), .ZN(n5446) );
  INV_X1 U5471 ( .A(n4829), .ZN(n4828) );
  OAI22_X1 U5472 ( .A1(n5438), .A2(n4831), .B1(n4833), .B2(n4830), .ZN(n4829)
         );
  INV_X1 U5473 ( .A(n4827), .ZN(n5442) );
  AOI21_X1 U5474 ( .B1(n5439), .B2(n4833), .A(n4830), .ZN(n4827) );
  NAND2_X1 U5475 ( .A1(n4400), .A2(n5312), .ZN(n4673) );
  AOI21_X1 U5476 ( .B1(n5313), .B2(n5315), .A(n4410), .ZN(n4672) );
  XNOR2_X1 U5477 ( .A(n5290), .B(SI_10_), .ZN(n5315) );
  NOR2_X2 U5478 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5119) );
  NOR2_X2 U5479 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5083) );
  OAI211_X1 U5480 ( .C1(n4651), .C2(n4649), .A(n4647), .B(n4646), .ZN(n5079)
         );
  NAND2_X1 U5481 ( .A1(n4648), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4647) );
  INV_X1 U5482 ( .A(n4650), .ZN(n4648) );
  NOR2_X1 U5483 ( .A1(n4699), .A2(n4701), .ZN(n4698) );
  INV_X1 U5484 ( .A(n6421), .ZN(n4699) );
  OR2_X1 U5485 ( .A1(n7957), .A2(n4701), .ZN(n4700) );
  NOR2_X1 U5486 ( .A1(n4655), .A2(n8932), .ZN(n4653) );
  INV_X1 U5487 ( .A(n4372), .ZN(n4655) );
  NAND2_X1 U5488 ( .A1(n7271), .A2(n4719), .ZN(n4721) );
  NAND2_X1 U5489 ( .A1(n4661), .A2(n4658), .ZN(n6446) );
  AND2_X1 U5490 ( .A1(n6456), .A2(n8492), .ZN(n8402) );
  OR2_X1 U5491 ( .A1(n6463), .A2(n6462), .ZN(n8403) );
  AND2_X1 U5492 ( .A1(n8492), .A2(n6441), .ZN(n8438) );
  AND2_X1 U5493 ( .A1(n8413), .A2(n6475), .ZN(n8446) );
  NAND2_X1 U5494 ( .A1(n8458), .A2(n4677), .ZN(n8397) );
  AND2_X1 U5495 ( .A1(n8388), .A2(n8458), .ZN(n8395) );
  AND2_X1 U5496 ( .A1(n8399), .A2(n6447), .ZN(n8458) );
  NAND2_X1 U5497 ( .A1(n4661), .A2(n4657), .ZN(n6447) );
  AND2_X1 U5498 ( .A1(n4658), .A2(n8951), .ZN(n4657) );
  XNOR2_X1 U5499 ( .A(n6404), .B(n6402), .ZN(n6403) );
  INV_X1 U5500 ( .A(n8883), .ZN(n8509) );
  AND4_X1 U5501 ( .A1(n8543), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n8772)
         );
  AND4_X1 U5502 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n6443)
         );
  NOR2_X1 U5503 ( .A1(n7479), .A2(n7478), .ZN(n7477) );
  NOR2_X1 U5504 ( .A1(n7489), .A2(n7490), .ZN(n7488) );
  NAND2_X1 U5505 ( .A1(n9990), .A2(n7349), .ZN(n7350) );
  AND2_X1 U5506 ( .A1(n4559), .A2(n4558), .ZN(n7410) );
  NAND2_X1 U5507 ( .A1(n7408), .A2(n10015), .ZN(n4558) );
  OAI21_X1 U5508 ( .B1(n4737), .B2(n7427), .A(n4736), .ZN(n7443) );
  AOI21_X1 U5509 ( .B1(n7429), .B2(n4739), .A(n4738), .ZN(n4736) );
  INV_X1 U5510 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4739) );
  NAND2_X1 U5511 ( .A1(n4448), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10008) );
  NAND2_X1 U5512 ( .A1(n7440), .A2(n7439), .ZN(n7744) );
  NAND2_X1 U5513 ( .A1(n7723), .A2(n10028), .ZN(n10033) );
  OR2_X1 U5514 ( .A1(n4741), .A2(n4740), .ZN(n10031) );
  INV_X1 U5515 ( .A(n10029), .ZN(n4740) );
  NAND2_X1 U5516 ( .A1(n4549), .A2(n4553), .ZN(n7801) );
  NAND2_X1 U5517 ( .A1(n7732), .A2(n4554), .ZN(n4549) );
  INV_X1 U5518 ( .A(n7740), .ZN(n4545) );
  INV_X1 U5519 ( .A(n7804), .ZN(n4546) );
  NAND2_X1 U5520 ( .A1(n4553), .A2(n7804), .ZN(n4548) );
  NAND2_X1 U5521 ( .A1(n4542), .A2(n4550), .ZN(n7800) );
  OR2_X1 U5522 ( .A1(n7732), .A2(n4552), .ZN(n4542) );
  NAND2_X1 U5523 ( .A1(n7789), .A2(n7751), .ZN(n7752) );
  NAND2_X1 U5524 ( .A1(n7983), .A2(n7984), .ZN(n7985) );
  NAND2_X1 U5525 ( .A1(n10043), .A2(n8832), .ZN(n10060) );
  AOI21_X1 U5526 ( .B1(n4534), .B2(n4537), .A(n4445), .ZN(n4533) );
  XNOR2_X1 U5527 ( .A(n4731), .B(n4730), .ZN(n10084) );
  NAND2_X1 U5528 ( .A1(n10077), .A2(n8803), .ZN(n10095) );
  NAND2_X1 U5529 ( .A1(n10095), .A2(n10096), .ZN(n10094) );
  INV_X1 U5530 ( .A(n4731), .ZN(n8789) );
  NAND2_X1 U5531 ( .A1(n10112), .A2(n10113), .ZN(n10111) );
  NAND2_X1 U5532 ( .A1(n10109), .A2(n8838), .ZN(n9790) );
  OAI21_X1 U5533 ( .B1(n8846), .B2(n8845), .A(n4526), .ZN(n4525) );
  INV_X1 U5534 ( .A(n8823), .ZN(n4526) );
  NAND2_X1 U5535 ( .A1(n9790), .A2(n9791), .ZN(n9789) );
  NAND2_X1 U5536 ( .A1(n8857), .A2(n6277), .ZN(n8532) );
  NAND2_X1 U5537 ( .A1(n6261), .A2(n7008), .ZN(n6271) );
  NOR2_X1 U5538 ( .A1(n6244), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U5539 ( .A1(n6219), .A2(n6218), .ZN(n6231) );
  OR2_X1 U5540 ( .A1(n6192), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U5541 ( .A1(n6179), .A2(n7070), .ZN(n6192) );
  AND2_X1 U5542 ( .A1(n6169), .A2(n6168), .ZN(n6179) );
  NOR2_X1 U5543 ( .A1(n6152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U5544 ( .A1(n6127), .A2(n7055), .ZN(n6138) );
  NOR3_X1 U5545 ( .A1(n4357), .A2(n7916), .A3(n4935), .ZN(n4934) );
  NOR2_X1 U5546 ( .A1(n4936), .A2(n7916), .ZN(n4933) );
  INV_X1 U5547 ( .A(n6317), .ZN(n4935) );
  AND4_X1 U5548 ( .A1(n6143), .A2(n6142), .A3(n6141), .A4(n6140), .ZN(n8366)
         );
  OR2_X1 U5549 ( .A1(n6109), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6117) );
  NOR2_X1 U5550 ( .A1(n6117), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6127) );
  OR2_X1 U5551 ( .A1(n6094), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U5552 ( .A1(n6086), .A2(n7754), .ZN(n6094) );
  NAND2_X1 U5553 ( .A1(n8641), .A2(n8632), .ZN(n8570) );
  NOR2_X1 U5554 ( .A1(n6061), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6071) );
  AND2_X1 U5555 ( .A1(n8639), .A2(n7516), .ZN(n8635) );
  AND4_X1 U5556 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n7595)
         );
  AND2_X1 U5557 ( .A1(n8623), .A2(n8619), .ZN(n8566) );
  OR2_X1 U5558 ( .A1(n8732), .A2(n8733), .ZN(n8871) );
  NAND2_X1 U5559 ( .A1(n4592), .A2(n8726), .ZN(n4591) );
  AND2_X1 U5560 ( .A1(n4589), .A2(n8727), .ZN(n4588) );
  INV_X1 U5561 ( .A(n8881), .ZN(n8879) );
  INV_X1 U5562 ( .A(n4567), .ZN(n8968) );
  AOI21_X1 U5563 ( .B1(n9016), .B2(n4570), .A(n4568), .ZN(n4567) );
  OAI21_X1 U5564 ( .B1(n4571), .B2(n4569), .A(n8986), .ZN(n4568) );
  AND2_X1 U5565 ( .A1(n6126), .A2(n6125), .ZN(n6429) );
  AOI21_X1 U5566 ( .B1(n4584), .B2(n8575), .A(n8664), .ZN(n4582) );
  NAND2_X1 U5567 ( .A1(n7719), .A2(n4584), .ZN(n4583) );
  NAND2_X1 U5568 ( .A1(n8597), .A2(n6928), .ZN(n10186) );
  OR2_X1 U5569 ( .A1(n6387), .A2(n8767), .ZN(n10192) );
  NAND2_X1 U5570 ( .A1(n4713), .A2(n4711), .ZN(n6346) );
  INV_X1 U5571 ( .A(n4712), .ZN(n4711) );
  OAI21_X1 U5572 ( .B1(n4714), .B2(n9166), .A(n6379), .ZN(n4712) );
  NOR2_X1 U5573 ( .A1(n4725), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n4722) );
  NOR3_X1 U5574 ( .A1(n6042), .A2(n4924), .A3(P2_IR_REG_8__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U5575 ( .A1(n7768), .A2(n7770), .ZN(n7769) );
  OAI21_X1 U5576 ( .B1(n5086), .B2(n5835), .A(n5037), .ZN(n5039) );
  OR2_X1 U5577 ( .A1(n5605), .A2(n5604), .ZN(n5624) );
  NAND2_X1 U5578 ( .A1(n4864), .A2(n4865), .ZN(n4861) );
  OR2_X1 U5579 ( .A1(n9225), .A2(n4862), .ZN(n4859) );
  NAND2_X1 U5580 ( .A1(n4865), .A2(n4866), .ZN(n4862) );
  INV_X1 U5581 ( .A(n5489), .ZN(n4844) );
  NOR2_X1 U5582 ( .A1(n4844), .A2(n4843), .ZN(n4842) );
  INV_X1 U5583 ( .A(n7770), .ZN(n4843) );
  OAI22_X1 U5584 ( .A1(n6910), .A2(n5061), .B1(n6837), .B2(n5086), .ZN(n5113)
         );
  NAND2_X1 U5585 ( .A1(n4471), .A2(n4874), .ZN(n4877) );
  NOR2_X1 U5586 ( .A1(n5636), .A2(n4875), .ZN(n4874) );
  INV_X1 U5587 ( .A(n5615), .ZN(n4875) );
  OR2_X1 U5588 ( .A1(n5090), .A2(n5088), .ZN(n5091) );
  INV_X1 U5589 ( .A(n5504), .ZN(n5502) );
  NAND2_X1 U5590 ( .A1(n4483), .A2(n5547), .ZN(n5548) );
  NAND2_X1 U5591 ( .A1(n4479), .A2(n4482), .ZN(n5552) );
  INV_X1 U5592 ( .A(n4483), .ZN(n4479) );
  NAND2_X1 U5593 ( .A1(n5142), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5168) );
  INV_X1 U5594 ( .A(n5144), .ZN(n5142) );
  INV_X2 U5595 ( .A(n5040), .ZN(n5754) );
  MUX2_X1 U5596 ( .A(n8209), .B(n8207), .S(n8176), .Z(n8168) );
  AND2_X1 U5597 ( .A1(n9734), .A2(n9461), .ZN(n8183) );
  INV_X1 U5598 ( .A(n8183), .ZN(n8315) );
  AND4_X1 U5599 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n7941)
         );
  OR2_X1 U5600 ( .A1(n9824), .A2(n9823), .ZN(n9826) );
  NOR3_X1 U5601 ( .A1(n9485), .A2(n9458), .A3(n4750), .ZN(n4748) );
  NAND2_X1 U5602 ( .A1(n4751), .A2(n9738), .ZN(n4750) );
  INV_X1 U5603 ( .A(n4751), .ZN(n4749) );
  NOR3_X1 U5604 ( .A1(n4944), .A2(n4756), .A3(n9486), .ZN(n5885) );
  NOR2_X1 U5605 ( .A1(n4944), .A2(n4755), .ZN(n9527) );
  INV_X1 U5606 ( .A(n4757), .ZN(n4755) );
  OR3_X1 U5607 ( .A1(n5669), .A2(n9228), .A3(n5668), .ZN(n5696) );
  NAND2_X1 U5608 ( .A1(n5622), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5669) );
  INV_X1 U5609 ( .A(n5624), .ZN(n5622) );
  NAND2_X1 U5610 ( .A1(n9606), .A2(n8058), .ZN(n9590) );
  NAND2_X1 U5611 ( .A1(n9590), .A2(n9591), .ZN(n9589) );
  NOR2_X1 U5612 ( .A1(n7824), .A2(n4760), .ZN(n9625) );
  INV_X1 U5613 ( .A(n4762), .ZN(n4760) );
  AND2_X1 U5614 ( .A1(n4460), .A2(n7688), .ZN(n4459) );
  OR2_X1 U5615 ( .A1(n4356), .A2(n4461), .ZN(n4460) );
  INV_X1 U5616 ( .A(n5852), .ZN(n4461) );
  INV_X1 U5617 ( .A(n4801), .ZN(n4800) );
  OAI21_X1 U5618 ( .B1(n8235), .B2(n4802), .A(n8291), .ZN(n4801) );
  INV_X1 U5619 ( .A(n4803), .ZN(n4802) );
  NAND2_X1 U5620 ( .A1(n5453), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5480) );
  OR2_X1 U5621 ( .A1(n5480), .A2(n5454), .ZN(n5504) );
  NOR2_X1 U5622 ( .A1(n7560), .A2(n9725), .ZN(n7643) );
  NAND2_X1 U5623 ( .A1(n7643), .A2(n7788), .ZN(n7682) );
  NAND2_X1 U5624 ( .A1(n7557), .A2(n8235), .ZN(n4805) );
  NAND2_X1 U5625 ( .A1(n4805), .A2(n4803), .ZN(n7687) );
  NAND2_X1 U5626 ( .A1(n4753), .A2(n4752), .ZN(n7560) );
  INV_X1 U5627 ( .A(n4753), .ZN(n7386) );
  NAND2_X1 U5628 ( .A1(n7384), .A2(n7390), .ZN(n7383) );
  OR2_X1 U5629 ( .A1(n5369), .A2(n5368), .ZN(n5390) );
  NAND2_X1 U5630 ( .A1(n5297), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5369) );
  INV_X1 U5631 ( .A(n5326), .ZN(n5297) );
  NAND2_X1 U5632 ( .A1(n5241), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U5633 ( .A1(n4807), .A2(n4806), .ZN(n8093) );
  AND2_X1 U5634 ( .A1(n9294), .A2(n5273), .ZN(n4806) );
  AND4_X1 U5635 ( .A1(n5249), .A2(n5248), .A3(n5247), .A4(n5246), .ZN(n7263)
         );
  NAND2_X1 U5636 ( .A1(n6939), .A2(n4766), .ZN(n6883) );
  AOI21_X1 U5637 ( .B1(n6937), .B2(n4465), .A(n4395), .ZN(n4464) );
  NAND2_X1 U5638 ( .A1(n4950), .A2(n6937), .ZN(n4463) );
  OAI21_X1 U5639 ( .B1(n6587), .B2(n5110), .A(n4521), .ZN(n6943) );
  AND2_X1 U5640 ( .A1(n5187), .A2(n4416), .ZN(n4521) );
  AND4_X1 U5641 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n6931)
         );
  NAND2_X1 U5642 ( .A1(n8080), .A2(n8275), .ZN(n8225) );
  NOR2_X1 U5643 ( .A1(n6707), .A2(n6818), .ZN(n6747) );
  INV_X1 U5644 ( .A(n5555), .ZN(n4485) );
  NAND2_X1 U5645 ( .A1(n8075), .A2(n8266), .ZN(n8218) );
  NAND2_X1 U5646 ( .A1(n8175), .A2(n8174), .ZN(n9467) );
  NAND2_X1 U5647 ( .A1(n8014), .A2(n8172), .ZN(n4838) );
  NAND2_X1 U5648 ( .A1(n5718), .A2(n5717), .ZN(n9665) );
  NAND2_X1 U5649 ( .A1(n5667), .A2(n5666), .ZN(n9676) );
  NAND2_X1 U5650 ( .A1(n5621), .A2(n5620), .ZN(n9688) );
  NOR2_X1 U5651 ( .A1(n5716), .A2(n4649), .ZN(n4878) );
  AND2_X1 U5652 ( .A1(n5916), .A2(n5915), .ZN(n6814) );
  NAND2_X1 U5653 ( .A1(n6806), .A2(n5882), .ZN(n9978) );
  INV_X1 U5654 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5001) );
  INV_X1 U5655 ( .A(n4984), .ZN(n4981) );
  NAND2_X1 U5656 ( .A1(n4973), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U5657 ( .A1(n4969), .A2(n4379), .ZN(n4869) );
  NAND2_X1 U5658 ( .A1(n5289), .A2(n5286), .ZN(n4639) );
  CLKBUF_X1 U5659 ( .A(n5994), .Z(n6563) );
  NAND2_X1 U5660 ( .A1(n7271), .A2(n4962), .ZN(n7505) );
  AND4_X1 U5661 ( .A1(n6276), .A2(n6275), .A3(n6274), .A4(n6273), .ZN(n8591)
         );
  AND2_X1 U5662 ( .A1(n6191), .A2(n6190), .ZN(n8394) );
  AND2_X1 U5663 ( .A1(n8396), .A2(n8388), .ZN(n8459) );
  AND2_X1 U5664 ( .A1(n4721), .A2(n4380), .ZN(n7630) );
  NAND2_X1 U5665 ( .A1(n7893), .A2(n6421), .ZN(n7958) );
  NAND2_X1 U5666 ( .A1(n7958), .A2(n7957), .ZN(n7956) );
  INV_X1 U5667 ( .A(n10132), .ZN(n7192) );
  AND2_X1 U5668 ( .A1(n4696), .A2(n4355), .ZN(n7188) );
  INV_X1 U5669 ( .A(n4717), .ZN(n4716) );
  OAI22_X1 U5670 ( .A1(n7629), .A2(n4380), .B1(n8780), .B2(n6415), .ZN(n4717)
         );
  AND4_X1 U5671 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n7908)
         );
  XNOR2_X1 U5672 ( .A(n6403), .B(n8782), .ZN(n6868) );
  AND4_X1 U5673 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n7656)
         );
  NAND2_X1 U5674 ( .A1(n6489), .A2(n6488), .ZN(n8507) );
  INV_X1 U5675 ( .A(n8524), .ZN(n8514) );
  AND2_X1 U5676 ( .A1(n6137), .A2(n6136), .ZN(n8560) );
  NAND2_X1 U5677 ( .A1(n8362), .A2(n4709), .ZN(n8521) );
  AND2_X1 U5678 ( .A1(n4710), .A2(n6435), .ZN(n4709) );
  INV_X1 U5679 ( .A(n8519), .ZN(n4710) );
  NAND2_X1 U5680 ( .A1(n8362), .A2(n6435), .ZN(n8520) );
  INV_X1 U5681 ( .A(n4353), .ZN(n8762) );
  INV_X1 U5682 ( .A(n8591), .ZN(n8873) );
  NAND4_X1 U5683 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n8775)
         );
  INV_X1 U5684 ( .A(n7908), .ZN(n8778) );
  NAND4_X1 U5685 ( .A1(n6076), .A2(n6075), .A3(n6074), .A4(n6073), .ZN(n8779)
         );
  INV_X1 U5686 ( .A(n7511), .ZN(n8780) );
  INV_X1 U5687 ( .A(n7656), .ZN(n7634) );
  INV_X1 U5688 ( .A(n7595), .ZN(n8781) );
  NAND2_X1 U5689 ( .A1(n4958), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5983) );
  NOR2_X1 U5690 ( .A1(n7457), .A2(n7456), .ZN(n7478) );
  AND2_X1 U5691 ( .A1(n7349), .A2(n4733), .ZN(n9991) );
  INV_X1 U5692 ( .A(n4561), .ZN(n7406) );
  INV_X1 U5693 ( .A(n4559), .ZN(n10003) );
  AOI21_X1 U5694 ( .B1(n7732), .B2(n7731), .A(n4365), .ZN(n10038) );
  AND2_X1 U5695 ( .A1(n4547), .A2(n4543), .ZN(n7871) );
  INV_X1 U5696 ( .A(n4544), .ZN(n4543) );
  OR2_X1 U5697 ( .A1(n7732), .A2(n4548), .ZN(n4547) );
  OAI21_X1 U5698 ( .B1(n4550), .B2(n4546), .A(n4545), .ZN(n4544) );
  INV_X1 U5699 ( .A(n4729), .ZN(n7725) );
  INV_X1 U5700 ( .A(n4606), .ZN(n7968) );
  OAI21_X1 U5701 ( .B1(n7881), .B2(n4604), .A(n4603), .ZN(n8785) );
  NAND2_X1 U5702 ( .A1(n4607), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4604) );
  NAND2_X1 U5703 ( .A1(n7969), .A2(n4607), .ZN(n4603) );
  INV_X1 U5704 ( .A(n7971), .ZN(n4607) );
  INV_X1 U5705 ( .A(n7969), .ZN(n4605) );
  AND2_X1 U5706 ( .A1(n4536), .A2(n4540), .ZN(n10046) );
  NAND2_X1 U5707 ( .A1(n4536), .A2(n4534), .ZN(n10045) );
  INV_X1 U5708 ( .A(n4614), .ZN(n10050) );
  INV_X1 U5709 ( .A(n8787), .ZN(n4613) );
  INV_X1 U5710 ( .A(n4617), .ZN(n10118) );
  INV_X1 U5711 ( .A(n9794), .ZN(n9797) );
  NAND2_X1 U5712 ( .A1(n4617), .A2(n4616), .ZN(n9796) );
  NOR2_X1 U5713 ( .A1(n8793), .A2(n4745), .ZN(n4616) );
  INV_X1 U5714 ( .A(n8840), .ZN(n10116) );
  OR2_X1 U5715 ( .A1(n9786), .A2(n9785), .ZN(n9787) );
  INV_X1 U5716 ( .A(n10004), .ZN(n10115) );
  XNOR2_X1 U5717 ( .A(n8532), .B(n8738), .ZN(n6525) );
  NAND2_X1 U5718 ( .A1(n6217), .A2(n6216), .ZN(n8938) );
  AOI21_X1 U5719 ( .B1(n9006), .B2(n4915), .A(n4912), .ZN(n8969) );
  INV_X1 U5720 ( .A(n6092), .ZN(n7711) );
  NAND2_X1 U5721 ( .A1(n10145), .A2(n7300), .ZN(n9026) );
  AND2_X1 U5722 ( .A1(n6686), .A2(n6539), .ZN(n10140) );
  NAND2_X1 U5723 ( .A1(n5994), .A2(n4926), .ZN(n4925) );
  OAI22_X1 U5724 ( .A1(n6580), .A2(n5716), .B1(n4652), .B2(n4840), .ZN(n4926)
         );
  INV_X1 U5725 ( .A(n10140), .ZN(n8977) );
  OR2_X1 U5726 ( .A1(n6388), .A2(n8899), .ZN(n8855) );
  INV_X1 U5727 ( .A(n4597), .ZN(n4596) );
  INV_X1 U5728 ( .A(n8855), .ZN(n10138) );
  NAND2_X1 U5729 ( .A1(n4585), .A2(n8656), .ZN(n7811) );
  OR2_X1 U5730 ( .A1(n7719), .A2(n8575), .ZN(n4585) );
  INV_X1 U5731 ( .A(n9048), .ZN(n9075) );
  INV_X1 U5732 ( .A(n8852), .ZN(n9080) );
  AND2_X1 U5733 ( .A1(n8536), .A2(n8535), .ZN(n9086) );
  NAND2_X1 U5734 ( .A1(n6270), .A2(n6269), .ZN(n9089) );
  NAND2_X1 U5735 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  NAND2_X1 U5736 ( .A1(n8883), .A2(n10129), .ZN(n8861) );
  NAND2_X1 U5737 ( .A1(n6260), .A2(n6259), .ZN(n9095) );
  NAND2_X1 U5738 ( .A1(n6250), .A2(n6249), .ZN(n9101) );
  NAND2_X1 U5739 ( .A1(n7762), .A2(n8544), .ZN(n6250) );
  NAND2_X1 U5740 ( .A1(n8891), .A2(n6327), .ZN(n8882) );
  NAND2_X1 U5741 ( .A1(n6243), .A2(n6242), .ZN(n9107) );
  NAND2_X1 U5742 ( .A1(n4587), .A2(n4592), .ZN(n8889) );
  NAND2_X1 U5743 ( .A1(n8941), .A2(n4594), .ZN(n4587) );
  NAND2_X1 U5744 ( .A1(n6237), .A2(n6236), .ZN(n9113) );
  NAND2_X1 U5745 ( .A1(n8941), .A2(n4595), .ZN(n8911) );
  AND2_X1 U5746 ( .A1(n6228), .A2(n6227), .ZN(n9119) );
  NAND2_X1 U5747 ( .A1(n8929), .A2(n6325), .ZN(n8918) );
  NAND2_X1 U5748 ( .A1(n6208), .A2(n6207), .ZN(n9126) );
  NAND2_X1 U5749 ( .A1(n6199), .A2(n6198), .ZN(n9132) );
  NAND2_X1 U5750 ( .A1(n6178), .A2(n6177), .ZN(n9142) );
  NAND2_X1 U5751 ( .A1(n4913), .A2(n4917), .ZN(n8990) );
  NAND2_X1 U5752 ( .A1(n9006), .A2(n4916), .ZN(n4913) );
  NAND2_X1 U5753 ( .A1(n4428), .A2(n4575), .ZN(n8985) );
  NAND2_X1 U5754 ( .A1(n6166), .A2(n6165), .ZN(n9148) );
  OAI21_X1 U5755 ( .B1(n9006), .B2(n9007), .A(n4921), .ZN(n8998) );
  INV_X1 U5756 ( .A(n4572), .ZN(n8997) );
  OAI21_X1 U5757 ( .B1(n9016), .B2(n4574), .A(n4573), .ZN(n4572) );
  INV_X1 U5758 ( .A(n4578), .ZN(n4574) );
  NAND2_X1 U5759 ( .A1(n6151), .A2(n6150), .ZN(n9154) );
  INV_X1 U5760 ( .A(n8560), .ZN(n9160) );
  INV_X1 U5761 ( .A(n6429), .ZN(n8372) );
  NAND2_X1 U5762 ( .A1(n6116), .A2(n6115), .ZN(n8479) );
  NOR2_X1 U5763 ( .A1(n7812), .A2(n4357), .ZN(n7917) );
  INV_X1 U5764 ( .A(n9118), .ZN(n9161) );
  NAND2_X1 U5765 ( .A1(n5972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5973) );
  AND2_X1 U5766 ( .A1(n5965), .A2(n5970), .ZN(n5971) );
  NOR2_X1 U5767 ( .A1(n4840), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9169) );
  NOR2_X1 U5768 ( .A1(n4349), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7850) );
  XNOR2_X1 U5769 ( .A(n6287), .B(n6286), .ZN(n8755) );
  NAND2_X1 U5770 ( .A1(n6007), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4618) );
  NOR2_X1 U5771 ( .A1(n5995), .A2(n9166), .ZN(n4727) );
  XNOR2_X1 U5772 ( .A(n5986), .B(n5985), .ZN(n7483) );
  NOR2_X1 U5773 ( .A1(n6796), .A2(n4873), .ZN(n4872) );
  INV_X1 U5774 ( .A(n5195), .ZN(n4873) );
  NAND2_X1 U5775 ( .A1(n6767), .A2(n5195), .ZN(n6795) );
  NAND2_X1 U5776 ( .A1(n4484), .A2(n4431), .ZN(n4474) );
  INV_X1 U5777 ( .A(n5515), .ZN(n4475) );
  NAND2_X1 U5778 ( .A1(n5559), .A2(n5558), .ZN(n9628) );
  NAND2_X1 U5779 ( .A1(n6658), .A2(n6657), .ZN(n5066) );
  NAND2_X1 U5780 ( .A1(n5601), .A2(n5600), .ZN(n9597) );
  NAND2_X1 U5781 ( .A1(n4859), .A2(n4861), .ZN(n9272) );
  OR2_X1 U5782 ( .A1(n9225), .A2(n9223), .ZN(n4860) );
  NAND2_X1 U5783 ( .A1(n5452), .A2(n5451), .ZN(n9720) );
  AND4_X1 U5784 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n6882)
         );
  NAND2_X1 U5785 ( .A1(n6720), .A2(n4847), .ZN(n6568) );
  NAND2_X1 U5786 ( .A1(n5500), .A2(n5499), .ZN(n7866) );
  AOI21_X1 U5787 ( .B1(n9225), .B2(n9224), .A(n9223), .ZN(n9227) );
  NAND2_X1 U5788 ( .A1(n6728), .A2(n6729), .ZN(n6727) );
  NOR2_X1 U5789 ( .A1(n4480), .A2(n4477), .ZN(n4476) );
  NAND2_X1 U5790 ( .A1(n7374), .A2(n7375), .ZN(n4854) );
  NAND2_X1 U5791 ( .A1(n5552), .A2(n5548), .ZN(n9257) );
  INV_X1 U5792 ( .A(n6943), .ZN(n9964) );
  AND2_X1 U5793 ( .A1(n5752), .A2(n5751), .ZN(n9280) );
  OR2_X1 U5794 ( .A1(n9488), .A2(n5069), .ZN(n5752) );
  INV_X1 U5795 ( .A(n9285), .ZN(n9265) );
  OR2_X1 U5796 ( .A1(n9276), .A2(n5069), .ZN(n5730) );
  NAND2_X1 U5797 ( .A1(n5118), .A2(n4385), .ZN(n6625) );
  NAND2_X1 U5798 ( .A1(n5100), .A2(n4690), .ZN(n9298) );
  AND2_X1 U5799 ( .A1(n5099), .A2(n4688), .ZN(n4690) );
  AND2_X1 U5800 ( .A1(n4689), .A2(n4691), .ZN(n4688) );
  NOR2_X1 U5801 ( .A1(n9459), .A2(n9682), .ZN(n9652) );
  INV_X1 U5802 ( .A(n4746), .ZN(n9459) );
  AOI211_X1 U5803 ( .C1(n9485), .C2(n9458), .A(n4748), .B(n4747), .ZN(n4746)
         );
  AND2_X1 U5804 ( .A1(n4750), .A2(n9458), .ZN(n4747) );
  NOR2_X1 U5805 ( .A1(n5932), .A2(n5871), .ZN(n5879) );
  AND2_X1 U5806 ( .A1(n8151), .A2(n6874), .ZN(n5871) );
  OR2_X1 U5807 ( .A1(n5903), .A2(n9546), .ZN(n5911) );
  NAND2_X1 U5808 ( .A1(n4682), .A2(n4683), .ZN(n9484) );
  NAND2_X1 U5809 ( .A1(n4881), .A2(n5865), .ZN(n9536) );
  NAND2_X1 U5810 ( .A1(n5864), .A2(n4885), .ZN(n4881) );
  NAND2_X1 U5811 ( .A1(n5864), .A2(n5863), .ZN(n9554) );
  OAI21_X1 U5812 ( .B1(n9606), .B2(n4778), .A(n4775), .ZN(n9581) );
  NAND2_X1 U5813 ( .A1(n4891), .A2(n4887), .ZN(n9605) );
  OAI21_X1 U5814 ( .B1(n7925), .B2(n4375), .A(n5856), .ZN(n9624) );
  NAND2_X1 U5815 ( .A1(n4458), .A2(n5852), .ZN(n7681) );
  NAND2_X1 U5816 ( .A1(n5851), .A2(n4356), .ZN(n4458) );
  NAND2_X1 U5817 ( .A1(n5851), .A2(n5850), .ZN(n7642) );
  OAI21_X1 U5818 ( .B1(n6950), .B2(n8230), .A(n4769), .ZN(n7281) );
  NAND2_X1 U5819 ( .A1(n7213), .A2(n7214), .ZN(n7212) );
  NAND2_X1 U5820 ( .A1(n6950), .A2(n8115), .ZN(n7213) );
  NAND2_X1 U5821 ( .A1(n6938), .A2(n6937), .ZN(n6936) );
  NAND2_X1 U5822 ( .A1(n6781), .A2(n5841), .ZN(n6938) );
  OR2_X1 U5823 ( .A1(n5917), .A2(n8325), .ZN(n9630) );
  NAND2_X1 U5824 ( .A1(n5948), .A2(n9988), .ZN(n4693) );
  INV_X1 U5825 ( .A(n9467), .ZN(n9738) );
  AND2_X1 U5826 ( .A1(n5162), .A2(n5161), .ZN(n6981) );
  AND2_X1 U5827 ( .A1(n5160), .A2(n4381), .ZN(n5161) );
  XNOR2_X1 U5828 ( .A(n8031), .B(n8030), .ZN(n9781) );
  OAI21_X1 U5829 ( .B1(n8171), .B2(n8170), .A(n8027), .ZN(n8031) );
  NAND2_X1 U5830 ( .A1(n5017), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U5831 ( .A1(n4948), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n5019) );
  XNOR2_X1 U5832 ( .A(n5873), .B(n5872), .ZN(n7854) );
  NAND2_X1 U5833 ( .A1(n5020), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U5834 ( .A1(n4992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4989) );
  NAND2_X1 U5835 ( .A1(n4984), .A2(n4900), .ZN(n4994) );
  XNOR2_X1 U5836 ( .A(n5598), .B(n5583), .ZN(n6827) );
  NOR2_X1 U5837 ( .A1(n4840), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9780) );
  CLKBUF_X1 U5838 ( .A(n5555), .Z(n8317) );
  INV_X1 U5839 ( .A(n6592), .ZN(n6079) );
  AOI21_X1 U5840 ( .B1(n4371), .B2(n4784), .A(n4780), .ZN(n4779) );
  INV_X1 U5841 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5210) );
  XNOR2_X1 U5842 ( .A(n5312), .B(n5224), .ZN(n6587) );
  AND2_X1 U5843 ( .A1(n4835), .A2(n4383), .ZN(n5130) );
  OAI21_X1 U5844 ( .B1(n4840), .B2(n5049), .A(n5048), .ZN(n5051) );
  INV_X1 U5845 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5006) );
  NAND2_X1 U5846 ( .A1(n4530), .A2(n8815), .ZN(n4529) );
  AOI21_X1 U5847 ( .B1(n4527), .B2(n9803), .A(n4523), .ZN(n4522) );
  OAI22_X1 U5848 ( .A1(n6545), .A2(n9048), .B1(n10225), .B2(n6544), .ZN(n6546)
         );
  NOR2_X1 U5849 ( .A1(n6537), .A2(n4952), .ZN(n6538) );
  NOR2_X1 U5850 ( .A1(n10205), .A2(n6535), .ZN(n6537) );
  AOI21_X1 U5851 ( .B1(n4486), .B2(n4382), .A(n5832), .ZN(n5833) );
  OR2_X1 U5852 ( .A1(n8328), .A2(n8327), .ZN(n4819) );
  INV_X1 U5853 ( .A(n5945), .ZN(n5946) );
  OAI22_X1 U5854 ( .A1(n8339), .A2(n9770), .B1(n9981), .B2(n5944), .ZN(n5945)
         );
  AND2_X1 U5855 ( .A1(n8456), .A2(n8894), .ZN(n8718) );
  INV_X1 U5856 ( .A(n8115), .ZN(n4771) );
  NAND2_X1 U5857 ( .A1(n4563), .A2(n5951), .ZN(n6017) );
  INV_X1 U5858 ( .A(n6404), .ZN(n6405) );
  NAND2_X2 U5859 ( .A1(n4996), .A2(n5036), .ZN(n5040) );
  INV_X1 U5860 ( .A(n9493), .ZN(n4796) );
  NAND2_X1 U5861 ( .A1(n4575), .A2(n8691), .ZN(n4571) );
  NAND2_X1 U5862 ( .A1(n6407), .A2(n10130), .ZN(n4355) );
  AND2_X1 U5863 ( .A1(n5850), .A2(n4399), .ZN(n4356) );
  INV_X1 U5864 ( .A(n8999), .ZN(n4919) );
  AND2_X1 U5865 ( .A1(n8663), .A2(n8776), .ZN(n4357) );
  AND2_X1 U5866 ( .A1(n5036), .A2(n5035), .ZN(n5175) );
  INV_X1 U5867 ( .A(n5175), .ZN(n5212) );
  INV_X2 U5868 ( .A(n5175), .ZN(n5061) );
  AND3_X1 U5869 ( .A1(n5954), .A2(n5956), .A3(n5955), .ZN(n4359) );
  AND2_X1 U5870 ( .A1(n5289), .A2(n5184), .ZN(n4360) );
  INV_X1 U5871 ( .A(n4922), .ZN(n4921) );
  NOR2_X1 U5872 ( .A1(n8436), .A2(n8774), .ZN(n4922) );
  AND2_X1 U5873 ( .A1(n6455), .A2(n6445), .ZN(n8400) );
  NAND2_X1 U5874 ( .A1(n4818), .A2(n8324), .ZN(n4361) );
  INV_X1 U5875 ( .A(n4880), .ZN(n4455) );
  NOR2_X1 U5876 ( .A1(n4832), .A2(n5358), .ZN(n4362) );
  AND2_X1 U5877 ( .A1(n4764), .A2(n4763), .ZN(n4363) );
  AND2_X1 U5878 ( .A1(n5757), .A2(n4823), .ZN(n4364) );
  AND2_X1 U5879 ( .A1(n7729), .A2(n7730), .ZN(n4365) );
  NAND2_X1 U5880 ( .A1(n8113), .A2(n8101), .ZN(n4366) );
  INV_X1 U5881 ( .A(n9795), .ZN(n4745) );
  NOR2_X1 U5882 ( .A1(n8317), .A2(n5818), .ZN(n4367) );
  INV_X1 U5883 ( .A(n5095), .ZN(n5626) );
  NAND2_X4 U5884 ( .A1(n8344), .A2(n5028), .ZN(n5095) );
  NAND2_X1 U5885 ( .A1(n5357), .A2(n5356), .ZN(n5439) );
  NAND2_X1 U5886 ( .A1(n5994), .A2(n5716), .ZN(n6008) );
  NAND2_X1 U5887 ( .A1(n8344), .A2(n8016), .ZN(n5097) );
  NAND2_X1 U5888 ( .A1(n4358), .A2(n5176), .ZN(n5293) );
  AND2_X1 U5889 ( .A1(n4983), .A2(n4901), .ZN(n4368) );
  AND2_X1 U5890 ( .A1(n4563), .A2(n4565), .ZN(n6028) );
  OR2_X1 U5891 ( .A1(n6042), .A2(n4924), .ZN(n4369) );
  NAND2_X1 U5892 ( .A1(n6291), .A2(n6289), .ZN(n4370) );
  AND2_X1 U5893 ( .A1(n4782), .A2(n5228), .ZN(n4371) );
  OR2_X1 U5894 ( .A1(n6467), .A2(n6466), .ZN(n4372) );
  NAND2_X1 U5895 ( .A1(n9529), .A2(n9512), .ZN(n4373) );
  OR2_X1 U5896 ( .A1(n5033), .A2(n5032), .ZN(n9300) );
  AND2_X2 U5897 ( .A1(n5040), .A2(n5038), .ZN(n5086) );
  NOR2_X1 U5898 ( .A1(n8669), .A2(n8775), .ZN(n4374) );
  AND2_X1 U5899 ( .A1(n6320), .A2(n8688), .ZN(n9007) );
  NOR2_X1 U5900 ( .A1(n9709), .A2(n9642), .ZN(n4375) );
  NOR2_X1 U5901 ( .A1(n5179), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5235) );
  AND2_X1 U5902 ( .A1(n5929), .A2(n5930), .ZN(n4376) );
  OR2_X1 U5903 ( .A1(n10201), .A2(n8777), .ZN(n4377) );
  AND2_X1 U5904 ( .A1(n4879), .A2(n4373), .ZN(n4378) );
  AND2_X1 U5905 ( .A1(n4871), .A2(n4870), .ZN(n4379) );
  OR2_X1 U5906 ( .A1(n6414), .A2(n7634), .ZN(n4380) );
  OR2_X1 U5907 ( .A1(n6611), .A2(n9370), .ZN(n4381) );
  INV_X1 U5908 ( .A(n8190), .ZN(n4795) );
  INV_X1 U5909 ( .A(n8668), .ZN(n4937) );
  INV_X1 U5910 ( .A(n5069), .ZN(n5763) );
  NAND2_X1 U5911 ( .A1(n5818), .A2(n8264), .ZN(n5034) );
  AND3_X1 U5912 ( .A1(n5828), .A2(n9274), .A3(n5827), .ZN(n4382) );
  XNOR2_X1 U5913 ( .A(n4618), .B(n5951), .ZN(n7348) );
  NAND2_X1 U5914 ( .A1(n4656), .A2(n6472), .ZN(n8375) );
  NAND2_X1 U5915 ( .A1(n8856), .A2(n8858), .ZN(n8857) );
  OR2_X1 U5916 ( .A1(n5126), .A2(n5125), .ZN(n4383) );
  NAND2_X1 U5917 ( .A1(n6028), .A2(n6029), .ZN(n6042) );
  NOR2_X1 U5918 ( .A1(n4481), .A2(n4478), .ZN(n4384) );
  NAND2_X1 U5919 ( .A1(n8167), .A2(n8166), .ZN(n8250) );
  INV_X1 U5920 ( .A(n8250), .ZN(n4797) );
  AND3_X1 U5921 ( .A1(n5117), .A2(n5116), .A3(n4466), .ZN(n4385) );
  OR2_X1 U5922 ( .A1(n4793), .A2(n4797), .ZN(n4386) );
  AND2_X1 U5923 ( .A1(n8090), .A2(n6846), .ZN(n4387) );
  NAND2_X1 U5924 ( .A1(n4853), .A2(n4852), .ZN(n5431) );
  OR2_X1 U5925 ( .A1(n8688), .A2(n8747), .ZN(n4388) );
  NAND2_X1 U5926 ( .A1(n5533), .A2(n5532), .ZN(n9709) );
  AND2_X1 U5927 ( .A1(n5988), .A2(n4925), .ZN(n10147) );
  INV_X1 U5928 ( .A(n10147), .ZN(n4927) );
  AND2_X1 U5929 ( .A1(n9676), .A2(n9560), .ZN(n4389) );
  INV_X1 U5930 ( .A(n9529), .ZN(n9747) );
  NAND2_X1 U5931 ( .A1(n5694), .A2(n5693), .ZN(n9529) );
  AND2_X1 U5932 ( .A1(n7724), .A2(n7796), .ZN(n4390) );
  NOR2_X1 U5933 ( .A1(n9119), .A2(n8488), .ZN(n4391) );
  INV_X1 U5934 ( .A(n4754), .ZN(n9504) );
  NOR2_X1 U5935 ( .A1(n4944), .A2(n4756), .ZN(n4754) );
  INV_X1 U5936 ( .A(n4514), .ZN(n4513) );
  NAND2_X1 U5937 ( .A1(n4517), .A2(n8200), .ZN(n4514) );
  NOR2_X1 U5938 ( .A1(n9485), .A2(n4750), .ZN(n4392) );
  INV_X1 U5939 ( .A(n4571), .ZN(n4570) );
  AND2_X1 U5940 ( .A1(n4767), .A2(n7282), .ZN(n4393) );
  AND2_X1 U5941 ( .A1(n5953), .A2(n4923), .ZN(n4394) );
  AND2_X1 U5942 ( .A1(n6882), .A2(n9964), .ZN(n4395) );
  AND2_X1 U5943 ( .A1(n4860), .A2(n4863), .ZN(n4396) );
  INV_X1 U5944 ( .A(n9223), .ZN(n4866) );
  AND2_X1 U5945 ( .A1(n4654), .A2(n4372), .ZN(n6472) );
  AND2_X1 U5946 ( .A1(n5402), .A2(n5401), .ZN(n4397) );
  NAND2_X1 U5947 ( .A1(n5225), .A2(n5224), .ZN(n5286) );
  AND2_X1 U5948 ( .A1(n8394), .A2(n8498), .ZN(n4398) );
  OR2_X1 U5949 ( .A1(n7947), .A2(n9288), .ZN(n4399) );
  NAND2_X1 U5950 ( .A1(n4807), .A2(n5273), .ZN(n6853) );
  INV_X1 U5951 ( .A(n6853), .ZN(n4765) );
  AND2_X1 U5952 ( .A1(n5311), .A2(n5315), .ZN(n4400) );
  OR2_X1 U5953 ( .A1(n6042), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n4401) );
  NAND2_X1 U5954 ( .A1(n4984), .A2(n4368), .ZN(n4402) );
  AND2_X1 U5955 ( .A1(n9101), .A2(n8895), .ZN(n4403) );
  AND2_X1 U5956 ( .A1(n9119), .A2(n8488), .ZN(n4404) );
  AND2_X1 U5957 ( .A1(n8941), .A2(n8702), .ZN(n4405) );
  AND2_X1 U5958 ( .A1(n8039), .A2(n8040), .ZN(n9582) );
  INV_X1 U5959 ( .A(n9582), .ZN(n4774) );
  INV_X1 U5960 ( .A(n8725), .ZN(n8892) );
  AND2_X1 U5961 ( .A1(n8727), .A2(n8726), .ZN(n8725) );
  AND2_X1 U5962 ( .A1(n4693), .A2(n4692), .ZN(n4406) );
  AND2_X1 U5963 ( .A1(n8517), .A2(n8420), .ZN(n4407) );
  AND2_X1 U5964 ( .A1(n7866), .A2(n9287), .ZN(n4408) );
  NOR2_X1 U5965 ( .A1(n6454), .A2(n6453), .ZN(n4409) );
  NAND2_X1 U5966 ( .A1(n5995), .A2(n5996), .ZN(n6007) );
  AND2_X1 U5967 ( .A1(n5995), .A2(n5996), .ZN(n4563) );
  AND2_X1 U5968 ( .A1(n5291), .A2(SI_10_), .ZN(n4410) );
  INV_X1 U5969 ( .A(n6320), .ZN(n8694) );
  OR2_X1 U5970 ( .A1(n9154), .A2(n8774), .ZN(n6320) );
  AND2_X1 U5971 ( .A1(n8746), .A2(n8537), .ZN(n8738) );
  INV_X1 U5972 ( .A(n4864), .ZN(n4863) );
  OAI21_X1 U5973 ( .B1(n9223), .B2(n9224), .A(n5687), .ZN(n4864) );
  OR2_X1 U5974 ( .A1(n8151), .A2(n9496), .ZN(n8143) );
  INV_X1 U5975 ( .A(n5965), .ZN(n4942) );
  OR2_X1 U5976 ( .A1(n4680), .A2(n4408), .ZN(n4411) );
  OR2_X1 U5977 ( .A1(n4917), .A2(n4914), .ZN(n4412) );
  OR2_X1 U5978 ( .A1(n8088), .A2(n8176), .ZN(n4413) );
  AND3_X1 U5979 ( .A1(n4978), .A2(n4979), .A3(n4977), .ZN(n4414) );
  AND2_X1 U5980 ( .A1(n9148), .A2(n9008), .ZN(n4415) );
  OR2_X1 U5981 ( .A1(n6611), .A2(n9368), .ZN(n4416) );
  AND3_X1 U5982 ( .A1(n6000), .A2(n5999), .A3(n5998), .ZN(n6402) );
  AND2_X1 U5983 ( .A1(n4719), .A2(n4718), .ZN(n4417) );
  AND2_X1 U5984 ( .A1(n8939), .A2(n4354), .ZN(n4418) );
  OR2_X1 U5985 ( .A1(n5041), .A2(n5040), .ZN(n4419) );
  NOR2_X1 U5986 ( .A1(n9270), .A2(n9271), .ZN(n4420) );
  INV_X1 U5987 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5236) );
  INV_X1 U5988 ( .A(n5184), .ZN(n4783) );
  NAND2_X1 U5989 ( .A1(n5437), .A2(n5355), .ZN(n5358) );
  AND2_X1 U5990 ( .A1(n6425), .A2(n4700), .ZN(n4421) );
  OR2_X1 U5991 ( .A1(n4816), .A2(n8329), .ZN(n4422) );
  INV_X1 U5992 ( .A(n4686), .ZN(n4685) );
  NOR2_X1 U5993 ( .A1(n5870), .A2(n4687), .ZN(n4686) );
  AND2_X1 U5994 ( .A1(n4796), .A2(n4683), .ZN(n4423) );
  AND2_X1 U5995 ( .A1(n5965), .A2(n4941), .ZN(n4424) );
  AND2_X1 U5996 ( .A1(n4722), .A2(n6028), .ZN(n4425) );
  INV_X1 U5997 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4649) );
  INV_X1 U5998 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4652) );
  OAI21_X1 U5999 ( .B1(n7579), .B2(n5283), .A(n5282), .ZN(n7599) );
  NAND2_X1 U6000 ( .A1(n7769), .A2(n5434), .ZN(n7938) );
  OR2_X1 U6001 ( .A1(n4869), .A2(n5179), .ZN(n4426) );
  NOR2_X1 U6002 ( .A1(n7973), .A2(n4541), .ZN(n4427) );
  NOR2_X1 U6003 ( .A1(n7682), .A2(n9720), .ZN(n5884) );
  OR2_X1 U6004 ( .A1(n9016), .A2(n4576), .ZN(n4428) );
  AND2_X1 U6005 ( .A1(n5815), .A2(n5814), .ZN(n5936) );
  INV_X1 U6006 ( .A(n5936), .ZN(n4837) );
  AOI21_X1 U6007 ( .B1(n7716), .B2(n4934), .A(n4933), .ZN(n7996) );
  OAI21_X1 U6008 ( .B1(n9016), .B2(n8681), .A(n8683), .ZN(n9005) );
  NAND2_X1 U6009 ( .A1(n4474), .A2(n4480), .ZN(n9187) );
  NAND2_X1 U6010 ( .A1(n4681), .A2(n5853), .ZN(n7823) );
  NAND2_X1 U6011 ( .A1(n4854), .A2(n5383), .ZN(n7542) );
  INV_X1 U6012 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4923) );
  OR2_X1 U6013 ( .A1(n9742), .A2(n9285), .ZN(n4429) );
  NOR3_X1 U6014 ( .A1(n7824), .A2(n9615), .A3(n4761), .ZN(n4758) );
  NOR2_X1 U6015 ( .A1(n10082), .A2(n8790), .ZN(n4430) );
  INV_X1 U6016 ( .A(n4555), .ZN(n4554) );
  OAI21_X1 U6017 ( .B1(n7731), .B2(n4365), .A(n4556), .ZN(n4555) );
  NOR2_X1 U6018 ( .A1(n4481), .A2(n4475), .ZN(n4431) );
  INV_X1 U6019 ( .A(n4759), .ZN(n9626) );
  NOR2_X1 U6020 ( .A1(n7824), .A2(n4761), .ZN(n4759) );
  AND2_X1 U6021 ( .A1(n4614), .A2(n4613), .ZN(n4432) );
  AND3_X1 U6022 ( .A1(n6235), .A2(n6234), .A3(n6233), .ZN(n8488) );
  AND2_X1 U6023 ( .A1(n4805), .A2(n8105), .ZN(n4433) );
  INV_X1 U6024 ( .A(n4553), .ZN(n4552) );
  AOI21_X1 U6025 ( .B1(n4554), .B2(n4365), .A(n4557), .ZN(n4553) );
  AND2_X1 U6026 ( .A1(n5496), .A2(n7147), .ZN(n4434) );
  INV_X1 U6027 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6029) );
  INV_X1 U6028 ( .A(n5868), .ZN(n4687) );
  AND2_X1 U6029 ( .A1(n5548), .A2(n5551), .ZN(n4435) );
  OR2_X1 U6030 ( .A1(n9570), .A2(n5862), .ZN(n4436) );
  OR2_X1 U6031 ( .A1(n5496), .A2(n7147), .ZN(n4437) );
  OR2_X1 U6032 ( .A1(n5617), .A2(n7110), .ZN(n4438) );
  AND2_X1 U6033 ( .A1(n4435), .A2(n5552), .ZN(n4439) );
  AND2_X1 U6034 ( .A1(n4940), .A2(n4377), .ZN(n4440) );
  XNOR2_X1 U6035 ( .A(n4989), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5779) );
  INV_X1 U6036 ( .A(n10074), .ZN(n4730) );
  NAND2_X1 U6037 ( .A1(n6816), .A2(n9630), .ZN(n9633) );
  NAND2_X1 U6038 ( .A1(n5388), .A2(n5387), .ZN(n7549) );
  INV_X1 U6039 ( .A(n7549), .ZN(n4752) );
  INV_X1 U6040 ( .A(n9988), .ZN(n9986) );
  NAND2_X1 U6041 ( .A1(n6939), .A2(n9964), .ZN(n4441) );
  OAI21_X1 U6042 ( .B1(n7518), .B2(n7698), .A(n6316), .ZN(n7716) );
  INV_X1 U6043 ( .A(n8437), .ZN(n4708) );
  AND2_X1 U6044 ( .A1(n4583), .A2(n4582), .ZN(n4442) );
  INV_X1 U6045 ( .A(n8457), .ZN(n4677) );
  INV_X1 U6046 ( .A(n8237), .ZN(n4804) );
  XNOR2_X1 U6047 ( .A(n6351), .B(n6354), .ZN(n6364) );
  NAND2_X1 U6048 ( .A1(n4846), .A2(n4845), .ZN(n6766) );
  OR2_X1 U6049 ( .A1(n6363), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6398) );
  INV_X1 U6050 ( .A(n8800), .ZN(n4540) );
  AND2_X1 U6051 ( .A1(n5840), .A2(n6912), .ZN(n4443) );
  AND2_X1 U6052 ( .A1(n4606), .A2(n4605), .ZN(n4444) );
  NOR2_X1 U6053 ( .A1(n8801), .A2(n8830), .ZN(n4445) );
  AND2_X1 U6054 ( .A1(n5760), .A2(n7144), .ZN(n4446) );
  NAND2_X1 U6055 ( .A1(n6353), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6378) );
  AND2_X1 U6056 ( .A1(n4585), .A2(n4584), .ZN(n4447) );
  NAND2_X1 U6057 ( .A1(n4597), .A2(n8595), .ZN(n7236) );
  NAND2_X1 U6058 ( .A1(n5060), .A2(n5064), .ZN(n6657) );
  AND2_X1 U6059 ( .A1(n7427), .A2(n7429), .ZN(n4448) );
  AND2_X1 U6060 ( .A1(n7977), .A2(n7988), .ZN(n4449) );
  INV_X1 U6061 ( .A(n9968), .ZN(n4763) );
  NAND2_X1 U6062 ( .A1(n5035), .A2(n4485), .ZN(n6805) );
  INV_X1 U6063 ( .A(n7428), .ZN(n4738) );
  AND2_X1 U6064 ( .A1(n8816), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n4450) );
  AND2_X1 U6065 ( .A1(n4596), .A2(n8595), .ZN(n4451) );
  NAND2_X1 U6066 ( .A1(n7445), .A2(n7743), .ZN(n10029) );
  INV_X1 U6067 ( .A(SI_13_), .ZN(n4834) );
  NAND2_X1 U6068 ( .A1(n4735), .A2(n7348), .ZN(n7349) );
  AND2_X1 U6069 ( .A1(n6612), .A2(n4367), .ZN(n4452) );
  NOR2_X2 U6070 ( .A1(n6515), .A2(n6514), .ZN(n8527) );
  OR2_X1 U6071 ( .A1(n6508), .A2(n6638), .ZN(n6515) );
  OR2_X2 U6072 ( .A1(n7248), .A2(n8324), .ZN(n9682) );
  NAND2_X1 U6073 ( .A1(n7876), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U6074 ( .A1(n10044), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U6075 ( .A1(n8844), .A2(n4524), .ZN(n4523) );
  NAND2_X1 U6076 ( .A1(n4529), .A2(n4522), .ZN(P2_U3201) );
  NAND3_X1 U6077 ( .A1(n4957), .A2(n4984), .A3(n4453), .ZN(n4679) );
  AND4_X2 U6078 ( .A1(n4358), .A2(n5176), .A3(n4980), .A4(n4414), .ZN(n4984)
         );
  AND3_X2 U6079 ( .A1(n4964), .A2(n5119), .A3(n5083), .ZN(n5176) );
  OAI21_X1 U6080 ( .B1(n5851), .B2(n4461), .A(n4459), .ZN(n4681) );
  NAND2_X1 U6081 ( .A1(n4457), .A2(n4456), .ZN(n5855) );
  NAND2_X1 U6082 ( .A1(n5851), .A2(n4459), .ZN(n4457) );
  NAND3_X1 U6083 ( .A1(n4463), .A2(n4464), .A3(n4462), .ZN(n6877) );
  NAND3_X1 U6084 ( .A1(n5840), .A2(n6937), .A3(n6912), .ZN(n4462) );
  NAND2_X1 U6085 ( .A1(n4891), .A2(n4468), .ZN(n4467) );
  OAI21_X2 U6086 ( .B1(n9242), .B2(n9246), .A(n9179), .ZN(n9225) );
  AND2_X2 U6087 ( .A1(n4470), .A2(n5636), .ZN(n9246) );
  INV_X1 U6088 ( .A(n5547), .ZN(n4482) );
  AND2_X2 U6089 ( .A1(n4859), .A2(n4858), .ZN(n9269) );
  NAND2_X1 U6090 ( .A1(n4488), .A2(n4413), .ZN(n8089) );
  AND2_X1 U6091 ( .A1(n8087), .A2(n8086), .ZN(n4489) );
  MUX2_X1 U6092 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5716), .Z(n5122) );
  INV_X1 U6093 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4493) );
  NAND4_X1 U6094 ( .A1(n4497), .A2(n4422), .A3(n4819), .A4(n4494), .ZN(
        P1_U3242) );
  OAI21_X1 U6095 ( .B1(n8255), .B2(n4496), .A(n4495), .ZN(n4494) );
  NAND2_X1 U6096 ( .A1(n4499), .A2(n4498), .ZN(n4497) );
  OAI21_X1 U6097 ( .B1(n8255), .B2(n8254), .A(n8264), .ZN(n4499) );
  NAND2_X1 U6098 ( .A1(n8112), .A2(n4503), .ZN(n4500) );
  NAND2_X1 U6099 ( .A1(n4500), .A2(n4501), .ZN(n8104) );
  NAND2_X1 U6100 ( .A1(n8136), .A2(n4516), .ZN(n4515) );
  NAND2_X1 U6101 ( .A1(n4510), .A2(n4511), .ZN(n8155) );
  AOI21_X1 U6102 ( .B1(n4512), .B2(n4513), .A(n8188), .ZN(n4511) );
  NAND3_X1 U6103 ( .A1(n8819), .A2(n8818), .A3(n4528), .ZN(n4527) );
  NAND2_X1 U6104 ( .A1(n4532), .A2(n4533), .ZN(n10063) );
  NAND2_X1 U6105 ( .A1(n7973), .A2(n4534), .ZN(n4532) );
  AND2_X1 U6106 ( .A1(n7974), .A2(n7975), .ZN(n4541) );
  NOR2_X1 U6107 ( .A1(n7733), .A2(n10026), .ZN(n4557) );
  AND3_X2 U6108 ( .A1(n6028), .A2(n4941), .A3(n4564), .ZN(n6288) );
  NAND4_X1 U6109 ( .A1(n6028), .A2(n4941), .A3(n4564), .A4(n5964), .ZN(n6359)
         );
  MUX2_X1 U6110 ( .A(P2_REG1_REG_0__SCAN_IN), .B(P2_REG2_REG_0__SCAN_IN), .S(
        n8811), .Z(n7457) );
  OAI21_X2 U6111 ( .B1(n8941), .B2(n4591), .A(n4588), .ZN(n8880) );
  NAND3_X1 U6112 ( .A1(n4590), .A2(n4592), .A3(n8726), .ZN(n4589) );
  NAND3_X1 U6113 ( .A1(n5980), .A2(n8599), .A3(n6821), .ZN(n4597) );
  NAND2_X1 U6114 ( .A1(n5980), .A2(n6821), .ZN(n8594) );
  NAND2_X1 U6115 ( .A1(n8595), .A2(n8599), .ZN(n7463) );
  NAND3_X1 U6116 ( .A1(n4733), .A2(n7349), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n9990) );
  NOR2_X1 U6117 ( .A1(n10084), .A2(n10083), .ZN(n10082) );
  OAI211_X1 U6118 ( .C1(n8790), .C2(P2_REG2_REG_15__SCAN_IN), .A(n4599), .B(
        n4602), .ZN(n4601) );
  NAND2_X1 U6119 ( .A1(n4600), .A2(n10084), .ZN(n4599) );
  INV_X1 U6120 ( .A(n8790), .ZN(n4600) );
  INV_X1 U6121 ( .A(n4601), .ZN(n10099) );
  INV_X1 U6122 ( .A(n10100), .ZN(n4602) );
  XNOR2_X1 U6123 ( .A(n7967), .B(n7975), .ZN(n7881) );
  OAI21_X1 U6124 ( .B1(n7723), .B2(n4610), .A(n4608), .ZN(n4729) );
  XNOR2_X1 U6125 ( .A(n8786), .B(n10042), .ZN(n10052) );
  OAI21_X1 U6126 ( .B1(n4612), .B2(n10052), .A(n4611), .ZN(n10067) );
  NAND2_X1 U6127 ( .A1(n8701), .A2(n4624), .ZN(n4627) );
  NAND3_X1 U6128 ( .A1(n4627), .A2(n8716), .A3(n8717), .ZN(n4626) );
  NAND2_X1 U6129 ( .A1(n4628), .A2(n8667), .ZN(n8672) );
  NAND2_X1 U6130 ( .A1(n4630), .A2(n8747), .ZN(n4629) );
  INV_X1 U6131 ( .A(n4631), .ZN(n4630) );
  AOI21_X1 U6132 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n4631) );
  AOI21_X1 U6133 ( .B1(n8659), .B2(n8653), .A(n8652), .ZN(n4632) );
  NOR2_X2 U6134 ( .A1(n8740), .A2(n4637), .ZN(n8749) );
  NAND2_X1 U6135 ( .A1(n10187), .A2(n8779), .ZN(n8632) );
  AOI21_X2 U6136 ( .B1(n6592), .B2(n8544), .A(n4638), .ZN(n10187) );
  NAND2_X1 U6137 ( .A1(n5185), .A2(n4360), .ZN(n4640) );
  NAND2_X1 U6138 ( .A1(n5185), .A2(n5184), .ZN(n5312) );
  NAND3_X1 U6139 ( .A1(n4640), .A2(n4639), .A3(n5285), .ZN(n5234) );
  NAND2_X1 U6140 ( .A1(n4645), .A2(n4641), .ZN(n8709) );
  NAND3_X1 U6141 ( .A1(n4643), .A2(n8697), .A3(n8987), .ZN(n4642) );
  NAND3_X1 U6142 ( .A1(n4651), .A2(n4650), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n4646) );
  NAND3_X1 U6143 ( .A1(n4654), .A2(n4653), .A3(n4656), .ZN(n8376) );
  OR2_X2 U6144 ( .A1(n6471), .A2(n6470), .ZN(n4656) );
  NAND2_X1 U6145 ( .A1(n5467), .A2(n4667), .ZN(n4666) );
  NAND3_X1 U6146 ( .A1(n4984), .A2(n4368), .A3(n4957), .ZN(n5020) );
  NAND2_X1 U6147 ( .A1(n4455), .A2(n4686), .ZN(n4682) );
  NAND2_X1 U6148 ( .A1(n4682), .A2(n4423), .ZN(n5931) );
  NAND2_X1 U6149 ( .A1(n4880), .A2(n4879), .ZN(n9518) );
  NAND2_X1 U6150 ( .A1(n5627), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4689) );
  NAND2_X1 U6151 ( .A1(n9986), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4692) );
  NAND2_X1 U6152 ( .A1(n4695), .A2(n4694), .ZN(n4696) );
  INV_X1 U6153 ( .A(n7200), .ZN(n4694) );
  INV_X1 U6154 ( .A(n4696), .ZN(n7199) );
  XNOR2_X1 U6155 ( .A(n6407), .B(n10130), .ZN(n7201) );
  OAI22_X1 U6156 ( .A1(n6868), .A2(n6869), .B1(n6403), .B2(n8782), .ZN(n7200)
         );
  NAND2_X1 U6157 ( .A1(n4697), .A2(n4421), .ZN(n6428) );
  NAND2_X1 U6158 ( .A1(n7893), .A2(n4698), .ZN(n4697) );
  NAND2_X1 U6159 ( .A1(n8425), .A2(n4702), .ZN(n4706) );
  NAND3_X1 U6160 ( .A1(n4704), .A2(n4706), .A3(n8481), .ZN(n8484) );
  NAND2_X1 U6162 ( .A1(n6291), .A2(n4714), .ZN(n6353) );
  NAND2_X1 U6163 ( .A1(n7271), .A2(n4417), .ZN(n4715) );
  NAND2_X1 U6164 ( .A1(n4715), .A2(n4716), .ZN(n7910) );
  INV_X1 U6165 ( .A(n4721), .ZN(n7504) );
  MUX2_X1 U6166 ( .A(n8634), .B(n8633), .S(n8747), .Z(n8645) );
  NAND2_X1 U6167 ( .A1(n5864), .A2(n4882), .ZN(n4880) );
  XNOR2_X2 U6168 ( .A(n4727), .B(P2_IR_REG_2__SCAN_IN), .ZN(n7487) );
  NOR2_X1 U6169 ( .A1(n7791), .A2(n7624), .ZN(n7792) );
  NAND2_X1 U6170 ( .A1(n7496), .A2(n7347), .ZN(n4735) );
  INV_X1 U6171 ( .A(n7348), .ZN(n4734) );
  INV_X1 U6172 ( .A(n7429), .ZN(n4737) );
  NAND2_X1 U6173 ( .A1(n4741), .A2(n10029), .ZN(n7723) );
  NAND2_X1 U6174 ( .A1(n7444), .A2(n7730), .ZN(n4742) );
  AND2_X1 U6175 ( .A1(n4742), .A2(n10029), .ZN(n7446) );
  NOR2_X1 U6176 ( .A1(n9485), .A2(n4749), .ZN(n9465) );
  NOR2_X1 U6177 ( .A1(n9485), .A2(n8151), .ZN(n5942) );
  INV_X1 U6178 ( .A(n4758), .ZN(n9614) );
  NAND2_X1 U6179 ( .A1(n9606), .A2(n4775), .ZN(n4772) );
  NAND2_X1 U6180 ( .A1(n4772), .A2(n4773), .ZN(n9580) );
  OAI21_X1 U6181 ( .B1(n5185), .B2(n4784), .A(n4371), .ZN(n5265) );
  NAND2_X1 U6182 ( .A1(n4781), .A2(n4779), .ZN(n5267) );
  NAND2_X1 U6183 ( .A1(n5185), .A2(n4371), .ZN(n4781) );
  NAND2_X1 U6184 ( .A1(n9509), .A2(n4786), .ZN(n4785) );
  OAI211_X1 U6185 ( .C1(n9509), .C2(n4791), .A(n4788), .B(n4785), .ZN(n5903)
         );
  NAND2_X1 U6186 ( .A1(n9509), .A2(n8190), .ZN(n9492) );
  AOI21_X1 U6187 ( .B1(n5893), .B2(n8095), .A(n4798), .ZN(n5892) );
  OAI21_X1 U6188 ( .B1(n7557), .B2(n4802), .A(n4800), .ZN(n7830) );
  INV_X1 U6189 ( .A(n4809), .ZN(n5638) );
  INV_X1 U6190 ( .A(n5597), .ZN(n4815) );
  NOR2_X1 U6191 ( .A1(n8257), .A2(n4485), .ZN(n4817) );
  NAND2_X1 U6192 ( .A1(n5357), .A2(n4362), .ZN(n4826) );
  NAND2_X1 U6193 ( .A1(n5128), .A2(n5127), .ZN(n4835) );
  NAND3_X1 U6194 ( .A1(n4835), .A2(n4383), .A3(n5151), .ZN(n5154) );
  NAND2_X1 U6195 ( .A1(n4838), .A2(n5878), .ZN(n5883) );
  NAND2_X1 U6196 ( .A1(n5206), .A2(SI_0_), .ZN(n5950) );
  MUX2_X1 U6197 ( .A(n8345), .B(n8534), .S(n4840), .Z(n8024) );
  MUX2_X1 U6198 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4840), .Z(n8029) );
  NAND2_X1 U6199 ( .A1(n7768), .A2(n4842), .ZN(n4841) );
  OAI21_X1 U6200 ( .B1(n4848), .B2(n4847), .A(n6720), .ZN(n4846) );
  INV_X1 U6201 ( .A(n5165), .ZN(n4850) );
  NAND2_X1 U6202 ( .A1(n4851), .A2(n5165), .ZN(n6567) );
  NAND2_X1 U6203 ( .A1(n7374), .A2(n4855), .ZN(n4853) );
  INV_X1 U6204 ( .A(n5179), .ZN(n4868) );
  NAND3_X1 U6205 ( .A1(n4868), .A2(n4969), .A3(n4867), .ZN(n4971) );
  NAND3_X1 U6206 ( .A1(n4868), .A2(n4969), .A3(n4871), .ZN(n5408) );
  NAND2_X1 U6207 ( .A1(n6767), .A2(n4872), .ZN(n6799) );
  INV_X1 U6208 ( .A(n4877), .ZN(n9244) );
  NAND2_X1 U6209 ( .A1(n7925), .A2(n4892), .ZN(n4891) );
  NAND2_X1 U6210 ( .A1(n4984), .A2(n4983), .ZN(n4986) );
  AND2_X2 U6211 ( .A1(n4984), .A2(n4898), .ZN(n4997) );
  NAND2_X1 U6212 ( .A1(n8930), .A2(n4904), .ZN(n4903) );
  NAND2_X1 U6213 ( .A1(n9006), .A2(n4910), .ZN(n4909) );
  INV_X1 U6214 ( .A(n8783), .ZN(n4928) );
  OAI21_X1 U6215 ( .B1(n8890), .B2(n4931), .A(n4929), .ZN(n8872) );
  OR2_X1 U6216 ( .A1(n8890), .A2(n8725), .ZN(n8891) );
  NAND2_X1 U6217 ( .A1(n6101), .A2(n4424), .ZN(n5966) );
  NAND2_X1 U6218 ( .A1(n6101), .A2(n5954), .ZN(n6105) );
  NAND2_X1 U6219 ( .A1(n6706), .A2(n6711), .ZN(n6705) );
  OAI21_X1 U6220 ( .B1(n5716), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n5220), .ZN(
        n5221) );
  OAI21_X1 U6221 ( .B1(n8856), .B2(n8858), .A(n8857), .ZN(n9092) );
  INV_X1 U6222 ( .A(n6472), .ZN(n8447) );
  OAI21_X1 U6223 ( .B1(n8958), .B2(n6206), .A(n8708), .ZN(n8944) );
  NOR2_X1 U6224 ( .A1(n8482), .A2(n8403), .ZN(n4943) );
  OR2_X2 U6225 ( .A1(n9574), .A2(n9562), .ZN(n4944) );
  AND2_X1 U6226 ( .A1(n6418), .A2(n7908), .ZN(n4945) );
  INV_X1 U6227 ( .A(n8570), .ZN(n6081) );
  NAND2_X1 U6228 ( .A1(n8398), .A2(n8397), .ZN(n4946) );
  NAND2_X1 U6229 ( .A1(n5576), .A2(n9188), .ZN(n9233) );
  NAND2_X1 U6230 ( .A1(n5970), .A2(n5968), .ZN(n4947) );
  NAND2_X1 U6231 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n4948) );
  AND2_X1 U6232 ( .A1(n5351), .A2(n5350), .ZN(n4949) );
  NOR2_X1 U6233 ( .A1(n5839), .A2(n6780), .ZN(n4950) );
  OR2_X1 U6234 ( .A1(n6611), .A2(n9316), .ZN(n4951) );
  NOR2_X1 U6235 ( .A1(n6545), .A2(n9118), .ZN(n4952) );
  NOR2_X1 U6236 ( .A1(n4947), .A2(n4942), .ZN(n4953) );
  OR2_X1 U6237 ( .A1(n5351), .A2(n5350), .ZN(n4954) );
  AND2_X1 U6238 ( .A1(n5445), .A2(n5468), .ZN(n4955) );
  AND2_X1 U6239 ( .A1(n5285), .A2(n5223), .ZN(n4956) );
  AND2_X1 U6240 ( .A1(n5004), .A2(n5003), .ZN(n4957) );
  INV_X1 U6241 ( .A(n5885), .ZN(n9485) );
  OR2_X1 U6242 ( .A1(n5036), .A2(n5058), .ZN(n4959) );
  OR2_X1 U6243 ( .A1(n6563), .A2(n10026), .ZN(n4960) );
  NAND2_X1 U6244 ( .A1(n5285), .A2(n5284), .ZN(n4961) );
  INV_X1 U6245 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6604) );
  OR2_X1 U6246 ( .A1(n6413), .A2(n7595), .ZN(n4962) );
  AND3_X1 U6247 ( .A1(n6494), .A2(n8507), .A3(n6493), .ZN(n4963) );
  INV_X2 U6248 ( .A(n10207), .ZN(n10205) );
  AND3_X2 U6249 ( .A1(n6543), .A2(n6542), .A3(n6541), .ZN(n10225) );
  AND2_X1 U6250 ( .A1(n6388), .A2(n8977), .ZN(n10146) );
  INV_X1 U6251 ( .A(n9770), .ZN(n5926) );
  INV_X1 U6252 ( .A(n9717), .ZN(n5919) );
  INV_X1 U6253 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4976) );
  INV_X1 U6254 ( .A(n5349), .ZN(n5351) );
  NAND2_X1 U6255 ( .A1(n8741), .A2(n8548), .ZN(n8549) );
  INV_X1 U6256 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5954) );
  OAI22_X1 U6257 ( .A1(n6750), .A2(n5061), .B1(n6735), .B2(n5086), .ZN(n5087)
         );
  NAND2_X1 U6258 ( .A1(n4349), .A2(n5219), .ZN(n5220) );
  AND2_X1 U6259 ( .A1(n7700), .A2(n6315), .ZN(n6316) );
  OAI22_X1 U6260 ( .A1(n8905), .A2(n6326), .B1(n8922), .B2(n8456), .ZN(n8890)
         );
  NAND2_X1 U6261 ( .A1(n6189), .A2(n5997), .ZN(n5998) );
  INV_X1 U6262 ( .A(n5562), .ZN(n5560) );
  INV_X1 U6263 ( .A(n5478), .ZN(n5453) );
  INV_X1 U6264 ( .A(n5258), .ZN(n5241) );
  NAND2_X1 U6265 ( .A1(n4971), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5498) );
  NOR2_X1 U6266 ( .A1(n5286), .A2(n4961), .ZN(n5311) );
  OR2_X1 U6267 ( .A1(n6049), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6061) );
  INV_X1 U6268 ( .A(n8552), .ZN(n8553) );
  AOI21_X1 U6269 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8827), .A(n8785), .ZN(
        n8786) );
  OR2_X1 U6270 ( .A1(n6138), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6152) );
  INV_X1 U6271 ( .A(n6340), .ZN(n6341) );
  OAI211_X1 U6272 ( .C1(n6605), .C2(n5993), .A(n6068), .B(n4960), .ZN(n7632)
         );
  NAND2_X1 U6273 ( .A1(n5166), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5198) );
  OR2_X1 U6274 ( .A1(n5696), .A2(n5695), .ZN(n5721) );
  OR2_X1 U6275 ( .A1(n5535), .A2(n5534), .ZN(n5562) );
  OR2_X1 U6276 ( .A1(n9819), .A2(n9818), .ZN(n9821) );
  INV_X1 U6277 ( .A(n9734), .ZN(n9458) );
  NAND2_X1 U6278 ( .A1(n5560), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U6279 ( .A1(n5502), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5535) );
  OR2_X1 U6280 ( .A1(n5390), .A2(n5389), .ZN(n5421) );
  OR2_X1 U6281 ( .A1(n5324), .A2(n5323), .ZN(n5326) );
  NAND2_X1 U6282 ( .A1(n9297), .A2(n6981), .ZN(n8275) );
  INV_X1 U6283 ( .A(n5358), .ZN(n5356) );
  NAND2_X1 U6284 ( .A1(n5221), .A2(n7028), .ZN(n5285) );
  OR2_X1 U6285 ( .A1(n6408), .A2(n8618), .ZN(n6409) );
  OR2_X1 U6286 ( .A1(n6238), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6244) );
  AND2_X1 U6287 ( .A1(n6071), .A2(n6070), .ZN(n6086) );
  AND2_X1 U6288 ( .A1(n9080), .A2(n8758), .ZN(n8759) );
  OR2_X1 U6289 ( .A1(n6281), .A2(n7306), .ZN(n6005) );
  XNOR2_X1 U6290 ( .A(n7487), .B(n7344), .ZN(n7498) );
  NAND2_X1 U6291 ( .A1(n7410), .A2(n7409), .ZN(n7437) );
  AOI21_X1 U6292 ( .B1(n8814), .B2(n8817), .A(n10004), .ZN(n8815) );
  NOR2_X1 U6293 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n6271), .ZN(n8849) );
  OR2_X1 U6294 ( .A1(n6231), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6238) );
  AND2_X1 U6295 ( .A1(n6209), .A2(n8406), .ZN(n6219) );
  INV_X1 U6296 ( .A(n8775), .ZN(n8670) );
  NAND2_X1 U6297 ( .A1(n7778), .A2(n8544), .ZN(n6260) );
  OR2_X1 U6298 ( .A1(n9062), .A2(n8498), .ZN(n8697) );
  AND2_X1 U6299 ( .A1(n9224), .A2(n5659), .ZN(n9179) );
  AND2_X1 U6300 ( .A1(n5738), .A2(n5737), .ZN(n6550) );
  INV_X1 U6301 ( .A(n8248), .ZN(n5929) );
  AND2_X1 U6302 ( .A1(n8303), .A2(n8156), .ZN(n9493) );
  AND2_X1 U6303 ( .A1(n8137), .A2(n9543), .ZN(n9558) );
  AND2_X1 U6304 ( .A1(n8195), .A2(n8131), .ZN(n9591) );
  INV_X1 U6305 ( .A(n9616), .ZN(n7290) );
  INV_X1 U6306 ( .A(n5883), .ZN(n9479) );
  OR2_X1 U6307 ( .A1(n6748), .A2(n6918), .ZN(n6913) );
  INV_X1 U6308 ( .A(n9644), .ZN(n9551) );
  INV_X1 U6309 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U6310 ( .A1(n5218), .A2(SI_7_), .ZN(n5266) );
  NAND2_X1 U6311 ( .A1(n5182), .A2(n5181), .ZN(n5185) );
  OR3_X1 U6312 ( .A1(n6364), .A2(n6361), .A3(n7764), .ZN(n6566) );
  NAND2_X1 U6313 ( .A1(n6520), .A2(n6519), .ZN(n6521) );
  NAND2_X1 U6314 ( .A1(n6498), .A2(n8977), .ZN(n8478) );
  OR2_X1 U6315 ( .A1(n6096), .A2(n6389), .ZN(n8543) );
  AND4_X1 U6316 ( .A1(n6226), .A2(n6225), .A3(n6224), .A4(n6223), .ZN(n8921)
         );
  AND4_X1 U6317 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n8662)
         );
  AOI21_X1 U6318 ( .B1(n9797), .B2(n9796), .A(n10122), .ZN(n9798) );
  OR2_X1 U6319 ( .A1(n6261), .A2(n6252), .ZN(n8886) );
  INV_X1 U6320 ( .A(n8394), .ZN(n9062) );
  INV_X1 U6321 ( .A(n9026), .ZN(n10142) );
  OR2_X1 U6322 ( .A1(n6487), .A2(n6639), .ZN(n6541) );
  INV_X1 U6323 ( .A(n10186), .ZN(n10200) );
  OR2_X1 U6324 ( .A1(n6530), .A2(n6529), .ZN(n6534) );
  INV_X1 U6325 ( .A(n9250), .ZN(n9279) );
  INV_X1 U6326 ( .A(n9280), .ZN(n9513) );
  OR2_X1 U6327 ( .A1(n5426), .A2(n5425), .ZN(n7943) );
  AND2_X1 U6328 ( .A1(n8153), .A2(n8190), .ZN(n9511) );
  AND2_X1 U6329 ( .A1(n8185), .A2(n8198), .ZN(n9545) );
  AND2_X1 U6330 ( .A1(n9636), .A2(n8051), .ZN(n7927) );
  AND2_X1 U6331 ( .A1(n8124), .A2(n8105), .ZN(n8235) );
  INV_X1 U6332 ( .A(n9469), .ZN(n7692) );
  AND2_X1 U6333 ( .A1(n5036), .A2(n6560), .ZN(n6613) );
  AND2_X1 U6334 ( .A1(n5272), .A2(n5271), .ZN(n9430) );
  NOR2_X1 U6335 ( .A1(n6566), .A2(n7318), .ZN(n7355) );
  INV_X1 U6336 ( .A(n8507), .ZN(n8518) );
  INV_X1 U6337 ( .A(n8478), .ZN(n8530) );
  INV_X1 U6338 ( .A(n8431), .ZN(n9008) );
  INV_X1 U6339 ( .A(n10010), .ZN(n10122) );
  INV_X1 U6340 ( .A(n6546), .ZN(n6547) );
  INV_X1 U6341 ( .A(n10225), .ZN(n10222) );
  NAND2_X1 U6342 ( .A1(n10205), .A2(n10198), .ZN(n9164) );
  AND2_X1 U6343 ( .A1(n6534), .A2(n6533), .ZN(n10207) );
  AND2_X1 U6344 ( .A1(n6565), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6764) );
  INV_X1 U6345 ( .A(n8592), .ZN(n6928) );
  AND2_X1 U6346 ( .A1(n5824), .A2(n8329), .ZN(n9260) );
  AND2_X1 U6347 ( .A1(n5807), .A2(n9630), .ZN(n9285) );
  INV_X1 U6348 ( .A(n9274), .ZN(n9267) );
  OR2_X1 U6349 ( .A1(n5566), .A2(n5565), .ZN(n9610) );
  INV_X1 U6350 ( .A(n6750), .ZN(n9299) );
  NAND2_X1 U6351 ( .A1(n5883), .A2(n5919), .ZN(n5920) );
  NAND2_X1 U6352 ( .A1(n5883), .A2(n5926), .ZN(n5927) );
  INV_X1 U6353 ( .A(n9981), .ZN(n9980) );
  INV_X1 U6354 ( .A(n9301), .ZN(P1_U3973) );
  NAND2_X1 U6355 ( .A1(n4406), .A2(n5949), .ZN(P1_U3550) );
  OAI21_X1 U6356 ( .B1(n5947), .B2(n9980), .A(n5946), .ZN(P1_U3518) );
  NOR2_X1 U6357 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4964) );
  NAND2_X1 U6358 ( .A1(n5176), .A2(n4965), .ZN(n5179) );
  NOR2_X1 U6359 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5409) );
  NOR2_X1 U6360 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4968) );
  NOR2_X1 U6361 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4967) );
  INV_X1 U6362 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4966) );
  AND4_X1 U6363 ( .A1(n5409), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n4969)
         );
  INV_X1 U6364 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U6365 ( .A1(n5498), .A2(n4972), .ZN(n4973) );
  INV_X1 U6366 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U6367 ( .A1(n5529), .A2(n5528), .ZN(n5531) );
  INV_X1 U6368 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4974) );
  NOR2_X2 U6369 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5317) );
  NOR2_X1 U6370 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4979) );
  NOR2_X1 U6371 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4978) );
  NOR2_X1 U6372 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4977) );
  NAND2_X1 U6373 ( .A1(n4981), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4982) );
  NAND2_X1 U6374 ( .A1(n4986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U6375 ( .A1(n4402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5799) );
  XNOR2_X1 U6376 ( .A(n5799), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U6377 ( .A1(n4987), .A2(n5880), .ZN(n4996) );
  NOR2_X1 U6378 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5004) );
  NAND2_X1 U6379 ( .A1(n4997), .A2(n4988), .ZN(n4992) );
  INV_X1 U6380 ( .A(n4997), .ZN(n4990) );
  NAND2_X1 U6381 ( .A1(n4990), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4991) );
  MUX2_X1 U6382 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4991), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n4993) );
  NAND2_X1 U6383 ( .A1(n4994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4995) );
  XNOR2_X1 U6384 ( .A(n4995), .B(P1_IR_REG_24__SCAN_IN), .ZN(n7552) );
  NOR2_X1 U6385 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5000) );
  NAND2_X1 U6386 ( .A1(n4997), .A2(n5000), .ZN(n4998) );
  NAND2_X1 U6387 ( .A1(n5001), .A2(n5000), .ZN(n5002) );
  NOR2_X1 U6388 ( .A1(n5002), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5003) );
  INV_X1 U6389 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5005) );
  INV_X1 U6390 ( .A(SI_1_), .ZN(n5007) );
  INV_X1 U6391 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5009) );
  AND2_X1 U6392 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6393 ( .A1(n5716), .A2(n5008), .ZN(n5050) );
  OAI21_X1 U6394 ( .B1(n5950), .B2(n5009), .A(n5050), .ZN(n5077) );
  XNOR2_X1 U6395 ( .A(n5078), .B(n5077), .ZN(n6580) );
  OR2_X1 U6396 ( .A1(n5110), .A2(n6580), .ZN(n5013) );
  INV_X1 U6397 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U6398 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5010) );
  XNOR2_X1 U6399 ( .A(n5011), .B(n5010), .ZN(n6668) );
  OR2_X1 U6400 ( .A1(n5052), .A2(n6668), .ZN(n5012) );
  NAND2_X1 U6401 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5015) );
  INV_X1 U6402 ( .A(n5020), .ZN(n5022) );
  NOR3_X1 U6403 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .A3(
        P1_IR_REG_30__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U6404 ( .A1(n5022), .A2(n5021), .ZN(n9778) );
  INV_X1 U6405 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5024) );
  INV_X1 U6406 ( .A(n5028), .ZN(n8016) );
  OR2_X2 U6407 ( .A1(n8344), .A2(n8016), .ZN(n5069) );
  INV_X1 U6408 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9303) );
  INV_X1 U6409 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5026) );
  OR2_X1 U6410 ( .A1(n5095), .A2(n5026), .ZN(n5027) );
  OAI21_X1 U6411 ( .B1(n5069), .B2(n9303), .A(n5027), .ZN(n5033) );
  OR2_X1 U6412 ( .A1(n8344), .A2(n5028), .ZN(n5094) );
  INV_X1 U6413 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5031) );
  INV_X1 U6414 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5029) );
  OR2_X1 U6415 ( .A1(n5097), .A2(n5029), .ZN(n5030) );
  OAI21_X1 U6416 ( .B1(n5094), .B2(n5031), .A(n5030), .ZN(n5032) );
  INV_X1 U6417 ( .A(n5034), .ZN(n5035) );
  NAND2_X1 U6418 ( .A1(n9300), .A2(n5175), .ZN(n5037) );
  XNOR2_X1 U6419 ( .A(n5039), .B(n5188), .ZN(n5046) );
  INV_X1 U6420 ( .A(n5046), .ZN(n5044) );
  INV_X1 U6421 ( .A(n9300), .ZN(n5041) );
  OR2_X1 U6422 ( .A1(n5835), .A2(n5212), .ZN(n5042) );
  AND2_X1 U6423 ( .A1(n4419), .A2(n5042), .ZN(n5045) );
  INV_X1 U6424 ( .A(n5045), .ZN(n5043) );
  NAND2_X1 U6425 ( .A1(n5044), .A2(n5043), .ZN(n5047) );
  NAND2_X1 U6426 ( .A1(n5046), .A2(n5045), .ZN(n6693) );
  NAND2_X1 U6427 ( .A1(n5047), .A2(n6693), .ZN(n6646) );
  INV_X1 U6428 ( .A(n6646), .ZN(n5068) );
  INV_X1 U6429 ( .A(SI_0_), .ZN(n5049) );
  INV_X1 U6430 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5048) );
  AND2_X1 U6431 ( .A1(n5051), .A2(n5050), .ZN(n9783) );
  MUX2_X1 U6432 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9783), .S(n6611), .Z(n6709) );
  INV_X1 U6433 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6434 ( .A1(n5907), .A2(n6644), .ZN(n5053) );
  OAI21_X1 U6435 ( .B1(n5094), .B2(n5054), .A(n5053), .ZN(n5057) );
  INV_X1 U6436 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7253) );
  INV_X1 U6437 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5058) );
  OR2_X1 U6438 ( .A1(n5095), .A2(n5058), .ZN(n5055) );
  OAI21_X1 U6439 ( .B1(n5069), .B2(n7253), .A(n5055), .ZN(n5056) );
  NAND2_X1 U6440 ( .A1(n9302), .A2(n4351), .ZN(n5059) );
  NAND2_X1 U6441 ( .A1(n9302), .A2(n5754), .ZN(n5063) );
  INV_X1 U6442 ( .A(n5036), .ZN(n5823) );
  AOI22_X1 U6443 ( .A1(n6709), .A2(n4351), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5823), .ZN(n5062) );
  NAND2_X1 U6444 ( .A1(n5063), .A2(n5062), .ZN(n6658) );
  NAND2_X1 U6445 ( .A1(n5064), .A2(n5188), .ZN(n5065) );
  NAND2_X1 U6446 ( .A1(n5066), .A2(n5065), .ZN(n6648) );
  INV_X1 U6447 ( .A(n6648), .ZN(n5067) );
  NAND2_X1 U6448 ( .A1(n6692), .A2(n6693), .ZN(n5092) );
  INV_X1 U6449 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9317) );
  OR2_X1 U6450 ( .A1(n5069), .A2(n9317), .ZN(n5076) );
  INV_X1 U6451 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5070) );
  OR2_X1 U6452 ( .A1(n5094), .A2(n5070), .ZN(n5075) );
  INV_X1 U6453 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5071) );
  OR2_X1 U6454 ( .A1(n5095), .A2(n5071), .ZN(n5074) );
  INV_X1 U6455 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5072) );
  OR2_X1 U6456 ( .A1(n5907), .A2(n5072), .ZN(n5073) );
  NAND2_X1 U6457 ( .A1(n5078), .A2(n5077), .ZN(n5081) );
  NAND2_X1 U6458 ( .A1(n5079), .A2(SI_1_), .ZN(n5080) );
  NAND2_X1 U6459 ( .A1(n5081), .A2(n5080), .ZN(n5106) );
  MUX2_X1 U6460 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4350), .Z(n5107) );
  INV_X1 U6461 ( .A(SI_2_), .ZN(n5082) );
  XNOR2_X1 U6462 ( .A(n5106), .B(n5105), .ZN(n6581) );
  OR2_X1 U6463 ( .A1(n5110), .A2(n6581), .ZN(n5085) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6582) );
  OR2_X1 U6465 ( .A1(n8173), .A2(n6582), .ZN(n5084) );
  OR2_X1 U6466 ( .A1(n5083), .A2(n5236), .ZN(n5121) );
  INV_X1 U6467 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5101) );
  XNOR2_X1 U6468 ( .A(n5121), .B(n5101), .ZN(n9316) );
  XNOR2_X1 U6469 ( .A(n5087), .B(n5188), .ZN(n5090) );
  OAI22_X1 U6470 ( .A1(n6750), .A2(n5040), .B1(n6735), .B2(n5212), .ZN(n5089)
         );
  INV_X1 U6471 ( .A(n5089), .ZN(n5088) );
  NAND2_X1 U6472 ( .A1(n5090), .A2(n5088), .ZN(n5093) );
  AND2_X1 U6473 ( .A1(n5093), .A2(n5091), .ZN(n6691) );
  NAND2_X1 U6474 ( .A1(n5092), .A2(n6691), .ZN(n6695) );
  NAND2_X1 U6475 ( .A1(n6695), .A2(n5093), .ZN(n6728) );
  OR2_X1 U6476 ( .A1(n5069), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5100) );
  INV_X1 U6477 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6835) );
  INV_X1 U6478 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5096) );
  INV_X1 U6479 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5098) );
  OR2_X1 U6480 ( .A1(n5907), .A2(n5098), .ZN(n5099) );
  NAND2_X1 U6481 ( .A1(n5121), .A2(n5101), .ZN(n5102) );
  NAND2_X1 U6482 ( .A1(n5102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5104) );
  INV_X1 U6483 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5103) );
  XNOR2_X1 U6484 ( .A(n5104), .B(n5103), .ZN(n6672) );
  NAND2_X1 U6485 ( .A1(n5106), .A2(n5105), .ZN(n5128) );
  NAND2_X1 U6486 ( .A1(n5107), .A2(SI_2_), .ZN(n5123) );
  NAND2_X1 U6487 ( .A1(n5128), .A2(n5123), .ZN(n5109) );
  INV_X1 U6488 ( .A(SI_3_), .ZN(n5108) );
  XNOR2_X1 U6489 ( .A(n5109), .B(n5126), .ZN(n6578) );
  OR2_X1 U6490 ( .A1(n5110), .A2(n6578), .ZN(n5112) );
  INV_X1 U6491 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6579) );
  OR2_X1 U6492 ( .A1(n8173), .A2(n6579), .ZN(n5111) );
  OAI211_X1 U6493 ( .C1(n6611), .C2(n6672), .A(n5112), .B(n5111), .ZN(n6754)
         );
  XNOR2_X1 U6494 ( .A(n5113), .B(n5188), .ZN(n5136) );
  OAI22_X1 U6495 ( .A1(n6910), .A2(n5040), .B1(n6837), .B2(n5061), .ZN(n5134)
         );
  XNOR2_X1 U6496 ( .A(n5136), .B(n5134), .ZN(n6729) );
  OAI21_X1 U6497 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n5144), .ZN(n6915) );
  OR2_X1 U6498 ( .A1(n5069), .A2(n6915), .ZN(n5118) );
  INV_X1 U6499 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6916) );
  INV_X1 U6500 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5114) );
  OR2_X1 U6501 ( .A1(n5095), .A2(n5114), .ZN(n5117) );
  INV_X1 U6502 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5115) );
  OR2_X1 U6503 ( .A1(n5907), .A2(n5115), .ZN(n5116) );
  OR2_X1 U6504 ( .A1(n5119), .A2(n5236), .ZN(n5120) );
  NAND2_X1 U6505 ( .A1(n5121), .A2(n5120), .ZN(n5157) );
  XNOR2_X1 U6506 ( .A(n5157), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6679) );
  INV_X1 U6507 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6584) );
  OR2_X1 U6508 ( .A1(n8173), .A2(n6584), .ZN(n5132) );
  NAND2_X1 U6509 ( .A1(n5122), .A2(SI_3_), .ZN(n5124) );
  AND2_X1 U6510 ( .A1(n5123), .A2(n5124), .ZN(n5127) );
  INV_X1 U6511 ( .A(n5124), .ZN(n5125) );
  MUX2_X1 U6512 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5716), .Z(n5152) );
  INV_X1 U6513 ( .A(SI_4_), .ZN(n5129) );
  XNOR2_X1 U6514 ( .A(n5130), .B(n5151), .ZN(n6583) );
  OR2_X1 U6515 ( .A1(n5110), .A2(n6583), .ZN(n5131) );
  OAI211_X1 U6516 ( .C1(n6679), .C2(n6611), .A(n5132), .B(n5131), .ZN(n6918)
         );
  INV_X1 U6517 ( .A(n6918), .ZN(n9959) );
  OAI22_X1 U6518 ( .A1(n6785), .A2(n5061), .B1(n9959), .B2(n5086), .ZN(n5133)
         );
  XNOR2_X1 U6519 ( .A(n5133), .B(n5188), .ZN(n5138) );
  OAI22_X1 U6520 ( .A1(n6785), .A2(n5040), .B1(n9959), .B2(n5212), .ZN(n5139)
         );
  XNOR2_X1 U6521 ( .A(n5138), .B(n5139), .ZN(n6721) );
  INV_X1 U6522 ( .A(n5134), .ZN(n5135) );
  NAND2_X1 U6523 ( .A1(n5136), .A2(n5135), .ZN(n6719) );
  AND2_X1 U6524 ( .A1(n6721), .A2(n6719), .ZN(n5137) );
  INV_X1 U6525 ( .A(n5138), .ZN(n5140) );
  NAND2_X1 U6526 ( .A1(n5140), .A2(n5139), .ZN(n5141) );
  INV_X1 U6527 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9363) );
  OR2_X1 U6528 ( .A1(n8035), .A2(n9363), .ZN(n5150) );
  INV_X1 U6529 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6530 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  NAND2_X1 U6531 ( .A1(n5168), .A2(n5145), .ZN(n6982) );
  OR2_X1 U6532 ( .A1(n5069), .A2(n6982), .ZN(n5149) );
  INV_X1 U6533 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9369) );
  OR2_X1 U6534 ( .A1(n5095), .A2(n9369), .ZN(n5148) );
  INV_X1 U6535 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5146) );
  OR2_X1 U6536 ( .A1(n5907), .A2(n5146), .ZN(n5147) );
  NAND2_X1 U6537 ( .A1(n5152), .A2(SI_4_), .ZN(n5153) );
  MUX2_X1 U6538 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5716), .Z(n5183) );
  INV_X1 U6539 ( .A(SI_5_), .ZN(n5155) );
  XNOR2_X1 U6540 ( .A(n5182), .B(n5181), .ZN(n6589) );
  OR2_X1 U6541 ( .A1(n5110), .A2(n6589), .ZN(n5162) );
  INV_X1 U6542 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5156) );
  OR2_X1 U6543 ( .A1(n8173), .A2(n5156), .ZN(n5160) );
  OAI21_X1 U6544 ( .B1(n5157), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5159) );
  INV_X1 U6545 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5158) );
  XNOR2_X1 U6546 ( .A(n5159), .B(n5158), .ZN(n9370) );
  OAI22_X1 U6547 ( .A1(n6932), .A2(n5212), .B1(n6981), .B2(n5086), .ZN(n5163)
         );
  XNOR2_X1 U6548 ( .A(n5163), .B(n5038), .ZN(n5165) );
  OAI22_X1 U6549 ( .A1(n6932), .A2(n5040), .B1(n6981), .B2(n5212), .ZN(n5164)
         );
  INV_X1 U6550 ( .A(n5164), .ZN(n6569) );
  INV_X1 U6551 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6552 ( .A1(n5168), .A2(n5167), .ZN(n5169) );
  NAND2_X1 U6553 ( .A1(n5198), .A2(n5169), .ZN(n6940) );
  OR2_X1 U6554 ( .A1(n5069), .A2(n6940), .ZN(n5174) );
  INV_X1 U6555 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6941) );
  OR2_X1 U6556 ( .A1(n8035), .A2(n6941), .ZN(n5173) );
  OR2_X1 U6557 ( .A1(n5095), .A2(n9983), .ZN(n5172) );
  INV_X1 U6558 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5170) );
  OR2_X1 U6559 ( .A1(n5907), .A2(n5170), .ZN(n5171) );
  INV_X1 U6560 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6561 ( .A1(n5177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5178) );
  MUX2_X1 U6562 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5178), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5180) );
  NAND2_X1 U6563 ( .A1(n5180), .A2(n5179), .ZN(n9368) );
  NAND2_X1 U6564 ( .A1(n5183), .A2(SI_5_), .ZN(n5184) );
  MUX2_X1 U6565 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5716), .Z(n5205) );
  INV_X1 U6566 ( .A(SI_6_), .ZN(n5186) );
  INV_X1 U6567 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6588) );
  OR2_X1 U6568 ( .A1(n8173), .A2(n6588), .ZN(n5187) );
  OAI22_X1 U6569 ( .A1(n6882), .A2(n5061), .B1(n9964), .B2(n5086), .ZN(n5189)
         );
  XNOR2_X1 U6570 ( .A(n5189), .B(n5188), .ZN(n5191) );
  OAI22_X1 U6571 ( .A1(n6882), .A2(n5040), .B1(n9964), .B2(n5061), .ZN(n5192)
         );
  INV_X1 U6572 ( .A(n5192), .ZN(n5190) );
  NAND2_X1 U6573 ( .A1(n5191), .A2(n5190), .ZN(n5195) );
  INV_X1 U6574 ( .A(n5191), .ZN(n5193) );
  NAND2_X1 U6575 ( .A1(n5193), .A2(n5192), .ZN(n5194) );
  AND2_X1 U6576 ( .A1(n5195), .A2(n5194), .ZN(n6768) );
  INV_X1 U6577 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9404) );
  OR2_X1 U6578 ( .A1(n8035), .A2(n9404), .ZN(n5204) );
  INV_X1 U6579 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6580 ( .A1(n5198), .A2(n5197), .ZN(n5199) );
  NAND2_X1 U6581 ( .A1(n5256), .A2(n5199), .ZN(n6885) );
  OR2_X1 U6582 ( .A1(n5069), .A2(n6885), .ZN(n5203) );
  INV_X1 U6583 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9398) );
  OR2_X1 U6584 ( .A1(n5095), .A2(n9398), .ZN(n5202) );
  INV_X1 U6585 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5200) );
  OR2_X1 U6586 ( .A1(n5907), .A2(n5200), .ZN(n5201) );
  NAND2_X1 U6587 ( .A1(n5205), .A2(SI_6_), .ZN(n5228) );
  INV_X1 U6588 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6590) );
  MUX2_X1 U6589 ( .A(n5210), .B(n6590), .S(n5206), .Z(n5217) );
  XNOR2_X1 U6590 ( .A(n5265), .B(n5264), .ZN(n6591) );
  OR2_X1 U6591 ( .A1(n6591), .A2(n5110), .ZN(n5209) );
  NAND2_X1 U6592 ( .A1(n5179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5207) );
  XNOR2_X1 U6593 ( .A(n5207), .B(n4871), .ZN(n9405) );
  OR2_X1 U6594 ( .A1(n6611), .A2(n9405), .ZN(n5208) );
  OAI211_X1 U6595 ( .C1(n8173), .C2(n5210), .A(n5209), .B(n5208), .ZN(n6902)
         );
  OAI22_X1 U6596 ( .A1(n6931), .A2(n5212), .B1(n6904), .B2(n5086), .ZN(n5211)
         );
  XNOR2_X1 U6597 ( .A(n5211), .B(n5188), .ZN(n5214) );
  OAI22_X1 U6598 ( .A1(n6931), .A2(n5040), .B1(n6904), .B2(n5212), .ZN(n5215)
         );
  INV_X1 U6599 ( .A(n5215), .ZN(n5213) );
  AND2_X1 U6600 ( .A1(n5214), .A2(n5213), .ZN(n6796) );
  INV_X1 U6601 ( .A(n5214), .ZN(n5216) );
  NAND2_X1 U6602 ( .A1(n5216), .A2(n5215), .ZN(n6794) );
  INV_X1 U6603 ( .A(n5217), .ZN(n5218) );
  INV_X1 U6604 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5219) );
  INV_X1 U6605 ( .A(n5221), .ZN(n5222) );
  NAND2_X1 U6606 ( .A1(n5222), .A2(SI_8_), .ZN(n5223) );
  NAND2_X1 U6607 ( .A1(n5266), .A2(n4956), .ZN(n5226) );
  INV_X1 U6608 ( .A(n5225), .ZN(n5230) );
  INV_X1 U6609 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6599) );
  INV_X1 U6610 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6593) );
  MUX2_X1 U6611 ( .A(n6599), .B(n6593), .S(n4349), .Z(n5231) );
  INV_X1 U6612 ( .A(SI_9_), .ZN(n7046) );
  NAND2_X1 U6613 ( .A1(n5231), .A2(n7046), .ZN(n5284) );
  INV_X1 U6614 ( .A(n5231), .ZN(n5232) );
  AND2_X1 U6615 ( .A1(n5284), .A2(n5288), .ZN(n5233) );
  XNOR2_X1 U6616 ( .A(n5234), .B(n5233), .ZN(n6592) );
  INV_X2 U6617 ( .A(n5110), .ZN(n8172) );
  NAND2_X1 U6618 ( .A1(n6592), .A2(n8172), .ZN(n5240) );
  OR2_X1 U6619 ( .A1(n5235), .A2(n5236), .ZN(n5269) );
  INV_X1 U6620 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6621 ( .A1(n5269), .A2(n5237), .ZN(n5271) );
  NAND2_X1 U6622 ( .A1(n5271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5238) );
  XNOR2_X1 U6623 ( .A(n5238), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9435) );
  AOI22_X1 U6624 ( .A1(n5557), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5556), .B2(
        n9435), .ZN(n5239) );
  NAND2_X1 U6625 ( .A1(n9968), .A2(n5774), .ZN(n5251) );
  INV_X1 U6626 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6969) );
  OR2_X1 U6627 ( .A1(n8035), .A2(n6969), .ZN(n5249) );
  INV_X1 U6628 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5255) );
  INV_X1 U6629 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6630 ( .A1(n5258), .A2(n5242), .ZN(n5243) );
  NAND2_X1 U6631 ( .A1(n5324), .A2(n5243), .ZN(n7577) );
  OR2_X1 U6632 ( .A1(n5069), .A2(n7577), .ZN(n5248) );
  INV_X1 U6633 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5244) );
  OR2_X1 U6634 ( .A1(n5095), .A2(n5244), .ZN(n5247) );
  INV_X1 U6635 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5245) );
  OR2_X1 U6636 ( .A1(n5907), .A2(n5245), .ZN(n5246) );
  INV_X1 U6637 ( .A(n7263), .ZN(n9293) );
  NAND2_X1 U6638 ( .A1(n9293), .A2(n4351), .ZN(n5250) );
  NAND2_X1 U6639 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  XNOR2_X1 U6640 ( .A(n5252), .B(n5188), .ZN(n7582) );
  NAND2_X1 U6641 ( .A1(n9968), .A2(n4351), .ZN(n5254) );
  NAND2_X1 U6642 ( .A1(n9293), .A2(n5754), .ZN(n5253) );
  AND2_X1 U6643 ( .A1(n5254), .A2(n5253), .ZN(n7581) );
  INV_X1 U6644 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9403) );
  OR2_X1 U6645 ( .A1(n8035), .A2(n9403), .ZN(n5263) );
  NAND2_X1 U6646 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  NAND2_X1 U6647 ( .A1(n5258), .A2(n5257), .ZN(n7264) );
  OR2_X1 U6648 ( .A1(n5069), .A2(n7264), .ZN(n5262) );
  INV_X1 U6649 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9397) );
  OR2_X1 U6650 ( .A1(n5095), .A2(n9397), .ZN(n5261) );
  INV_X1 U6651 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5259) );
  OR2_X1 U6652 ( .A1(n5907), .A2(n5259), .ZN(n5260) );
  NAND2_X1 U6653 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  XNOR2_X1 U6654 ( .A(n5268), .B(n4956), .ZN(n6605) );
  INV_X1 U6655 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6656 ( .A1(n5270), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5272) );
  AOI22_X1 U6657 ( .A1(n5557), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5556), .B2(
        n9430), .ZN(n5273) );
  NAND2_X1 U6658 ( .A1(n6853), .A2(n5774), .ZN(n5274) );
  OAI21_X1 U6659 ( .B1(n6881), .B2(n5212), .A(n5274), .ZN(n5275) );
  XNOR2_X1 U6660 ( .A(n5275), .B(n5188), .ZN(n7259) );
  INV_X1 U6661 ( .A(n6881), .ZN(n9294) );
  NAND2_X1 U6662 ( .A1(n9294), .A2(n5754), .ZN(n5277) );
  NAND2_X1 U6663 ( .A1(n6853), .A2(n4351), .ZN(n5276) );
  AND2_X1 U6664 ( .A1(n5277), .A2(n5276), .ZN(n7261) );
  OAI22_X1 U6665 ( .A1(n7582), .A2(n7581), .B1(n7259), .B2(n7261), .ZN(n5283)
         );
  INV_X1 U6666 ( .A(n7259), .ZN(n7580) );
  INV_X1 U6667 ( .A(n7261), .ZN(n5278) );
  INV_X1 U6668 ( .A(n7581), .ZN(n5279) );
  OAI21_X1 U6669 ( .B1(n7580), .B2(n5278), .A(n5279), .ZN(n5281) );
  NOR2_X1 U6670 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  AOI22_X1 U6671 ( .A1(n5281), .A2(n7582), .B1(n7259), .B2(n5280), .ZN(n5282)
         );
  INV_X1 U6672 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6600) );
  INV_X1 U6673 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5287) );
  MUX2_X1 U6674 ( .A(n6600), .B(n5287), .S(n4350), .Z(n5290) );
  INV_X1 U6675 ( .A(n5290), .ZN(n5291) );
  MUX2_X1 U6676 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5716), .Z(n5349) );
  XNOR2_X1 U6677 ( .A(n5349), .B(SI_11_), .ZN(n5292) );
  XNOR2_X1 U6678 ( .A(n5348), .B(n5292), .ZN(n6597) );
  NAND2_X1 U6679 ( .A1(n6597), .A2(n8172), .ZN(n5296) );
  NAND2_X1 U6680 ( .A1(n5293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5294) );
  XNOR2_X1 U6681 ( .A(n5294), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U6682 ( .A1(n5557), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5556), .B2(
        n9836), .ZN(n5295) );
  NAND2_X1 U6683 ( .A1(n5296), .A2(n5295), .ZN(n7610) );
  NAND2_X1 U6684 ( .A1(n7610), .A2(n5774), .ZN(n5307) );
  INV_X1 U6685 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7221) );
  OR2_X1 U6686 ( .A1(n8035), .A2(n7221), .ZN(n5305) );
  INV_X1 U6687 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5323) );
  INV_X1 U6688 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6689 ( .A1(n5326), .A2(n5298), .ZN(n5299) );
  NAND2_X1 U6690 ( .A1(n5369), .A2(n5299), .ZN(n7608) );
  OR2_X1 U6691 ( .A1(n5069), .A2(n7608), .ZN(n5304) );
  INV_X1 U6692 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5300) );
  OR2_X1 U6693 ( .A1(n5095), .A2(n5300), .ZN(n5303) );
  INV_X1 U6694 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5301) );
  OR2_X1 U6695 ( .A1(n5907), .A2(n5301), .ZN(n5302) );
  INV_X1 U6696 ( .A(n6952), .ZN(n9291) );
  NAND2_X1 U6697 ( .A1(n9291), .A2(n4351), .ZN(n5306) );
  NAND2_X1 U6698 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  XNOR2_X1 U6699 ( .A(n5308), .B(n5038), .ZN(n7602) );
  NAND2_X1 U6700 ( .A1(n7610), .A2(n4351), .ZN(n5310) );
  NAND2_X1 U6701 ( .A1(n9291), .A2(n5754), .ZN(n5309) );
  NAND2_X1 U6702 ( .A1(n5310), .A2(n5309), .ZN(n5342) );
  AND2_X1 U6703 ( .A1(n5312), .A2(n5311), .ZN(n5314) );
  NOR2_X1 U6704 ( .A1(n5314), .A2(n5313), .ZN(n5316) );
  XNOR2_X1 U6705 ( .A(n5316), .B(n5315), .ZN(n6594) );
  NAND2_X1 U6706 ( .A1(n6594), .A2(n8172), .ZN(n5322) );
  NAND2_X1 U6707 ( .A1(n5235), .A2(n5317), .ZN(n5318) );
  NAND2_X1 U6708 ( .A1(n5318), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5319) );
  MUX2_X1 U6709 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5319), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5320) );
  AND2_X1 U6710 ( .A1(n5320), .A2(n5293), .ZN(n9814) );
  AOI22_X1 U6711 ( .A1(n5557), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5556), .B2(
        n9814), .ZN(n5321) );
  NAND2_X1 U6712 ( .A1(n5322), .A2(n5321), .ZN(n7679) );
  NAND2_X1 U6713 ( .A1(n7679), .A2(n4351), .ZN(n5334) );
  NAND2_X1 U6714 ( .A1(n5324), .A2(n5323), .ZN(n5325) );
  NAND2_X1 U6715 ( .A1(n5326), .A2(n5325), .ZN(n7672) );
  OR2_X1 U6716 ( .A1(n5069), .A2(n7672), .ZN(n5332) );
  INV_X1 U6717 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6958) );
  OR2_X1 U6718 ( .A1(n8035), .A2(n6958), .ZN(n5331) );
  INV_X1 U6719 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5327) );
  OR2_X1 U6720 ( .A1(n5095), .A2(n5327), .ZN(n5330) );
  INV_X1 U6721 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6722 ( .A1(n5907), .A2(n5328), .ZN(n5329) );
  INV_X1 U6723 ( .A(n7605), .ZN(n9292) );
  NAND2_X1 U6724 ( .A1(n9292), .A2(n5754), .ZN(n5333) );
  NAND2_X1 U6725 ( .A1(n5334), .A2(n5333), .ZN(n7674) );
  NAND2_X1 U6726 ( .A1(n7679), .A2(n5774), .ZN(n5336) );
  NAND2_X1 U6727 ( .A1(n9292), .A2(n4351), .ZN(n5335) );
  NAND2_X1 U6728 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  XNOR2_X1 U6729 ( .A(n5337), .B(n5038), .ZN(n5339) );
  AOI22_X1 U6730 ( .A1(n7602), .A2(n5342), .B1(n7674), .B2(n5339), .ZN(n5338)
         );
  NAND2_X1 U6731 ( .A1(n7599), .A2(n5338), .ZN(n5347) );
  INV_X1 U6732 ( .A(n7602), .ZN(n5345) );
  INV_X1 U6733 ( .A(n5339), .ZN(n7600) );
  INV_X1 U6734 ( .A(n7674), .ZN(n5340) );
  NAND2_X1 U6735 ( .A1(n7600), .A2(n5340), .ZN(n5341) );
  NAND2_X1 U6736 ( .A1(n5341), .A2(n5342), .ZN(n5344) );
  INV_X1 U6737 ( .A(n5341), .ZN(n5343) );
  INV_X1 U6738 ( .A(n5342), .ZN(n7601) );
  AOI22_X1 U6739 ( .A1(n5345), .A2(n5344), .B1(n5343), .B2(n7601), .ZN(n5346)
         );
  NAND2_X1 U6740 ( .A1(n5347), .A2(n5346), .ZN(n7374) );
  INV_X1 U6741 ( .A(SI_11_), .ZN(n5350) );
  MUX2_X1 U6742 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5716), .Z(n5353) );
  INV_X1 U6743 ( .A(n5353), .ZN(n5354) );
  INV_X1 U6744 ( .A(SI_12_), .ZN(n7135) );
  NAND2_X1 U6745 ( .A1(n5354), .A2(n7135), .ZN(n5355) );
  INV_X1 U6746 ( .A(n5357), .ZN(n5359) );
  NAND2_X1 U6747 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  AND2_X1 U6748 ( .A1(n5439), .A2(n5360), .ZN(n6619) );
  NAND2_X1 U6749 ( .A1(n6619), .A2(n8172), .ZN(n5367) );
  INV_X1 U6750 ( .A(n5293), .ZN(n5362) );
  INV_X1 U6751 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6752 ( .A1(n5362), .A2(n5361), .ZN(n5411) );
  NAND2_X1 U6753 ( .A1(n5411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5364) );
  INV_X1 U6754 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5363) );
  OR2_X1 U6755 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  NAND2_X1 U6756 ( .A1(n5364), .A2(n5363), .ZN(n5385) );
  AND2_X1 U6757 ( .A1(n5365), .A2(n5385), .ZN(n9852) );
  AOI22_X1 U6758 ( .A1(n5557), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5556), .B2(
        n9852), .ZN(n5366) );
  NAND2_X1 U6759 ( .A1(n7380), .A2(n5774), .ZN(n5377) );
  INV_X1 U6760 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7287) );
  OR2_X1 U6761 ( .A1(n8035), .A2(n7287), .ZN(n5375) );
  INV_X1 U6762 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6763 ( .A1(n5369), .A2(n5368), .ZN(n5370) );
  NAND2_X1 U6764 ( .A1(n5390), .A2(n5370), .ZN(n7378) );
  OR2_X1 U6765 ( .A1(n5069), .A2(n7378), .ZN(n5374) );
  INV_X1 U6766 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9419) );
  OR2_X1 U6767 ( .A1(n5095), .A2(n9419), .ZN(n5373) );
  INV_X1 U6768 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5371) );
  OR2_X1 U6769 ( .A1(n5907), .A2(n5371), .ZN(n5372) );
  INV_X1 U6770 ( .A(n7546), .ZN(n9290) );
  NAND2_X1 U6771 ( .A1(n9290), .A2(n4351), .ZN(n5376) );
  NAND2_X1 U6772 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  XNOR2_X1 U6773 ( .A(n5378), .B(n5038), .ZN(n5380) );
  NOR2_X1 U6774 ( .A1(n7546), .A2(n5040), .ZN(n5379) );
  AOI21_X1 U6775 ( .B1(n7380), .B2(n4351), .A(n5379), .ZN(n5381) );
  XNOR2_X1 U6776 ( .A(n5380), .B(n5381), .ZN(n7375) );
  INV_X1 U6777 ( .A(n5380), .ZN(n5382) );
  NAND2_X1 U6778 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  MUX2_X1 U6779 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4350), .Z(n5403) );
  XNOR2_X1 U6780 ( .A(n5403), .B(SI_13_), .ZN(n5384) );
  XNOR2_X1 U6781 ( .A(n5404), .B(n5384), .ZN(n6627) );
  NAND2_X1 U6782 ( .A1(n6627), .A2(n8172), .ZN(n5388) );
  NAND2_X1 U6783 ( .A1(n5385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5386) );
  XNOR2_X1 U6784 ( .A(n5386), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9437) );
  AOI22_X1 U6785 ( .A1(n5557), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5556), .B2(
        n9437), .ZN(n5387) );
  NAND2_X1 U6786 ( .A1(n7549), .A2(n5774), .ZN(n5397) );
  INV_X1 U6787 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7387) );
  OR2_X1 U6788 ( .A1(n8035), .A2(n7387), .ZN(n5395) );
  INV_X1 U6789 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6790 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  NAND2_X1 U6791 ( .A1(n5421), .A2(n5391), .ZN(n7544) );
  OR2_X1 U6792 ( .A1(n5069), .A2(n7544), .ZN(n5394) );
  INV_X1 U6793 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7572) );
  OR2_X1 U6794 ( .A1(n5095), .A2(n7572), .ZN(n5393) );
  INV_X1 U6795 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7569) );
  OR2_X1 U6796 ( .A1(n5907), .A2(n7569), .ZN(n5392) );
  INV_X1 U6797 ( .A(n7559), .ZN(n9289) );
  NAND2_X1 U6798 ( .A1(n9289), .A2(n4351), .ZN(n5396) );
  NAND2_X1 U6799 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  XNOR2_X1 U6800 ( .A(n5398), .B(n5038), .ZN(n5400) );
  NOR2_X1 U6801 ( .A1(n7559), .A2(n5040), .ZN(n5399) );
  AOI21_X1 U6802 ( .B1(n7549), .B2(n4351), .A(n5399), .ZN(n5401) );
  XNOR2_X1 U6803 ( .A(n5400), .B(n5401), .ZN(n7543) );
  INV_X1 U6804 ( .A(n5400), .ZN(n5402) );
  NAND2_X1 U6805 ( .A1(n5404), .A2(SI_13_), .ZN(n5405) );
  NAND2_X1 U6806 ( .A1(n5442), .A2(n5405), .ZN(n5407) );
  MUX2_X1 U6807 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4350), .Z(n5435) );
  XNOR2_X1 U6808 ( .A(n5435), .B(SI_14_), .ZN(n5406) );
  XNOR2_X1 U6809 ( .A(n5407), .B(n5406), .ZN(n6631) );
  NAND2_X1 U6810 ( .A1(n6631), .A2(n8172), .ZN(n5415) );
  INV_X1 U6811 ( .A(n5409), .ZN(n5410) );
  OAI21_X1 U6812 ( .B1(n5411), .B2(n5410), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5412) );
  MUX2_X1 U6813 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5412), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5413) );
  AND2_X1 U6814 ( .A1(n5408), .A2(n5413), .ZN(n9883) );
  AOI22_X1 U6815 ( .A1(n5557), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5556), .B2(
        n9883), .ZN(n5414) );
  NAND2_X1 U6816 ( .A1(n9725), .A2(n5774), .ZN(n5428) );
  INV_X1 U6817 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5418) );
  INV_X1 U6818 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5416) );
  OR2_X1 U6819 ( .A1(n5095), .A2(n5416), .ZN(n5417) );
  OAI21_X1 U6820 ( .B1(n8035), .B2(n5418), .A(n5417), .ZN(n5426) );
  INV_X1 U6821 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6822 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  NAND2_X1 U6823 ( .A1(n5478), .A2(n5422), .ZN(n7561) );
  INV_X1 U6824 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5423) );
  OR2_X1 U6825 ( .A1(n5907), .A2(n5423), .ZN(n5424) );
  OAI21_X1 U6826 ( .B1(n5069), .B2(n7561), .A(n5424), .ZN(n5425) );
  NAND2_X1 U6827 ( .A1(n7943), .A2(n4351), .ZN(n5427) );
  NAND2_X1 U6828 ( .A1(n5428), .A2(n5427), .ZN(n5429) );
  XNOR2_X1 U6829 ( .A(n5429), .B(n5038), .ZN(n5432) );
  XNOR2_X1 U6830 ( .A(n5431), .B(n5432), .ZN(n7768) );
  AND2_X1 U6831 ( .A1(n7943), .A2(n5754), .ZN(n5430) );
  AOI21_X1 U6832 ( .B1(n9725), .B2(n4351), .A(n5430), .ZN(n7770) );
  INV_X1 U6833 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U6834 ( .A1(n5431), .A2(n5433), .ZN(n5434) );
  INV_X1 U6835 ( .A(SI_14_), .ZN(n5443) );
  INV_X1 U6836 ( .A(n5440), .ZN(n5436) );
  NAND2_X1 U6837 ( .A1(n5444), .A2(n5443), .ZN(n5466) );
  MUX2_X1 U6838 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4350), .Z(n5469) );
  INV_X1 U6839 ( .A(n5469), .ZN(n5445) );
  INV_X1 U6840 ( .A(SI_15_), .ZN(n5468) );
  NAND2_X1 U6841 ( .A1(n5469), .A2(SI_15_), .ZN(n5448) );
  MUX2_X1 U6842 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4349), .Z(n5495) );
  XNOR2_X1 U6843 ( .A(n5495), .B(SI_16_), .ZN(n5449) );
  XNOR2_X1 U6844 ( .A(n5497), .B(n5449), .ZN(n6653) );
  NAND2_X1 U6845 ( .A1(n6653), .A2(n8172), .ZN(n5452) );
  NAND2_X1 U6846 ( .A1(n4426), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5450) );
  XNOR2_X1 U6847 ( .A(n5450), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9443) );
  AOI22_X1 U6848 ( .A1(n5557), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5556), .B2(
        n9443), .ZN(n5451) );
  NAND2_X1 U6849 ( .A1(n9720), .A2(n5774), .ZN(n5462) );
  INV_X1 U6850 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6851 ( .A1(n5480), .A2(n5454), .ZN(n5455) );
  NAND2_X1 U6852 ( .A1(n5504), .A2(n5455), .ZN(n9216) );
  OR2_X1 U6853 ( .A1(n5069), .A2(n9216), .ZN(n5460) );
  INV_X1 U6854 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7683) );
  OR2_X1 U6855 ( .A1(n8035), .A2(n7683), .ZN(n5459) );
  INV_X1 U6856 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9413) );
  OR2_X1 U6857 ( .A1(n5095), .A2(n9413), .ZN(n5458) );
  INV_X1 U6858 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5456) );
  OR2_X1 U6859 ( .A1(n5907), .A2(n5456), .ZN(n5457) );
  INV_X1 U6860 ( .A(n7941), .ZN(n7831) );
  NAND2_X1 U6861 ( .A1(n7831), .A2(n4351), .ZN(n5461) );
  NAND2_X1 U6862 ( .A1(n5462), .A2(n5461), .ZN(n5463) );
  XNOR2_X1 U6863 ( .A(n5463), .B(n5038), .ZN(n5490) );
  NAND2_X1 U6864 ( .A1(n9720), .A2(n4351), .ZN(n5465) );
  NAND2_X1 U6865 ( .A1(n7831), .A2(n5754), .ZN(n5464) );
  NAND2_X1 U6866 ( .A1(n5465), .A2(n5464), .ZN(n9212) );
  NAND2_X1 U6867 ( .A1(n5467), .A2(n5466), .ZN(n5471) );
  XNOR2_X1 U6868 ( .A(n5469), .B(n5468), .ZN(n5470) );
  XNOR2_X1 U6869 ( .A(n5471), .B(n5470), .ZN(n6635) );
  NAND2_X1 U6870 ( .A1(n6635), .A2(n8172), .ZN(n5475) );
  NAND2_X1 U6871 ( .A1(n5408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5472) );
  MUX2_X1 U6872 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5472), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5473) );
  NAND2_X1 U6873 ( .A1(n5473), .A2(n4426), .ZN(n9440) );
  INV_X1 U6874 ( .A(n9440), .ZN(n9907) );
  AOI22_X1 U6875 ( .A1(n5557), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5556), .B2(
        n9907), .ZN(n5474) );
  NAND2_X1 U6876 ( .A1(n7947), .A2(n4351), .ZN(n5485) );
  INV_X1 U6877 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7646) );
  INV_X1 U6878 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9901) );
  OR2_X1 U6879 ( .A1(n5095), .A2(n9901), .ZN(n5476) );
  OAI21_X1 U6880 ( .B1(n8035), .B2(n7646), .A(n5476), .ZN(n5483) );
  INV_X1 U6881 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6882 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  NAND2_X1 U6883 ( .A1(n5480), .A2(n5479), .ZN(n7945) );
  INV_X1 U6884 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7784) );
  OR2_X1 U6885 ( .A1(n5907), .A2(n7784), .ZN(n5481) );
  OAI21_X1 U6886 ( .B1(n5069), .B2(n7945), .A(n5481), .ZN(n5482) );
  OR2_X1 U6887 ( .A1(n5483), .A2(n5482), .ZN(n9288) );
  NAND2_X1 U6888 ( .A1(n9288), .A2(n5754), .ZN(n5484) );
  NAND2_X1 U6889 ( .A1(n5485), .A2(n5484), .ZN(n7939) );
  NAND2_X1 U6890 ( .A1(n7947), .A2(n5774), .ZN(n5487) );
  NAND2_X1 U6891 ( .A1(n9288), .A2(n4351), .ZN(n5486) );
  NAND2_X1 U6892 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  XNOR2_X1 U6893 ( .A(n5488), .B(n5038), .ZN(n5491) );
  AOI22_X1 U6894 ( .A1(n5490), .A2(n9212), .B1(n7939), .B2(n5491), .ZN(n5489)
         );
  INV_X1 U6895 ( .A(n5490), .ZN(n9213) );
  OAI21_X1 U6896 ( .B1(n5491), .B2(n7939), .A(n9212), .ZN(n5493) );
  NOR2_X1 U6897 ( .A1(n9212), .A2(n7939), .ZN(n5492) );
  INV_X1 U6898 ( .A(n5491), .ZN(n9211) );
  AOI22_X1 U6899 ( .A1(n9213), .A2(n5493), .B1(n5492), .B2(n9211), .ZN(n5494)
         );
  INV_X1 U6900 ( .A(SI_16_), .ZN(n7147) );
  MUX2_X1 U6901 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4349), .Z(n5519) );
  INV_X1 U6902 ( .A(SI_17_), .ZN(n5520) );
  XNOR2_X1 U6903 ( .A(n5519), .B(n5520), .ZN(n5517) );
  XNOR2_X1 U6904 ( .A(n5518), .B(n5517), .ZN(n6715) );
  NAND2_X1 U6905 ( .A1(n6715), .A2(n8172), .ZN(n5500) );
  XNOR2_X1 U6906 ( .A(n5498), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U6907 ( .A1(n5557), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5556), .B2(
        n9926), .ZN(n5499) );
  NAND2_X1 U6908 ( .A1(n7866), .A2(n5774), .ZN(n5510) );
  INV_X1 U6909 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9427) );
  INV_X1 U6910 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9715) );
  OR2_X1 U6911 ( .A1(n5095), .A2(n9715), .ZN(n5501) );
  OAI21_X1 U6912 ( .B1(n8035), .B2(n9427), .A(n5501), .ZN(n5508) );
  INV_X1 U6913 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U6914 ( .A1(n5504), .A2(n5503), .ZN(n5505) );
  NAND2_X1 U6915 ( .A1(n5535), .A2(n5505), .ZN(n7864) );
  INV_X1 U6916 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9768) );
  OR2_X1 U6917 ( .A1(n5907), .A2(n9768), .ZN(n5506) );
  OAI21_X1 U6918 ( .B1(n5069), .B2(n7864), .A(n5506), .ZN(n5507) );
  OR2_X1 U6919 ( .A1(n5508), .A2(n5507), .ZN(n9287) );
  NAND2_X1 U6920 ( .A1(n9287), .A2(n4351), .ZN(n5509) );
  NAND2_X1 U6921 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  XNOR2_X1 U6922 ( .A(n5511), .B(n5188), .ZN(n7859) );
  AND2_X1 U6923 ( .A1(n9287), .A2(n5754), .ZN(n5512) );
  AOI21_X1 U6924 ( .B1(n7866), .B2(n4351), .A(n5512), .ZN(n7858) );
  AND2_X1 U6925 ( .A1(n7859), .A2(n7858), .ZN(n5516) );
  INV_X1 U6926 ( .A(n7859), .ZN(n5514) );
  INV_X1 U6927 ( .A(n7858), .ZN(n5513) );
  NAND2_X1 U6928 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  INV_X1 U6929 ( .A(n5519), .ZN(n5521) );
  NAND2_X1 U6930 ( .A1(n5521), .A2(n5520), .ZN(n5522) );
  NAND2_X1 U6931 ( .A1(n5523), .A2(n5522), .ZN(n5526) );
  MUX2_X1 U6932 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5716), .Z(n5524) );
  NAND2_X1 U6933 ( .A1(n5524), .A2(SI_18_), .ZN(n5553) );
  OAI21_X1 U6934 ( .B1(n5524), .B2(SI_18_), .A(n5553), .ZN(n5525) );
  NAND2_X1 U6935 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  AND2_X1 U6936 ( .A1(n5554), .A2(n5527), .ZN(n6739) );
  NAND2_X1 U6937 ( .A1(n6739), .A2(n8172), .ZN(n5533) );
  OR2_X1 U6938 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  AND2_X1 U6939 ( .A1(n5531), .A2(n5530), .ZN(n9940) );
  AOI22_X1 U6940 ( .A1(n5557), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5556), .B2(
        n9940), .ZN(n5532) );
  NAND2_X1 U6941 ( .A1(n9709), .A2(n5774), .ZN(n5545) );
  INV_X1 U6942 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U6943 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  NAND2_X1 U6944 ( .A1(n5562), .A2(n5536), .ZN(n9259) );
  OR2_X1 U6945 ( .A1(n5069), .A2(n9259), .ZN(n5543) );
  INV_X1 U6946 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5537) );
  OR2_X1 U6947 ( .A1(n8035), .A2(n5537), .ZN(n5542) );
  INV_X1 U6948 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n5538) );
  OR2_X1 U6949 ( .A1(n5095), .A2(n5538), .ZN(n5541) );
  INV_X1 U6950 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5539) );
  OR2_X1 U6951 ( .A1(n5907), .A2(n5539), .ZN(n5540) );
  NAND4_X1 U6952 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(n9642)
         );
  NAND2_X1 U6953 ( .A1(n9642), .A2(n4351), .ZN(n5544) );
  NAND2_X1 U6954 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  XNOR2_X1 U6955 ( .A(n5546), .B(n5038), .ZN(n5547) );
  NAND2_X1 U6956 ( .A1(n9709), .A2(n4351), .ZN(n5550) );
  NAND2_X1 U6957 ( .A1(n9642), .A2(n5754), .ZN(n5549) );
  NAND2_X1 U6958 ( .A1(n5550), .A2(n5549), .ZN(n9258) );
  INV_X1 U6959 ( .A(n9258), .ZN(n5551) );
  MUX2_X1 U6960 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4350), .Z(n5580) );
  XNOR2_X1 U6961 ( .A(n5580), .B(SI_19_), .ZN(n5578) );
  XNOR2_X1 U6962 ( .A(n5577), .B(n5578), .ZN(n6776) );
  NAND2_X1 U6963 ( .A1(n6776), .A2(n8172), .ZN(n5559) );
  AOI22_X1 U6964 ( .A1(n5557), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4485), .B2(
        n5556), .ZN(n5558) );
  NAND2_X1 U6965 ( .A1(n9628), .A2(n5774), .ZN(n5568) );
  INV_X1 U6966 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6967 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  NAND2_X1 U6968 ( .A1(n5605), .A2(n5563), .ZN(n9631) );
  INV_X1 U6969 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9763) );
  OAI22_X1 U6970 ( .A1(n9631), .A2(n5069), .B1(n5907), .B2(n9763), .ZN(n5566)
         );
  INV_X1 U6971 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9632) );
  INV_X1 U6972 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9705) );
  OR2_X1 U6973 ( .A1(n5095), .A2(n9705), .ZN(n5564) );
  OAI21_X1 U6974 ( .B1(n8035), .B2(n9632), .A(n5564), .ZN(n5565) );
  NAND2_X1 U6975 ( .A1(n9610), .A2(n4351), .ZN(n5567) );
  NAND2_X1 U6976 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  XNOR2_X1 U6977 ( .A(n5569), .B(n5038), .ZN(n5572) );
  NAND2_X1 U6978 ( .A1(n9628), .A2(n4351), .ZN(n5571) );
  NAND2_X1 U6979 ( .A1(n9610), .A2(n5754), .ZN(n5570) );
  NAND2_X1 U6980 ( .A1(n5571), .A2(n5570), .ZN(n5573) );
  NAND2_X1 U6981 ( .A1(n5572), .A2(n5573), .ZN(n9189) );
  INV_X1 U6982 ( .A(n5572), .ZN(n5575) );
  INV_X1 U6983 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U6984 ( .A1(n5575), .A2(n5574), .ZN(n9188) );
  INV_X1 U6985 ( .A(n5578), .ZN(n5579) );
  INV_X1 U6986 ( .A(n5580), .ZN(n5581) );
  INV_X1 U6987 ( .A(SI_19_), .ZN(n7090) );
  NAND2_X1 U6988 ( .A1(n5581), .A2(n7090), .ZN(n5582) );
  MUX2_X1 U6989 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4349), .Z(n5597) );
  INV_X1 U6990 ( .A(SI_20_), .ZN(n5596) );
  XNOR2_X1 U6991 ( .A(n5597), .B(n5596), .ZN(n5583) );
  NAND2_X1 U6992 ( .A1(n6827), .A2(n8172), .ZN(n5585) );
  INV_X1 U6993 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6793) );
  OR2_X1 U6994 ( .A1(n8173), .A2(n6793), .ZN(n5584) );
  NAND2_X1 U6995 ( .A1(n9615), .A2(n5774), .ZN(n5592) );
  INV_X1 U6996 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9759) );
  XNOR2_X1 U6997 ( .A(n5605), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U6998 ( .A1(n9618), .A2(n5763), .ZN(n5590) );
  INV_X1 U6999 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5587) );
  INV_X1 U7000 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9700) );
  OR2_X1 U7001 ( .A1(n5095), .A2(n9700), .ZN(n5586) );
  OAI21_X1 U7002 ( .B1(n8035), .B2(n5587), .A(n5586), .ZN(n5588) );
  INV_X1 U7003 ( .A(n5588), .ZN(n5589) );
  OAI211_X1 U7004 ( .C1(n5907), .C2(n9759), .A(n5590), .B(n5589), .ZN(n9645)
         );
  NAND2_X1 U7005 ( .A1(n9645), .A2(n4351), .ZN(n5591) );
  NAND2_X1 U7006 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  XNOR2_X1 U7007 ( .A(n5593), .B(n5188), .ZN(n9235) );
  AND2_X1 U7008 ( .A1(n9645), .A2(n5754), .ZN(n5594) );
  AOI21_X1 U7009 ( .B1(n9615), .B2(n4351), .A(n5594), .ZN(n9234) );
  AND2_X1 U7010 ( .A1(n9235), .A2(n9234), .ZN(n5595) );
  OAI22_X1 U7011 ( .A1(n9233), .A2(n5595), .B1(n9235), .B2(n9234), .ZN(n9196)
         );
  MUX2_X1 U7012 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n5716), .Z(n5616) );
  XNOR2_X1 U7013 ( .A(n5616), .B(SI_21_), .ZN(n5599) );
  XNOR2_X1 U7014 ( .A(n5619), .B(n5599), .ZN(n6923) );
  NAND2_X1 U7015 ( .A1(n6923), .A2(n8172), .ZN(n5601) );
  INV_X1 U7016 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6925) );
  OR2_X1 U7017 ( .A1(n8173), .A2(n6925), .ZN(n5600) );
  NAND2_X1 U7018 ( .A1(n9597), .A2(n5774), .ZN(n5610) );
  INV_X1 U7019 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9755) );
  INV_X1 U7020 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5603) );
  INV_X1 U7021 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5602) );
  OAI21_X1 U7022 ( .B1(n5605), .B2(n5603), .A(n5602), .ZN(n5606) );
  NAND2_X1 U7023 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n5604) );
  NAND2_X1 U7024 ( .A1(n5606), .A2(n5624), .ZN(n9598) );
  OR2_X1 U7025 ( .A1(n9598), .A2(n5069), .ZN(n5608) );
  AOI22_X1 U7026 ( .A1(n5627), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5626), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n5607) );
  OAI211_X1 U7027 ( .C1(n5907), .C2(n9755), .A(n5608), .B(n5607), .ZN(n9611)
         );
  NAND2_X1 U7028 ( .A1(n9611), .A2(n4351), .ZN(n5609) );
  NAND2_X1 U7029 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  XNOR2_X1 U7030 ( .A(n5611), .B(n5188), .ZN(n5614) );
  AND2_X1 U7031 ( .A1(n9611), .A2(n5754), .ZN(n5612) );
  AOI21_X1 U7032 ( .B1(n9597), .B2(n4351), .A(n5612), .ZN(n5613) );
  XNOR2_X1 U7033 ( .A(n5614), .B(n5613), .ZN(n9197) );
  NAND2_X1 U7034 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  INV_X1 U7035 ( .A(n5616), .ZN(n5617) );
  INV_X1 U7036 ( .A(SI_21_), .ZN(n7110) );
  NAND2_X1 U7037 ( .A1(n5617), .A2(n7110), .ZN(n5618) );
  MUX2_X1 U7038 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n4350), .Z(n5639) );
  INV_X1 U7039 ( .A(SI_22_), .ZN(n5640) );
  XNOR2_X1 U7040 ( .A(n5639), .B(n5640), .ZN(n5637) );
  XNOR2_X1 U7041 ( .A(n5638), .B(n5637), .ZN(n7257) );
  NAND2_X1 U7042 ( .A1(n7257), .A2(n8172), .ZN(n5621) );
  INV_X1 U7043 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7270) );
  OR2_X1 U7044 ( .A1(n8173), .A2(n7270), .ZN(n5620) );
  NAND2_X1 U7045 ( .A1(n9688), .A2(n5774), .ZN(n5632) );
  INV_X1 U7046 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5630) );
  INV_X1 U7047 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7048 ( .A1(n5624), .A2(n5623), .ZN(n5625) );
  NAND2_X1 U7049 ( .A1(n5669), .A2(n5625), .ZN(n9249) );
  OR2_X1 U7050 ( .A1(n9249), .A2(n5069), .ZN(n5629) );
  AOI22_X1 U7051 ( .A1(n5627), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n5626), .B2(
        P1_REG1_REG_22__SCAN_IN), .ZN(n5628) );
  OAI211_X1 U7052 ( .C1(n5907), .C2(n5630), .A(n5629), .B(n5628), .ZN(n9593)
         );
  NAND2_X1 U7053 ( .A1(n9593), .A2(n4351), .ZN(n5631) );
  NAND2_X1 U7054 ( .A1(n5632), .A2(n5631), .ZN(n5633) );
  XNOR2_X1 U7055 ( .A(n5633), .B(n5188), .ZN(n5636) );
  NAND2_X1 U7056 ( .A1(n9688), .A2(n5175), .ZN(n5635) );
  NAND2_X1 U7057 ( .A1(n9593), .A2(n5754), .ZN(n5634) );
  NAND2_X1 U7058 ( .A1(n5635), .A2(n5634), .ZN(n9243) );
  NAND2_X1 U7059 ( .A1(n5638), .A2(n5637), .ZN(n5643) );
  INV_X1 U7060 ( .A(n5639), .ZN(n5641) );
  NAND2_X1 U7061 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  NAND2_X1 U7062 ( .A1(n5643), .A2(n5642), .ZN(n5661) );
  MUX2_X1 U7063 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n5716), .Z(n5662) );
  INV_X1 U7064 ( .A(SI_23_), .ZN(n7122) );
  XNOR2_X1 U7065 ( .A(n5662), .B(n7122), .ZN(n5660) );
  XNOR2_X1 U7066 ( .A(n5661), .B(n5660), .ZN(n7321) );
  NAND2_X1 U7067 ( .A1(n7321), .A2(n8172), .ZN(n5645) );
  INV_X1 U7068 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7323) );
  OR2_X1 U7069 ( .A1(n8173), .A2(n7323), .ZN(n5644) );
  NAND2_X1 U7070 ( .A1(n9562), .A2(n5774), .ZN(n5652) );
  XNOR2_X1 U7071 ( .A(n5669), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U7072 ( .A1(n9555), .A2(n5763), .ZN(n5650) );
  INV_X1 U7073 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9564) );
  INV_X1 U7074 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9685) );
  OR2_X1 U7075 ( .A1(n5095), .A2(n9685), .ZN(n5647) );
  INV_X1 U7076 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9750) );
  OR2_X1 U7077 ( .A1(n5907), .A2(n9750), .ZN(n5646) );
  OAI211_X1 U7078 ( .C1(n8035), .C2(n9564), .A(n5647), .B(n5646), .ZN(n5648)
         );
  INV_X1 U7079 ( .A(n5648), .ZN(n5649) );
  NAND2_X1 U7080 ( .A1(n5650), .A2(n5649), .ZN(n9583) );
  NAND2_X1 U7081 ( .A1(n9583), .A2(n5175), .ZN(n5651) );
  NAND2_X1 U7082 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  XNOR2_X1 U7083 ( .A(n5653), .B(n5188), .ZN(n5655) );
  AND2_X1 U7084 ( .A1(n9583), .A2(n5754), .ZN(n5654) );
  AOI21_X1 U7085 ( .B1(n9562), .B2(n4351), .A(n5654), .ZN(n5656) );
  NAND2_X1 U7086 ( .A1(n5655), .A2(n5656), .ZN(n9224) );
  INV_X1 U7087 ( .A(n5655), .ZN(n5658) );
  INV_X1 U7088 ( .A(n5656), .ZN(n5657) );
  NAND2_X1 U7089 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  NAND2_X1 U7090 ( .A1(n5661), .A2(n5660), .ZN(n5665) );
  INV_X1 U7091 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U7092 ( .A1(n5663), .A2(n7122), .ZN(n5664) );
  MUX2_X1 U7093 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4349), .Z(n5690) );
  INV_X1 U7094 ( .A(SI_24_), .ZN(n7112) );
  XNOR2_X1 U7095 ( .A(n5690), .B(n7112), .ZN(n5688) );
  NAND2_X1 U7096 ( .A1(n7553), .A2(n8172), .ZN(n5667) );
  INV_X1 U7097 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7555) );
  OR2_X1 U7098 ( .A1(n8173), .A2(n7555), .ZN(n5666) );
  NAND2_X1 U7099 ( .A1(n9676), .A2(n5774), .ZN(n5679) );
  INV_X1 U7100 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5668) );
  INV_X1 U7101 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9228) );
  OAI21_X1 U7102 ( .B1(n5669), .B2(n5668), .A(n9228), .ZN(n5670) );
  NAND2_X1 U7103 ( .A1(n5670), .A2(n5696), .ZN(n9540) );
  OR2_X1 U7104 ( .A1(n9540), .A2(n5069), .ZN(n5677) );
  INV_X1 U7105 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9539) );
  INV_X1 U7106 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5671) );
  OR2_X1 U7107 ( .A1(n5907), .A2(n5671), .ZN(n5674) );
  INV_X1 U7108 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5672) );
  OR2_X1 U7109 ( .A1(n5095), .A2(n5672), .ZN(n5673) );
  OAI211_X1 U7110 ( .C1(n8035), .C2(n9539), .A(n5674), .B(n5673), .ZN(n5675)
         );
  INV_X1 U7111 ( .A(n5675), .ZN(n5676) );
  NAND2_X1 U7112 ( .A1(n5677), .A2(n5676), .ZN(n9560) );
  NAND2_X1 U7113 ( .A1(n9560), .A2(n4351), .ZN(n5678) );
  NAND2_X1 U7114 ( .A1(n5679), .A2(n5678), .ZN(n5680) );
  XNOR2_X1 U7115 ( .A(n5680), .B(n5188), .ZN(n5682) );
  AND2_X1 U7116 ( .A1(n9560), .A2(n5754), .ZN(n5681) );
  AOI21_X1 U7117 ( .B1(n9676), .B2(n4351), .A(n5681), .ZN(n5683) );
  NAND2_X1 U7118 ( .A1(n5682), .A2(n5683), .ZN(n5687) );
  INV_X1 U7119 ( .A(n5682), .ZN(n5685) );
  INV_X1 U7120 ( .A(n5683), .ZN(n5684) );
  NAND2_X1 U7121 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  NAND2_X1 U7122 ( .A1(n5687), .A2(n5686), .ZN(n9223) );
  INV_X1 U7123 ( .A(n5690), .ZN(n5691) );
  NAND2_X1 U7124 ( .A1(n5691), .A2(n7112), .ZN(n5692) );
  MUX2_X1 U7125 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n4350), .Z(n5711) );
  INV_X1 U7126 ( .A(SI_25_), .ZN(n5712) );
  XNOR2_X1 U7127 ( .A(n5711), .B(n5712), .ZN(n5709) );
  XNOR2_X1 U7128 ( .A(n5710), .B(n5709), .ZN(n7666) );
  NAND2_X1 U7129 ( .A1(n7666), .A2(n8172), .ZN(n5694) );
  INV_X1 U7130 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7668) );
  OR2_X1 U7131 ( .A1(n8173), .A2(n7668), .ZN(n5693) );
  NAND2_X1 U7132 ( .A1(n9529), .A2(n5774), .ZN(n5705) );
  INV_X1 U7133 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U7134 ( .A1(n5696), .A2(n5695), .ZN(n5697) );
  AND2_X1 U7135 ( .A1(n5721), .A2(n5697), .ZN(n9530) );
  NAND2_X1 U7136 ( .A1(n9530), .A2(n5763), .ZN(n5703) );
  INV_X1 U7137 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5700) );
  INV_X1 U7138 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9672) );
  OR2_X1 U7139 ( .A1(n5095), .A2(n9672), .ZN(n5699) );
  INV_X1 U7140 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9745) );
  OR2_X1 U7141 ( .A1(n5907), .A2(n9745), .ZN(n5698) );
  OAI211_X1 U7142 ( .C1(n8035), .C2(n5700), .A(n5699), .B(n5698), .ZN(n5701)
         );
  INV_X1 U7143 ( .A(n5701), .ZN(n5702) );
  NAND2_X1 U7144 ( .A1(n5703), .A2(n5702), .ZN(n9512) );
  NAND2_X1 U7145 ( .A1(n9512), .A2(n5175), .ZN(n5704) );
  NAND2_X1 U7146 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  XNOR2_X1 U7147 ( .A(n5706), .B(n5038), .ZN(n5708) );
  INV_X1 U7148 ( .A(n9512), .ZN(n9550) );
  OAI22_X1 U7149 ( .A1(n9747), .A2(n5061), .B1(n9550), .B2(n5040), .ZN(n5707)
         );
  XNOR2_X1 U7150 ( .A(n5708), .B(n5707), .ZN(n9203) );
  NOR2_X1 U7151 ( .A1(n5708), .A2(n5707), .ZN(n9271) );
  INV_X1 U7152 ( .A(n5711), .ZN(n5713) );
  NAND2_X1 U7153 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  MUX2_X1 U7154 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n5716), .Z(n5741) );
  INV_X1 U7155 ( .A(SI_26_), .ZN(n7082) );
  XNOR2_X1 U7156 ( .A(n5741), .B(n7082), .ZN(n5739) );
  NAND2_X1 U7157 ( .A1(n7762), .A2(n8172), .ZN(n5718) );
  INV_X1 U7158 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7767) );
  OR2_X1 U7159 ( .A1(n8173), .A2(n7767), .ZN(n5717) );
  NAND2_X1 U7160 ( .A1(n9665), .A2(n5774), .ZN(n5732) );
  INV_X1 U7161 ( .A(n5721), .ZN(n5719) );
  NAND2_X1 U7162 ( .A1(n5719), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5746) );
  INV_X1 U7163 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7164 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  NAND2_X1 U7165 ( .A1(n5746), .A2(n5722), .ZN(n9276) );
  INV_X1 U7166 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5727) );
  INV_X1 U7167 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5723) );
  OR2_X1 U7168 ( .A1(n5907), .A2(n5723), .ZN(n5726) );
  INV_X1 U7169 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5724) );
  OR2_X1 U7170 ( .A1(n5095), .A2(n5724), .ZN(n5725) );
  OAI211_X1 U7171 ( .C1(n8035), .C2(n5727), .A(n5726), .B(n5725), .ZN(n5728)
         );
  INV_X1 U7172 ( .A(n5728), .ZN(n5729) );
  NAND2_X1 U7173 ( .A1(n5730), .A2(n5729), .ZN(n9524) );
  NAND2_X1 U7174 ( .A1(n9524), .A2(n5175), .ZN(n5731) );
  NAND2_X1 U7175 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  XNOR2_X1 U7176 ( .A(n5733), .B(n5188), .ZN(n5735) );
  AND2_X1 U7177 ( .A1(n9524), .A2(n5754), .ZN(n5734) );
  AOI21_X1 U7178 ( .B1(n9665), .B2(n4351), .A(n5734), .ZN(n5736) );
  XNOR2_X1 U7179 ( .A(n5735), .B(n5736), .ZN(n9270) );
  INV_X1 U7180 ( .A(n5735), .ZN(n5738) );
  INV_X1 U7181 ( .A(n5736), .ZN(n5737) );
  INV_X1 U7182 ( .A(n5741), .ZN(n5742) );
  NAND2_X1 U7183 ( .A1(n5742), .A2(n7082), .ZN(n5743) );
  MUX2_X1 U7184 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n4349), .Z(n5759) );
  INV_X1 U7185 ( .A(SI_27_), .ZN(n7144) );
  XNOR2_X1 U7186 ( .A(n5759), .B(n7144), .ZN(n5757) );
  NAND2_X1 U7187 ( .A1(n7778), .A2(n8172), .ZN(n5745) );
  INV_X1 U7188 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8330) );
  OR2_X1 U7189 ( .A1(n8173), .A2(n8330), .ZN(n5744) );
  INV_X1 U7190 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U7191 ( .A1(n5746), .A2(n6554), .ZN(n5747) );
  NAND2_X1 U7192 ( .A1(n9475), .A2(n5747), .ZN(n9488) );
  INV_X1 U7193 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9487) );
  INV_X1 U7194 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9662) );
  OR2_X1 U7195 ( .A1(n5095), .A2(n9662), .ZN(n5749) );
  INV_X1 U7196 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9740) );
  OR2_X1 U7197 ( .A1(n5907), .A2(n9740), .ZN(n5748) );
  OAI211_X1 U7198 ( .C1(n8035), .C2(n9487), .A(n5749), .B(n5748), .ZN(n5750)
         );
  INV_X1 U7199 ( .A(n5750), .ZN(n5751) );
  AOI22_X1 U7200 ( .A1(n9486), .A2(n5774), .B1(n4351), .B2(n9513), .ZN(n5753)
         );
  XNOR2_X1 U7201 ( .A(n5753), .B(n5038), .ZN(n5756) );
  AOI22_X1 U7202 ( .A1(n9486), .A2(n4351), .B1(n5754), .B2(n9513), .ZN(n5755)
         );
  NAND2_X1 U7203 ( .A1(n5756), .A2(n5755), .ZN(n5827) );
  OAI21_X1 U7204 ( .B1(n5756), .B2(n5755), .A(n5827), .ZN(n6549) );
  INV_X1 U7205 ( .A(n5759), .ZN(n5760) );
  MUX2_X1 U7206 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4350), .Z(n5874) );
  INV_X1 U7207 ( .A(SI_28_), .ZN(n7151) );
  XNOR2_X1 U7208 ( .A(n5874), .B(n7151), .ZN(n5872) );
  NAND2_X1 U7209 ( .A1(n7854), .A2(n8172), .ZN(n5762) );
  INV_X1 U7210 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7855) );
  OR2_X1 U7211 ( .A1(n8173), .A2(n7855), .ZN(n5761) );
  NAND2_X1 U7212 ( .A1(n8151), .A2(n4351), .ZN(n5772) );
  XNOR2_X1 U7213 ( .A(n9475), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U7214 ( .A1(n8336), .A2(n5763), .ZN(n5770) );
  INV_X1 U7215 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5767) );
  INV_X1 U7216 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7217 ( .A1(n5907), .A2(n5944), .ZN(n5766) );
  INV_X1 U7218 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5764) );
  OR2_X1 U7219 ( .A1(n5095), .A2(n5764), .ZN(n5765) );
  OAI211_X1 U7220 ( .C1(n8035), .C2(n5767), .A(n5766), .B(n5765), .ZN(n5768)
         );
  INV_X1 U7221 ( .A(n5768), .ZN(n5769) );
  OR2_X1 U7222 ( .A1(n9496), .A2(n5040), .ZN(n5771) );
  NAND2_X1 U7223 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  XNOR2_X1 U7224 ( .A(n5773), .B(n5188), .ZN(n5777) );
  NAND2_X1 U7225 ( .A1(n8151), .A2(n5774), .ZN(n5775) );
  OAI21_X1 U7226 ( .B1(n9496), .B2(n5061), .A(n5775), .ZN(n5776) );
  XNOR2_X1 U7227 ( .A(n5777), .B(n5776), .ZN(n5804) );
  INV_X1 U7228 ( .A(n5781), .ZN(n7667) );
  NAND2_X1 U7229 ( .A1(n7667), .A2(P1_B_REG_SCAN_IN), .ZN(n5778) );
  MUX2_X1 U7230 ( .A(n5778), .B(P1_B_REG_SCAN_IN), .S(n7552), .Z(n5780) );
  NAND2_X1 U7231 ( .A1(n5780), .A2(n5779), .ZN(n5912) );
  OR2_X1 U7232 ( .A1(n5781), .A2(n5779), .ZN(n9774) );
  OAI21_X1 U7233 ( .B1(n5912), .B2(P1_D_REG_1__SCAN_IN), .A(n9774), .ZN(n6812)
         );
  NOR2_X1 U7234 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5785) );
  NOR4_X1 U7235 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5784) );
  NOR4_X1 U7236 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5783) );
  NOR4_X1 U7237 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5782) );
  NAND4_X1 U7238 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n5791)
         );
  NOR4_X1 U7239 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5789) );
  NOR4_X1 U7240 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5788) );
  NOR4_X1 U7241 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5787) );
  NOR4_X1 U7242 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5786) );
  NAND4_X1 U7243 ( .A1(n5789), .A2(n5788), .A3(n5787), .A4(n5786), .ZN(n5790)
         );
  NOR2_X1 U7244 ( .A1(n5791), .A2(n5790), .ZN(n5913) );
  NOR2_X1 U7245 ( .A1(n5912), .A2(n5913), .ZN(n5792) );
  NOR2_X1 U7246 ( .A1(n6812), .A2(n5792), .ZN(n5795) );
  INV_X1 U7247 ( .A(n5912), .ZN(n5794) );
  INV_X1 U7248 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5793) );
  NOR2_X1 U7249 ( .A1(n5779), .A2(n7552), .ZN(n6603) );
  AOI21_X1 U7250 ( .B1(n5794), .B2(n5793), .A(n6603), .ZN(n5922) );
  AND2_X1 U7251 ( .A1(n5795), .A2(n5922), .ZN(n5805) );
  INV_X1 U7252 ( .A(n8326), .ZN(n8254) );
  INV_X1 U7253 ( .A(n8264), .ZN(n6924) );
  NAND2_X1 U7254 ( .A1(n8254), .A2(n6924), .ZN(n7248) );
  INV_X1 U7255 ( .A(n7248), .ZN(n5797) );
  AND2_X1 U7256 ( .A1(n5796), .A2(n5797), .ZN(n9726) );
  AND2_X1 U7257 ( .A1(n8326), .A2(n8264), .ZN(n8213) );
  OR2_X1 U7258 ( .A1(n9726), .A2(n8213), .ZN(n5819) );
  INV_X1 U7259 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7260 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  NAND2_X1 U7261 ( .A1(n5800), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5802) );
  INV_X1 U7262 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5801) );
  XNOR2_X1 U7263 ( .A(n5802), .B(n5801), .ZN(n6609) );
  AND2_X1 U7264 ( .A1(n6609), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6560) );
  INV_X1 U7265 ( .A(n6613), .ZN(n8325) );
  NOR2_X1 U7266 ( .A1(n5819), .A2(n8325), .ZN(n5803) );
  NAND3_X1 U7267 ( .A1(n6553), .A2(n5804), .A3(n9274), .ZN(n5834) );
  INV_X1 U7268 ( .A(n5804), .ZN(n5828) );
  INV_X1 U7269 ( .A(n5805), .ZN(n5821) );
  NOR2_X1 U7270 ( .A1(n7248), .A2(n5818), .ZN(n6817) );
  NAND2_X1 U7271 ( .A1(n6613), .A2(n6817), .ZN(n5806) );
  OR2_X1 U7272 ( .A1(n5821), .A2(n5806), .ZN(n5807) );
  INV_X1 U7273 ( .A(n5818), .ZN(n8324) );
  OR2_X1 U7274 ( .A1(n5882), .A2(n8264), .ZN(n5917) );
  INV_X1 U7275 ( .A(n5796), .ZN(n8319) );
  NAND2_X1 U7276 ( .A1(n6613), .A2(n8319), .ZN(n5808) );
  OR2_X1 U7277 ( .A1(n5821), .A2(n5808), .ZN(n5816) );
  INV_X1 U7278 ( .A(n7856), .ZN(n6677) );
  AND2_X1 U7279 ( .A1(n6677), .A2(n8213), .ZN(n9643) );
  INV_X1 U7280 ( .A(n9643), .ZN(n9549) );
  NOR2_X2 U7281 ( .A1(n5816), .A2(n9549), .ZN(n9277) );
  INV_X1 U7282 ( .A(n9277), .ZN(n9252) );
  INV_X1 U7283 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9474) );
  OR2_X1 U7284 ( .A1(n5069), .A2(n9474), .ZN(n5809) );
  OR2_X1 U7285 ( .A1(n9475), .A2(n5809), .ZN(n5815) );
  INV_X1 U7286 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5812) );
  INV_X1 U7287 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5925) );
  OR2_X1 U7288 ( .A1(n5907), .A2(n5925), .ZN(n5811) );
  INV_X1 U7289 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7290 ( .A1(n5095), .A2(n5918), .ZN(n5810) );
  OAI211_X1 U7291 ( .C1(n8035), .C2(n5812), .A(n5811), .B(n5810), .ZN(n5813)
         );
  INV_X1 U7292 ( .A(n5813), .ZN(n5814) );
  AND2_X1 U7293 ( .A1(n7856), .A2(n8213), .ZN(n9644) );
  NOR2_X2 U7294 ( .A1(n5816), .A2(n9551), .ZN(n9250) );
  AOI22_X1 U7295 ( .A1(n4837), .A2(n9250), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5826) );
  INV_X1 U7296 ( .A(n8213), .ZN(n5817) );
  OR2_X1 U7297 ( .A1(n5796), .A2(n5817), .ZN(n7249) );
  OR2_X1 U7298 ( .A1(n5818), .A2(P1_U3086), .ZN(n6791) );
  NAND3_X1 U7299 ( .A1(n5819), .A2(n7249), .A3(n6791), .ZN(n5820) );
  NAND2_X1 U7300 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  NAND2_X1 U7301 ( .A1(n5796), .A2(n8213), .ZN(n5915) );
  NAND2_X1 U7302 ( .A1(n5822), .A2(n5915), .ZN(n6649) );
  OAI21_X1 U7303 ( .B1(n6649), .B2(n5823), .A(P1_STATE_REG_SCAN_IN), .ZN(n5824) );
  OR2_X1 U7304 ( .A1(n6609), .A2(P1_U3086), .ZN(n8329) );
  INV_X1 U7305 ( .A(n9260), .ZN(n9282) );
  NAND2_X1 U7306 ( .A1(n8336), .A2(n9282), .ZN(n5825) );
  OAI211_X1 U7307 ( .C1(n9280), .C2(n9252), .A(n5826), .B(n5825), .ZN(n5830)
         );
  NOR3_X1 U7308 ( .A1(n5828), .A2(n5827), .A3(n9267), .ZN(n5829) );
  AOI211_X1 U7309 ( .C1(n8151), .C2(n9265), .A(n5830), .B(n5829), .ZN(n5831)
         );
  INV_X1 U7310 ( .A(n5831), .ZN(n5832) );
  NAND2_X1 U7311 ( .A1(n5834), .A2(n5833), .ZN(P1_U3220) );
  NAND2_X1 U7312 ( .A1(n9302), .A2(n6709), .ZN(n6706) );
  XNOR2_X1 U7313 ( .A(n9300), .B(n5835), .ZN(n6711) );
  NAND2_X1 U7314 ( .A1(n5041), .A2(n5835), .ZN(n5836) );
  NAND2_X1 U7315 ( .A1(n6705), .A2(n5836), .ZN(n6702) );
  NAND2_X1 U7316 ( .A1(n6750), .A2(n6818), .ZN(n8075) );
  NAND2_X1 U7317 ( .A1(n6702), .A2(n8218), .ZN(n6701) );
  NAND2_X1 U7318 ( .A1(n6750), .A2(n6735), .ZN(n5837) );
  NAND2_X1 U7319 ( .A1(n6701), .A2(n5837), .ZN(n6746) );
  NAND2_X1 U7320 ( .A1(n6910), .A2(n6754), .ZN(n8268) );
  NAND2_X1 U7321 ( .A1(n9298), .A2(n6837), .ZN(n8071) );
  NAND2_X1 U7322 ( .A1(n8268), .A2(n8071), .ZN(n8219) );
  NAND2_X1 U7323 ( .A1(n6746), .A2(n8219), .ZN(n6745) );
  NAND2_X1 U7324 ( .A1(n6910), .A2(n6837), .ZN(n5838) );
  NAND2_X1 U7325 ( .A1(n6745), .A2(n5838), .ZN(n6912) );
  NAND2_X1 U7326 ( .A1(n6785), .A2(n6918), .ZN(n8068) );
  NAND2_X1 U7327 ( .A1(n6625), .A2(n9959), .ZN(n8070) );
  NAND2_X1 U7328 ( .A1(n8068), .A2(n8070), .ZN(n8220) );
  NAND2_X1 U7329 ( .A1(n6932), .A2(n6786), .ZN(n8080) );
  INV_X1 U7330 ( .A(n6932), .ZN(n9297) );
  AND2_X1 U7331 ( .A1(n8220), .A2(n8225), .ZN(n5840) );
  INV_X1 U7332 ( .A(n8225), .ZN(n5839) );
  NAND2_X1 U7333 ( .A1(n6785), .A2(n9959), .ZN(n6780) );
  NAND2_X1 U7334 ( .A1(n6932), .A2(n6981), .ZN(n5841) );
  NAND2_X1 U7335 ( .A1(n6882), .A2(n6943), .ZN(n8082) );
  INV_X1 U7336 ( .A(n6882), .ZN(n9296) );
  NAND2_X1 U7337 ( .A1(n9296), .A2(n9964), .ZN(n6846) );
  NAND2_X1 U7338 ( .A1(n8082), .A2(n6846), .ZN(n6937) );
  NAND2_X1 U7339 ( .A1(n6931), .A2(n6902), .ZN(n8091) );
  INV_X1 U7340 ( .A(n6931), .ZN(n9295) );
  NAND2_X1 U7341 ( .A1(n9295), .A2(n6904), .ZN(n8090) );
  NAND2_X1 U7342 ( .A1(n8091), .A2(n8090), .ZN(n6879) );
  NAND2_X1 U7343 ( .A1(n6877), .A2(n6879), .ZN(n6876) );
  NAND2_X1 U7344 ( .A1(n6931), .A2(n6904), .ZN(n5842) );
  NAND2_X1 U7345 ( .A1(n6876), .A2(n5842), .ZN(n6844) );
  NAND2_X1 U7346 ( .A1(n6881), .A2(n6853), .ZN(n8101) );
  NAND2_X1 U7347 ( .A1(n8101), .A2(n8093), .ZN(n6850) );
  NAND2_X1 U7348 ( .A1(n6844), .A2(n6850), .ZN(n6843) );
  NAND2_X1 U7349 ( .A1(n6881), .A2(n4765), .ZN(n5843) );
  NAND2_X1 U7350 ( .A1(n6843), .A2(n5843), .ZN(n6976) );
  OR2_X1 U7351 ( .A1(n7263), .A2(n9968), .ZN(n8102) );
  NAND2_X1 U7352 ( .A1(n9968), .A2(n7263), .ZN(n8113) );
  NAND2_X1 U7353 ( .A1(n8102), .A2(n8113), .ZN(n6975) );
  NAND2_X1 U7354 ( .A1(n6976), .A2(n6975), .ZN(n6974) );
  OR2_X1 U7355 ( .A1(n9968), .A2(n9293), .ZN(n5844) );
  NAND2_X1 U7356 ( .A1(n6974), .A2(n5844), .ZN(n6957) );
  OR2_X1 U7357 ( .A1(n7679), .A2(n7605), .ZN(n8279) );
  NAND2_X1 U7358 ( .A1(n7679), .A2(n7605), .ZN(n8115) );
  NAND2_X1 U7359 ( .A1(n8279), .A2(n8115), .ZN(n6956) );
  NAND2_X1 U7360 ( .A1(n6957), .A2(n6956), .ZN(n6955) );
  OR2_X1 U7361 ( .A1(n7679), .A2(n9292), .ZN(n5845) );
  NAND2_X1 U7362 ( .A1(n6955), .A2(n5845), .ZN(n7217) );
  OR2_X1 U7363 ( .A1(n7610), .A2(n6952), .ZN(n8118) );
  NAND2_X1 U7364 ( .A1(n7610), .A2(n6952), .ZN(n8116) );
  NAND2_X1 U7365 ( .A1(n8118), .A2(n8116), .ZN(n8230) );
  NAND2_X1 U7366 ( .A1(n7217), .A2(n8230), .ZN(n7216) );
  OR2_X1 U7367 ( .A1(n7610), .A2(n9291), .ZN(n5846) );
  NAND2_X1 U7368 ( .A1(n7216), .A2(n5846), .ZN(n7285) );
  OR2_X1 U7369 ( .A1(n7380), .A2(n7546), .ZN(n8119) );
  NAND2_X1 U7370 ( .A1(n7380), .A2(n7546), .ZN(n8284) );
  NAND2_X1 U7371 ( .A1(n8119), .A2(n8284), .ZN(n8232) );
  NAND2_X1 U7372 ( .A1(n7285), .A2(n8232), .ZN(n7284) );
  INV_X1 U7373 ( .A(n7380), .ZN(n7400) );
  NAND2_X1 U7374 ( .A1(n7400), .A2(n7546), .ZN(n5847) );
  NAND2_X1 U7375 ( .A1(n7284), .A2(n5847), .ZN(n7384) );
  OR2_X1 U7376 ( .A1(n7549), .A2(n7559), .ZN(n8121) );
  NAND2_X1 U7377 ( .A1(n7549), .A2(n7559), .ZN(n8261) );
  NAND2_X1 U7378 ( .A1(n8121), .A2(n8261), .ZN(n7390) );
  OR2_X1 U7379 ( .A1(n7549), .A2(n9289), .ZN(n5848) );
  NAND2_X1 U7380 ( .A1(n7383), .A2(n5848), .ZN(n7556) );
  NAND2_X1 U7381 ( .A1(n9725), .A2(n7943), .ZN(n5849) );
  NAND2_X1 U7382 ( .A1(n7556), .A2(n5849), .ZN(n5851) );
  OR2_X1 U7383 ( .A1(n9725), .A2(n7943), .ZN(n5850) );
  NAND2_X1 U7384 ( .A1(n7947), .A2(n9288), .ZN(n5852) );
  OR2_X1 U7385 ( .A1(n9720), .A2(n7941), .ZN(n8063) );
  NAND2_X1 U7386 ( .A1(n9720), .A2(n7941), .ZN(n8108) );
  NAND2_X1 U7387 ( .A1(n8063), .A2(n8108), .ZN(n7688) );
  NAND2_X1 U7388 ( .A1(n9720), .A2(n7831), .ZN(n5853) );
  OR2_X1 U7389 ( .A1(n7866), .A2(n9287), .ZN(n5854) );
  NAND2_X1 U7390 ( .A1(n5855), .A2(n5854), .ZN(n7925) );
  NAND2_X1 U7391 ( .A1(n9709), .A2(n9642), .ZN(n5856) );
  AND2_X1 U7392 ( .A1(n9628), .A2(n9610), .ZN(n5857) );
  NOR2_X1 U7393 ( .A1(n9615), .A2(n9645), .ZN(n5858) );
  NAND2_X1 U7394 ( .A1(n9615), .A2(n9645), .ZN(n5859) );
  AND2_X1 U7395 ( .A1(n9597), .A2(n9611), .ZN(n9570) );
  AND2_X1 U7396 ( .A1(n9688), .A2(n9593), .ZN(n5862) );
  OR2_X1 U7397 ( .A1(n9597), .A2(n9611), .ZN(n9571) );
  OR2_X1 U7398 ( .A1(n9688), .A2(n9593), .ZN(n5860) );
  AND2_X1 U7399 ( .A1(n9571), .A2(n5860), .ZN(n5861) );
  OR2_X1 U7400 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  NOR2_X1 U7401 ( .A1(n9562), .A2(n9583), .ZN(n5866) );
  NAND2_X1 U7402 ( .A1(n9562), .A2(n9583), .ZN(n5865) );
  OR2_X1 U7403 ( .A1(n9676), .A2(n9560), .ZN(n5867) );
  OR2_X1 U7404 ( .A1(n9529), .A2(n9512), .ZN(n5868) );
  NOR2_X1 U7405 ( .A1(n9665), .A2(n9524), .ZN(n5870) );
  NAND2_X1 U7406 ( .A1(n9665), .A2(n9524), .ZN(n5869) );
  NAND2_X1 U7407 ( .A1(n9486), .A2(n9280), .ZN(n8156) );
  NAND2_X1 U7408 ( .A1(n8151), .A2(n9496), .ZN(n8158) );
  OR2_X1 U7409 ( .A1(n9486), .A2(n9513), .ZN(n5930) );
  NAND2_X1 U7410 ( .A1(n5873), .A2(n5872), .ZN(n5877) );
  INV_X1 U7411 ( .A(n5874), .ZN(n5875) );
  NAND2_X1 U7412 ( .A1(n5875), .A2(n7151), .ZN(n5876) );
  INV_X1 U7413 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9173) );
  INV_X1 U7414 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8015) );
  MUX2_X1 U7415 ( .A(n9173), .B(n8015), .S(n5716), .Z(n8020) );
  OR2_X1 U7416 ( .A1(n8173), .A2(n8015), .ZN(n5878) );
  NAND2_X1 U7417 ( .A1(n5883), .A2(n5936), .ZN(n8166) );
  XNOR2_X1 U7418 ( .A(n5879), .B(n8250), .ZN(n9472) );
  NAND2_X1 U7419 ( .A1(n5796), .A2(n5880), .ZN(n5881) );
  NAND3_X1 U7420 ( .A1(n7249), .A2(n7248), .A3(n5881), .ZN(n6806) );
  INV_X1 U7421 ( .A(n9665), .ZN(n9508) );
  INV_X1 U7422 ( .A(n9688), .ZN(n9579) );
  INV_X1 U7423 ( .A(n5835), .ZN(n5887) );
  OR2_X1 U7424 ( .A1(n5887), .A2(n6709), .ZN(n6707) );
  NAND2_X1 U7425 ( .A1(n6747), .A2(n6837), .ZN(n6748) );
  INV_X1 U7426 ( .A(n7679), .ZN(n9976) );
  INV_X1 U7427 ( .A(n7610), .ZN(n7220) );
  NAND2_X1 U7428 ( .A1(n6959), .A2(n7220), .ZN(n7218) );
  INV_X1 U7429 ( .A(n7947), .ZN(n7788) );
  INV_X1 U7430 ( .A(n5884), .ZN(n7824) );
  INV_X1 U7431 ( .A(n9709), .ZN(n7935) );
  INV_X1 U7432 ( .A(n9628), .ZN(n9765) );
  NOR2_X2 U7433 ( .A1(n9597), .A2(n9614), .ZN(n9596) );
  NAND2_X1 U7434 ( .A1(n9579), .A2(n9596), .ZN(n9574) );
  INV_X1 U7435 ( .A(n5942), .ZN(n5886) );
  AOI211_X1 U7436 ( .C1(n5883), .C2(n5886), .A(n9682), .B(n9465), .ZN(n9473)
         );
  INV_X1 U7437 ( .A(n6711), .ZN(n8221) );
  INV_X1 U7438 ( .A(n6709), .ZN(n7252) );
  NAND2_X1 U7439 ( .A1(n8221), .A2(n6710), .ZN(n5889) );
  NAND2_X1 U7440 ( .A1(n5041), .A2(n5887), .ZN(n5888) );
  NAND2_X1 U7441 ( .A1(n5889), .A2(n5888), .ZN(n8074) );
  INV_X1 U7442 ( .A(n8075), .ZN(n5890) );
  OR2_X1 U7443 ( .A1(n8074), .A2(n5890), .ZN(n8067) );
  NAND2_X1 U7444 ( .A1(n8067), .A2(n8266), .ZN(n8269) );
  OAI21_X1 U7445 ( .B1(n8269), .B2(n8219), .A(n8268), .ZN(n6908) );
  NAND2_X1 U7446 ( .A1(n6908), .A2(n8070), .ZN(n6845) );
  AND2_X1 U7447 ( .A1(n8080), .A2(n8068), .ZN(n8271) );
  NAND2_X1 U7448 ( .A1(n6845), .A2(n8271), .ZN(n5891) );
  NAND2_X1 U7449 ( .A1(n5891), .A2(n8275), .ZN(n6929) );
  AND2_X1 U7450 ( .A1(n8102), .A2(n8093), .ZN(n5893) );
  NAND2_X1 U7451 ( .A1(n8091), .A2(n8101), .ZN(n8095) );
  AND2_X1 U7452 ( .A1(n5892), .A2(n8082), .ZN(n8276) );
  NAND2_X1 U7453 ( .A1(n6929), .A2(n8276), .ZN(n6948) );
  INV_X1 U7454 ( .A(n6956), .ZN(n8228) );
  NAND2_X1 U7455 ( .A1(n6948), .A2(n5894), .ZN(n6950) );
  INV_X1 U7456 ( .A(n8230), .ZN(n7214) );
  INV_X1 U7457 ( .A(n8232), .ZN(n7282) );
  NAND2_X1 U7458 ( .A1(n7280), .A2(n8284), .ZN(n7391) );
  NAND2_X1 U7459 ( .A1(n7391), .A2(n8121), .ZN(n5895) );
  NAND2_X1 U7460 ( .A1(n5895), .A2(n8261), .ZN(n7557) );
  INV_X1 U7461 ( .A(n7943), .ZN(n5896) );
  OR2_X1 U7462 ( .A1(n9725), .A2(n5896), .ZN(n8124) );
  NAND2_X1 U7463 ( .A1(n9725), .A2(n5896), .ZN(n8105) );
  INV_X1 U7464 ( .A(n9288), .ZN(n9218) );
  OR2_X1 U7465 ( .A1(n7947), .A2(n9218), .ZN(n7686) );
  NAND2_X1 U7466 ( .A1(n7947), .A2(n9218), .ZN(n8106) );
  NAND2_X1 U7467 ( .A1(n7686), .A2(n8106), .ZN(n8237) );
  AND2_X1 U7468 ( .A1(n8063), .A2(n7686), .ZN(n8291) );
  INV_X1 U7469 ( .A(n9287), .ZN(n7691) );
  OR2_X1 U7470 ( .A1(n7866), .A2(n7691), .ZN(n8046) );
  NAND2_X1 U7471 ( .A1(n7866), .A2(n7691), .ZN(n8129) );
  NAND2_X1 U7472 ( .A1(n8046), .A2(n8129), .ZN(n7828) );
  INV_X1 U7473 ( .A(n8108), .ZN(n8298) );
  NOR2_X1 U7474 ( .A1(n7828), .A2(n8298), .ZN(n5897) );
  NAND2_X1 U7475 ( .A1(n7830), .A2(n5897), .ZN(n7827) );
  NAND2_X1 U7476 ( .A1(n7827), .A2(n8046), .ZN(n7926) );
  NAND2_X1 U7477 ( .A1(n7935), .A2(n9642), .ZN(n9636) );
  INV_X1 U7478 ( .A(n9642), .ZN(n5898) );
  NAND2_X1 U7479 ( .A1(n9709), .A2(n5898), .ZN(n8051) );
  NAND2_X1 U7480 ( .A1(n7926), .A2(n7927), .ZN(n9637) );
  INV_X1 U7481 ( .A(n9610), .ZN(n9262) );
  OR2_X1 U7482 ( .A1(n9628), .A2(n9262), .ZN(n8242) );
  AND2_X1 U7483 ( .A1(n8242), .A2(n9636), .ZN(n8296) );
  NAND2_X1 U7484 ( .A1(n9637), .A2(n8296), .ZN(n5899) );
  NAND2_X1 U7485 ( .A1(n9628), .A2(n9262), .ZN(n8241) );
  NAND2_X1 U7486 ( .A1(n5899), .A2(n8241), .ZN(n9608) );
  XNOR2_X1 U7487 ( .A(n9615), .B(n9645), .ZN(n9607) );
  NAND2_X1 U7488 ( .A1(n9608), .A2(n9607), .ZN(n9606) );
  INV_X1 U7489 ( .A(n9645), .ZN(n8041) );
  NAND2_X1 U7490 ( .A1(n9615), .A2(n8041), .ZN(n8058) );
  INV_X1 U7491 ( .A(n9611), .ZN(n9253) );
  OR2_X1 U7492 ( .A1(n9597), .A2(n9253), .ZN(n8195) );
  NAND2_X1 U7493 ( .A1(n9597), .A2(n9253), .ZN(n8131) );
  INV_X1 U7494 ( .A(n9593), .ZN(n9183) );
  OR2_X1 U7495 ( .A1(n9688), .A2(n9183), .ZN(n8039) );
  NAND2_X1 U7496 ( .A1(n9688), .A2(n9183), .ZN(n8040) );
  NAND2_X1 U7497 ( .A1(n9580), .A2(n8040), .ZN(n9557) );
  INV_X1 U7498 ( .A(n9583), .ZN(n9548) );
  OR2_X1 U7499 ( .A1(n9562), .A2(n9548), .ZN(n8137) );
  NAND2_X1 U7500 ( .A1(n9562), .A2(n9548), .ZN(n9543) );
  NAND2_X1 U7501 ( .A1(n9557), .A2(n9558), .ZN(n9556) );
  INV_X1 U7502 ( .A(n9560), .ZN(n9206) );
  OR2_X1 U7503 ( .A1(n9676), .A2(n9206), .ZN(n8185) );
  NAND2_X1 U7504 ( .A1(n9676), .A2(n9206), .ZN(n8198) );
  NAND3_X1 U7505 ( .A1(n9556), .A2(n9545), .A3(n9543), .ZN(n5900) );
  NAND2_X1 U7506 ( .A1(n5900), .A2(n8185), .ZN(n9520) );
  OR2_X1 U7507 ( .A1(n9529), .A2(n9550), .ZN(n8152) );
  NAND2_X1 U7508 ( .A1(n9529), .A2(n9550), .ZN(n8200) );
  NAND2_X1 U7509 ( .A1(n8152), .A2(n8200), .ZN(n9519) );
  NAND2_X1 U7510 ( .A1(n9522), .A2(n8200), .ZN(n9510) );
  INV_X1 U7511 ( .A(n9524), .ZN(n9495) );
  OR2_X1 U7512 ( .A1(n9665), .A2(n9495), .ZN(n8153) );
  NAND2_X1 U7513 ( .A1(n9665), .A2(n9495), .ZN(n8190) );
  NAND2_X1 U7514 ( .A1(n9510), .A2(n9511), .ZN(n9509) );
  AND2_X1 U7515 ( .A1(n8158), .A2(n8156), .ZN(n8205) );
  INV_X1 U7516 ( .A(n8143), .ZN(n8206) );
  NAND2_X1 U7517 ( .A1(n4485), .A2(n8326), .ZN(n5902) );
  NAND2_X1 U7518 ( .A1(n8264), .A2(n8324), .ZN(n5901) );
  INV_X1 U7519 ( .A(n5904), .ZN(n6665) );
  NAND2_X1 U7520 ( .A1(n6665), .A2(P1_B_REG_SCAN_IN), .ZN(n5905) );
  AND2_X1 U7521 ( .A1(n9644), .A2(n5905), .ZN(n9460) );
  INV_X1 U7522 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9657) );
  INV_X1 U7523 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5906) );
  OR2_X1 U7524 ( .A1(n8035), .A2(n5906), .ZN(n5909) );
  INV_X1 U7525 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9736) );
  OR2_X1 U7526 ( .A1(n5907), .A2(n9736), .ZN(n5908) );
  OAI211_X1 U7527 ( .C1(n5095), .C2(n9657), .A(n5909), .B(n5908), .ZN(n9286)
         );
  AOI22_X1 U7528 ( .A1(n6874), .A2(n9643), .B1(n9460), .B2(n9286), .ZN(n5910)
         );
  NAND2_X1 U7529 ( .A1(n5911), .A2(n5910), .ZN(n9481) );
  AOI211_X1 U7530 ( .C1(n9472), .C2(n9978), .A(n9473), .B(n9481), .ZN(n5924)
         );
  NAND2_X2 U7531 ( .A1(n6613), .A2(n5912), .ZN(n9957) );
  NAND2_X1 U7532 ( .A1(n6613), .A2(n5913), .ZN(n5914) );
  NAND2_X1 U7533 ( .A1(n9957), .A2(n5914), .ZN(n5916) );
  AND2_X1 U7534 ( .A1(n6812), .A2(n5917), .ZN(n5923) );
  AND3_X2 U7535 ( .A1(n6814), .A2(n5923), .A3(n5922), .ZN(n9988) );
  MUX2_X1 U7536 ( .A(n5918), .B(n5924), .S(n9988), .Z(n5921) );
  NAND2_X1 U7537 ( .A1(n9988), .A2(n9726), .ZN(n9717) );
  NAND2_X1 U7538 ( .A1(n5921), .A2(n5920), .ZN(P1_U3551) );
  INV_X1 U7539 ( .A(n5922), .ZN(n6815) );
  AND3_X2 U7540 ( .A1(n6815), .A2(n6814), .A3(n5923), .ZN(n9981) );
  MUX2_X1 U7541 ( .A(n5925), .B(n5924), .S(n9981), .Z(n5928) );
  NAND2_X1 U7542 ( .A1(n9981), .A2(n9726), .ZN(n9770) );
  NAND2_X1 U7543 ( .A1(n5928), .A2(n5927), .ZN(P1_U3519) );
  AOI21_X1 U7544 ( .B1(n5931), .B2(n5930), .A(n5929), .ZN(n5933) );
  INV_X1 U7545 ( .A(n9978), .ZN(n9728) );
  NAND2_X1 U7546 ( .A1(n9491), .A2(n8156), .ZN(n5934) );
  XNOR2_X1 U7547 ( .A(n5934), .B(n8248), .ZN(n5935) );
  NAND2_X1 U7548 ( .A1(n5935), .A2(n9640), .ZN(n5939) );
  OAI22_X1 U7549 ( .A1(n9280), .A2(n9549), .B1(n5936), .B2(n9551), .ZN(n5937)
         );
  INV_X1 U7550 ( .A(n5937), .ZN(n5938) );
  NAND2_X1 U7551 ( .A1(n5939), .A2(n5938), .ZN(n8341) );
  NAND2_X1 U7552 ( .A1(n8151), .A2(n9485), .ZN(n5940) );
  INV_X1 U7553 ( .A(n9682), .ZN(n7288) );
  NAND2_X1 U7554 ( .A1(n5940), .A2(n7288), .ZN(n5941) );
  NOR2_X1 U7555 ( .A1(n5942), .A2(n5941), .ZN(n8335) );
  NOR2_X1 U7556 ( .A1(n8341), .A2(n8335), .ZN(n5943) );
  INV_X1 U7557 ( .A(n5948), .ZN(n5947) );
  INV_X1 U7558 ( .A(n8151), .ZN(n8339) );
  NAND2_X1 U7559 ( .A1(n8151), .A2(n5919), .ZN(n5949) );
  XNOR2_X1 U7560 ( .A(n5950), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9178) );
  INV_X1 U7561 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5996) );
  INV_X1 U7562 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5953) );
  NOR2_X1 U7563 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5958) );
  NOR2_X1 U7564 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5957) );
  NOR2_X1 U7565 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5956) );
  NOR2_X1 U7566 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5955) );
  NOR2_X1 U7567 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5961) );
  NOR2_X1 U7568 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5960) );
  NOR2_X1 U7569 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5959) );
  INV_X1 U7570 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6344) );
  INV_X1 U7571 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5963) );
  AND2_X1 U7572 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  INV_X1 U7573 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5970) );
  XNOR2_X2 U7574 ( .A(n5967), .B(n5970), .ZN(n6334) );
  MUX2_X1 U7575 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9178), .S(n5994), .Z(n6821) );
  INV_X1 U7576 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7577 ( .A1(n6288), .A2(n4953), .ZN(n9167) );
  NAND2_X1 U7578 ( .A1(n6288), .A2(n5971), .ZN(n5972) );
  NAND2_X1 U7579 ( .A1(n6263), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7580 ( .A1(n4958), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7581 ( .A1(n8539), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5977) );
  INV_X1 U7582 ( .A(n5974), .ZN(n8358) );
  NAND2_X1 U7583 ( .A1(n6012), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5976) );
  NAND4_X1 U7584 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n8784)
         );
  INV_X1 U7585 ( .A(n8784), .ZN(n5980) );
  NAND2_X1 U7586 ( .A1(n6263), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7587 ( .A1(n8539), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5982) );
  INV_X1 U7588 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7589 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5985) );
  INV_X1 U7590 ( .A(n7483), .ZN(n5987) );
  NAND2_X1 U7591 ( .A1(n6189), .A2(n5987), .ZN(n5988) );
  NAND2_X1 U7592 ( .A1(n8783), .A2(n10147), .ZN(n8599) );
  NAND2_X1 U7593 ( .A1(n4958), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7594 ( .A1(n6012), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7595 ( .A1(n8539), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7596 ( .A1(n6263), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7597 ( .A1(n5993), .A2(n6581), .ZN(n6000) );
  INV_X1 U7598 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6576) );
  OR2_X1 U7599 ( .A1(n6008), .A2(n6576), .ZN(n5999) );
  INV_X1 U7600 ( .A(n7487), .ZN(n5997) );
  OR2_X1 U7601 ( .A1(n8782), .A2(n6402), .ZN(n8604) );
  NAND2_X1 U7602 ( .A1(n8782), .A2(n6402), .ZN(n8605) );
  NAND2_X2 U7603 ( .A1(n8604), .A2(n8605), .ZN(n8563) );
  INV_X1 U7604 ( .A(n8563), .ZN(n7238) );
  NAND2_X1 U7605 ( .A1(n7236), .A2(n7238), .ZN(n6001) );
  NAND2_X1 U7606 ( .A1(n6001), .A2(n8604), .ZN(n7296) );
  INV_X1 U7607 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6002) );
  OR2_X1 U7608 ( .A1(n6167), .A2(n6002), .ZN(n6006) );
  INV_X1 U7609 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7306) );
  NAND2_X1 U7610 ( .A1(n4958), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6004) );
  OR2_X1 U7611 ( .A1(n6096), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6003) );
  OR2_X1 U7612 ( .A1(n5993), .A2(n6578), .ZN(n6010) );
  INV_X1 U7613 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6577) );
  OR2_X1 U7614 ( .A1(n6008), .A2(n6577), .ZN(n6009) );
  NAND2_X1 U7615 ( .A1(n6300), .A2(n10156), .ZN(n8617) );
  INV_X1 U7616 ( .A(n8562), .ZN(n7302) );
  NAND2_X1 U7617 ( .A1(n7296), .A2(n7302), .ZN(n7297) );
  NAND2_X1 U7618 ( .A1(n7297), .A2(n8617), .ZN(n10135) );
  AND2_X1 U7619 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6011) );
  NOR2_X1 U7620 ( .A1(n6035), .A2(n6011), .ZN(n10137) );
  OR2_X1 U7621 ( .A1(n6096), .A2(n10137), .ZN(n6016) );
  NAND2_X1 U7622 ( .A1(n4958), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7623 ( .A1(n8539), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7624 ( .A1(n6012), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6013) );
  NAND4_X1 U7625 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n8618)
         );
  NAND2_X1 U7626 ( .A1(n6017), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6019) );
  INV_X1 U7627 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6018) );
  XNOR2_X1 U7628 ( .A(n6019), .B(n6018), .ZN(n7413) );
  INV_X1 U7629 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6020) );
  OR2_X1 U7630 ( .A1(n6008), .A2(n6020), .ZN(n6022) );
  OR2_X1 U7631 ( .A1(n5993), .A2(n6583), .ZN(n6021) );
  XNOR2_X1 U7632 ( .A(n8618), .B(n10139), .ZN(n10136) );
  NAND2_X1 U7633 ( .A1(n10135), .A2(n10136), .ZN(n6023) );
  NAND2_X1 U7634 ( .A1(n7594), .A2(n10139), .ZN(n8613) );
  NAND2_X1 U7635 ( .A1(n6023), .A2(n8613), .ZN(n7589) );
  NAND2_X1 U7636 ( .A1(n6012), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6027) );
  XNOR2_X1 U7637 ( .A(n6035), .B(P2_REG3_REG_5__SCAN_IN), .ZN(n7591) );
  OR2_X1 U7638 ( .A1(n6096), .A2(n7591), .ZN(n6026) );
  NAND2_X1 U7639 ( .A1(n4958), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U7640 ( .A1(n8539), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6024) );
  NAND4_X1 U7641 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n10132)
         );
  OR2_X1 U7642 ( .A1(n6028), .A2(n9166), .ZN(n6030) );
  XNOR2_X1 U7643 ( .A(n6030), .B(n6029), .ZN(n10015) );
  OR2_X1 U7644 ( .A1(n5993), .A2(n6589), .ZN(n6032) );
  INV_X1 U7645 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6585) );
  OR2_X1 U7646 ( .A1(n6008), .A2(n6585), .ZN(n6031) );
  OAI211_X1 U7647 ( .C1(n6563), .C2(n10015), .A(n6032), .B(n6031), .ZN(n7228)
         );
  NAND2_X1 U7648 ( .A1(n7192), .A2(n7228), .ZN(n8623) );
  INV_X1 U7649 ( .A(n7228), .ZN(n10166) );
  NAND2_X1 U7650 ( .A1(n10132), .A2(n10166), .ZN(n8619) );
  NAND2_X1 U7651 ( .A1(n7589), .A2(n8566), .ZN(n7590) );
  NAND2_X1 U7652 ( .A1(n7590), .A2(n8623), .ZN(n7660) );
  NAND2_X1 U7653 ( .A1(n4958), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6041) );
  INV_X1 U7654 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7412) );
  OR2_X1 U7655 ( .A1(n6167), .A2(n7412), .ZN(n6040) );
  INV_X1 U7656 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7229) );
  NAND2_X1 U7657 ( .A1(n6035), .A2(n7229), .ZN(n6033) );
  NAND2_X1 U7658 ( .A1(n6033), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6036) );
  NOR2_X1 U7659 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .ZN(n6034) );
  NAND2_X1 U7660 ( .A1(n6035), .A2(n6034), .ZN(n6049) );
  AND2_X1 U7661 ( .A1(n6036), .A2(n6049), .ZN(n7661) );
  OR2_X1 U7662 ( .A1(n6096), .A2(n7661), .ZN(n6039) );
  INV_X1 U7663 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6037) );
  OR2_X1 U7664 ( .A1(n6281), .A2(n6037), .ZN(n6038) );
  NAND2_X1 U7665 ( .A1(n6042), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6044) );
  INV_X1 U7666 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6043) );
  XNOR2_X1 U7667 ( .A(n6044), .B(n6043), .ZN(n7441) );
  OR2_X1 U7668 ( .A1(n5993), .A2(n6587), .ZN(n6046) );
  INV_X1 U7669 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6586) );
  OR2_X1 U7670 ( .A1(n6008), .A2(n6586), .ZN(n6045) );
  OAI211_X1 U7671 ( .C1(n6563), .C2(n7441), .A(n6046), .B(n6045), .ZN(n10172)
         );
  NAND2_X1 U7672 ( .A1(n7595), .A2(n10172), .ZN(n8624) );
  INV_X1 U7673 ( .A(n8624), .ZN(n6047) );
  INV_X1 U7674 ( .A(n10172), .ZN(n7662) );
  NAND2_X1 U7675 ( .A1(n8781), .A2(n7662), .ZN(n8625) );
  OAI21_X1 U7676 ( .B1(n7660), .B2(n6047), .A(n8625), .ZN(n7531) );
  NAND2_X1 U7677 ( .A1(n6012), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6055) );
  INV_X1 U7678 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7679 ( .A1(n6280), .A2(n6048), .ZN(n6054) );
  NAND2_X1 U7680 ( .A1(n6049), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6050) );
  AND2_X1 U7681 ( .A1(n6061), .A2(n6050), .ZN(n7507) );
  OR2_X1 U7682 ( .A1(n6096), .A2(n7507), .ZN(n6053) );
  INV_X1 U7683 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6051) );
  OR2_X1 U7684 ( .A1(n6281), .A2(n6051), .ZN(n6052) );
  NAND2_X1 U7685 ( .A1(n4401), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6056) );
  MUX2_X1 U7686 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6056), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n6057) );
  NAND2_X1 U7687 ( .A1(n6057), .A2(n4369), .ZN(n7743) );
  OR2_X1 U7688 ( .A1(n5993), .A2(n6591), .ZN(n6059) );
  OR2_X1 U7689 ( .A1(n6008), .A2(n6590), .ZN(n6058) );
  OAI211_X1 U7690 ( .C1(n6563), .C2(n7743), .A(n6059), .B(n6058), .ZN(n7537)
         );
  NAND2_X1 U7691 ( .A1(n7656), .A2(n7537), .ZN(n8639) );
  INV_X1 U7692 ( .A(n7537), .ZN(n10178) );
  NAND2_X1 U7693 ( .A1(n7634), .A2(n10178), .ZN(n7516) );
  NAND2_X1 U7694 ( .A1(n7531), .A2(n8635), .ZN(n7515) );
  NAND2_X1 U7695 ( .A1(n6012), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6066) );
  INV_X1 U7696 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6060) );
  OR2_X1 U7697 ( .A1(n6280), .A2(n6060), .ZN(n6065) );
  AND2_X1 U7698 ( .A1(n6061), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6062) );
  NOR2_X1 U7699 ( .A1(n6071), .A2(n6062), .ZN(n7631) );
  OR2_X1 U7700 ( .A1(n6096), .A2(n7631), .ZN(n6064) );
  INV_X1 U7701 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7524) );
  OR2_X1 U7702 ( .A1(n6281), .A2(n7524), .ZN(n6063) );
  OR2_X1 U7703 ( .A1(n6008), .A2(n6604), .ZN(n6068) );
  NAND2_X1 U7704 ( .A1(n4369), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7705 ( .A(n6067), .B(n4923), .ZN(n10026) );
  INV_X1 U7706 ( .A(n7632), .ZN(n10182) );
  NAND2_X1 U7707 ( .A1(n8780), .A2(n10182), .ZN(n8631) );
  AND2_X1 U7708 ( .A1(n7516), .A2(n8631), .ZN(n8644) );
  NAND2_X1 U7709 ( .A1(n7515), .A2(n8644), .ZN(n6069) );
  NAND2_X1 U7710 ( .A1(n7511), .A2(n7632), .ZN(n8640) );
  NAND2_X1 U7711 ( .A1(n6069), .A2(n8640), .ZN(n7613) );
  INV_X1 U7712 ( .A(n7613), .ZN(n6082) );
  NAND2_X1 U7713 ( .A1(n6012), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7714 ( .A1(n4958), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6075) );
  INV_X1 U7715 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6070) );
  NOR2_X1 U7716 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  OR2_X1 U7717 ( .A1(n6086), .A2(n6072), .ZN(n7914) );
  NAND2_X1 U7718 ( .A1(n6263), .A2(n7914), .ZN(n6074) );
  NAND2_X1 U7719 ( .A1(n8539), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7720 ( .A1(n6077), .A2(n9166), .ZN(n6078) );
  XNOR2_X1 U7721 ( .A(n6078), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7796) );
  AOI22_X1 U7722 ( .A1(n6188), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6189), .B2(
        n7796), .ZN(n6080) );
  NAND2_X1 U7723 ( .A1(n6594), .A2(n8544), .ZN(n6085) );
  OR2_X1 U7724 ( .A1(n4425), .A2(n9166), .ZN(n6083) );
  XNOR2_X1 U7725 ( .A(n6083), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7875) );
  AOI22_X1 U7726 ( .A1(n6188), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6189), .B2(
        n7875), .ZN(n6084) );
  NAND2_X1 U7727 ( .A1(n6085), .A2(n6084), .ZN(n6092) );
  NAND2_X1 U7728 ( .A1(n4958), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6091) );
  INV_X1 U7729 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7735) );
  OR2_X1 U7730 ( .A1(n6167), .A2(n7735), .ZN(n6090) );
  INV_X1 U7731 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7754) );
  OR2_X1 U7732 ( .A1(n6086), .A2(n7754), .ZN(n6087) );
  AND2_X1 U7733 ( .A1(n6094), .A2(n6087), .ZN(n7846) );
  OR2_X1 U7734 ( .A1(n6096), .A2(n7846), .ZN(n6089) );
  INV_X1 U7735 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7736) );
  OR2_X1 U7736 ( .A1(n6281), .A2(n7736), .ZN(n6088) );
  NAND2_X1 U7737 ( .A1(n7711), .A2(n8778), .ZN(n8654) );
  AND2_X1 U7738 ( .A1(n8654), .A2(n8632), .ZN(n8643) );
  NAND2_X1 U7739 ( .A1(n7908), .A2(n6092), .ZN(n8651) );
  INV_X1 U7740 ( .A(n8651), .ZN(n6093) );
  NAND2_X1 U7741 ( .A1(n6012), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7742 ( .A1(n6094), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6095) );
  AND2_X1 U7743 ( .A1(n6109), .A2(n6095), .ZN(n7896) );
  OR2_X1 U7744 ( .A1(n6096), .A2(n7896), .ZN(n6099) );
  NAND2_X1 U7745 ( .A1(n4958), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7746 ( .A1(n8539), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6097) );
  NAND4_X1 U7747 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n8777)
         );
  NAND2_X1 U7748 ( .A1(n6597), .A2(n8544), .ZN(n6104) );
  OR2_X1 U7749 ( .A1(n6101), .A2(n9166), .ZN(n6102) );
  XNOR2_X1 U7750 ( .A(n6102), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7975) );
  AOI22_X1 U7751 ( .A1(n6188), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6189), .B2(
        n7975), .ZN(n6103) );
  NAND2_X1 U7752 ( .A1(n10201), .A2(n7961), .ZN(n8656) );
  NAND2_X1 U7753 ( .A1(n6619), .A2(n8544), .ZN(n6108) );
  NAND2_X1 U7754 ( .A1(n6105), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6106) );
  XNOR2_X1 U7755 ( .A(n6106), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7988) );
  AOI22_X1 U7756 ( .A1(n6188), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6189), .B2(
        n7988), .ZN(n6107) );
  NAND2_X1 U7757 ( .A1(n4958), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6114) );
  INV_X1 U7758 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7980) );
  OR2_X1 U7759 ( .A1(n6167), .A2(n7980), .ZN(n6113) );
  NAND2_X1 U7760 ( .A1(n6109), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6110) );
  AND2_X1 U7761 ( .A1(n6117), .A2(n6110), .ZN(n7819) );
  OR2_X1 U7762 ( .A1(n6096), .A2(n7819), .ZN(n6112) );
  INV_X1 U7763 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7976) );
  OR2_X1 U7764 ( .A1(n6281), .A2(n7976), .ZN(n6111) );
  NOR2_X1 U7765 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  NAND2_X1 U7766 ( .A1(n6627), .A2(n8544), .ZN(n6116) );
  OR2_X1 U7767 ( .A1(n6105), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7768 ( .A1(n6148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6123) );
  XNOR2_X1 U7769 ( .A(n6123), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U7770 ( .A1(n6188), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6189), .B2(
        n10042), .ZN(n6115) );
  INV_X1 U7771 ( .A(n8479), .ZN(n8669) );
  NAND2_X1 U7772 ( .A1(n4958), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6122) );
  AND2_X1 U7773 ( .A1(n6117), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6118) );
  NOR2_X1 U7774 ( .A1(n6127), .A2(n6118), .ZN(n8471) );
  OR2_X1 U7775 ( .A1(n6096), .A2(n8471), .ZN(n6121) );
  NAND2_X1 U7776 ( .A1(n8539), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7777 ( .A1(n6012), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7778 ( .A1(n6631), .A2(n8544), .ZN(n6126) );
  INV_X1 U7779 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7780 ( .A1(n6123), .A2(n6145), .ZN(n6124) );
  NAND2_X1 U7781 ( .A1(n6124), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6133) );
  XNOR2_X1 U7782 ( .A(n6133), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10058) );
  AOI22_X1 U7783 ( .A1(n6188), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6189), .B2(
        n10058), .ZN(n6125) );
  NAND2_X1 U7784 ( .A1(n4958), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6132) );
  INV_X1 U7785 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8825) );
  OR2_X1 U7786 ( .A1(n6167), .A2(n8825), .ZN(n6131) );
  INV_X1 U7787 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7055) );
  OR2_X1 U7788 ( .A1(n6127), .A2(n7055), .ZN(n6128) );
  AND2_X1 U7789 ( .A1(n6128), .A2(n6138), .ZN(n8370) );
  OR2_X1 U7790 ( .A1(n6096), .A2(n8370), .ZN(n6130) );
  INV_X1 U7791 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8009) );
  OR2_X1 U7792 ( .A1(n6281), .A2(n8009), .ZN(n6129) );
  NOR2_X1 U7793 ( .A1(n8372), .A2(n6433), .ZN(n8678) );
  NAND2_X1 U7794 ( .A1(n8372), .A2(n6433), .ZN(n7997) );
  NAND2_X1 U7795 ( .A1(n6635), .A2(n8544), .ZN(n6137) );
  INV_X1 U7796 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7797 ( .A1(n6133), .A2(n6146), .ZN(n6134) );
  NAND2_X1 U7798 ( .A1(n6134), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6135) );
  XNOR2_X1 U7799 ( .A(n6135), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10074) );
  AOI22_X1 U7800 ( .A1(n6188), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6189), .B2(
        n10074), .ZN(n6136) );
  NAND2_X1 U7801 ( .A1(n4958), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6143) );
  INV_X1 U7802 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9074) );
  OR2_X1 U7803 ( .A1(n6167), .A2(n9074), .ZN(n6142) );
  NAND2_X1 U7804 ( .A1(n6138), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6139) );
  AND2_X1 U7805 ( .A1(n6152), .A2(n6139), .ZN(n9022) );
  OR2_X1 U7806 ( .A1(n6096), .A2(n9022), .ZN(n6141) );
  INV_X1 U7807 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10083) );
  OR2_X1 U7808 ( .A1(n6281), .A2(n10083), .ZN(n6140) );
  OR2_X1 U7809 ( .A1(n9160), .A2(n8366), .ZN(n8683) );
  NAND2_X1 U7810 ( .A1(n6653), .A2(n8544), .ZN(n6151) );
  INV_X1 U7811 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6144) );
  NAND3_X1 U7812 ( .A1(n6146), .A2(n6145), .A3(n6144), .ZN(n6147) );
  OR2_X1 U7813 ( .A1(n6159), .A2(n9166), .ZN(n6149) );
  XNOR2_X1 U7814 ( .A(n6149), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U7815 ( .A1(n6188), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6189), .B2(
        n10090), .ZN(n6150) );
  NAND2_X1 U7816 ( .A1(n4958), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6157) );
  INV_X1 U7817 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9071) );
  OR2_X1 U7818 ( .A1(n6167), .A2(n9071), .ZN(n6156) );
  AND2_X1 U7819 ( .A1(n6152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6153) );
  NOR2_X1 U7820 ( .A1(n6169), .A2(n6153), .ZN(n9012) );
  OR2_X1 U7821 ( .A1(n6096), .A2(n9012), .ZN(n6155) );
  INV_X1 U7822 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9011) );
  OR2_X1 U7823 ( .A1(n6281), .A2(n9011), .ZN(n6154) );
  NAND2_X1 U7824 ( .A1(n9154), .A2(n8774), .ZN(n8688) );
  NAND2_X1 U7825 ( .A1(n6715), .A2(n8544), .ZN(n6166) );
  INV_X1 U7826 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6158) );
  NOR2_X1 U7827 ( .A1(n6163), .A2(n9166), .ZN(n6160) );
  MUX2_X1 U7828 ( .A(n9166), .B(n6160), .S(P2_IR_REG_17__SCAN_IN), .Z(n6161)
         );
  INV_X1 U7829 ( .A(n6161), .ZN(n6164) );
  INV_X1 U7830 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6162) );
  AND2_X1 U7831 ( .A1(n6164), .A2(n6185), .ZN(n10108) );
  AOI22_X1 U7832 ( .A1(n6189), .A2(n10108), .B1(n6188), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7833 ( .A1(n4958), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6175) );
  INV_X1 U7834 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9068) );
  OR2_X1 U7835 ( .A1(n6167), .A2(n9068), .ZN(n6174) );
  INV_X1 U7836 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6168) );
  NOR2_X1 U7837 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  OR2_X1 U7838 ( .A1(n6179), .A2(n6170), .ZN(n9002) );
  INV_X1 U7839 ( .A(n9002), .ZN(n6171) );
  OR2_X1 U7840 ( .A1(n6096), .A2(n6171), .ZN(n6173) );
  INV_X1 U7841 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10119) );
  OR2_X1 U7842 ( .A1(n6281), .A2(n10119), .ZN(n6172) );
  NAND2_X1 U7843 ( .A1(n9148), .A2(n8431), .ZN(n8559) );
  NAND2_X1 U7844 ( .A1(n6739), .A2(n8544), .ZN(n6178) );
  NAND2_X1 U7845 ( .A1(n6185), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6176) );
  XNOR2_X1 U7846 ( .A(n6176), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U7847 ( .A1(n6188), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9805), .B2(
        n6189), .ZN(n6177) );
  INV_X1 U7848 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9065) );
  OR2_X1 U7849 ( .A1(n6167), .A2(n9065), .ZN(n6184) );
  INV_X1 U7850 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7070) );
  OR2_X1 U7851 ( .A1(n6179), .A2(n7070), .ZN(n6180) );
  AND2_X1 U7852 ( .A1(n6192), .A2(n6180), .ZN(n8993) );
  OR2_X1 U7853 ( .A1(n6096), .A2(n8993), .ZN(n6183) );
  NAND2_X1 U7854 ( .A1(n4958), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7855 ( .A1(n8539), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6181) );
  NAND4_X1 U7856 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n9000)
         );
  NAND2_X1 U7857 ( .A1(n8503), .A2(n9000), .ZN(n8987) );
  NAND2_X1 U7858 ( .A1(n8987), .A2(n8983), .ZN(n8690) );
  NAND2_X1 U7859 ( .A1(n9142), .A2(n8973), .ZN(n8986) );
  NAND2_X1 U7860 ( .A1(n6776), .A2(n8544), .ZN(n6191) );
  INV_X1 U7861 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6186) );
  AOI22_X1 U7862 ( .A1(n8762), .A2(n6189), .B1(n6188), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7863 ( .A1(n4958), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6197) );
  INV_X1 U7864 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9063) );
  OR2_X1 U7865 ( .A1(n6167), .A2(n9063), .ZN(n6196) );
  NAND2_X1 U7866 ( .A1(n6192), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6193) );
  AND2_X1 U7867 ( .A1(n6200), .A2(n6193), .ZN(n8978) );
  OR2_X1 U7868 ( .A1(n6096), .A2(n8978), .ZN(n6195) );
  INV_X1 U7869 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8979) );
  OR2_X1 U7870 ( .A1(n6281), .A2(n8979), .ZN(n6194) );
  NAND2_X1 U7871 ( .A1(n9062), .A2(n8498), .ZN(n8707) );
  INV_X1 U7872 ( .A(n8707), .ZN(n8698) );
  NAND2_X1 U7873 ( .A1(n6827), .A2(n8544), .ZN(n6199) );
  INV_X1 U7874 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6828) );
  OR2_X1 U7875 ( .A1(n6008), .A2(n6828), .ZN(n6198) );
  NAND2_X1 U7876 ( .A1(n6012), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6205) );
  INV_X1 U7877 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9131) );
  OR2_X1 U7878 ( .A1(n6280), .A2(n9131), .ZN(n6204) );
  AND2_X1 U7879 ( .A1(n6200), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6201) );
  NOR2_X1 U7880 ( .A1(n6209), .A2(n6201), .ZN(n8461) );
  OR2_X1 U7881 ( .A1(n6096), .A2(n8461), .ZN(n6203) );
  INV_X1 U7882 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8964) );
  OR2_X1 U7883 ( .A1(n6281), .A2(n8964), .ZN(n6202) );
  INV_X1 U7884 ( .A(n8710), .ZN(n6206) );
  NAND2_X1 U7885 ( .A1(n9132), .A2(n8975), .ZN(n8708) );
  NAND2_X1 U7886 ( .A1(n6923), .A2(n8544), .ZN(n6208) );
  INV_X1 U7887 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6926) );
  OR2_X1 U7888 ( .A1(n6008), .A2(n6926), .ZN(n6207) );
  INV_X1 U7889 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8406) );
  NOR2_X1 U7890 ( .A1(n6209), .A2(n8406), .ZN(n6210) );
  OR2_X1 U7891 ( .A1(n6219), .A2(n6210), .ZN(n8954) );
  NAND2_X1 U7892 ( .A1(n6263), .A2(n8954), .ZN(n6214) );
  INV_X1 U7893 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9055) );
  OR2_X1 U7894 ( .A1(n6167), .A2(n9055), .ZN(n6213) );
  INV_X1 U7895 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9125) );
  OR2_X1 U7896 ( .A1(n6280), .A2(n9125), .ZN(n6212) );
  INV_X1 U7897 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8953) );
  OR2_X1 U7898 ( .A1(n6281), .A2(n8953), .ZN(n6211) );
  NAND2_X1 U7899 ( .A1(n9126), .A2(n6443), .ZN(n8713) );
  INV_X1 U7900 ( .A(n8713), .ZN(n6215) );
  OAI21_X1 U7901 ( .B1(n8944), .B2(n6215), .A(n8711), .ZN(n8940) );
  NAND2_X1 U7902 ( .A1(n7257), .A2(n8544), .ZN(n6217) );
  INV_X1 U7903 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7258) );
  OR2_X1 U7904 ( .A1(n6008), .A2(n7258), .ZN(n6216) );
  INV_X1 U7905 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6218) );
  OR2_X1 U7906 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  NAND2_X1 U7907 ( .A1(n6231), .A2(n6220), .ZN(n8934) );
  NAND2_X1 U7908 ( .A1(n6263), .A2(n8934), .ZN(n6226) );
  INV_X1 U7909 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6221) );
  OR2_X1 U7910 ( .A1(n6167), .A2(n6221), .ZN(n6225) );
  INV_X1 U7911 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6222) );
  OR2_X1 U7912 ( .A1(n6280), .A2(n6222), .ZN(n6224) );
  INV_X1 U7913 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8936) );
  OR2_X1 U7914 ( .A1(n6281), .A2(n8936), .ZN(n6223) );
  NAND2_X1 U7915 ( .A1(n8940), .A2(n8939), .ZN(n8941) );
  OR2_X1 U7916 ( .A1(n8938), .A2(n8921), .ZN(n8702) );
  NAND2_X1 U7917 ( .A1(n7321), .A2(n8544), .ZN(n6228) );
  INV_X1 U7918 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7320) );
  OR2_X1 U7919 ( .A1(n6008), .A2(n7320), .ZN(n6227) );
  NAND2_X1 U7920 ( .A1(n6012), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7921 ( .A1(n4958), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6229) );
  AND2_X1 U7922 ( .A1(n6230), .A2(n6229), .ZN(n6235) );
  NAND2_X1 U7923 ( .A1(n6231), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7924 ( .A1(n6238), .A2(n6232), .ZN(n8925) );
  NAND2_X1 U7925 ( .A1(n8925), .A2(n6263), .ZN(n6234) );
  NAND2_X1 U7926 ( .A1(n8539), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7927 ( .A1(n7553), .A2(n8544), .ZN(n6237) );
  INV_X1 U7928 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8360) );
  OR2_X1 U7929 ( .A1(n6008), .A2(n8360), .ZN(n6236) );
  INV_X1 U7930 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U7931 ( .A1(n6238), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7932 ( .A1(n6244), .A2(n6239), .ZN(n8908) );
  NAND2_X1 U7933 ( .A1(n8908), .A2(n6263), .ZN(n6241) );
  AOI22_X1 U7934 ( .A1(n6012), .A2(P2_REG1_REG_24__SCAN_IN), .B1(n4958), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n6240) );
  OAI211_X1 U7935 ( .C1(n6281), .C2(n8915), .A(n6241), .B(n6240), .ZN(n8894)
         );
  INV_X1 U7936 ( .A(n8894), .ZN(n8922) );
  NAND2_X1 U7937 ( .A1(n9113), .A2(n8922), .ZN(n8557) );
  NAND2_X1 U7938 ( .A1(n8926), .A2(n8488), .ZN(n8912) );
  NAND2_X1 U7939 ( .A1(n7666), .A2(n8544), .ZN(n6243) );
  INV_X1 U7940 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8356) );
  OR2_X1 U7941 ( .A1(n6008), .A2(n8356), .ZN(n6242) );
  AND2_X1 U7942 ( .A1(n6244), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6245) );
  OR2_X1 U7943 ( .A1(n6245), .A2(n6251), .ZN(n8897) );
  NAND2_X1 U7944 ( .A1(n8897), .A2(n6263), .ZN(n6248) );
  AOI22_X1 U7945 ( .A1(n6012), .A2(P2_REG1_REG_25__SCAN_IN), .B1(n4958), .B2(
        P2_REG0_REG_25__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7946 ( .A1(n8539), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7947 ( .A1(n9107), .A2(n8773), .ZN(n8726) );
  INV_X1 U7948 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7763) );
  OR2_X1 U7949 ( .A1(n6008), .A2(n7763), .ZN(n6249) );
  INV_X1 U7950 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8510) );
  NOR2_X1 U7951 ( .A1(n6251), .A2(n8510), .ZN(n6252) );
  NAND2_X1 U7952 ( .A1(n8886), .A2(n6263), .ZN(n6257) );
  INV_X1 U7953 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U7954 ( .A1(n8539), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7955 ( .A1(n4958), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6253) );
  OAI211_X1 U7956 ( .C1(n6167), .C2(n9039), .A(n6254), .B(n6253), .ZN(n6255)
         );
  INV_X1 U7957 ( .A(n6255), .ZN(n6256) );
  NAND2_X1 U7958 ( .A1(n9101), .A2(n8420), .ZN(n8556) );
  INV_X1 U7959 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6258) );
  OR2_X1 U7960 ( .A1(n6008), .A2(n6258), .ZN(n6259) );
  INV_X1 U7961 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7008) );
  OR2_X1 U7962 ( .A1(n6261), .A2(n7008), .ZN(n6262) );
  NAND2_X1 U7963 ( .A1(n6262), .A2(n6271), .ZN(n8876) );
  NAND2_X1 U7964 ( .A1(n8876), .A2(n6263), .ZN(n6268) );
  INV_X1 U7965 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U7966 ( .A1(n8539), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7967 ( .A1(n4958), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6264) );
  OAI211_X1 U7968 ( .C1(n6167), .C2(n9036), .A(n6265), .B(n6264), .ZN(n6266)
         );
  INV_X1 U7969 ( .A(n6266), .ZN(n6267) );
  OAI21_X2 U7970 ( .B1(n8870), .B2(n8733), .A(n8555), .ZN(n8856) );
  NAND2_X1 U7971 ( .A1(n7854), .A2(n8544), .ZN(n6270) );
  INV_X1 U7972 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7853) );
  OR2_X1 U7973 ( .A1(n6008), .A2(n7853), .ZN(n6269) );
  NAND2_X1 U7974 ( .A1(n6012), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6276) );
  INV_X1 U7975 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9088) );
  OR2_X1 U7976 ( .A1(n6280), .A2(n9088), .ZN(n6275) );
  AND2_X1 U7977 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n6271), .ZN(n6272) );
  NOR2_X1 U7978 ( .A1(n8849), .A2(n6272), .ZN(n8866) );
  OR2_X1 U7979 ( .A1(n6096), .A2(n8866), .ZN(n6274) );
  INV_X1 U7980 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8865) );
  OR2_X1 U7981 ( .A1(n6281), .A2(n8865), .ZN(n6273) );
  INV_X1 U7982 ( .A(n9089), .ZN(n8752) );
  NAND2_X1 U7983 ( .A1(n8752), .A2(n8873), .ZN(n6277) );
  NAND2_X1 U7984 ( .A1(n8014), .A2(n8544), .ZN(n6279) );
  OR2_X1 U7985 ( .A1(n6008), .A2(n9173), .ZN(n6278) );
  INV_X1 U7986 ( .A(n8849), .ZN(n6389) );
  INV_X1 U7987 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6535) );
  OR2_X1 U7988 ( .A1(n6280), .A2(n6535), .ZN(n6284) );
  INV_X1 U7989 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6390) );
  OR2_X1 U7990 ( .A1(n6281), .A2(n6390), .ZN(n6283) );
  INV_X1 U7991 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6544) );
  OR2_X1 U7992 ( .A1(n6167), .A2(n6544), .ZN(n6282) );
  NAND2_X1 U7993 ( .A1(n6536), .A2(n8772), .ZN(n8537) );
  INV_X1 U7994 ( .A(n6288), .ZN(n6285) );
  NAND2_X1 U7995 ( .A1(n6285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6287) );
  INV_X1 U7996 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6286) );
  INV_X1 U7997 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7998 ( .A1(n4370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6290) );
  INV_X1 U7999 ( .A(n6291), .ZN(n6292) );
  NAND2_X1 U8000 ( .A1(n6292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6293) );
  MUX2_X1 U8001 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6293), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6294) );
  OR2_X1 U8002 ( .A1(n6399), .A2(n4354), .ZN(n7367) );
  INV_X1 U8003 ( .A(n8767), .ZN(n8597) );
  OAI21_X1 U8004 ( .B1(n8767), .B2(n8755), .A(n10186), .ZN(n6295) );
  NOR2_X1 U8005 ( .A1(n8762), .A2(n6295), .ZN(n6296) );
  NAND2_X1 U8006 ( .A1(n7367), .A2(n6296), .ZN(n7622) );
  NAND2_X1 U8007 ( .A1(n8784), .A2(n6821), .ZN(n7465) );
  NAND2_X1 U8008 ( .A1(n7463), .A2(n7465), .ZN(n7239) );
  NAND2_X1 U8009 ( .A1(n10147), .A2(n4928), .ZN(n7240) );
  NAND2_X1 U8010 ( .A1(n7239), .A2(n7240), .ZN(n6297) );
  NAND2_X1 U8011 ( .A1(n6297), .A2(n8563), .ZN(n7237) );
  INV_X1 U8012 ( .A(n6402), .ZN(n6298) );
  OR2_X1 U8013 ( .A1(n8782), .A2(n6298), .ZN(n7301) );
  NAND2_X1 U8014 ( .A1(n7237), .A2(n7301), .ZN(n6299) );
  NAND2_X1 U8015 ( .A1(n6299), .A2(n8562), .ZN(n7304) );
  NAND2_X1 U8016 ( .A1(n6300), .A2(n6406), .ZN(n6301) );
  NAND2_X1 U8017 ( .A1(n7304), .A2(n6301), .ZN(n10128) );
  NAND2_X1 U8018 ( .A1(n8618), .A2(n10139), .ZN(n6302) );
  NAND2_X1 U8019 ( .A1(n10128), .A2(n6302), .ZN(n6304) );
  INV_X1 U8020 ( .A(n10139), .ZN(n10162) );
  NAND2_X1 U8021 ( .A1(n7594), .A2(n10162), .ZN(n6303) );
  NAND2_X1 U8022 ( .A1(n6304), .A2(n6303), .ZN(n7592) );
  NOR2_X1 U8023 ( .A1(n10132), .A2(n7228), .ZN(n6306) );
  NAND2_X1 U8024 ( .A1(n10132), .A2(n7228), .ZN(n6305) );
  OAI21_X1 U8025 ( .B1(n7592), .B2(n6306), .A(n6305), .ZN(n7654) );
  NAND2_X1 U8026 ( .A1(n8624), .A2(n8625), .ZN(n8568) );
  NAND2_X1 U8027 ( .A1(n7654), .A2(n8568), .ZN(n6308) );
  NAND2_X1 U8028 ( .A1(n8781), .A2(n10172), .ZN(n6307) );
  NAND2_X1 U8029 ( .A1(n6308), .A2(n6307), .ZN(n7518) );
  NAND2_X1 U8030 ( .A1(n8651), .A2(n8654), .ZN(n8574) );
  INV_X1 U8031 ( .A(n10187), .ZN(n7904) );
  INV_X1 U8032 ( .A(n7701), .ZN(n6309) );
  NAND2_X1 U8033 ( .A1(n8574), .A2(n6309), .ZN(n6312) );
  INV_X1 U8034 ( .A(n6312), .ZN(n6311) );
  NAND2_X1 U8035 ( .A1(n8780), .A2(n7632), .ZN(n7616) );
  AND2_X1 U8036 ( .A1(n7615), .A2(n8574), .ZN(n6310) );
  NAND2_X1 U8037 ( .A1(n8640), .A2(n8631), .ZN(n8571) );
  NAND2_X1 U8038 ( .A1(n7656), .A2(n10178), .ZN(n7520) );
  AND2_X1 U8039 ( .A1(n8571), .A2(n7520), .ZN(n7519) );
  AND2_X1 U8040 ( .A1(n7519), .A2(n6312), .ZN(n6313) );
  NAND2_X1 U8041 ( .A1(n7908), .A2(n7711), .ZN(n6315) );
  NAND2_X1 U8042 ( .A1(n10201), .A2(n8777), .ZN(n6317) );
  NOR2_X1 U8043 ( .A1(n8479), .A2(n8775), .ZN(n8668) );
  NAND2_X1 U8044 ( .A1(n8479), .A2(n8775), .ZN(n8674) );
  NOR2_X1 U8045 ( .A1(n6429), .A2(n6433), .ZN(n6318) );
  OAI22_X1 U8046 ( .A1(n7996), .A2(n6318), .B1(n8372), .B2(n9019), .ZN(n9018)
         );
  AOI21_X1 U8047 ( .B1(n8560), .B2(n8366), .A(n9018), .ZN(n6319) );
  INV_X1 U8048 ( .A(n9154), .ZN(n8436) );
  NAND2_X1 U8049 ( .A1(n8983), .A2(n8559), .ZN(n8999) );
  NAND2_X1 U8050 ( .A1(n9142), .A2(n9000), .ZN(n6321) );
  INV_X1 U8051 ( .A(n8498), .ZN(n8991) );
  NAND2_X1 U8052 ( .A1(n8710), .A2(n8708), .ZN(n8960) );
  NAND2_X1 U8053 ( .A1(n8961), .A2(n8960), .ZN(n8959) );
  INV_X1 U8054 ( .A(n9132), .ZN(n8466) );
  NAND2_X1 U8055 ( .A1(n8466), .A2(n8975), .ZN(n8946) );
  NAND2_X1 U8056 ( .A1(n8959), .A2(n8946), .ZN(n6323) );
  NAND2_X1 U8057 ( .A1(n8711), .A2(n8713), .ZN(n8945) );
  NAND2_X1 U8058 ( .A1(n6323), .A2(n8945), .ZN(n8949) );
  INV_X1 U8059 ( .A(n9126), .ZN(n8411) );
  NAND2_X1 U8060 ( .A1(n8411), .A2(n6443), .ZN(n6324) );
  NAND2_X1 U8061 ( .A1(n8949), .A2(n6324), .ZN(n8930) );
  INV_X1 U8062 ( .A(n8938), .ZN(n9054) );
  NAND2_X1 U8063 ( .A1(n9054), .A2(n8921), .ZN(n6325) );
  NOR2_X1 U8064 ( .A1(n9113), .A2(n8894), .ZN(n6326) );
  INV_X1 U8065 ( .A(n9107), .ZN(n8900) );
  NAND2_X1 U8066 ( .A1(n8900), .A2(n8773), .ZN(n6327) );
  INV_X1 U8067 ( .A(n9101), .ZN(n8517) );
  NOR2_X1 U8068 ( .A1(n9095), .A2(n8883), .ZN(n6329) );
  NAND2_X1 U8069 ( .A1(n9095), .A2(n8883), .ZN(n6328) );
  NAND2_X1 U8070 ( .A1(n8859), .A2(n8585), .ZN(n6331) );
  NAND2_X1 U8071 ( .A1(n9089), .A2(n8873), .ZN(n6330) );
  NAND2_X1 U8072 ( .A1(n6331), .A2(n6330), .ZN(n6332) );
  XNOR2_X1 U8073 ( .A(n6332), .B(n8738), .ZN(n6342) );
  NAND2_X1 U8074 ( .A1(n8762), .A2(n8767), .ZN(n6333) );
  INV_X1 U8075 ( .A(n8755), .ZN(n6483) );
  NAND2_X1 U8076 ( .A1(n8592), .A2(n6483), .ZN(n8550) );
  INV_X1 U8077 ( .A(n6334), .ZN(n8764) );
  INV_X1 U8078 ( .A(n8806), .ZN(n8811) );
  NAND2_X1 U8079 ( .A1(n8764), .A2(n8811), .ZN(n6335) );
  NAND2_X1 U8080 ( .A1(n6563), .A2(n6335), .ZN(n6513) );
  NAND2_X1 U8081 ( .A1(n6513), .A2(n8747), .ZN(n8976) );
  AND2_X1 U8082 ( .A1(n6563), .A2(P2_B_REG_SCAN_IN), .ZN(n6336) );
  NOR2_X1 U8083 ( .A1(n8976), .A2(n6336), .ZN(n8847) );
  NAND2_X1 U8084 ( .A1(n6012), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U8085 ( .A1(n4958), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8086 ( .A1(n8539), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6337) );
  NAND4_X1 U8087 ( .A1(n8543), .A2(n6339), .A3(n6338), .A4(n6337), .ZN(n8771)
         );
  INV_X1 U8088 ( .A(n6513), .ZN(n6511) );
  AND2_X2 U8089 ( .A1(n6511), .A2(n8747), .ZN(n10129) );
  AOI22_X1 U8090 ( .A1(n8847), .A2(n8771), .B1(n8873), .B2(n10129), .ZN(n6340)
         );
  AOI21_X1 U8091 ( .B1(n6342), .B2(n10134), .A(n6341), .ZN(n6343) );
  INV_X1 U8092 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6379) );
  INV_X1 U8093 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8094 ( .A1(n6350), .A2(n6355), .ZN(n6348) );
  OR2_X1 U8095 ( .A1(n9166), .A2(n6355), .ZN(n6349) );
  INV_X1 U8096 ( .A(n6349), .ZN(n6345) );
  NAND2_X1 U8097 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  NAND2_X1 U8098 ( .A1(n6348), .A2(n6347), .ZN(n6361) );
  XNOR2_X1 U8099 ( .A(n6361), .B(P2_B_REG_SCAN_IN), .ZN(n6352) );
  INV_X1 U8100 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U8101 ( .A1(n6352), .A2(n6364), .ZN(n6360) );
  NAND3_X1 U8102 ( .A1(n6355), .A2(n6379), .A3(n6354), .ZN(n6356) );
  OAI21_X1 U8103 ( .B1(n6353), .B2(n6356), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6357) );
  MUX2_X1 U8104 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6357), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6358) );
  AND2_X1 U8105 ( .A1(n6359), .A2(n6358), .ZN(n6362) );
  NAND2_X1 U8106 ( .A1(n6360), .A2(n6362), .ZN(n6363) );
  INV_X1 U8107 ( .A(n6362), .ZN(n7764) );
  NAND2_X1 U8108 ( .A1(n6361), .A2(n7764), .ZN(n6762) );
  NAND2_X1 U8109 ( .A1(n6398), .A2(n6762), .ZN(n6487) );
  OR2_X1 U8110 ( .A1(n6363), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U8111 ( .A1(n6364), .A2(n7764), .ZN(n6365) );
  NAND2_X1 U8112 ( .A1(n6366), .A2(n6365), .ZN(n6639) );
  NOR2_X1 U8113 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6370) );
  NOR4_X1 U8114 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6369) );
  NOR4_X1 U8115 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6368) );
  NOR4_X1 U8116 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6367) );
  NAND4_X1 U8117 ( .A1(n6370), .A2(n6369), .A3(n6368), .A4(n6367), .ZN(n6376)
         );
  NOR4_X1 U8118 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6374) );
  NOR4_X1 U8119 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6373) );
  NOR4_X1 U8120 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6372) );
  NOR4_X1 U8121 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6371) );
  NAND4_X1 U8122 ( .A1(n6374), .A2(n6373), .A3(n6372), .A4(n6371), .ZN(n6375)
         );
  NOR2_X1 U8123 ( .A1(n6376), .A2(n6375), .ZN(n6377) );
  XNOR2_X1 U8124 ( .A(n6378), .B(n6379), .ZN(n6565) );
  NAND2_X1 U8125 ( .A1(n6399), .A2(n8747), .ZN(n6502) );
  NAND3_X1 U8126 ( .A1(n6486), .A2(n6686), .A3(n6502), .ZN(n6540) );
  AOI21_X1 U8127 ( .B1(n6487), .B2(n6639), .A(n6540), .ZN(n6386) );
  NAND3_X1 U8128 ( .A1(n4353), .A2(n8767), .A3(n6483), .ZN(n6380) );
  NAND2_X1 U8129 ( .A1(n6380), .A2(n4354), .ZN(n6381) );
  OR2_X1 U8130 ( .A1(n6487), .A2(n6381), .ZN(n6384) );
  INV_X1 U8131 ( .A(n6381), .ZN(n6382) );
  OR2_X1 U8132 ( .A1(n6639), .A2(n6382), .ZN(n6383) );
  NAND2_X1 U8133 ( .A1(n6384), .A2(n6383), .ZN(n6543) );
  INV_X1 U8134 ( .A(n6543), .ZN(n6385) );
  NAND2_X1 U8135 ( .A1(n6386), .A2(n6385), .ZN(n6388) );
  NAND2_X1 U8136 ( .A1(n8762), .A2(n8755), .ZN(n6387) );
  NOR2_X1 U8137 ( .A1(n10192), .A2(n8592), .ZN(n6539) );
  INV_X2 U8138 ( .A(n10146), .ZN(n10145) );
  NAND2_X1 U8139 ( .A1(n6527), .A2(n10145), .ZN(n6395) );
  NOR2_X1 U8140 ( .A1(n6387), .A2(n6928), .ZN(n7298) );
  NAND2_X1 U8141 ( .A1(n10145), .A2(n7298), .ZN(n7628) );
  NAND2_X1 U8142 ( .A1(n6387), .A2(n10200), .ZN(n8899) );
  OAI22_X1 U8143 ( .A1(n10145), .A2(n6390), .B1(n6389), .B2(n8977), .ZN(n6391)
         );
  AOI21_X1 U8144 ( .B1(n6536), .B2(n10138), .A(n6391), .ZN(n6392) );
  OAI21_X1 U8145 ( .B1(n6525), .B2(n7628), .A(n6392), .ZN(n6393) );
  INV_X1 U8146 ( .A(n6393), .ZN(n6394) );
  NAND2_X1 U8147 ( .A1(n6395), .A2(n6394), .ZN(P2_U3204) );
  XNOR2_X1 U8148 ( .A(n8592), .B(n8755), .ZN(n6396) );
  AND2_X1 U8149 ( .A1(n6762), .A2(n6396), .ZN(n6397) );
  NAND2_X1 U8150 ( .A1(n6398), .A2(n6397), .ZN(n6400) );
  OAI21_X1 U8151 ( .B1(n6404), .B2(n6821), .A(n8594), .ZN(n7205) );
  AOI22_X1 U8152 ( .A1(n7206), .A2(n7205), .B1(n4928), .B2(n6401), .ZN(n6869)
         );
  XNOR2_X1 U8153 ( .A(n6404), .B(n6406), .ZN(n6407) );
  XNOR2_X1 U8154 ( .A(n6404), .B(n10162), .ZN(n6408) );
  XNOR2_X1 U8155 ( .A(n6408), .B(n7594), .ZN(n7187) );
  XNOR2_X1 U8156 ( .A(n6404), .B(n10166), .ZN(n6410) );
  XNOR2_X1 U8157 ( .A(n6410), .B(n7192), .ZN(n7227) );
  INV_X1 U8158 ( .A(n6410), .ZN(n6411) );
  XNOR2_X1 U8159 ( .A(n6404), .B(n7662), .ZN(n6412) );
  XNOR2_X1 U8160 ( .A(n6412), .B(n7595), .ZN(n7272) );
  NAND2_X1 U8161 ( .A1(n7273), .A2(n7272), .ZN(n7271) );
  INV_X1 U8162 ( .A(n6412), .ZN(n6413) );
  XNOR2_X1 U8163 ( .A(n6404), .B(n10178), .ZN(n6414) );
  XNOR2_X1 U8164 ( .A(n6414), .B(n7634), .ZN(n7506) );
  XNOR2_X1 U8165 ( .A(n10182), .B(n6404), .ZN(n6415) );
  XNOR2_X1 U8166 ( .A(n6415), .B(n8780), .ZN(n7629) );
  XNOR2_X1 U8167 ( .A(n6404), .B(n10187), .ZN(n6416) );
  XNOR2_X1 U8168 ( .A(n6416), .B(n8779), .ZN(n7911) );
  OR2_X2 U8169 ( .A1(n7910), .A2(n7911), .ZN(n7838) );
  XNOR2_X1 U8170 ( .A(n6404), .B(n7711), .ZN(n7840) );
  INV_X1 U8171 ( .A(n6416), .ZN(n6417) );
  INV_X1 U8172 ( .A(n8779), .ZN(n7637) );
  NOR2_X1 U8173 ( .A1(n6417), .A2(n7637), .ZN(n7839) );
  AOI21_X1 U8174 ( .B1(n7840), .B2(n8778), .A(n7839), .ZN(n6419) );
  INV_X1 U8175 ( .A(n7840), .ZN(n6418) );
  XNOR2_X1 U8176 ( .A(n8575), .B(n6405), .ZN(n7894) );
  NAND2_X1 U8177 ( .A1(n7895), .A2(n7894), .ZN(n7893) );
  INV_X1 U8178 ( .A(n7894), .ZN(n6420) );
  NAND2_X1 U8179 ( .A1(n6420), .A2(n8777), .ZN(n6421) );
  XNOR2_X1 U8180 ( .A(n8663), .B(n6404), .ZN(n6422) );
  XNOR2_X1 U8181 ( .A(n6422), .B(n8776), .ZN(n7957) );
  INV_X1 U8182 ( .A(n6422), .ZN(n6423) );
  NAND2_X1 U8183 ( .A1(n6423), .A2(n8776), .ZN(n6424) );
  XNOR2_X1 U8184 ( .A(n8479), .B(n6404), .ZN(n8472) );
  NAND2_X1 U8185 ( .A1(n8472), .A2(n8670), .ZN(n6425) );
  INV_X1 U8186 ( .A(n8472), .ZN(n6426) );
  NAND2_X1 U8187 ( .A1(n6426), .A2(n8775), .ZN(n6427) );
  NAND2_X1 U8188 ( .A1(n6428), .A2(n6427), .ZN(n8364) );
  INV_X1 U8189 ( .A(n8364), .ZN(n6431) );
  XNOR2_X1 U8190 ( .A(n6429), .B(n6404), .ZN(n6432) );
  XNOR2_X1 U8191 ( .A(n6432), .B(n9019), .ZN(n8365) );
  INV_X1 U8192 ( .A(n8365), .ZN(n6430) );
  INV_X1 U8193 ( .A(n6432), .ZN(n6434) );
  NAND2_X1 U8194 ( .A1(n6434), .A2(n6433), .ZN(n6435) );
  XNOR2_X1 U8195 ( .A(n8560), .B(n6404), .ZN(n6437) );
  XNOR2_X1 U8196 ( .A(n6437), .B(n9009), .ZN(n8519) );
  XNOR2_X1 U8197 ( .A(n9154), .B(n6404), .ZN(n6436) );
  NAND2_X1 U8198 ( .A1(n6436), .A2(n8774), .ZN(n8437) );
  OAI21_X1 U8199 ( .B1(n6436), .B2(n8774), .A(n8437), .ZN(n8427) );
  AND2_X1 U8200 ( .A1(n6437), .A2(n9009), .ZN(n8426) );
  NOR2_X1 U8201 ( .A1(n8427), .A2(n8426), .ZN(n6438) );
  NAND2_X1 U8202 ( .A1(n8521), .A2(n6438), .ZN(n8425) );
  XNOR2_X1 U8203 ( .A(n9148), .B(n6404), .ZN(n6439) );
  NAND2_X1 U8204 ( .A1(n6439), .A2(n8431), .ZN(n8492) );
  INV_X1 U8205 ( .A(n6439), .ZN(n6440) );
  NAND2_X1 U8206 ( .A1(n6440), .A2(n9008), .ZN(n6441) );
  XNOR2_X1 U8207 ( .A(n9126), .B(n6404), .ZN(n6442) );
  NAND2_X1 U8208 ( .A1(n6442), .A2(n6443), .ZN(n6455) );
  INV_X1 U8209 ( .A(n6442), .ZN(n6444) );
  INV_X1 U8210 ( .A(n6443), .ZN(n8962) );
  NAND2_X1 U8211 ( .A1(n6444), .A2(n8962), .ZN(n6445) );
  NAND2_X1 U8212 ( .A1(n6446), .A2(n8975), .ZN(n8399) );
  INV_X1 U8213 ( .A(n8975), .ZN(n8951) );
  XNOR2_X1 U8214 ( .A(n8394), .B(n6405), .ZN(n6448) );
  NAND2_X1 U8215 ( .A1(n6448), .A2(n8498), .ZN(n8457) );
  INV_X1 U8216 ( .A(n6448), .ZN(n6449) );
  NAND2_X1 U8217 ( .A1(n6449), .A2(n8991), .ZN(n6450) );
  AND2_X1 U8218 ( .A1(n8457), .A2(n6450), .ZN(n8388) );
  INV_X1 U8219 ( .A(n6460), .ZN(n6454) );
  XNOR2_X1 U8220 ( .A(n9142), .B(n6404), .ZN(n6457) );
  NAND2_X1 U8221 ( .A1(n6457), .A2(n8973), .ZN(n8386) );
  AND2_X1 U8222 ( .A1(n8386), .A2(n6452), .ZN(n6453) );
  INV_X1 U8223 ( .A(n6455), .ZN(n8482) );
  INV_X1 U8224 ( .A(n6456), .ZN(n6463) );
  INV_X1 U8225 ( .A(n6457), .ZN(n6458) );
  NAND2_X1 U8226 ( .A1(n6458), .A2(n9000), .ZN(n6459) );
  AND2_X1 U8227 ( .A1(n8386), .A2(n6459), .ZN(n8493) );
  AND2_X1 U8228 ( .A1(n8493), .A2(n6460), .ZN(n6461) );
  AND2_X1 U8229 ( .A1(n6461), .A2(n8400), .ZN(n6462) );
  XNOR2_X1 U8230 ( .A(n8938), .B(n6405), .ZN(n6464) );
  XNOR2_X1 U8231 ( .A(n6464), .B(n8921), .ZN(n8481) );
  INV_X1 U8232 ( .A(n6464), .ZN(n6465) );
  NAND2_X1 U8233 ( .A1(n6465), .A2(n8921), .ZN(n6466) );
  NAND2_X1 U8234 ( .A1(n8484), .A2(n6466), .ZN(n6471) );
  XNOR2_X1 U8235 ( .A(n8926), .B(n6404), .ZN(n6470) );
  AND2_X1 U8236 ( .A1(n8481), .A2(n6470), .ZN(n6468) );
  INV_X1 U8237 ( .A(n6470), .ZN(n6467) );
  INV_X1 U8238 ( .A(n8488), .ZN(n8932) );
  NAND2_X1 U8239 ( .A1(n8376), .A2(n6472), .ZN(n6476) );
  XNOR2_X1 U8240 ( .A(n9113), .B(n6404), .ZN(n6473) );
  NAND2_X1 U8241 ( .A1(n6473), .A2(n8922), .ZN(n8413) );
  INV_X1 U8242 ( .A(n6473), .ZN(n6474) );
  NAND2_X1 U8243 ( .A1(n6474), .A2(n8894), .ZN(n6475) );
  NAND2_X1 U8244 ( .A1(n6476), .A2(n8446), .ZN(n8412) );
  NAND2_X1 U8245 ( .A1(n8412), .A2(n8413), .ZN(n6477) );
  XNOR2_X1 U8246 ( .A(n9107), .B(n6405), .ZN(n6478) );
  XNOR2_X1 U8247 ( .A(n6478), .B(n8773), .ZN(n8414) );
  NAND2_X1 U8248 ( .A1(n6477), .A2(n8414), .ZN(n8416) );
  INV_X1 U8249 ( .A(n6478), .ZN(n6479) );
  NAND2_X1 U8250 ( .A1(n6479), .A2(n8773), .ZN(n6480) );
  NAND2_X1 U8251 ( .A1(n8416), .A2(n6480), .ZN(n8504) );
  NAND2_X1 U8252 ( .A1(n8504), .A2(n8420), .ZN(n8347) );
  XNOR2_X1 U8253 ( .A(n9095), .B(n6404), .ZN(n6495) );
  NOR2_X1 U8254 ( .A1(n6495), .A2(n8509), .ZN(n6492) );
  AOI21_X1 U8255 ( .B1(n8509), .B2(n6495), .A(n6492), .ZN(n8348) );
  XNOR2_X1 U8256 ( .A(n9101), .B(n6404), .ZN(n8505) );
  XNOR2_X1 U8257 ( .A(n6404), .B(n8591), .ZN(n6481) );
  XNOR2_X1 U8258 ( .A(n9089), .B(n6481), .ZN(n6497) );
  INV_X1 U8259 ( .A(n6486), .ZN(n6482) );
  NOR2_X1 U8260 ( .A1(n6541), .A2(n6482), .ZN(n6501) );
  NAND2_X1 U8261 ( .A1(n6501), .A2(n6686), .ZN(n6530) );
  NAND3_X1 U8262 ( .A1(n6928), .A2(n8767), .A3(n6483), .ZN(n6484) );
  OR2_X1 U8263 ( .A1(n4353), .A2(n6484), .ZN(n6528) );
  NOR2_X1 U8264 ( .A1(n10200), .A2(n8747), .ZN(n6485) );
  NAND2_X1 U8265 ( .A1(n6528), .A2(n6485), .ZN(n6499) );
  OR2_X1 U8266 ( .A1(n6530), .A2(n6499), .ZN(n6489) );
  NAND3_X1 U8267 ( .A1(n6487), .A2(n6639), .A3(n6486), .ZN(n6508) );
  INV_X1 U8268 ( .A(n6686), .ZN(n6638) );
  INV_X1 U8269 ( .A(n6528), .ZN(n6504) );
  NAND2_X1 U8270 ( .A1(n6532), .A2(n6504), .ZN(n6488) );
  AND2_X1 U8271 ( .A1(n6497), .A2(n8507), .ZN(n6490) );
  NAND2_X1 U8272 ( .A1(n8354), .A2(n6490), .ZN(n6524) );
  NAND2_X1 U8273 ( .A1(n8346), .A2(n6491), .ZN(n6522) );
  INV_X1 U8274 ( .A(n6497), .ZN(n6494) );
  INV_X1 U8275 ( .A(n6492), .ZN(n6493) );
  INV_X1 U8276 ( .A(n6495), .ZN(n6496) );
  NAND4_X1 U8277 ( .A1(n6497), .A2(n6496), .A3(n8883), .A4(n8507), .ZN(n6520)
         );
  OR2_X1 U8278 ( .A1(n6530), .A2(n10186), .ZN(n6498) );
  NAND2_X1 U8279 ( .A1(n6499), .A2(n8899), .ZN(n6531) );
  INV_X1 U8280 ( .A(n6531), .ZN(n6500) );
  OR2_X1 U8281 ( .A1(n6501), .A2(n6500), .ZN(n6506) );
  NAND3_X1 U8282 ( .A1(n6566), .A2(n6565), .A3(n6502), .ZN(n6503) );
  AOI21_X1 U8283 ( .B1(n6508), .B2(n6504), .A(n6503), .ZN(n6505) );
  NAND2_X1 U8284 ( .A1(n6506), .A2(n6505), .ZN(n6510) );
  INV_X1 U8285 ( .A(n7367), .ZN(n6507) );
  AND2_X1 U8286 ( .A1(n6686), .A2(n6507), .ZN(n8765) );
  AND2_X1 U8287 ( .A1(n6508), .A2(n8765), .ZN(n6509) );
  AOI21_X2 U8288 ( .B1(n6510), .B2(P2_STATE_REG_SCAN_IN), .A(n6509), .ZN(n8524) );
  NOR2_X1 U8289 ( .A1(n8524), .A2(n8866), .ZN(n6518) );
  NOR2_X1 U8290 ( .A1(n7367), .A2(n6511), .ZN(n6512) );
  NAND2_X1 U8291 ( .A1(n6532), .A2(n6512), .ZN(n8523) );
  OR2_X1 U8292 ( .A1(n7367), .A2(n6513), .ZN(n6514) );
  AOI22_X1 U8293 ( .A1(n8527), .A2(n8883), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n6516) );
  OAI21_X1 U8294 ( .B1(n8772), .B2(n8523), .A(n6516), .ZN(n6517) );
  AOI211_X1 U8295 ( .C1(n9089), .C2(n8478), .A(n6518), .B(n6517), .ZN(n6519)
         );
  NAND2_X1 U8296 ( .A1(n6524), .A2(n6523), .ZN(P2_U3160) );
  NOR2_X1 U8297 ( .A1(n6525), .A2(n10192), .ZN(n6526) );
  AND2_X1 U8298 ( .A1(n7367), .A2(n6528), .ZN(n6529) );
  NAND2_X1 U8299 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  INV_X1 U8300 ( .A(n6536), .ZN(n6545) );
  NAND2_X1 U8301 ( .A1(n10205), .A2(n10200), .ZN(n9118) );
  OAI21_X1 U8302 ( .B1(n6548), .B2(n10207), .A(n6538), .ZN(P2_U3456) );
  NOR2_X1 U8303 ( .A1(n6540), .A2(n6539), .ZN(n6542) );
  NAND2_X1 U8304 ( .A1(n10225), .A2(n10200), .ZN(n9048) );
  OAI21_X1 U8305 ( .B1(n6548), .B2(n10222), .A(n6547), .ZN(P2_U3488) );
  OAI21_X1 U8306 ( .B1(n9269), .B2(n6550), .A(n6549), .ZN(n6551) );
  INV_X1 U8307 ( .A(n6551), .ZN(n6552) );
  OAI21_X1 U8308 ( .B1(n6553), .B2(n6552), .A(n9274), .ZN(n6559) );
  NOR2_X1 U8309 ( .A1(n6554), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6555) );
  AOI21_X1 U8310 ( .B1(n9524), .B2(n9277), .A(n6555), .ZN(n6556) );
  OAI21_X1 U8311 ( .B1(n9260), .B2(n9488), .A(n6556), .ZN(n6557) );
  AOI21_X1 U8312 ( .B1(n6874), .B2(n9250), .A(n6557), .ZN(n6558) );
  INV_X1 U8313 ( .A(n9486), .ZN(n9742) );
  NAND3_X1 U8314 ( .A1(n6559), .A2(n6558), .A3(n4429), .ZN(P1_U3214) );
  INV_X1 U8315 ( .A(n6560), .ZN(n6561) );
  OR2_X2 U8316 ( .A1(n5036), .A2(n6561), .ZN(n9301) );
  NAND2_X1 U8317 ( .A1(n6566), .A2(n4354), .ZN(n6562) );
  NAND2_X1 U8318 ( .A1(n6562), .A2(n6565), .ZN(n7356) );
  NAND2_X1 U8319 ( .A1(n7356), .A2(n6563), .ZN(n6564) );
  NAND2_X1 U8320 ( .A1(n6564), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8321 ( .A(n6565), .ZN(n7318) );
  NAND2_X1 U8322 ( .A1(n6568), .A2(n6567), .ZN(n6570) );
  XNOR2_X1 U8323 ( .A(n6570), .B(n6569), .ZN(n6571) );
  NOR2_X1 U8324 ( .A1(n6571), .A2(n9267), .ZN(n6575) );
  NOR2_X1 U8325 ( .A1(n9260), .A2(n6982), .ZN(n6574) );
  NAND2_X1 U8326 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9344) );
  OAI21_X1 U8327 ( .B1(n9279), .B2(n6882), .A(n9344), .ZN(n6573) );
  OAI22_X1 U8328 ( .A1(n9252), .A2(n6785), .B1(n6981), .B2(n9285), .ZN(n6572)
         );
  OR4_X1 U8329 ( .A1(n6575), .A2(n6574), .A3(n6573), .A4(n6572), .ZN(P1_U3227)
         );
  INV_X2 U8330 ( .A(n7850), .ZN(n9175) );
  INV_X2 U8331 ( .A(n9169), .ZN(n9172) );
  OAI222_X1 U8332 ( .A1(n7483), .A2(P2_U3151), .B1(n9175), .B2(n6580), .C1(
        n4652), .C2(n9172), .ZN(P2_U3294) );
  OAI222_X1 U8333 ( .A1(n7487), .A2(P2_U3151), .B1(n9175), .B2(n6581), .C1(
        n6576), .C2(n9172), .ZN(P2_U3293) );
  OAI222_X1 U8334 ( .A1(n7348), .A2(P2_U3151), .B1(n9175), .B2(n6578), .C1(
        n6577), .C2(n9172), .ZN(P2_U3292) );
  OAI222_X1 U8335 ( .A1(n9775), .A2(n6579), .B1(n8017), .B2(n6578), .C1(
        P1_U3086), .C2(n6672), .ZN(P1_U3352) );
  OAI222_X1 U8336 ( .A1(n9775), .A2(n4649), .B1(n8017), .B2(n6580), .C1(
        P1_U3086), .C2(n6668), .ZN(P1_U3354) );
  OAI222_X1 U8337 ( .A1(n9775), .A2(n6582), .B1(n8017), .B2(n6581), .C1(
        P1_U3086), .C2(n9316), .ZN(P1_U3353) );
  OAI222_X1 U8338 ( .A1(n7413), .A2(P2_U3151), .B1(n9175), .B2(n6583), .C1(
        n9172), .C2(n6020), .ZN(P2_U3291) );
  OAI222_X1 U8339 ( .A1(n9775), .A2(n6584), .B1(P1_U3086), .B2(n6679), .C1(
        n8017), .C2(n6583), .ZN(P1_U3351) );
  OAI222_X1 U8340 ( .A1(n10015), .A2(P2_U3151), .B1(n9175), .B2(n6589), .C1(
        n6585), .C2(n9172), .ZN(P2_U3290) );
  OAI222_X1 U8341 ( .A1(n7441), .A2(P2_U3151), .B1(n9175), .B2(n6587), .C1(
        n6586), .C2(n9172), .ZN(P2_U3289) );
  OAI222_X1 U8342 ( .A1(n9775), .A2(n6588), .B1(n8017), .B2(n6587), .C1(
        P1_U3086), .C2(n9368), .ZN(P1_U3349) );
  OAI222_X1 U8343 ( .A1(n9370), .A2(P1_U3086), .B1(n8017), .B2(n6589), .C1(
        n9775), .C2(n5156), .ZN(P1_U3350) );
  OAI222_X1 U8344 ( .A1(n7743), .A2(P2_U3151), .B1(n9175), .B2(n6591), .C1(
        n6590), .C2(n9172), .ZN(P2_U3288) );
  OAI222_X1 U8345 ( .A1(n9405), .A2(P1_U3086), .B1(n8017), .B2(n6591), .C1(
        n9775), .C2(n5210), .ZN(P1_U3348) );
  INV_X1 U8346 ( .A(n9435), .ZN(n9830) );
  OAI222_X1 U8347 ( .A1(n8017), .A2(n6079), .B1(n9830), .B2(P1_U3086), .C1(
        n6593), .C2(n9775), .ZN(P1_U3346) );
  INV_X1 U8348 ( .A(n6594), .ZN(n6601) );
  INV_X1 U8349 ( .A(n9775), .ZN(n6740) );
  AOI22_X1 U8350 ( .A1(n9814), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n6740), .ZN(n6595) );
  OAI21_X1 U8351 ( .B1(n6601), .B2(n8017), .A(n6595), .ZN(P1_U3345) );
  AOI22_X1 U8352 ( .A1(n9430), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n6740), .ZN(n6596) );
  OAI21_X1 U8353 ( .B1(n6605), .B2(n8017), .A(n6596), .ZN(P1_U3347) );
  INV_X1 U8354 ( .A(n6597), .ZN(n6607) );
  AOI22_X1 U8355 ( .A1(n9836), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n6740), .ZN(n6598) );
  OAI21_X1 U8356 ( .B1(n6607), .B2(n8017), .A(n6598), .ZN(P1_U3344) );
  INV_X1 U8357 ( .A(n7796), .ZN(n7749) );
  OAI222_X1 U8358 ( .A1(P2_U3151), .A2(n7749), .B1(n9175), .B2(n6079), .C1(
        n6599), .C2(n9172), .ZN(P2_U3286) );
  INV_X1 U8359 ( .A(n7875), .ZN(n7880) );
  OAI222_X1 U8360 ( .A1(P2_U3151), .A2(n7880), .B1(n9175), .B2(n6601), .C1(
        n6600), .C2(n9172), .ZN(P2_U3285) );
  NAND2_X1 U8361 ( .A1(n9957), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6602) );
  OAI21_X1 U8362 ( .B1(n9957), .B2(n6603), .A(n6602), .ZN(P1_U3439) );
  OAI222_X1 U8363 ( .A1(n10026), .A2(P2_U3151), .B1(n9175), .B2(n6605), .C1(
        n6604), .C2(n9172), .ZN(P2_U3287) );
  INV_X1 U8364 ( .A(n7975), .ZN(n7982) );
  INV_X1 U8365 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6606) );
  OAI222_X1 U8366 ( .A1(n7982), .A2(P2_U3151), .B1(n9175), .B2(n6607), .C1(
        n6606), .C2(n9172), .ZN(P2_U3284) );
  AOI21_X1 U8367 ( .B1(n6665), .B2(n5054), .A(n7856), .ZN(n6661) );
  OAI21_X1 U8368 ( .B1(n6665), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6661), .ZN(
        n6608) );
  XOR2_X1 U8369 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6608), .Z(n6618) );
  NAND2_X1 U8370 ( .A1(n8213), .A2(n6609), .ZN(n6610) );
  NAND2_X1 U8371 ( .A1(n6611), .A2(n6610), .ZN(n6615) );
  INV_X1 U8372 ( .A(n8329), .ZN(n6612) );
  NOR2_X1 U8373 ( .A1(n6613), .A2(n6612), .ZN(n6614) );
  OR2_X1 U8374 ( .A1(n6615), .A2(n6614), .ZN(n6678) );
  INV_X1 U8375 ( .A(n6614), .ZN(n6616) );
  NAND2_X1 U8376 ( .A1(n6616), .A2(n6615), .ZN(n9956) );
  INV_X1 U8377 ( .A(n9956), .ZN(n9456) );
  AOI22_X1 U8378 ( .A1(n9456), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6617) );
  OAI21_X1 U8379 ( .B1(n6618), .B2(n6678), .A(n6617), .ZN(P1_U3243) );
  INV_X1 U8380 ( .A(n6619), .ZN(n6622) );
  AOI22_X1 U8381 ( .A1(n9852), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n6740), .ZN(n6620) );
  OAI21_X1 U8382 ( .B1(n6622), .B2(n8017), .A(n6620), .ZN(P1_U3343) );
  INV_X1 U8383 ( .A(n7988), .ZN(n8827) );
  INV_X1 U8384 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6621) );
  OAI222_X1 U8385 ( .A1(P2_U3151), .A2(n8827), .B1(n9175), .B2(n6622), .C1(
        n6621), .C2(n9172), .ZN(P2_U3283) );
  NOR2_X1 U8386 ( .A1(n9456), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8387 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U8388 ( .A1(n7831), .A2(P1_U3973), .ZN(n6623) );
  OAI21_X1 U8389 ( .B1(n6655), .B2(P1_U3973), .A(n6623), .ZN(P1_U3570) );
  INV_X1 U8390 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8391 ( .A1(n7943), .A2(P1_U3973), .ZN(n6624) );
  OAI21_X1 U8392 ( .B1(n6633), .B2(P1_U3973), .A(n6624), .ZN(P1_U3568) );
  NAND2_X1 U8393 ( .A1(n6625), .A2(P1_U3973), .ZN(n6626) );
  OAI21_X1 U8394 ( .B1(P1_U3973), .B2(n6020), .A(n6626), .ZN(P1_U3558) );
  INV_X1 U8395 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6628) );
  INV_X1 U8396 ( .A(n6627), .ZN(n6630) );
  INV_X1 U8397 ( .A(n9437), .ZN(n9878) );
  OAI222_X1 U8398 ( .A1(n9775), .A2(n6628), .B1(n8017), .B2(n6630), .C1(
        P1_U3086), .C2(n9878), .ZN(P1_U3342) );
  INV_X1 U8399 ( .A(n10042), .ZN(n8830) );
  INV_X1 U8400 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6629) );
  OAI222_X1 U8401 ( .A1(n8830), .A2(P2_U3151), .B1(n9175), .B2(n6630), .C1(
        n6629), .C2(n9172), .ZN(P2_U3282) );
  INV_X1 U8402 ( .A(n6631), .ZN(n6634) );
  AOI22_X1 U8403 ( .A1(n9883), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n6740), .ZN(n6632) );
  OAI21_X1 U8404 ( .B1(n6634), .B2(n8017), .A(n6632), .ZN(P1_U3341) );
  INV_X1 U8405 ( .A(n10058), .ZN(n8826) );
  OAI222_X1 U8406 ( .A1(n8826), .A2(P2_U3151), .B1(n9175), .B2(n6634), .C1(
        n9172), .C2(n6633), .ZN(P2_U3281) );
  INV_X1 U8407 ( .A(n6635), .ZN(n6641) );
  INV_X1 U8408 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6636) );
  OAI222_X1 U8409 ( .A1(n8017), .A2(n6641), .B1(n9440), .B2(P1_U3086), .C1(
        n6636), .C2(n9775), .ZN(P1_U3340) );
  NAND2_X1 U8410 ( .A1(n6638), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6637) );
  OAI21_X1 U8411 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(P2_U3377) );
  INV_X1 U8412 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6640) );
  OAI222_X1 U8413 ( .A1(P2_U3151), .A2(n4730), .B1(n9175), .B2(n6641), .C1(
        n6640), .C2(n9172), .ZN(P2_U3280) );
  INV_X1 U8414 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6644) );
  AND2_X1 U8415 ( .A1(n9302), .A2(n7252), .ZN(n8262) );
  OR2_X1 U8416 ( .A1(n8262), .A2(n6710), .ZN(n8217) );
  OAI21_X1 U8417 ( .B1(n9978), .B2(n9640), .A(n8217), .ZN(n6642) );
  NAND2_X1 U8418 ( .A1(n9300), .A2(n9644), .ZN(n7250) );
  OAI211_X1 U8419 ( .C1(n7248), .C2(n7252), .A(n6642), .B(n7250), .ZN(n9730)
         );
  NAND2_X1 U8420 ( .A1(n9730), .A2(n9981), .ZN(n6643) );
  OAI21_X1 U8421 ( .B1(n9981), .B2(n6644), .A(n6643), .ZN(P1_U3453) );
  NAND2_X1 U8422 ( .A1(n9583), .A2(P1_U3973), .ZN(n6645) );
  OAI21_X1 U8423 ( .B1(P1_U3973), .B2(n7320), .A(n6645), .ZN(P1_U3577) );
  INV_X1 U8424 ( .A(n6692), .ZN(n6647) );
  AOI21_X1 U8425 ( .B1(n6648), .B2(n6646), .A(n6647), .ZN(n6652) );
  AOI22_X1 U8426 ( .A1(n5887), .A2(n9265), .B1(n9277), .B2(n9302), .ZN(n6651)
         );
  NOR2_X1 U8427 ( .A1(n6649), .A2(n8325), .ZN(n6697) );
  INV_X1 U8428 ( .A(n6697), .ZN(n6688) );
  AOI22_X1 U8429 ( .A1(n6688), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9299), .B2(
        n9250), .ZN(n6650) );
  OAI211_X1 U8430 ( .C1(n6652), .C2(n9267), .A(n6651), .B(n6650), .ZN(P1_U3222) );
  INV_X1 U8431 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6654) );
  INV_X1 U8432 ( .A(n6653), .ZN(n6656) );
  INV_X1 U8433 ( .A(n9443), .ZN(n9915) );
  OAI222_X1 U8434 ( .A1(n9775), .A2(n6654), .B1(n8017), .B2(n6656), .C1(
        P1_U3086), .C2(n9915), .ZN(P1_U3339) );
  INV_X1 U8435 ( .A(n10090), .ZN(n8824) );
  OAI222_X1 U8436 ( .A1(n8824), .A2(P2_U3151), .B1(n9175), .B2(n6656), .C1(
        n9172), .C2(n6655), .ZN(P2_U3279) );
  XNOR2_X1 U8437 ( .A(n6657), .B(n6658), .ZN(n6690) );
  AND2_X1 U8438 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9312) );
  MUX2_X1 U8439 ( .A(n6690), .B(n9312), .S(n6665), .Z(n6659) );
  NAND2_X1 U8440 ( .A1(n6659), .A2(n6677), .ZN(n6660) );
  OAI211_X1 U8441 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6661), .A(n6660), .B(
        P1_U3973), .ZN(n9330) );
  INV_X1 U8442 ( .A(n9330), .ZN(n6685) );
  MUX2_X1 U8443 ( .A(n5071), .B(P1_REG1_REG_2__SCAN_IN), .S(n9316), .Z(n9326)
         );
  MUX2_X1 U8444 ( .A(n5026), .B(P1_REG1_REG_1__SCAN_IN), .S(n6668), .Z(n9309)
         );
  AND2_X1 U8445 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9308) );
  NAND2_X1 U8446 ( .A1(n9309), .A2(n9308), .ZN(n9307) );
  INV_X1 U8447 ( .A(n6668), .ZN(n9306) );
  NAND2_X1 U8448 ( .A1(n9306), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U8449 ( .A1(n9307), .A2(n6662), .ZN(n9325) );
  NAND2_X1 U8450 ( .A1(n9326), .A2(n9325), .ZN(n9324) );
  INV_X1 U8451 ( .A(n9316), .ZN(n6670) );
  NAND2_X1 U8452 ( .A1(n6670), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U8453 ( .A1(n9324), .A2(n6663), .ZN(n9339) );
  MUX2_X1 U8454 ( .A(n5096), .B(P1_REG1_REG_3__SCAN_IN), .S(n6672), .Z(n9340)
         );
  NAND2_X1 U8455 ( .A1(n9339), .A2(n9340), .ZN(n9338) );
  INV_X1 U8456 ( .A(n6672), .ZN(n9334) );
  NAND2_X1 U8457 ( .A1(n9334), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U8458 ( .A1(n9338), .A2(n6664), .ZN(n6667) );
  XNOR2_X1 U8459 ( .A(n6679), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n6666) );
  OR2_X1 U8460 ( .A1(n6678), .A2(n6665), .ZN(n9899) );
  INV_X1 U8461 ( .A(n9899), .ZN(n9946) );
  NAND2_X1 U8462 ( .A1(n6667), .A2(n6666), .ZN(n9354) );
  OAI211_X1 U8463 ( .C1(n6667), .C2(n6666), .A(n9946), .B(n9354), .ZN(n6683)
         );
  XNOR2_X1 U8464 ( .A(n6679), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6676) );
  MUX2_X1 U8465 ( .A(n5070), .B(P1_REG2_REG_2__SCAN_IN), .S(n9316), .Z(n9323)
         );
  MUX2_X1 U8466 ( .A(n5031), .B(P1_REG2_REG_1__SCAN_IN), .S(n6668), .Z(n9311)
         );
  NAND2_X1 U8467 ( .A1(n9311), .A2(n9312), .ZN(n9310) );
  NAND2_X1 U8468 ( .A1(n9306), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8469 ( .A1(n9310), .A2(n6669), .ZN(n9322) );
  NAND2_X1 U8470 ( .A1(n9323), .A2(n9322), .ZN(n9321) );
  NAND2_X1 U8471 ( .A1(n6670), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8472 ( .A1(n9321), .A2(n6671), .ZN(n9336) );
  MUX2_X1 U8473 ( .A(n6835), .B(P1_REG2_REG_3__SCAN_IN), .S(n6672), .Z(n9337)
         );
  NAND2_X1 U8474 ( .A1(n9336), .A2(n9337), .ZN(n9335) );
  NAND2_X1 U8475 ( .A1(n9334), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8476 ( .A1(n9335), .A2(n6673), .ZN(n6675) );
  OR2_X1 U8477 ( .A1(n7856), .A2(n5904), .ZN(n6674) );
  OR2_X1 U8478 ( .A1(n6678), .A2(n6674), .ZN(n9916) );
  INV_X1 U8479 ( .A(n9916), .ZN(n9942) );
  NAND2_X1 U8480 ( .A1(n6675), .A2(n6676), .ZN(n9349) );
  OAI211_X1 U8481 ( .C1(n6676), .C2(n6675), .A(n9942), .B(n9349), .ZN(n6682)
         );
  AND2_X1 U8482 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6724) );
  AOI21_X1 U8483 ( .B1(n9456), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6724), .ZN(
        n6681) );
  OR2_X1 U8484 ( .A1(n6678), .A2(n6677), .ZN(n9952) );
  INV_X1 U8485 ( .A(n9952), .ZN(n9908) );
  INV_X1 U8486 ( .A(n6679), .ZN(n9352) );
  NAND2_X1 U8487 ( .A1(n9908), .A2(n9352), .ZN(n6680) );
  NAND4_X1 U8488 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6684)
         );
  OR2_X1 U8489 ( .A1(n6685), .A2(n6684), .ZN(P1_U3247) );
  NAND2_X1 U8490 ( .A1(n6686), .A2(n6363), .ZN(n6761) );
  AND2_X1 U8491 ( .A1(n6761), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8492 ( .A1(n6761), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8493 ( .A1(n6761), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8494 ( .A1(n6761), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8495 ( .A1(n6761), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8496 ( .A1(n6761), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8497 ( .A1(n6761), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8498 ( .A1(n6761), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8499 ( .A1(n6761), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8500 ( .A1(n6761), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8501 ( .A1(n6761), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  OAI22_X1 U8502 ( .A1(n9279), .A2(n5041), .B1(n9285), .B2(n7252), .ZN(n6687)
         );
  AOI21_X1 U8503 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6688), .A(n6687), .ZN(
        n6689) );
  OAI21_X1 U8504 ( .B1(n9267), .B2(n6690), .A(n6689), .ZN(P1_U3232) );
  INV_X1 U8505 ( .A(n6691), .ZN(n6694) );
  NAND3_X1 U8506 ( .A1(n6694), .A2(n6693), .A3(n6692), .ZN(n6696) );
  AOI21_X1 U8507 ( .B1(n6696), .B2(n6695), .A(n9267), .ZN(n6700) );
  OAI22_X1 U8508 ( .A1(n9252), .A2(n5041), .B1(n6735), .B2(n9285), .ZN(n6699)
         );
  OAI22_X1 U8509 ( .A1(n9279), .A2(n6910), .B1(n6697), .B2(n9317), .ZN(n6698)
         );
  OR3_X1 U8510 ( .A1(n6700), .A2(n6699), .A3(n6698), .ZN(P1_U3237) );
  OAI21_X1 U8511 ( .B1(n6702), .B2(n8218), .A(n6701), .ZN(n6811) );
  AOI211_X1 U8512 ( .C1(n6818), .C2(n6707), .A(n9682), .B(n6747), .ZN(n6807)
         );
  XNOR2_X1 U8513 ( .A(n8074), .B(n8218), .ZN(n6703) );
  OAI222_X1 U8514 ( .A1(n9549), .A2(n5041), .B1(n9551), .B2(n6910), .C1(n6703), 
        .C2(n9546), .ZN(n6809) );
  AOI211_X1 U8515 ( .C1(n9978), .C2(n6811), .A(n6807), .B(n6809), .ZN(n6738)
         );
  AOI22_X1 U8516 ( .A1(n5919), .A2(n6818), .B1(n9986), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6704) );
  OAI21_X1 U8517 ( .B1(n6738), .B2(n9986), .A(n6704), .ZN(P1_U3524) );
  OAI21_X1 U8518 ( .B1(n6711), .B2(n6706), .A(n6705), .ZN(n6860) );
  INV_X1 U8519 ( .A(n6707), .ZN(n6708) );
  AOI211_X1 U8520 ( .C1(n6709), .C2(n5887), .A(n9682), .B(n6708), .ZN(n6864)
         );
  INV_X1 U8521 ( .A(n9302), .ZN(n6713) );
  XNOR2_X1 U8522 ( .A(n6711), .B(n6710), .ZN(n6712) );
  OAI222_X1 U8523 ( .A1(n9551), .A2(n6750), .B1(n9549), .B2(n6713), .C1(n6712), 
        .C2(n9546), .ZN(n6861) );
  AOI211_X1 U8524 ( .C1(n9978), .C2(n6860), .A(n6864), .B(n6861), .ZN(n6744)
         );
  AOI22_X1 U8525 ( .A1(n5919), .A2(n5887), .B1(n9986), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6714) );
  OAI21_X1 U8526 ( .B1(n6744), .B2(n9986), .A(n6714), .ZN(P1_U3523) );
  INV_X1 U8527 ( .A(n6715), .ZN(n6718) );
  AOI22_X1 U8528 ( .A1(n9926), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6740), .ZN(n6716) );
  OAI21_X1 U8529 ( .B1(n6718), .B2(n8017), .A(n6716), .ZN(P1_U3338) );
  INV_X1 U8530 ( .A(n10108), .ZN(n8836) );
  INV_X1 U8531 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6717) );
  OAI222_X1 U8532 ( .A1(P2_U3151), .A2(n8836), .B1(n9175), .B2(n6718), .C1(
        n6717), .C2(n9172), .ZN(P2_U3278) );
  AND2_X1 U8533 ( .A1(n6727), .A2(n6719), .ZN(n6722) );
  OAI211_X1 U8534 ( .C1(n6722), .C2(n6721), .A(n9274), .B(n6720), .ZN(n6726)
         );
  OAI22_X1 U8535 ( .A1(n6910), .A2(n9252), .B1(n9279), .B2(n6932), .ZN(n6723)
         );
  AOI211_X1 U8536 ( .C1(n6918), .C2(n9265), .A(n6724), .B(n6723), .ZN(n6725)
         );
  OAI211_X1 U8537 ( .C1(n9260), .C2(n6915), .A(n6726), .B(n6725), .ZN(P1_U3230) );
  OAI21_X1 U8538 ( .B1(n6729), .B2(n6728), .A(n6727), .ZN(n6730) );
  NAND2_X1 U8539 ( .A1(n6730), .A2(n9274), .ZN(n6734) );
  NAND2_X1 U8540 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9331) );
  INV_X1 U8541 ( .A(n9331), .ZN(n6732) );
  OAI22_X1 U8542 ( .A1(n6750), .A2(n9252), .B1(n9279), .B2(n6785), .ZN(n6731)
         );
  AOI211_X1 U8543 ( .C1(n6754), .C2(n9265), .A(n6732), .B(n6731), .ZN(n6733)
         );
  OAI211_X1 U8544 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9260), .A(n6734), .B(
        n6733), .ZN(P1_U3218) );
  OAI22_X1 U8545 ( .A1(n9770), .A2(n6735), .B1(n9981), .B2(n5072), .ZN(n6736)
         );
  INV_X1 U8546 ( .A(n6736), .ZN(n6737) );
  OAI21_X1 U8547 ( .B1(n6738), .B2(n9980), .A(n6737), .ZN(P1_U3459) );
  INV_X1 U8548 ( .A(n6739), .ZN(n6760) );
  AOI22_X1 U8549 ( .A1(n9940), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n6740), .ZN(n6741) );
  OAI21_X1 U8550 ( .B1(n6760), .B2(n8017), .A(n6741), .ZN(P1_U3337) );
  OAI22_X1 U8551 ( .A1(n9770), .A2(n5835), .B1(n9981), .B2(n5029), .ZN(n6742)
         );
  INV_X1 U8552 ( .A(n6742), .ZN(n6743) );
  OAI21_X1 U8553 ( .B1(n6744), .B2(n9980), .A(n6743), .ZN(P1_U3456) );
  OAI21_X1 U8554 ( .B1(n6746), .B2(n8219), .A(n6745), .ZN(n6833) );
  INV_X1 U8555 ( .A(n6747), .ZN(n6749) );
  INV_X1 U8556 ( .A(n6748), .ZN(n6914) );
  AOI211_X1 U8557 ( .C1(n6754), .C2(n6749), .A(n9682), .B(n6914), .ZN(n6839)
         );
  XNOR2_X1 U8558 ( .A(n8269), .B(n8219), .ZN(n6752) );
  OAI22_X1 U8559 ( .A1(n6750), .A2(n9549), .B1(n6785), .B2(n9551), .ZN(n6751)
         );
  AOI21_X1 U8560 ( .B1(n6752), .B2(n9640), .A(n6751), .ZN(n6836) );
  INV_X1 U8561 ( .A(n6836), .ZN(n6753) );
  AOI211_X1 U8562 ( .C1(n9978), .C2(n6833), .A(n6839), .B(n6753), .ZN(n6758)
         );
  AOI22_X1 U8563 ( .A1(n5919), .A2(n6754), .B1(n9986), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6755) );
  OAI21_X1 U8564 ( .B1(n6758), .B2(n9986), .A(n6755), .ZN(P1_U3525) );
  OAI22_X1 U8565 ( .A1(n9770), .A2(n6837), .B1(n9981), .B2(n5098), .ZN(n6756)
         );
  INV_X1 U8566 ( .A(n6756), .ZN(n6757) );
  OAI21_X1 U8567 ( .B1(n6758), .B2(n9980), .A(n6757), .ZN(P1_U3462) );
  INV_X1 U8568 ( .A(n9805), .ZN(n9803) );
  INV_X1 U8569 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6759) );
  OAI222_X1 U8570 ( .A1(P2_U3151), .A2(n9803), .B1(n9175), .B2(n6760), .C1(
        n6759), .C2(n9172), .ZN(P2_U3277) );
  INV_X1 U8571 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6765) );
  INV_X1 U8572 ( .A(n6762), .ZN(n6763) );
  AOI22_X1 U8573 ( .A1(n6761), .A2(n6765), .B1(n6764), .B2(n6763), .ZN(
        P2_U3376) );
  AND2_X1 U8574 ( .A1(n6761), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8575 ( .A1(n6761), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8576 ( .A1(n6761), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8577 ( .A1(n6761), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8578 ( .A1(n6761), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8579 ( .A1(n6761), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8580 ( .A1(n6761), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8581 ( .A1(n6761), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8582 ( .A1(n6761), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8583 ( .A1(n6761), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8584 ( .A1(n6761), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8585 ( .A1(n6761), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8586 ( .A1(n6761), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8587 ( .A1(n6761), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8588 ( .A1(n6761), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8589 ( .A1(n6761), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8590 ( .A1(n6761), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8591 ( .A1(n6761), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8592 ( .A1(n6761), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  OAI21_X1 U8593 ( .B1(n6768), .B2(n6766), .A(n6767), .ZN(n6774) );
  NOR2_X1 U8594 ( .A1(n9285), .A2(n9964), .ZN(n6773) );
  NAND2_X1 U8595 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9360) );
  INV_X1 U8596 ( .A(n9360), .ZN(n6769) );
  AOI21_X1 U8597 ( .B1(n9297), .B2(n9277), .A(n6769), .ZN(n6771) );
  NAND2_X1 U8598 ( .A1(n9295), .A2(n9250), .ZN(n6770) );
  OAI211_X1 U8599 ( .C1(n9260), .C2(n6940), .A(n6771), .B(n6770), .ZN(n6772)
         );
  AOI211_X1 U8600 ( .C1(n6774), .C2(n9274), .A(n6773), .B(n6772), .ZN(n6775)
         );
  INV_X1 U8601 ( .A(n6775), .ZN(P1_U3239) );
  INV_X1 U8602 ( .A(n6776), .ZN(n8333) );
  INV_X1 U8603 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6777) );
  OAI222_X1 U8604 ( .A1(P2_U3151), .A2(n4353), .B1(n9175), .B2(n8333), .C1(
        n6777), .C2(n9172), .ZN(P2_U3276) );
  INV_X1 U8605 ( .A(n6821), .ZN(n7366) );
  NAND2_X1 U8606 ( .A1(n8784), .A2(n7366), .ZN(n8593) );
  AND2_X1 U8607 ( .A1(n8594), .A2(n8593), .ZN(n8565) );
  NAND2_X1 U8608 ( .A1(n8524), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7209) );
  NAND2_X1 U8609 ( .A1(n7209), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6779) );
  INV_X1 U8610 ( .A(n8523), .ZN(n8468) );
  AOI22_X1 U8611 ( .A1(n8478), .A2(n6821), .B1(n8468), .B2(n8783), .ZN(n6778)
         );
  OAI211_X1 U8612 ( .C1(n8565), .C2(n8518), .A(n6779), .B(n6778), .ZN(P2_U3172) );
  NAND2_X1 U8613 ( .A1(n6912), .A2(n8220), .ZN(n6911) );
  NAND2_X1 U8614 ( .A1(n6911), .A2(n6780), .ZN(n6782) );
  OAI21_X1 U8615 ( .B1(n6782), .B2(n8225), .A(n6781), .ZN(n6979) );
  AOI211_X1 U8616 ( .C1(n6786), .C2(n6913), .A(n9682), .B(n6939), .ZN(n6985)
         );
  NAND2_X1 U8617 ( .A1(n6845), .A2(n8068), .ZN(n6783) );
  XNOR2_X1 U8618 ( .A(n6783), .B(n8225), .ZN(n6784) );
  OAI222_X1 U8619 ( .A1(n9551), .A2(n6882), .B1(n9549), .B2(n6785), .C1(n6784), 
        .C2(n9546), .ZN(n6980) );
  AOI211_X1 U8620 ( .C1(n9978), .C2(n6979), .A(n6985), .B(n6980), .ZN(n6790)
         );
  AOI22_X1 U8621 ( .A1(n5919), .A2(n6786), .B1(n9986), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n6787) );
  OAI21_X1 U8622 ( .B1(n6790), .B2(n9986), .A(n6787), .ZN(P1_U3527) );
  OAI22_X1 U8623 ( .A1(n9770), .A2(n6981), .B1(n9981), .B2(n5146), .ZN(n6788)
         );
  INV_X1 U8624 ( .A(n6788), .ZN(n6789) );
  OAI21_X1 U8625 ( .B1(n6790), .B2(n9980), .A(n6789), .ZN(P1_U3468) );
  NAND2_X1 U8626 ( .A1(n6827), .A2(n9780), .ZN(n6792) );
  OAI211_X1 U8627 ( .C1(n6793), .C2(n9775), .A(n6792), .B(n6791), .ZN(P1_U3335) );
  INV_X1 U8628 ( .A(n6794), .ZN(n6798) );
  OAI21_X1 U8629 ( .B1(n6798), .B2(n6796), .A(n6795), .ZN(n6797) );
  OAI211_X1 U8630 ( .C1(n6799), .C2(n6798), .A(n9274), .B(n6797), .ZN(n6804)
         );
  NAND2_X1 U8631 ( .A1(n9294), .A2(n9250), .ZN(n6800) );
  NAND2_X1 U8632 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9378) );
  OAI211_X1 U8633 ( .C1(n9252), .C2(n6882), .A(n6800), .B(n9378), .ZN(n6802)
         );
  NOR2_X1 U8634 ( .A1(n9260), .A2(n6885), .ZN(n6801) );
  AOI211_X1 U8635 ( .C1(n6902), .C2(n9265), .A(n6802), .B(n6801), .ZN(n6803)
         );
  NAND2_X1 U8636 ( .A1(n6804), .A2(n6803), .ZN(P1_U3213) );
  NAND2_X1 U8637 ( .A1(n6806), .A2(n6805), .ZN(n6834) );
  INV_X1 U8638 ( .A(n6807), .ZN(n6808) );
  OAI22_X1 U8639 ( .A1(n6808), .A2(n4485), .B1(n9630), .B2(n9317), .ZN(n6810)
         );
  AOI211_X1 U8640 ( .C1(n6834), .C2(n6811), .A(n6810), .B(n6809), .ZN(n6820)
         );
  INV_X1 U8641 ( .A(n6812), .ZN(n6813) );
  NAND3_X1 U8642 ( .A1(n6815), .A2(n6814), .A3(n6813), .ZN(n6816) );
  INV_X2 U8643 ( .A(n9633), .ZN(n9469) );
  INV_X1 U8644 ( .A(n9629), .ZN(n7293) );
  AOI22_X1 U8645 ( .A1(n7293), .A2(n6818), .B1(n9469), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n6819) );
  OAI21_X1 U8646 ( .B1(n6820), .B2(n9469), .A(n6819), .ZN(P1_U3291) );
  INV_X1 U8647 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8648 ( .A1(n7622), .A2(n10192), .ZN(n10198) );
  NOR2_X1 U8649 ( .A1(n10198), .A2(n10134), .ZN(n6823) );
  NAND2_X1 U8650 ( .A1(n6821), .A2(n10200), .ZN(n6822) );
  NAND2_X1 U8651 ( .A1(n8783), .A2(n10131), .ZN(n7369) );
  OAI211_X1 U8652 ( .C1(n8565), .C2(n6823), .A(n6822), .B(n7369), .ZN(n9079)
         );
  NAND2_X1 U8653 ( .A1(n10205), .A2(n9079), .ZN(n6824) );
  OAI21_X1 U8654 ( .B1(n10205), .B2(n6825), .A(n6824), .ZN(P2_U3390) );
  NAND2_X1 U8655 ( .A1(n9513), .A2(P1_U3973), .ZN(n6826) );
  OAI21_X1 U8656 ( .B1(P1_U3973), .B2(n6258), .A(n6826), .ZN(P1_U3581) );
  INV_X1 U8657 ( .A(n6827), .ZN(n6829) );
  OAI222_X1 U8658 ( .A1(n8755), .A2(P2_U3151), .B1(n9175), .B2(n6829), .C1(
        n6828), .C2(n9172), .ZN(P2_U3275) );
  NAND2_X1 U8659 ( .A1(P2_U3893), .A2(n7634), .ZN(n6830) );
  OAI21_X1 U8660 ( .B1(P2_U3893), .B2(n5210), .A(n6830), .ZN(P2_U3498) );
  NAND2_X1 U8661 ( .A1(P2_U3893), .A2(n8618), .ZN(n6831) );
  OAI21_X1 U8662 ( .B1(P2_U3893), .B2(n6584), .A(n6831), .ZN(P2_U3495) );
  NAND2_X1 U8663 ( .A1(P2_U3893), .A2(n10132), .ZN(n6832) );
  OAI21_X1 U8664 ( .B1(P2_U3893), .B2(n5156), .A(n6832), .ZN(P2_U3496) );
  INV_X1 U8665 ( .A(n6833), .ZN(n6842) );
  NAND2_X1 U8666 ( .A1(n7692), .A2(n6834), .ZN(n9650) );
  MUX2_X1 U8667 ( .A(n6836), .B(n6835), .S(n9469), .Z(n6841) );
  AND2_X2 U8668 ( .A1(n7692), .A2(n8317), .ZN(n9616) );
  OAI22_X1 U8669 ( .A1(n9629), .A2(n6837), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9630), .ZN(n6838) );
  AOI21_X1 U8670 ( .B1(n6839), .B2(n9616), .A(n6838), .ZN(n6840) );
  OAI211_X1 U8671 ( .C1(n6842), .C2(n9650), .A(n6841), .B(n6840), .ZN(P1_U3290) );
  OAI21_X1 U8672 ( .B1(n6844), .B2(n6850), .A(n6843), .ZN(n6893) );
  INV_X1 U8673 ( .A(n6893), .ZN(n6859) );
  INV_X1 U8674 ( .A(n6845), .ZN(n6849) );
  AND2_X1 U8675 ( .A1(n8275), .A2(n6846), .ZN(n8086) );
  INV_X1 U8676 ( .A(n8086), .ZN(n6847) );
  OR2_X1 U8677 ( .A1(n8271), .A2(n6847), .ZN(n6848) );
  AOI21_X1 U8678 ( .B1(n6849), .B2(n8086), .A(n8085), .ZN(n6878) );
  OAI21_X1 U8679 ( .B1(n6878), .B2(n6879), .A(n8091), .ZN(n6966) );
  XNOR2_X1 U8680 ( .A(n6966), .B(n6850), .ZN(n6851) );
  OAI222_X1 U8681 ( .A1(n9551), .A2(n7263), .B1(n9549), .B2(n6931), .C1(n6851), 
        .C2(n9546), .ZN(n6891) );
  INV_X1 U8682 ( .A(n6970), .ZN(n6852) );
  AOI211_X1 U8683 ( .C1(n6853), .C2(n6883), .A(n9682), .B(n6852), .ZN(n6892)
         );
  NAND2_X1 U8684 ( .A1(n6892), .A2(n9616), .ZN(n6856) );
  INV_X1 U8685 ( .A(n7264), .ZN(n6854) );
  INV_X1 U8686 ( .A(n9630), .ZN(n9617) );
  AOI22_X1 U8687 ( .A1(n9469), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6854), .B2(
        n9617), .ZN(n6855) );
  OAI211_X1 U8688 ( .C1(n4765), .C2(n9629), .A(n6856), .B(n6855), .ZN(n6857)
         );
  AOI21_X1 U8689 ( .B1(n6891), .B2(n9633), .A(n6857), .ZN(n6858) );
  OAI21_X1 U8690 ( .B1(n6859), .B2(n9650), .A(n6858), .ZN(P1_U3285) );
  INV_X1 U8691 ( .A(n6860), .ZN(n6867) );
  NAND2_X1 U8692 ( .A1(n6861), .A2(n7692), .ZN(n6866) );
  NOR2_X1 U8693 ( .A1(n9629), .A2(n5835), .ZN(n6863) );
  OAI22_X1 U8694 ( .A1(n7692), .A2(n5031), .B1(n9303), .B2(n9630), .ZN(n6862)
         );
  AOI211_X1 U8695 ( .C1(n6864), .C2(n9616), .A(n6863), .B(n6862), .ZN(n6865)
         );
  OAI211_X1 U8696 ( .C1(n6867), .C2(n9650), .A(n6866), .B(n6865), .ZN(P1_U3292) );
  XOR2_X1 U8697 ( .A(n6869), .B(n6868), .Z(n6873) );
  AOI22_X1 U8698 ( .A1(n8468), .A2(n10130), .B1(n8527), .B2(n8783), .ZN(n6870)
         );
  OAI21_X1 U8699 ( .B1(n8530), .B2(n6402), .A(n6870), .ZN(n6871) );
  AOI21_X1 U8700 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7209), .A(n6871), .ZN(
        n6872) );
  OAI21_X1 U8701 ( .B1(n6873), .B2(n8518), .A(n6872), .ZN(P2_U3177) );
  NAND2_X1 U8702 ( .A1(n6874), .A2(P1_U3973), .ZN(n6875) );
  OAI21_X1 U8703 ( .B1(P1_U3973), .B2(n7853), .A(n6875), .ZN(P1_U3582) );
  OAI21_X1 U8704 ( .B1(n6877), .B2(n6879), .A(n6876), .ZN(n6901) );
  INV_X1 U8705 ( .A(n6901), .ZN(n6890) );
  XOR2_X1 U8706 ( .A(n6879), .B(n6878), .Z(n6880) );
  OAI222_X1 U8707 ( .A1(n9549), .A2(n6882), .B1(n9551), .B2(n6881), .C1(n6880), 
        .C2(n9546), .ZN(n6899) );
  NAND2_X1 U8708 ( .A1(n6899), .A2(n7692), .ZN(n6889) );
  INV_X1 U8709 ( .A(n6883), .ZN(n6884) );
  AOI211_X1 U8710 ( .C1(n6902), .C2(n4441), .A(n9682), .B(n6884), .ZN(n6900)
         );
  NOR2_X1 U8711 ( .A1(n9629), .A2(n6904), .ZN(n6887) );
  OAI22_X1 U8712 ( .A1(n7692), .A2(n9404), .B1(n6885), .B2(n9630), .ZN(n6886)
         );
  AOI211_X1 U8713 ( .C1(n6900), .C2(n9616), .A(n6887), .B(n6886), .ZN(n6888)
         );
  OAI211_X1 U8714 ( .C1(n6890), .C2(n9650), .A(n6889), .B(n6888), .ZN(P1_U3286) );
  AOI211_X1 U8715 ( .C1(n9978), .C2(n6893), .A(n6892), .B(n6891), .ZN(n6898)
         );
  OAI22_X1 U8716 ( .A1(n4765), .A2(n9717), .B1(n9988), .B2(n9397), .ZN(n6894)
         );
  INV_X1 U8717 ( .A(n6894), .ZN(n6895) );
  OAI21_X1 U8718 ( .B1(n6898), .B2(n9986), .A(n6895), .ZN(P1_U3530) );
  OAI22_X1 U8719 ( .A1(n4765), .A2(n9770), .B1(n9981), .B2(n5259), .ZN(n6896)
         );
  INV_X1 U8720 ( .A(n6896), .ZN(n6897) );
  OAI21_X1 U8721 ( .B1(n6898), .B2(n9980), .A(n6897), .ZN(P1_U3477) );
  AOI211_X1 U8722 ( .C1(n9978), .C2(n6901), .A(n6900), .B(n6899), .ZN(n6907)
         );
  AOI22_X1 U8723 ( .A1(n5919), .A2(n6902), .B1(n9986), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n6903) );
  OAI21_X1 U8724 ( .B1(n6907), .B2(n9986), .A(n6903), .ZN(P1_U3529) );
  OAI22_X1 U8725 ( .A1(n9770), .A2(n6904), .B1(n9981), .B2(n5200), .ZN(n6905)
         );
  INV_X1 U8726 ( .A(n6905), .ZN(n6906) );
  OAI21_X1 U8727 ( .B1(n6907), .B2(n9980), .A(n6906), .ZN(P1_U3474) );
  XNOR2_X1 U8728 ( .A(n6908), .B(n8220), .ZN(n6909) );
  OAI222_X1 U8729 ( .A1(n9551), .A2(n6932), .B1(n9549), .B2(n6910), .C1(n6909), 
        .C2(n9546), .ZN(n9960) );
  INV_X1 U8730 ( .A(n9960), .ZN(n6922) );
  OAI21_X1 U8731 ( .B1(n6912), .B2(n8220), .A(n6911), .ZN(n9962) );
  INV_X1 U8732 ( .A(n9650), .ZN(n7286) );
  OAI211_X1 U8733 ( .C1(n6914), .C2(n9959), .A(n7288), .B(n6913), .ZN(n9958)
         );
  OAI22_X1 U8734 ( .A1(n7692), .A2(n6916), .B1(n6915), .B2(n9630), .ZN(n6917)
         );
  AOI21_X1 U8735 ( .B1(n7293), .B2(n6918), .A(n6917), .ZN(n6919) );
  OAI21_X1 U8736 ( .B1(n9958), .B2(n7290), .A(n6919), .ZN(n6920) );
  AOI21_X1 U8737 ( .B1(n9962), .B2(n7286), .A(n6920), .ZN(n6921) );
  OAI21_X1 U8738 ( .B1(n6922), .B2(n9469), .A(n6921), .ZN(P1_U3289) );
  INV_X1 U8739 ( .A(n6923), .ZN(n6927) );
  OAI222_X1 U8740 ( .A1(n9775), .A2(n6925), .B1(n8017), .B2(n6927), .C1(
        P1_U3086), .C2(n6924), .ZN(P1_U3334) );
  OAI222_X1 U8741 ( .A1(P2_U3151), .A2(n6928), .B1(n9175), .B2(n6927), .C1(
        n6926), .C2(n9172), .ZN(P2_U3274) );
  XNOR2_X1 U8742 ( .A(n6929), .B(n6937), .ZN(n6930) );
  NAND2_X1 U8743 ( .A1(n6930), .A2(n9640), .ZN(n6935) );
  OAI22_X1 U8744 ( .A1(n6932), .A2(n9549), .B1(n6931), .B2(n9551), .ZN(n6933)
         );
  INV_X1 U8745 ( .A(n6933), .ZN(n6934) );
  NAND2_X1 U8746 ( .A1(n6935), .A2(n6934), .ZN(n9965) );
  INV_X1 U8747 ( .A(n9965), .ZN(n6947) );
  OAI21_X1 U8748 ( .B1(n6938), .B2(n6937), .A(n6936), .ZN(n9967) );
  OAI211_X1 U8749 ( .C1(n9964), .C2(n6939), .A(n4441), .B(n7288), .ZN(n9963)
         );
  OAI22_X1 U8750 ( .A1(n7692), .A2(n6941), .B1(n6940), .B2(n9630), .ZN(n6942)
         );
  AOI21_X1 U8751 ( .B1(n7293), .B2(n6943), .A(n6942), .ZN(n6944) );
  OAI21_X1 U8752 ( .B1(n9963), .B2(n7290), .A(n6944), .ZN(n6945) );
  AOI21_X1 U8753 ( .B1(n9967), .B2(n7286), .A(n6945), .ZN(n6946) );
  OAI21_X1 U8754 ( .B1(n6947), .B2(n9469), .A(n6946), .ZN(P1_U3287) );
  NAND2_X1 U8755 ( .A1(n6948), .A2(n8280), .ZN(n6949) );
  NAND2_X1 U8756 ( .A1(n6949), .A2(n6956), .ZN(n6951) );
  NAND2_X1 U8757 ( .A1(n6951), .A2(n6950), .ZN(n6954) );
  OAI22_X1 U8758 ( .A1(n6952), .A2(n9551), .B1(n7263), .B2(n9549), .ZN(n6953)
         );
  AOI21_X1 U8759 ( .B1(n6954), .B2(n9640), .A(n6953), .ZN(n9974) );
  OAI21_X1 U8760 ( .B1(n6957), .B2(n6956), .A(n6955), .ZN(n9979) );
  NAND2_X1 U8761 ( .A1(n9979), .A2(n7286), .ZN(n6964) );
  OAI22_X1 U8762 ( .A1(n7692), .A2(n6958), .B1(n7672), .B2(n9630), .ZN(n6962)
         );
  INV_X1 U8763 ( .A(n6959), .ZN(n7219) );
  OAI211_X1 U8764 ( .C1(n9976), .C2(n6960), .A(n7219), .B(n7288), .ZN(n9973)
         );
  NOR2_X1 U8765 ( .A1(n9973), .A2(n7290), .ZN(n6961) );
  AOI211_X1 U8766 ( .C1(n7293), .C2(n7679), .A(n6962), .B(n6961), .ZN(n6963)
         );
  OAI211_X1 U8767 ( .C1(n9469), .C2(n9974), .A(n6964), .B(n6963), .ZN(P1_U3283) );
  INV_X1 U8768 ( .A(n8101), .ZN(n6965) );
  AOI21_X1 U8769 ( .B1(n6966), .B2(n8093), .A(n6965), .ZN(n6967) );
  XNOR2_X1 U8770 ( .A(n6967), .B(n6975), .ZN(n6968) );
  AOI22_X1 U8771 ( .A1(n6968), .A2(n9640), .B1(n9643), .B2(n9294), .ZN(n9970)
         );
  OAI22_X1 U8772 ( .A1(n7692), .A2(n6969), .B1(n7577), .B2(n9630), .ZN(n6973)
         );
  XOR2_X1 U8773 ( .A(n9968), .B(n6970), .Z(n6971) );
  AOI22_X1 U8774 ( .A1(n6971), .A2(n7288), .B1(n9644), .B2(n9292), .ZN(n9969)
         );
  NOR2_X1 U8775 ( .A1(n9969), .A2(n7290), .ZN(n6972) );
  AOI211_X1 U8776 ( .C1(n7293), .C2(n9968), .A(n6973), .B(n6972), .ZN(n6978)
         );
  OAI21_X1 U8777 ( .B1(n6976), .B2(n6975), .A(n6974), .ZN(n9972) );
  NAND2_X1 U8778 ( .A1(n9972), .A2(n7286), .ZN(n6977) );
  OAI211_X1 U8779 ( .C1(n9970), .C2(n9469), .A(n6978), .B(n6977), .ZN(P1_U3284) );
  INV_X1 U8780 ( .A(n6979), .ZN(n6988) );
  NAND2_X1 U8781 ( .A1(n6980), .A2(n7692), .ZN(n6987) );
  NOR2_X1 U8782 ( .A1(n9629), .A2(n6981), .ZN(n6984) );
  OAI22_X1 U8783 ( .A1(n7692), .A2(n9363), .B1(n6982), .B2(n9630), .ZN(n6983)
         );
  AOI211_X1 U8784 ( .C1(n6985), .C2(n9616), .A(n6984), .B(n6983), .ZN(n6986)
         );
  OAI211_X1 U8785 ( .C1(n6988), .C2(n9650), .A(n6987), .B(n6986), .ZN(P1_U3288) );
  AOI22_X1 U8786 ( .A1(SI_22_), .A2(keyinput_f10), .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n6989) );
  OAI221_X1 U8787 ( .B1(SI_22_), .B2(keyinput_f10), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n6989), .ZN(n6996) );
  AOI22_X1 U8788 ( .A1(SI_11_), .A2(keyinput_f21), .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n6990) );
  OAI221_X1 U8789 ( .B1(SI_11_), .B2(keyinput_f21), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n6990), .ZN(n6995) );
  AOI22_X1 U8790 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n6991) );
  OAI221_X1 U8791 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n6991), .ZN(n6994) );
  AOI22_X1 U8792 ( .A1(SI_25_), .A2(keyinput_f7), .B1(SI_28_), .B2(keyinput_f4), .ZN(n6992) );
  OAI221_X1 U8793 ( .B1(SI_25_), .B2(keyinput_f7), .C1(SI_28_), .C2(
        keyinput_f4), .A(n6992), .ZN(n6993) );
  NOR4_X1 U8794 ( .A1(n6996), .A2(n6995), .A3(n6994), .A4(n6993), .ZN(n7024)
         );
  XOR2_X1 U8795 ( .A(n7122), .B(keyinput_f9), .Z(n7003) );
  AOI22_X1 U8796 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_f41), .B1(n8406), 
        .B2(keyinput_f45), .ZN(n6997) );
  OAI221_X1 U8797 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .C1(n8406), .C2(keyinput_f45), .A(n6997), .ZN(n7002) );
  AOI22_X1 U8798 ( .A1(SI_26_), .A2(keyinput_f6), .B1(P2_REG3_REG_10__SCAN_IN), 
        .B2(keyinput_f39), .ZN(n6998) );
  OAI221_X1 U8799 ( .B1(SI_26_), .B2(keyinput_f6), .C1(P2_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n6998), .ZN(n7001) );
  AOI22_X1 U8800 ( .A1(SI_15_), .A2(keyinput_f17), .B1(SI_17_), .B2(
        keyinput_f15), .ZN(n6999) );
  OAI221_X1 U8801 ( .B1(SI_15_), .B2(keyinput_f17), .C1(SI_17_), .C2(
        keyinput_f15), .A(n6999), .ZN(n7000) );
  NOR4_X1 U8802 ( .A1(n7003), .A2(n7002), .A3(n7001), .A4(n7000), .ZN(n7023)
         );
  AOI22_X1 U8803 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(SI_3_), 
        .B2(keyinput_f29), .ZN(n7004) );
  OAI221_X1 U8804 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(SI_3_), 
        .C2(keyinput_f29), .A(n7004), .ZN(n7012) );
  AOI22_X1 U8805 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(keyinput_f42), .ZN(n7005) );
  OAI221_X1 U8806 ( .B1(SI_2_), .B2(keyinput_f30), .C1(P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n7005), .ZN(n7011) );
  AOI22_X1 U8807 ( .A1(n6168), .A2(keyinput_f50), .B1(keyinput_f33), .B2(n5006), .ZN(n7006) );
  OAI221_X1 U8808 ( .B1(n6168), .B2(keyinput_f50), .C1(n5006), .C2(
        keyinput_f33), .A(n7006), .ZN(n7010) );
  INV_X1 U8809 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8451) );
  AOI22_X1 U8810 ( .A1(n8451), .A2(keyinput_f51), .B1(n7008), .B2(keyinput_f36), .ZN(n7007) );
  OAI221_X1 U8811 ( .B1(n8451), .B2(keyinput_f51), .C1(n7008), .C2(
        keyinput_f36), .A(n7007), .ZN(n7009) );
  NOR4_X1 U8812 ( .A1(n7012), .A2(n7011), .A3(n7010), .A4(n7009), .ZN(n7022)
         );
  AOI22_X1 U8813 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(
        P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .ZN(n7013) );
  OAI221_X1 U8814 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n7013), .ZN(n7020) );
  AOI22_X1 U8815 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(keyinput_f47), .ZN(n7014) );
  OAI221_X1 U8816 ( .B1(SI_30_), .B2(keyinput_f2), .C1(P2_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n7014), .ZN(n7019) );
  AOI22_X1 U8817 ( .A1(SI_14_), .A2(keyinput_f18), .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n7015) );
  OAI221_X1 U8818 ( .B1(SI_14_), .B2(keyinput_f18), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n7015), .ZN(n7018) );
  AOI22_X1 U8819 ( .A1(SI_12_), .A2(keyinput_f20), .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n7016) );
  OAI221_X1 U8820 ( .B1(SI_12_), .B2(keyinput_f20), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n7016), .ZN(n7017) );
  NOR4_X1 U8821 ( .A1(n7020), .A2(n7019), .A3(n7018), .A4(n7017), .ZN(n7021)
         );
  NAND4_X1 U8822 ( .A1(n7024), .A2(n7023), .A3(n7022), .A4(n7021), .ZN(n7068)
         );
  INV_X1 U8823 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7189) );
  AOI22_X1 U8824 ( .A1(n7090), .A2(keyinput_f13), .B1(n7189), .B2(keyinput_f52), .ZN(n7025) );
  OAI221_X1 U8825 ( .B1(n7090), .B2(keyinput_f13), .C1(n7189), .C2(
        keyinput_f52), .A(n7025), .ZN(n7034) );
  INV_X1 U8826 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7448) );
  AOI22_X1 U8827 ( .A1(n5596), .A2(keyinput_f12), .B1(n7448), .B2(keyinput_f35), .ZN(n7026) );
  OAI221_X1 U8828 ( .B1(n5596), .B2(keyinput_f12), .C1(n7448), .C2(
        keyinput_f35), .A(n7026), .ZN(n7033) );
  INV_X1 U8829 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7124) );
  AOI22_X1 U8830 ( .A1(n7028), .A2(keyinput_f24), .B1(n7124), .B2(keyinput_f48), .ZN(n7027) );
  OAI221_X1 U8831 ( .B1(n7028), .B2(keyinput_f24), .C1(n7124), .C2(
        keyinput_f48), .A(n7027), .ZN(n7032) );
  XNOR2_X1 U8832 ( .A(SI_0_), .B(keyinput_f32), .ZN(n7030) );
  XNOR2_X1 U8833 ( .A(SI_6_), .B(keyinput_f26), .ZN(n7029) );
  NAND2_X1 U8834 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  NOR4_X1 U8835 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .ZN(n7066)
         );
  INV_X1 U8836 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7633) );
  AOI22_X1 U8837 ( .A1(n7633), .A2(keyinput_f43), .B1(P2_U3151), .B2(
        keyinput_f34), .ZN(n7035) );
  OAI221_X1 U8838 ( .B1(n7633), .B2(keyinput_f43), .C1(P2_U3151), .C2(
        keyinput_f34), .A(n7035), .ZN(n7043) );
  INV_X1 U8839 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8377) );
  AOI22_X1 U8840 ( .A1(n7144), .A2(keyinput_f5), .B1(n8377), .B2(keyinput_f38), 
        .ZN(n7036) );
  OAI221_X1 U8841 ( .B1(n7144), .B2(keyinput_f5), .C1(n8377), .C2(keyinput_f38), .A(n7036), .ZN(n7042) );
  INV_X1 U8842 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7877) );
  XOR2_X1 U8843 ( .A(n7877), .B(keyinput_f58), .Z(n7040) );
  XNOR2_X1 U8844 ( .A(SI_4_), .B(keyinput_f28), .ZN(n7039) );
  XNOR2_X1 U8845 ( .A(SI_5_), .B(keyinput_f27), .ZN(n7038) );
  XNOR2_X1 U8846 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n7037) );
  NAND4_X1 U8847 ( .A1(n7040), .A2(n7039), .A3(n7038), .A4(n7037), .ZN(n7041)
         );
  NOR3_X1 U8848 ( .A1(n7043), .A2(n7042), .A3(n7041), .ZN(n7065) );
  INV_X1 U8849 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7149) );
  AOI22_X1 U8850 ( .A1(n7149), .A2(keyinput_f56), .B1(keyinput_f53), .B2(n6070), .ZN(n7044) );
  OAI221_X1 U8851 ( .B1(n7149), .B2(keyinput_f56), .C1(n6070), .C2(
        keyinput_f53), .A(n7044), .ZN(n7053) );
  INV_X1 U8852 ( .A(SI_7_), .ZN(n7113) );
  AOI22_X1 U8853 ( .A1(n7113), .A2(keyinput_f25), .B1(n7046), .B2(keyinput_f23), .ZN(n7045) );
  OAI221_X1 U8854 ( .B1(n7113), .B2(keyinput_f25), .C1(n7046), .C2(
        keyinput_f23), .A(n7045), .ZN(n7052) );
  XNOR2_X1 U8855 ( .A(SI_21_), .B(keyinput_f11), .ZN(n7050) );
  XNOR2_X1 U8856 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_f59), .ZN(n7049) );
  XNOR2_X1 U8857 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_f44), .ZN(n7048) );
  XNOR2_X1 U8858 ( .A(SI_1_), .B(keyinput_f31), .ZN(n7047) );
  NAND4_X1 U8859 ( .A1(n7050), .A2(n7049), .A3(n7048), .A4(n7047), .ZN(n7051)
         );
  NOR3_X1 U8860 ( .A1(n7053), .A2(n7052), .A3(n7051), .ZN(n7064) );
  AOI22_X1 U8861 ( .A1(n4834), .A2(keyinput_f19), .B1(n7055), .B2(keyinput_f37), .ZN(n7054) );
  OAI221_X1 U8862 ( .B1(n4834), .B2(keyinput_f19), .C1(n7055), .C2(
        keyinput_f37), .A(n7054), .ZN(n7062) );
  INV_X1 U8863 ( .A(SI_18_), .ZN(n7127) );
  INV_X1 U8864 ( .A(SI_31_), .ZN(n8028) );
  AOI22_X1 U8865 ( .A1(n7127), .A2(keyinput_f14), .B1(keyinput_f1), .B2(n8028), 
        .ZN(n7056) );
  OAI221_X1 U8866 ( .B1(n7127), .B2(keyinput_f14), .C1(n8028), .C2(keyinput_f1), .A(n7056), .ZN(n7061) );
  INV_X1 U8867 ( .A(SI_29_), .ZN(n8018) );
  INV_X1 U8868 ( .A(SI_10_), .ZN(n7146) );
  AOI22_X1 U8869 ( .A1(n8018), .A2(keyinput_f3), .B1(keyinput_f22), .B2(n7146), 
        .ZN(n7057) );
  OAI221_X1 U8870 ( .B1(n8018), .B2(keyinput_f3), .C1(n7146), .C2(keyinput_f22), .A(n7057), .ZN(n7060) );
  AOI22_X1 U8871 ( .A1(n7112), .A2(keyinput_f8), .B1(keyinput_f16), .B2(n7147), 
        .ZN(n7058) );
  OAI221_X1 U8872 ( .B1(n7112), .B2(keyinput_f8), .C1(n7147), .C2(keyinput_f16), .A(n7058), .ZN(n7059) );
  NOR4_X1 U8873 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .ZN(n7063)
         );
  NAND4_X1 U8874 ( .A1(n7066), .A2(n7065), .A3(n7064), .A4(n7063), .ZN(n7067)
         );
  OAI22_X1 U8875 ( .A1(keyinput_f60), .A2(n7070), .B1(n7068), .B2(n7067), .ZN(
        n7069) );
  AOI21_X1 U8876 ( .B1(keyinput_f60), .B2(n7070), .A(n7069), .ZN(n7163) );
  AOI22_X1 U8877 ( .A1(SI_2_), .A2(keyinput_g30), .B1(SI_17_), .B2(
        keyinput_g15), .ZN(n7071) );
  OAI221_X1 U8878 ( .B1(SI_2_), .B2(keyinput_g30), .C1(SI_17_), .C2(
        keyinput_g15), .A(n7071), .ZN(n7078) );
  AOI22_X1 U8879 ( .A1(SI_13_), .A2(keyinput_g19), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_g33), .ZN(n7072) );
  OAI221_X1 U8880 ( .B1(SI_13_), .B2(keyinput_g19), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_g33), .A(n7072), .ZN(n7077) );
  AOI22_X1 U8881 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n7073) );
  OAI221_X1 U8882 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n7073), .ZN(n7076) );
  AOI22_X1 U8883 ( .A1(SI_20_), .A2(keyinput_g12), .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n7074) );
  OAI221_X1 U8884 ( .B1(SI_20_), .B2(keyinput_g12), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n7074), .ZN(n7075) );
  NOR4_X1 U8885 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n7108)
         );
  AOI22_X1 U8886 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_5_), 
        .B2(keyinput_g27), .ZN(n7079) );
  OAI221_X1 U8887 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(SI_5_), 
        .C2(keyinput_g27), .A(n7079), .ZN(n7086) );
  AOI22_X1 U8888 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(keyinput_g62), .ZN(n7080) );
  OAI221_X1 U8889 ( .B1(SI_4_), .B2(keyinput_g28), .C1(P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n7080), .ZN(n7085) );
  AOI22_X1 U8890 ( .A1(SI_8_), .A2(keyinput_g24), .B1(n7082), .B2(keyinput_g6), 
        .ZN(n7081) );
  OAI221_X1 U8891 ( .B1(SI_8_), .B2(keyinput_g24), .C1(n7082), .C2(keyinput_g6), .A(n7081), .ZN(n7084) );
  XNOR2_X1 U8892 ( .A(SI_0_), .B(keyinput_g32), .ZN(n7083) );
  NOR4_X1 U8893 ( .A1(n7086), .A2(n7085), .A3(n7084), .A4(n7083), .ZN(n7107)
         );
  AOI22_X1 U8894 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_14_), .B2(
        keyinput_g18), .ZN(n7087) );
  OAI221_X1 U8895 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_14_), .C2(
        keyinput_g18), .A(n7087), .ZN(n7096) );
  AOI22_X1 U8896 ( .A1(SI_22_), .A2(keyinput_g10), .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n7088) );
  OAI221_X1 U8897 ( .B1(SI_22_), .B2(keyinput_g10), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n7088), .ZN(n7095) );
  AOI22_X1 U8898 ( .A1(n8377), .A2(keyinput_g38), .B1(keyinput_g13), .B2(n7090), .ZN(n7089) );
  OAI221_X1 U8899 ( .B1(n8377), .B2(keyinput_g38), .C1(n7090), .C2(
        keyinput_g13), .A(n7089), .ZN(n7094) );
  INV_X1 U8900 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7274) );
  INV_X1 U8901 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7092) );
  AOI22_X1 U8902 ( .A1(n7274), .A2(keyinput_g61), .B1(keyinput_g54), .B2(n7092), .ZN(n7091) );
  OAI221_X1 U8903 ( .B1(n7274), .B2(keyinput_g61), .C1(n7092), .C2(
        keyinput_g54), .A(n7091), .ZN(n7093) );
  NOR4_X1 U8904 ( .A1(n7096), .A2(n7095), .A3(n7094), .A4(n7093), .ZN(n7106)
         );
  AOI22_X1 U8905 ( .A1(SI_25_), .A2(keyinput_g7), .B1(P2_STATE_REG_SCAN_IN), 
        .B2(keyinput_g34), .ZN(n7097) );
  OAI221_X1 U8906 ( .B1(SI_25_), .B2(keyinput_g7), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_g34), .A(n7097), .ZN(n7104) );
  AOI22_X1 U8907 ( .A1(SI_11_), .A2(keyinput_g21), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n7098) );
  OAI221_X1 U8908 ( .B1(SI_11_), .B2(keyinput_g21), .C1(SI_15_), .C2(
        keyinput_g17), .A(n7098), .ZN(n7103) );
  AOI22_X1 U8909 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(keyinput_g37), .ZN(n7099) );
  OAI221_X1 U8910 ( .B1(SI_29_), .B2(keyinput_g3), .C1(P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n7099), .ZN(n7102) );
  AOI22_X1 U8911 ( .A1(SI_9_), .A2(keyinput_g23), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n7100) );
  OAI221_X1 U8912 ( .B1(SI_9_), .B2(keyinput_g23), .C1(P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n7100), .ZN(n7101) );
  NOR4_X1 U8913 ( .A1(n7104), .A2(n7103), .A3(n7102), .A4(n7101), .ZN(n7105)
         );
  NAND4_X1 U8914 ( .A1(n7108), .A2(n7107), .A3(n7106), .A4(n7105), .ZN(n7161)
         );
  AOI22_X1 U8915 ( .A1(n7189), .A2(keyinput_g52), .B1(keyinput_g11), .B2(n7110), .ZN(n7109) );
  OAI221_X1 U8916 ( .B1(n7189), .B2(keyinput_g52), .C1(n7110), .C2(
        keyinput_g11), .A(n7109), .ZN(n7120) );
  AOI22_X1 U8917 ( .A1(n7113), .A2(keyinput_g25), .B1(n7112), .B2(keyinput_g8), 
        .ZN(n7111) );
  OAI221_X1 U8918 ( .B1(n7113), .B2(keyinput_g25), .C1(n7112), .C2(keyinput_g8), .A(n7111), .ZN(n7119) );
  XNOR2_X1 U8919 ( .A(SI_6_), .B(keyinput_g26), .ZN(n7117) );
  XNOR2_X1 U8920 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_g45), .ZN(n7116)
         );
  XNOR2_X1 U8921 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_g55), .ZN(n7115)
         );
  XNOR2_X1 U8922 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_g44), .ZN(n7114) );
  NAND4_X1 U8923 ( .A1(n7117), .A2(n7116), .A3(n7115), .A4(n7114), .ZN(n7118)
         );
  NOR3_X1 U8924 ( .A1(n7120), .A2(n7119), .A3(n7118), .ZN(n7159) );
  INV_X1 U8925 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9835) );
  AOI22_X1 U8926 ( .A1(n9835), .A2(keyinput_g0), .B1(n7122), .B2(keyinput_g9), 
        .ZN(n7121) );
  OAI221_X1 U8927 ( .B1(n9835), .B2(keyinput_g0), .C1(n7122), .C2(keyinput_g9), 
        .A(n7121), .ZN(n7131) );
  AOI22_X1 U8928 ( .A1(n7124), .A2(keyinput_g48), .B1(keyinput_g49), .B2(n7229), .ZN(n7123) );
  OAI221_X1 U8929 ( .B1(n7124), .B2(keyinput_g48), .C1(n7229), .C2(
        keyinput_g49), .A(n7123), .ZN(n7130) );
  INV_X1 U8930 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8419) );
  AOI22_X1 U8931 ( .A1(n8419), .A2(keyinput_g47), .B1(keyinput_g1), .B2(n8028), 
        .ZN(n7125) );
  OAI221_X1 U8932 ( .B1(n8419), .B2(keyinput_g47), .C1(n8028), .C2(keyinput_g1), .A(n7125), .ZN(n7129) );
  AOI22_X1 U8933 ( .A1(n7127), .A2(keyinput_g14), .B1(n6070), .B2(keyinput_g53), .ZN(n7126) );
  OAI221_X1 U8934 ( .B1(n7127), .B2(keyinput_g14), .C1(n6070), .C2(
        keyinput_g53), .A(n7126), .ZN(n7128) );
  NOR4_X1 U8935 ( .A1(n7131), .A2(n7130), .A3(n7129), .A4(n7128), .ZN(n7158)
         );
  INV_X1 U8936 ( .A(SI_30_), .ZN(n7133) );
  AOI22_X1 U8937 ( .A1(n6168), .A2(keyinput_g50), .B1(keyinput_g2), .B2(n7133), 
        .ZN(n7132) );
  OAI221_X1 U8938 ( .B1(n6168), .B2(keyinput_g50), .C1(n7133), .C2(keyinput_g2), .A(n7132), .ZN(n7142) );
  INV_X1 U8939 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7307) );
  AOI22_X1 U8940 ( .A1(n7307), .A2(keyinput_g40), .B1(keyinput_g20), .B2(n7135), .ZN(n7134) );
  OAI221_X1 U8941 ( .B1(n7307), .B2(keyinput_g40), .C1(n7135), .C2(
        keyinput_g20), .A(n7134), .ZN(n7141) );
  AOI22_X1 U8942 ( .A1(n7633), .A2(keyinput_g43), .B1(n8451), .B2(keyinput_g51), .ZN(n7136) );
  OAI221_X1 U8943 ( .B1(n7633), .B2(keyinput_g43), .C1(n8451), .C2(
        keyinput_g51), .A(n7136), .ZN(n7140) );
  XNOR2_X1 U8944 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_g36), .ZN(n7138)
         );
  XNOR2_X1 U8945 ( .A(SI_1_), .B(keyinput_g31), .ZN(n7137) );
  NAND2_X1 U8946 ( .A1(n7138), .A2(n7137), .ZN(n7139) );
  NOR4_X1 U8947 ( .A1(n7142), .A2(n7141), .A3(n7140), .A4(n7139), .ZN(n7157)
         );
  AOI22_X1 U8948 ( .A1(n7754), .A2(keyinput_g39), .B1(keyinput_g5), .B2(n7144), 
        .ZN(n7143) );
  OAI221_X1 U8949 ( .B1(n7754), .B2(keyinput_g39), .C1(n7144), .C2(keyinput_g5), .A(n7143), .ZN(n7155) );
  AOI22_X1 U8950 ( .A1(n7147), .A2(keyinput_g16), .B1(keyinput_g22), .B2(n7146), .ZN(n7145) );
  OAI221_X1 U8951 ( .B1(n7147), .B2(keyinput_g16), .C1(n7146), .C2(
        keyinput_g22), .A(n7145), .ZN(n7154) );
  AOI22_X1 U8952 ( .A1(n7149), .A2(keyinput_g56), .B1(keyinput_g35), .B2(n7448), .ZN(n7148) );
  OAI221_X1 U8953 ( .B1(n7149), .B2(keyinput_g56), .C1(n7448), .C2(
        keyinput_g35), .A(n7148), .ZN(n7153) );
  AOI22_X1 U8954 ( .A1(n7151), .A2(keyinput_g4), .B1(n7877), .B2(keyinput_g58), 
        .ZN(n7150) );
  OAI221_X1 U8955 ( .B1(n7151), .B2(keyinput_g4), .C1(n7877), .C2(keyinput_g58), .A(n7150), .ZN(n7152) );
  NOR4_X1 U8956 ( .A1(n7155), .A2(n7154), .A3(n7153), .A4(n7152), .ZN(n7156)
         );
  NAND4_X1 U8957 ( .A1(n7159), .A2(n7158), .A3(n7157), .A4(n7156), .ZN(n7160)
         );
  OAI22_X1 U8958 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(n7161), 
        .B2(n7160), .ZN(n7162) );
  AOI211_X1 U8959 ( .C1(P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n7163), 
        .B(n7162), .ZN(n7183) );
  INV_X1 U8960 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10232) );
  NOR2_X1 U8961 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7164) );
  AOI21_X1 U8962 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7164), .ZN(n10237) );
  NOR2_X1 U8963 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7165) );
  AOI21_X1 U8964 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7165), .ZN(n10240) );
  NOR2_X1 U8965 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7166) );
  AOI21_X1 U8966 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7166), .ZN(n10243) );
  NOR2_X1 U8967 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7167) );
  AOI21_X1 U8968 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7167), .ZN(n10246) );
  NOR2_X1 U8969 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7168) );
  AOI21_X1 U8970 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7168), .ZN(n10249) );
  NOR2_X1 U8971 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7169) );
  AOI21_X1 U8972 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7169), .ZN(n10252) );
  NOR2_X1 U8973 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7170) );
  AOI21_X1 U8974 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7170), .ZN(n10255) );
  NOR2_X1 U8975 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7171) );
  AOI21_X1 U8976 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7171), .ZN(n10258) );
  NOR2_X1 U8977 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7172) );
  AOI21_X1 U8978 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7172), .ZN(n10264) );
  NOR2_X1 U8979 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7173) );
  AOI21_X1 U8980 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7173), .ZN(n10267) );
  NOR2_X1 U8981 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7174) );
  AOI21_X1 U8982 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7174), .ZN(n10270) );
  NOR2_X1 U8983 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7175) );
  AOI21_X1 U8984 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7175), .ZN(n10273) );
  NOR2_X1 U8985 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n7176) );
  AOI21_X1 U8986 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n7176), .ZN(n10276) );
  AND2_X1 U8987 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7177) );
  NOR2_X1 U8988 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7177), .ZN(n10227) );
  INV_X1 U8989 ( .A(n10227), .ZN(n10228) );
  INV_X1 U8990 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10230) );
  NAND3_X1 U8991 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10229) );
  NAND2_X1 U8992 ( .A1(n10230), .A2(n10229), .ZN(n10226) );
  NAND2_X1 U8993 ( .A1(n10228), .A2(n10226), .ZN(n10261) );
  NAND2_X1 U8994 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7178) );
  OAI21_X1 U8995 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7178), .ZN(n10260) );
  NOR2_X1 U8996 ( .A1(n10261), .A2(n10260), .ZN(n10259) );
  AOI21_X1 U8997 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10259), .ZN(n10279) );
  NAND2_X1 U8998 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7179) );
  OAI21_X1 U8999 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7179), .ZN(n10278) );
  NOR2_X1 U9000 ( .A1(n10279), .A2(n10278), .ZN(n10277) );
  AOI21_X1 U9001 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10277), .ZN(n10282) );
  NOR2_X1 U9002 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7180) );
  AOI21_X1 U9003 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7180), .ZN(n10281) );
  NAND2_X1 U9004 ( .A1(n10282), .A2(n10281), .ZN(n10280) );
  OAI21_X1 U9005 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10280), .ZN(n10275) );
  NAND2_X1 U9006 ( .A1(n10276), .A2(n10275), .ZN(n10274) );
  OAI21_X1 U9007 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10274), .ZN(n10272) );
  NAND2_X1 U9008 ( .A1(n10273), .A2(n10272), .ZN(n10271) );
  OAI21_X1 U9009 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10271), .ZN(n10269) );
  NAND2_X1 U9010 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  OAI21_X1 U9011 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10268), .ZN(n10266) );
  NAND2_X1 U9012 ( .A1(n10267), .A2(n10266), .ZN(n10265) );
  OAI21_X1 U9013 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10265), .ZN(n10263) );
  NAND2_X1 U9014 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  OAI21_X1 U9015 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10262), .ZN(n10257) );
  NAND2_X1 U9016 ( .A1(n10258), .A2(n10257), .ZN(n10256) );
  OAI21_X1 U9017 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10256), .ZN(n10254) );
  NAND2_X1 U9018 ( .A1(n10255), .A2(n10254), .ZN(n10253) );
  OAI21_X1 U9019 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10253), .ZN(n10251) );
  NAND2_X1 U9020 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  OAI21_X1 U9021 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10250), .ZN(n10248) );
  NAND2_X1 U9022 ( .A1(n10249), .A2(n10248), .ZN(n10247) );
  OAI21_X1 U9023 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10247), .ZN(n10245) );
  NAND2_X1 U9024 ( .A1(n10246), .A2(n10245), .ZN(n10244) );
  OAI21_X1 U9025 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10244), .ZN(n10242) );
  NAND2_X1 U9026 ( .A1(n10243), .A2(n10242), .ZN(n10241) );
  OAI21_X1 U9027 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10241), .ZN(n10239) );
  NAND2_X1 U9028 ( .A1(n10240), .A2(n10239), .ZN(n10238) );
  OAI21_X1 U9029 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10238), .ZN(n10236) );
  NAND2_X1 U9030 ( .A1(n10237), .A2(n10236), .ZN(n10235) );
  OAI21_X1 U9031 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10235), .ZN(n10233) );
  NAND2_X1 U9032 ( .A1(n10232), .A2(n10233), .ZN(n7181) );
  NOR2_X1 U9033 ( .A1(n10232), .A2(n10233), .ZN(n10231) );
  AOI21_X1 U9034 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7181), .A(n10231), .ZN(
        n7182) );
  XOR2_X1 U9035 ( .A(n7183), .B(n7182), .Z(n7185) );
  XNOR2_X1 U9036 ( .A(n4492), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7184) );
  XNOR2_X1 U9037 ( .A(n7185), .B(n7184), .ZN(ADD_1068_U4) );
  OAI21_X1 U9038 ( .B1(n7188), .B2(n7187), .A(n7186), .ZN(n7195) );
  NOR2_X1 U9039 ( .A1(n8524), .A2(n10137), .ZN(n7194) );
  NAND2_X1 U9040 ( .A1(n8478), .A2(n10139), .ZN(n7191) );
  NOR2_X1 U9041 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7189), .ZN(n7359) );
  AOI21_X1 U9042 ( .B1(n8527), .B2(n10130), .A(n7359), .ZN(n7190) );
  OAI211_X1 U9043 ( .C1(n7192), .C2(n8523), .A(n7191), .B(n7190), .ZN(n7193)
         );
  AOI211_X1 U9044 ( .C1(n7195), .C2(n8507), .A(n7194), .B(n7193), .ZN(n7196)
         );
  INV_X1 U9045 ( .A(n7196), .ZN(P2_U3170) );
  NAND2_X1 U9046 ( .A1(n8478), .A2(n10156), .ZN(n7198) );
  NOR2_X1 U9047 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7307), .ZN(n9996) );
  AOI21_X1 U9048 ( .B1(n8527), .B2(n8782), .A(n9996), .ZN(n7197) );
  OAI211_X1 U9049 ( .C1(n7594), .C2(n8523), .A(n7198), .B(n7197), .ZN(n7203)
         );
  AOI211_X1 U9050 ( .C1(n7201), .C2(n7200), .A(n8518), .B(n7199), .ZN(n7202)
         );
  AOI211_X1 U9051 ( .C1(n7307), .C2(n8514), .A(n7203), .B(n7202), .ZN(n7204)
         );
  INV_X1 U9052 ( .A(n7204), .ZN(P2_U3158) );
  XOR2_X1 U9053 ( .A(n7206), .B(n7205), .Z(n7211) );
  AOI22_X1 U9054 ( .A1(n8468), .A2(n8782), .B1(n8527), .B2(n8784), .ZN(n7207)
         );
  OAI21_X1 U9055 ( .B1(n8530), .B2(n10147), .A(n7207), .ZN(n7208) );
  AOI21_X1 U9056 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7209), .A(n7208), .ZN(
        n7210) );
  OAI21_X1 U9057 ( .B1(n8518), .B2(n7211), .A(n7210), .ZN(P2_U3162) );
  OAI21_X1 U9058 ( .B1(n7214), .B2(n7213), .A(n7212), .ZN(n7215) );
  AOI222_X1 U9059 ( .A1(n9640), .A2(n7215), .B1(n9290), .B2(n9644), .C1(n9292), 
        .C2(n9643), .ZN(n7311) );
  OAI21_X1 U9060 ( .B1(n7217), .B2(n8230), .A(n7216), .ZN(n7314) );
  NAND2_X1 U9061 ( .A1(n7314), .A2(n7286), .ZN(n7225) );
  INV_X1 U9062 ( .A(n7218), .ZN(n7289) );
  AOI211_X1 U9063 ( .C1(n7610), .C2(n7219), .A(n9682), .B(n7289), .ZN(n7313)
         );
  NOR2_X1 U9064 ( .A1(n7220), .A2(n9629), .ZN(n7223) );
  OAI22_X1 U9065 ( .A1(n9633), .A2(n7221), .B1(n7608), .B2(n9630), .ZN(n7222)
         );
  AOI211_X1 U9066 ( .C1(n7313), .C2(n9616), .A(n7223), .B(n7222), .ZN(n7224)
         );
  OAI211_X1 U9067 ( .C1(n9469), .C2(n7311), .A(n7225), .B(n7224), .ZN(P1_U3282) );
  XOR2_X1 U9068 ( .A(n7227), .B(n7226), .Z(n7235) );
  INV_X1 U9069 ( .A(n7591), .ZN(n7233) );
  NAND2_X1 U9070 ( .A1(n8478), .A2(n7228), .ZN(n7231) );
  NOR2_X1 U9071 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7229), .ZN(n10012) );
  AOI21_X1 U9072 ( .B1(n8527), .B2(n8618), .A(n10012), .ZN(n7230) );
  OAI211_X1 U9073 ( .C1(n7595), .C2(n8523), .A(n7231), .B(n7230), .ZN(n7232)
         );
  AOI21_X1 U9074 ( .B1(n7233), .B2(n8514), .A(n7232), .ZN(n7234) );
  OAI21_X1 U9075 ( .B1(n7235), .B2(n8518), .A(n7234), .ZN(P2_U3167) );
  XNOR2_X1 U9076 ( .A(n8563), .B(n7236), .ZN(n10152) );
  INV_X1 U9077 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7344) );
  NOR2_X1 U9078 ( .A1(n6402), .A2(n8899), .ZN(n7245) );
  AOI22_X1 U9079 ( .A1(n10130), .A2(n10131), .B1(n10129), .B2(n8783), .ZN(
        n7244) );
  INV_X1 U9080 ( .A(n7237), .ZN(n7242) );
  AND3_X1 U9081 ( .A1(n7238), .A2(n7239), .A3(n7240), .ZN(n7241) );
  OAI21_X1 U9082 ( .B1(n7242), .B2(n7241), .A(n10134), .ZN(n7243) );
  OAI211_X1 U9083 ( .C1(n10152), .C2(n7622), .A(n7244), .B(n7243), .ZN(n10154)
         );
  AOI211_X1 U9084 ( .C1(n10140), .C2(P2_REG3_REG_2__SCAN_IN), .A(n7245), .B(
        n10154), .ZN(n7246) );
  MUX2_X1 U9085 ( .A(n7344), .B(n7246), .S(n10145), .Z(n7247) );
  OAI21_X1 U9086 ( .B1(n10152), .B2(n7628), .A(n7247), .ZN(P2_U3231) );
  NAND3_X1 U9087 ( .A1(n8217), .A2(n7249), .A3(n7248), .ZN(n7251) );
  AOI21_X1 U9088 ( .B1(n7251), .B2(n7250), .A(n9469), .ZN(n7256) );
  NAND2_X1 U9089 ( .A1(n9616), .A2(n7288), .ZN(n9563) );
  AOI21_X1 U9090 ( .B1(n9563), .B2(n9629), .A(n7252), .ZN(n7255) );
  OAI22_X1 U9091 ( .A1(n9633), .A2(n5054), .B1(n7253), .B2(n9630), .ZN(n7254)
         );
  OR3_X1 U9092 ( .A1(n7256), .A2(n7255), .A3(n7254), .ZN(P1_U3293) );
  INV_X1 U9093 ( .A(n7257), .ZN(n7269) );
  OAI222_X1 U9094 ( .A1(n8597), .A2(P2_U3151), .B1(n9175), .B2(n7269), .C1(
        n7258), .C2(n9172), .ZN(P2_U3273) );
  XNOR2_X1 U9095 ( .A(n7579), .B(n7259), .ZN(n7260) );
  NAND2_X1 U9096 ( .A1(n7260), .A2(n7261), .ZN(n7578) );
  OAI21_X1 U9097 ( .B1(n7261), .B2(n7260), .A(n7578), .ZN(n7262) );
  NAND2_X1 U9098 ( .A1(n7262), .A2(n9274), .ZN(n7268) );
  NAND2_X1 U9099 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9394) );
  OAI21_X1 U9100 ( .B1(n9279), .B2(n7263), .A(n9394), .ZN(n7266) );
  NOR2_X1 U9101 ( .A1(n9260), .A2(n7264), .ZN(n7265) );
  AOI211_X1 U9102 ( .C1(n9277), .C2(n9295), .A(n7266), .B(n7265), .ZN(n7267)
         );
  OAI211_X1 U9103 ( .C1(n4765), .C2(n9285), .A(n7268), .B(n7267), .ZN(P1_U3221) );
  OAI222_X1 U9104 ( .A1(n9775), .A2(n7270), .B1(n8254), .B2(P1_U3086), .C1(
        n8017), .C2(n7269), .ZN(P1_U3333) );
  OAI211_X1 U9105 ( .C1(n7273), .C2(n7272), .A(n7271), .B(n8507), .ZN(n7279)
         );
  NAND2_X1 U9106 ( .A1(n8478), .A2(n10172), .ZN(n7276) );
  NOR2_X1 U9107 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7274), .ZN(n7422) );
  AOI21_X1 U9108 ( .B1(n8527), .B2(n10132), .A(n7422), .ZN(n7275) );
  OAI211_X1 U9109 ( .C1(n7656), .C2(n8523), .A(n7276), .B(n7275), .ZN(n7277)
         );
  INV_X1 U9110 ( .A(n7277), .ZN(n7278) );
  OAI211_X1 U9111 ( .C1(n7661), .C2(n8524), .A(n7279), .B(n7278), .ZN(P2_U3179) );
  OAI21_X1 U9112 ( .B1(n7282), .B2(n7281), .A(n7280), .ZN(n7283) );
  AOI222_X1 U9113 ( .A1(n9640), .A2(n7283), .B1(n9289), .B2(n9644), .C1(n9291), 
        .C2(n9643), .ZN(n7399) );
  OAI21_X1 U9114 ( .B1(n7285), .B2(n8232), .A(n7284), .ZN(n7402) );
  NAND2_X1 U9115 ( .A1(n7402), .A2(n7286), .ZN(n7295) );
  OAI22_X1 U9116 ( .A1(n7692), .A2(n7287), .B1(n7378), .B2(n9630), .ZN(n7292)
         );
  OAI211_X1 U9117 ( .C1(n7289), .C2(n7400), .A(n7288), .B(n7386), .ZN(n7398)
         );
  NOR2_X1 U9118 ( .A1(n7398), .A2(n7290), .ZN(n7291) );
  AOI211_X1 U9119 ( .C1(n7293), .C2(n7380), .A(n7292), .B(n7291), .ZN(n7294)
         );
  OAI211_X1 U9120 ( .C1(n9469), .C2(n7399), .A(n7295), .B(n7294), .ZN(P1_U3281) );
  OAI21_X1 U9121 ( .B1(n7296), .B2(n7302), .A(n7297), .ZN(n10157) );
  INV_X1 U9122 ( .A(n10157), .ZN(n7310) );
  INV_X1 U9123 ( .A(n7298), .ZN(n7299) );
  NAND2_X1 U9124 ( .A1(n7299), .A2(n7622), .ZN(n7300) );
  NAND3_X1 U9125 ( .A1(n7237), .A2(n7302), .A3(n7301), .ZN(n7303) );
  NAND2_X1 U9126 ( .A1(n7304), .A2(n7303), .ZN(n7305) );
  AOI222_X1 U9127 ( .A1(n10134), .A2(n7305), .B1(n8782), .B2(n10129), .C1(
        n8618), .C2(n10131), .ZN(n10159) );
  MUX2_X1 U9128 ( .A(n7306), .B(n10159), .S(n10145), .Z(n7309) );
  AOI22_X1 U9129 ( .A1(n10138), .A2(n10156), .B1(n7307), .B2(n10140), .ZN(
        n7308) );
  OAI211_X1 U9130 ( .C1(n7310), .C2(n9026), .A(n7309), .B(n7308), .ZN(P2_U3230) );
  INV_X1 U9131 ( .A(n7311), .ZN(n7312) );
  AOI211_X1 U9132 ( .C1(n7314), .C2(n9978), .A(n7313), .B(n7312), .ZN(n7317)
         );
  AOI22_X1 U9133 ( .A1(n7610), .A2(n5926), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n9980), .ZN(n7315) );
  OAI21_X1 U9134 ( .B1(n7317), .B2(n9980), .A(n7315), .ZN(P1_U3486) );
  AOI22_X1 U9135 ( .A1(n7610), .A2(n5919), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n9986), .ZN(n7316) );
  OAI21_X1 U9136 ( .B1(n7317), .B2(n9986), .A(n7316), .ZN(P1_U3533) );
  NAND2_X1 U9137 ( .A1(n7321), .A2(n7850), .ZN(n7319) );
  NAND2_X1 U9138 ( .A1(n7318), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8769) );
  OAI211_X1 U9139 ( .C1(n7320), .C2(n9172), .A(n7319), .B(n8769), .ZN(P2_U3272) );
  NAND2_X1 U9140 ( .A1(n7321), .A2(n9780), .ZN(n7322) );
  OAI211_X1 U9141 ( .C1(n7323), .C2(n9775), .A(n7322), .B(n8329), .ZN(P1_U3332) );
  MUX2_X1 U9142 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8799), .Z(n7407) );
  XNOR2_X1 U9143 ( .A(n7407), .B(n7413), .ZN(n7328) );
  MUX2_X1 U9144 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8799), .Z(n7326) );
  MUX2_X1 U9145 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8799), .Z(n7325) );
  MUX2_X1 U9146 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8806), .Z(n7324) );
  XNOR2_X1 U9147 ( .A(n7324), .B(n7483), .ZN(n7479) );
  INV_X1 U9148 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7456) );
  AOI21_X1 U9149 ( .B1(n7324), .B2(n7483), .A(n7477), .ZN(n7489) );
  XNOR2_X1 U9150 ( .A(n7325), .B(n7487), .ZN(n7490) );
  AOI21_X1 U9151 ( .B1(n7325), .B2(n7487), .A(n7488), .ZN(n9999) );
  XOR2_X1 U9152 ( .A(n7348), .B(n7326), .Z(n9998) );
  NAND2_X1 U9153 ( .A1(n9999), .A2(n9998), .ZN(n9997) );
  OAI21_X1 U9154 ( .B1(n7326), .B2(n7348), .A(n9997), .ZN(n7327) );
  NAND2_X1 U9155 ( .A1(P2_U3893), .A2(n6334), .ZN(n10004) );
  AOI211_X1 U9156 ( .C1(n7328), .C2(n7327), .A(n10004), .B(n7406), .ZN(n7365)
         );
  INV_X1 U9157 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7363) );
  OR2_X1 U9158 ( .A1(P2_U3150), .A2(n7355), .ZN(n10020) );
  OR2_X1 U9159 ( .A1(n6334), .A2(P2_U3151), .ZN(n7851) );
  INV_X1 U9160 ( .A(n7851), .ZN(n7354) );
  AND2_X1 U9161 ( .A1(n7356), .A2(n7354), .ZN(n7459) );
  INV_X1 U9162 ( .A(n7459), .ZN(n7329) );
  OR2_X1 U9163 ( .A1(n7329), .A2(n8811), .ZN(n8840) );
  INV_X1 U9164 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7330) );
  MUX2_X1 U9165 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7330), .S(n7413), .Z(n7342)
         );
  INV_X1 U9166 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7331) );
  MUX2_X1 U9167 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7331), .S(n7487), .Z(n7495)
         );
  NAND2_X1 U9168 ( .A1(n5995), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7335) );
  NAND2_X1 U9169 ( .A1(n7483), .A2(n7335), .ZN(n7334) );
  NAND2_X1 U9170 ( .A1(n7456), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7332) );
  OR2_X1 U9171 ( .A1(n7332), .A2(n5995), .ZN(n7333) );
  NAND2_X1 U9172 ( .A1(n7334), .A2(n7333), .ZN(n7482) );
  NAND2_X1 U9173 ( .A1(n7482), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7336) );
  NAND2_X1 U9174 ( .A1(n7336), .A2(n7335), .ZN(n7494) );
  NAND2_X1 U9175 ( .A1(n7495), .A2(n7494), .ZN(n7493) );
  NAND2_X1 U9176 ( .A1(n7487), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7337) );
  NAND2_X1 U9177 ( .A1(n7493), .A2(n7337), .ZN(n7338) );
  NAND2_X1 U9178 ( .A1(n9989), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U9179 ( .A1(n7338), .A2(n7348), .ZN(n7339) );
  NAND2_X1 U9180 ( .A1(n7340), .A2(n7339), .ZN(n7341) );
  NAND2_X1 U9181 ( .A1(n7341), .A2(n7342), .ZN(n7415) );
  OAI21_X1 U9182 ( .B1(n7342), .B2(n7341), .A(n7415), .ZN(n7353) );
  AND2_X1 U9183 ( .A1(n7459), .A2(n8811), .ZN(n10010) );
  OR2_X1 U9184 ( .A1(n7413), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7343) );
  NAND2_X1 U9185 ( .A1(n7413), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7424) );
  AND2_X1 U9186 ( .A1(n7343), .A2(n7424), .ZN(n7351) );
  AND2_X1 U9187 ( .A1(n7456), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7345) );
  NAND2_X1 U9188 ( .A1(n5995), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7346) );
  OAI21_X1 U9189 ( .B1(n7483), .B2(n7345), .A(n7346), .ZN(n7474) );
  INV_X1 U9190 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7473) );
  OR2_X1 U9191 ( .A1(n7474), .A2(n7473), .ZN(n7476) );
  NAND2_X1 U9192 ( .A1(n7476), .A2(n7346), .ZN(n7497) );
  NAND2_X1 U9193 ( .A1(n7498), .A2(n7497), .ZN(n7496) );
  NAND2_X1 U9194 ( .A1(n7487), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U9195 ( .A1(n7350), .A2(n7351), .ZN(n7425) );
  OAI21_X1 U9196 ( .B1(n7351), .B2(n7350), .A(n7425), .ZN(n7352) );
  AOI22_X1 U9197 ( .A1(n10116), .A2(n7353), .B1(n10010), .B2(n7352), .ZN(n7362) );
  NAND2_X1 U9198 ( .A1(n7355), .A2(n7354), .ZN(n7358) );
  NOR2_X1 U9199 ( .A1(n8806), .A2(P2_U3151), .ZN(n7779) );
  NAND3_X1 U9200 ( .A1(n7356), .A2(n7779), .A3(n6334), .ZN(n7357) );
  NAND2_X1 U9201 ( .A1(n7358), .A2(n7357), .ZN(n10107) );
  INV_X1 U9202 ( .A(n7413), .ZN(n7360) );
  AOI21_X1 U9203 ( .B1(n10107), .B2(n7360), .A(n7359), .ZN(n7361) );
  OAI211_X1 U9204 ( .C1(n7363), .C2(n10020), .A(n7362), .B(n7361), .ZN(n7364)
         );
  OR2_X1 U9205 ( .A1(n7365), .A2(n7364), .ZN(P2_U3186) );
  NAND2_X1 U9206 ( .A1(n7367), .A2(n10186), .ZN(n7370) );
  NAND2_X1 U9207 ( .A1(n10140), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7368) );
  OAI211_X1 U9208 ( .C1(n8565), .C2(n7370), .A(n7369), .B(n7368), .ZN(n7371)
         );
  MUX2_X1 U9209 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n7371), .S(n10145), .Z(n7372)
         );
  AOI21_X1 U9210 ( .B1(n10138), .B2(n6821), .A(n7372), .ZN(n7373) );
  INV_X1 U9211 ( .A(n7373), .ZN(P2_U3233) );
  XOR2_X1 U9212 ( .A(n7374), .B(n7375), .Z(n7382) );
  NAND2_X1 U9213 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9865) );
  OAI21_X1 U9214 ( .B1(n9279), .B2(n7559), .A(n9865), .ZN(n7376) );
  AOI21_X1 U9215 ( .B1(n9277), .B2(n9291), .A(n7376), .ZN(n7377) );
  OAI21_X1 U9216 ( .B1(n9260), .B2(n7378), .A(n7377), .ZN(n7379) );
  AOI21_X1 U9217 ( .B1(n7380), .B2(n9265), .A(n7379), .ZN(n7381) );
  OAI21_X1 U9218 ( .B1(n7382), .B2(n9267), .A(n7381), .ZN(P1_U3224) );
  OAI21_X1 U9219 ( .B1(n7384), .B2(n7390), .A(n7383), .ZN(n7568) );
  INV_X1 U9220 ( .A(n7568), .ZN(n7397) );
  INV_X1 U9221 ( .A(n7560), .ZN(n7385) );
  AOI211_X1 U9222 ( .C1(n7549), .C2(n7386), .A(n9682), .B(n7385), .ZN(n7567)
         );
  NOR2_X1 U9223 ( .A1(n4752), .A2(n9629), .ZN(n7389) );
  OAI22_X1 U9224 ( .A1(n9633), .A2(n7387), .B1(n7544), .B2(n9630), .ZN(n7388)
         );
  AOI211_X1 U9225 ( .C1(n7567), .C2(n9616), .A(n7389), .B(n7388), .ZN(n7396)
         );
  INV_X1 U9226 ( .A(n7390), .ZN(n8234) );
  XNOR2_X1 U9227 ( .A(n7391), .B(n8234), .ZN(n7392) );
  NAND2_X1 U9228 ( .A1(n7392), .A2(n9640), .ZN(n7394) );
  AOI22_X1 U9229 ( .A1(n9290), .A2(n9643), .B1(n9644), .B2(n7943), .ZN(n7393)
         );
  NAND2_X1 U9230 ( .A1(n7394), .A2(n7393), .ZN(n7566) );
  NAND2_X1 U9231 ( .A1(n7566), .A2(n9633), .ZN(n7395) );
  OAI211_X1 U9232 ( .C1(n7397), .C2(n9650), .A(n7396), .B(n7395), .ZN(P1_U3280) );
  INV_X1 U9233 ( .A(n9726), .ZN(n9975) );
  OAI211_X1 U9234 ( .C1(n7400), .C2(n9975), .A(n7399), .B(n7398), .ZN(n7401)
         );
  AOI21_X1 U9235 ( .B1(n7402), .B2(n9978), .A(n7401), .ZN(n7405) );
  NAND2_X1 U9236 ( .A1(n9986), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7403) );
  OAI21_X1 U9237 ( .B1(n7405), .B2(n9986), .A(n7403), .ZN(P1_U3534) );
  NAND2_X1 U9238 ( .A1(n9980), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7404) );
  OAI21_X1 U9239 ( .B1(n7405), .B2(n9980), .A(n7404), .ZN(P1_U3489) );
  INV_X1 U9240 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7436) );
  MUX2_X1 U9241 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8799), .Z(n7408) );
  XNOR2_X1 U9242 ( .A(n7408), .B(n10015), .ZN(n10006) );
  MUX2_X1 U9243 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8799), .Z(n7438) );
  XOR2_X1 U9244 ( .A(n7441), .B(n7438), .Z(n7409) );
  OAI21_X1 U9245 ( .B1(n7410), .B2(n7409), .A(n7437), .ZN(n7411) );
  NAND2_X1 U9246 ( .A1(n7411), .A2(n10115), .ZN(n7435) );
  MUX2_X1 U9247 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7412), .S(n7441), .Z(n7421)
         );
  NAND2_X1 U9248 ( .A1(n7413), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7414) );
  INV_X1 U9249 ( .A(n10015), .ZN(n7416) );
  XNOR2_X1 U9250 ( .A(n7417), .B(n7416), .ZN(n10007) );
  NAND2_X1 U9251 ( .A1(n10007), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7419) );
  NAND2_X1 U9252 ( .A1(n7417), .A2(n10015), .ZN(n7418) );
  NAND2_X1 U9253 ( .A1(n7419), .A2(n7418), .ZN(n7420) );
  NAND2_X1 U9254 ( .A1(n7420), .A2(n7421), .ZN(n7440) );
  OAI21_X1 U9255 ( .B1(n7421), .B2(n7420), .A(n7440), .ZN(n7433) );
  INV_X1 U9256 ( .A(n10107), .ZN(n10027) );
  INV_X1 U9257 ( .A(n7422), .ZN(n7423) );
  OAI21_X1 U9258 ( .B1(n10027), .B2(n7441), .A(n7423), .ZN(n7432) );
  NAND2_X1 U9259 ( .A1(n7425), .A2(n7424), .ZN(n7426) );
  NAND2_X1 U9260 ( .A1(n7426), .A2(n10015), .ZN(n7429) );
  MUX2_X1 U9261 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6037), .S(n7441), .Z(n7428)
         );
  NAND3_X1 U9262 ( .A1(n10008), .A2(n4738), .A3(n7429), .ZN(n7430) );
  AOI21_X1 U9263 ( .B1(n7443), .B2(n7430), .A(n10122), .ZN(n7431) );
  AOI211_X1 U9264 ( .C1(n10116), .C2(n7433), .A(n7432), .B(n7431), .ZN(n7434)
         );
  OAI211_X1 U9265 ( .C1(n10020), .C2(n7436), .A(n7435), .B(n7434), .ZN(
        P2_U3188) );
  MUX2_X1 U9266 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8799), .Z(n7728) );
  XOR2_X1 U9267 ( .A(n7743), .B(n7728), .Z(n7731) );
  OAI21_X1 U9268 ( .B1(n7438), .B2(n7441), .A(n7437), .ZN(n7732) );
  XOR2_X1 U9269 ( .A(n7731), .B(n7732), .Z(n7455) );
  NAND2_X1 U9270 ( .A1(n7441), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7439) );
  INV_X1 U9271 ( .A(n7743), .ZN(n7730) );
  XNOR2_X1 U9272 ( .A(n7744), .B(n7730), .ZN(n7742) );
  XNOR2_X1 U9273 ( .A(n7742), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7453) );
  INV_X1 U9274 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7451) );
  NAND2_X1 U9275 ( .A1(n7441), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9276 ( .A1(n7443), .A2(n7442), .ZN(n7445) );
  INV_X1 U9277 ( .A(n7445), .ZN(n7444) );
  OAI21_X1 U9278 ( .B1(n7446), .B2(P2_REG2_REG_7__SCAN_IN), .A(n10031), .ZN(
        n7447) );
  NAND2_X1 U9279 ( .A1(n10010), .A2(n7447), .ZN(n7450) );
  NOR2_X1 U9280 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7448), .ZN(n7508) );
  AOI21_X1 U9281 ( .B1(n10107), .B2(n7730), .A(n7508), .ZN(n7449) );
  OAI211_X1 U9282 ( .C1(n10020), .C2(n7451), .A(n7450), .B(n7449), .ZN(n7452)
         );
  AOI21_X1 U9283 ( .B1(n10116), .B2(n7453), .A(n7452), .ZN(n7454) );
  OAI21_X1 U9284 ( .B1(n7455), .B2(n10004), .A(n7454), .ZN(P2_U3189) );
  INV_X1 U9285 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7462) );
  AND2_X1 U9286 ( .A1(n7457), .A2(n7456), .ZN(n7458) );
  OAI22_X1 U9287 ( .A1(n10115), .A2(n7459), .B1(n7478), .B2(n7458), .ZN(n7461)
         );
  AOI22_X1 U9288 ( .A1(n10107), .A2(P2_IR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n7460) );
  OAI211_X1 U9289 ( .C1(n7462), .C2(n10020), .A(n7461), .B(n7460), .ZN(
        P2_U3182) );
  INV_X1 U9290 ( .A(n7628), .ZN(n7714) );
  AOI21_X1 U9291 ( .B1(n7463), .B2(n8594), .A(n4451), .ZN(n10148) );
  INV_X1 U9292 ( .A(n10148), .ZN(n7471) );
  INV_X1 U9293 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7464) );
  OAI22_X1 U9294 ( .A1(n8855), .A2(n10147), .B1(n8977), .B2(n7464), .ZN(n7470)
         );
  AOI22_X1 U9295 ( .A1(n10129), .A2(n8784), .B1(n8782), .B2(n10131), .ZN(n7468) );
  OAI21_X1 U9296 ( .B1(n7465), .B2(n7463), .A(n7239), .ZN(n7466) );
  NAND2_X1 U9297 ( .A1(n7466), .A2(n10134), .ZN(n7467) );
  OAI211_X1 U9298 ( .C1(n10148), .C2(n7622), .A(n7468), .B(n7467), .ZN(n10150)
         );
  MUX2_X1 U9299 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10150), .S(n10145), .Z(n7469) );
  AOI211_X1 U9300 ( .C1(n7714), .C2(n7471), .A(n7470), .B(n7469), .ZN(n7472)
         );
  INV_X1 U9301 ( .A(n7472), .ZN(P2_U3232) );
  NAND2_X1 U9302 ( .A1(n7474), .A2(n7473), .ZN(n7475) );
  AOI21_X1 U9303 ( .B1(n7476), .B2(n7475), .A(n10122), .ZN(n7481) );
  AOI211_X1 U9304 ( .C1(n7479), .C2(n7478), .A(n7477), .B(n10004), .ZN(n7480)
         );
  AOI211_X1 U9305 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3151), .A(n7481), .B(
        n7480), .ZN(n7486) );
  XNOR2_X1 U9306 ( .A(n7482), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7484) );
  AOI22_X1 U9307 ( .A1(n10116), .A2(n7484), .B1(n10107), .B2(n5987), .ZN(n7485) );
  OAI211_X1 U9308 ( .C1(n10230), .C2(n10020), .A(n7486), .B(n7485), .ZN(
        P2_U3183) );
  INV_X1 U9309 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7503) );
  NOR2_X1 U9310 ( .A1(n10027), .A2(n7487), .ZN(n7492) );
  AOI211_X1 U9311 ( .C1(n7490), .C2(n7489), .A(n10004), .B(n7488), .ZN(n7491)
         );
  AOI211_X1 U9312 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(P2_U3151), .A(n7492), .B(
        n7491), .ZN(n7502) );
  OAI21_X1 U9313 ( .B1(n7495), .B2(n7494), .A(n7493), .ZN(n7500) );
  OAI21_X1 U9314 ( .B1(n7498), .B2(n7497), .A(n7496), .ZN(n7499) );
  AOI22_X1 U9315 ( .A1(n10116), .A2(n7500), .B1(n10010), .B2(n7499), .ZN(n7501) );
  OAI211_X1 U9316 ( .C1(n10020), .C2(n7503), .A(n7502), .B(n7501), .ZN(
        P2_U3184) );
  AOI21_X1 U9317 ( .B1(n7506), .B2(n7505), .A(n7504), .ZN(n7514) );
  INV_X1 U9318 ( .A(n7507), .ZN(n7536) );
  NAND2_X1 U9319 ( .A1(n8478), .A2(n7537), .ZN(n7510) );
  AOI21_X1 U9320 ( .B1(n8527), .B2(n8781), .A(n7508), .ZN(n7509) );
  OAI211_X1 U9321 ( .C1(n7511), .C2(n8523), .A(n7510), .B(n7509), .ZN(n7512)
         );
  AOI21_X1 U9322 ( .B1(n7536), .B2(n8514), .A(n7512), .ZN(n7513) );
  OAI21_X1 U9323 ( .B1(n7514), .B2(n8518), .A(n7513), .ZN(P2_U3153) );
  NAND2_X1 U9324 ( .A1(n7515), .A2(n7516), .ZN(n7517) );
  XNOR2_X1 U9325 ( .A(n7517), .B(n8571), .ZN(n10185) );
  INV_X1 U9326 ( .A(n10185), .ZN(n7528) );
  OR2_X1 U9327 ( .A1(n7518), .A2(n8635), .ZN(n7529) );
  NAND2_X1 U9328 ( .A1(n7529), .A2(n7519), .ZN(n7617) );
  NAND2_X1 U9329 ( .A1(n7617), .A2(n10134), .ZN(n7523) );
  AOI21_X1 U9330 ( .B1(n7529), .B2(n7520), .A(n8571), .ZN(n7522) );
  AOI22_X1 U9331 ( .A1(n7634), .A2(n10129), .B1(n10131), .B2(n8779), .ZN(n7521) );
  OAI21_X1 U9332 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n10183) );
  NOR2_X1 U9333 ( .A1(n10145), .A2(n7524), .ZN(n7526) );
  OAI22_X1 U9334 ( .A1(n8855), .A2(n10182), .B1(n7631), .B2(n8977), .ZN(n7525)
         );
  AOI211_X1 U9335 ( .C1(n10183), .C2(n10145), .A(n7526), .B(n7525), .ZN(n7527)
         );
  OAI21_X1 U9336 ( .B1(n7528), .B2(n9026), .A(n7527), .ZN(P2_U3225) );
  INV_X1 U9337 ( .A(n7529), .ZN(n7530) );
  AOI21_X1 U9338 ( .B1(n8635), .B2(n7518), .A(n7530), .ZN(n7535) );
  INV_X1 U9339 ( .A(n10134), .ZN(n8972) );
  AOI22_X1 U9340 ( .A1(n10129), .A2(n8781), .B1(n8780), .B2(n10131), .ZN(n7534) );
  OR2_X1 U9341 ( .A1(n7531), .A2(n8635), .ZN(n7532) );
  AND2_X1 U9342 ( .A1(n7515), .A2(n7532), .ZN(n10177) );
  INV_X1 U9343 ( .A(n7622), .ZN(n7710) );
  NAND2_X1 U9344 ( .A1(n10177), .A2(n7710), .ZN(n7533) );
  OAI211_X1 U9345 ( .C1(n7535), .C2(n8972), .A(n7534), .B(n7533), .ZN(n10181)
         );
  INV_X1 U9346 ( .A(n10181), .ZN(n7541) );
  AOI22_X1 U9347 ( .A1(n10138), .A2(n7537), .B1(n10140), .B2(n7536), .ZN(n7538) );
  OAI21_X1 U9348 ( .B1(n6051), .B2(n10145), .A(n7538), .ZN(n7539) );
  AOI21_X1 U9349 ( .B1(n10177), .B2(n7714), .A(n7539), .ZN(n7540) );
  OAI21_X1 U9350 ( .B1(n7541), .B2(n10146), .A(n7540), .ZN(P2_U3226) );
  XOR2_X1 U9351 ( .A(n7542), .B(n7543), .Z(n7551) );
  NOR2_X1 U9352 ( .A1(n9260), .A2(n7544), .ZN(n7548) );
  NAND2_X1 U9353 ( .A1(n9250), .A2(n7943), .ZN(n7545) );
  NAND2_X1 U9354 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9880) );
  OAI211_X1 U9355 ( .C1(n9252), .C2(n7546), .A(n7545), .B(n9880), .ZN(n7547)
         );
  AOI211_X1 U9356 ( .C1(n7549), .C2(n9265), .A(n7548), .B(n7547), .ZN(n7550)
         );
  OAI21_X1 U9357 ( .B1(n7551), .B2(n9267), .A(n7550), .ZN(P1_U3234) );
  INV_X1 U9358 ( .A(n7552), .ZN(n7554) );
  INV_X1 U9359 ( .A(n7553), .ZN(n8361) );
  OAI222_X1 U9360 ( .A1(n9775), .A2(n7555), .B1(n7554), .B2(P1_U3086), .C1(
        n8017), .C2(n8361), .ZN(P1_U3331) );
  XNOR2_X1 U9361 ( .A(n7556), .B(n8235), .ZN(n9729) );
  XOR2_X1 U9362 ( .A(n8235), .B(n7557), .Z(n7558) );
  OAI222_X1 U9363 ( .A1(n9551), .A2(n9218), .B1(n9549), .B2(n7559), .C1(n7558), 
        .C2(n9546), .ZN(n9723) );
  INV_X1 U9364 ( .A(n9725), .ZN(n7777) );
  AOI211_X1 U9365 ( .C1(n9725), .C2(n7560), .A(n9682), .B(n7643), .ZN(n9724)
         );
  NAND2_X1 U9366 ( .A1(n9724), .A2(n9616), .ZN(n7563) );
  INV_X1 U9367 ( .A(n7561), .ZN(n7774) );
  AOI22_X1 U9368 ( .A1(n9469), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7774), .B2(
        n9617), .ZN(n7562) );
  OAI211_X1 U9369 ( .C1(n7777), .C2(n9629), .A(n7563), .B(n7562), .ZN(n7564)
         );
  AOI21_X1 U9370 ( .B1(n9723), .B2(n9633), .A(n7564), .ZN(n7565) );
  OAI21_X1 U9371 ( .B1(n9729), .B2(n9650), .A(n7565), .ZN(P1_U3279) );
  AOI211_X1 U9372 ( .C1(n7568), .C2(n9978), .A(n7567), .B(n7566), .ZN(n7571)
         );
  MUX2_X1 U9373 ( .A(n7569), .B(n7571), .S(n9981), .Z(n7570) );
  OAI21_X1 U9374 ( .B1(n4752), .B2(n9770), .A(n7570), .ZN(P1_U3492) );
  MUX2_X1 U9375 ( .A(n7572), .B(n7571), .S(n9988), .Z(n7573) );
  OAI21_X1 U9376 ( .B1(n4752), .B2(n9717), .A(n7573), .ZN(P1_U3535) );
  NAND2_X1 U9377 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9832) );
  INV_X1 U9378 ( .A(n9832), .ZN(n7574) );
  AOI21_X1 U9379 ( .B1(n9292), .B2(n9250), .A(n7574), .ZN(n7576) );
  NAND2_X1 U9380 ( .A1(n9294), .A2(n9277), .ZN(n7575) );
  OAI211_X1 U9381 ( .C1(n9260), .C2(n7577), .A(n7576), .B(n7575), .ZN(n7587)
         );
  OAI21_X1 U9382 ( .B1(n7580), .B2(n7579), .A(n7578), .ZN(n7584) );
  XNOR2_X1 U9383 ( .A(n7582), .B(n7581), .ZN(n7583) );
  XNOR2_X1 U9384 ( .A(n7584), .B(n7583), .ZN(n7585) );
  NOR2_X1 U9385 ( .A1(n7585), .A2(n9267), .ZN(n7586) );
  AOI211_X1 U9386 ( .C1(n9968), .C2(n9265), .A(n7587), .B(n7586), .ZN(n7588)
         );
  INV_X1 U9387 ( .A(n7588), .ZN(P1_U3231) );
  OAI21_X1 U9388 ( .B1(n7589), .B2(n8566), .A(n7590), .ZN(n10169) );
  OAI22_X1 U9389 ( .A1(n8855), .A2(n10166), .B1(n8977), .B2(n7591), .ZN(n7597)
         );
  INV_X1 U9390 ( .A(n10129), .ZN(n8974) );
  XNOR2_X1 U9391 ( .A(n7592), .B(n8566), .ZN(n7593) );
  OAI222_X1 U9392 ( .A1(n8976), .A2(n7595), .B1(n8974), .B2(n7594), .C1(n8972), 
        .C2(n7593), .ZN(n10167) );
  MUX2_X1 U9393 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10167), .S(n10145), .Z(n7596) );
  AOI211_X1 U9394 ( .C1(n10169), .C2(n10142), .A(n7597), .B(n7596), .ZN(n7598)
         );
  INV_X1 U9395 ( .A(n7598), .ZN(P2_U3228) );
  XNOR2_X1 U9396 ( .A(n7599), .B(n7600), .ZN(n7675) );
  NOR2_X1 U9397 ( .A1(n7675), .A2(n7674), .ZN(n7673) );
  AOI21_X1 U9398 ( .B1(n7600), .B2(n7599), .A(n7673), .ZN(n7604) );
  XNOR2_X1 U9399 ( .A(n7602), .B(n7601), .ZN(n7603) );
  XNOR2_X1 U9400 ( .A(n7604), .B(n7603), .ZN(n7612) );
  NAND2_X1 U9401 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9849) );
  OAI21_X1 U9402 ( .B1(n9252), .B2(n7605), .A(n9849), .ZN(n7606) );
  AOI21_X1 U9403 ( .B1(n9250), .B2(n9290), .A(n7606), .ZN(n7607) );
  OAI21_X1 U9404 ( .B1(n9260), .B2(n7608), .A(n7607), .ZN(n7609) );
  AOI21_X1 U9405 ( .B1(n7610), .B2(n9265), .A(n7609), .ZN(n7611) );
  OAI21_X1 U9406 ( .B1(n7612), .B2(n9267), .A(n7611), .ZN(P1_U3236) );
  NAND2_X1 U9407 ( .A1(n7613), .A2(n8570), .ZN(n7614) );
  NAND2_X1 U9408 ( .A1(n7696), .A2(n7614), .ZN(n10188) );
  AOI22_X1 U9409 ( .A1(n10129), .A2(n8780), .B1(n8778), .B2(n10131), .ZN(n7621) );
  NAND2_X1 U9410 ( .A1(n7617), .A2(n7615), .ZN(n7703) );
  INV_X1 U9411 ( .A(n7703), .ZN(n7619) );
  AOI21_X1 U9412 ( .B1(n7617), .B2(n7616), .A(n8570), .ZN(n7618) );
  OAI21_X1 U9413 ( .B1(n7619), .B2(n7618), .A(n10134), .ZN(n7620) );
  OAI211_X1 U9414 ( .C1(n10188), .C2(n7622), .A(n7621), .B(n7620), .ZN(n10190)
         );
  NAND2_X1 U9415 ( .A1(n10190), .A2(n10145), .ZN(n7627) );
  INV_X1 U9416 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7624) );
  INV_X1 U9417 ( .A(n7914), .ZN(n7623) );
  OAI22_X1 U9418 ( .A1(n10145), .A2(n7624), .B1(n7623), .B2(n8977), .ZN(n7625)
         );
  AOI21_X1 U9419 ( .B1(n10138), .B2(n7904), .A(n7625), .ZN(n7626) );
  OAI211_X1 U9420 ( .C1(n10188), .C2(n7628), .A(n7627), .B(n7626), .ZN(
        P2_U3224) );
  XOR2_X1 U9421 ( .A(n7630), .B(n7629), .Z(n7641) );
  INV_X1 U9422 ( .A(n7631), .ZN(n7639) );
  NAND2_X1 U9423 ( .A1(n8478), .A2(n7632), .ZN(n7636) );
  NOR2_X1 U9424 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7633), .ZN(n10024) );
  AOI21_X1 U9425 ( .B1(n8527), .B2(n7634), .A(n10024), .ZN(n7635) );
  OAI211_X1 U9426 ( .C1(n7637), .C2(n8523), .A(n7636), .B(n7635), .ZN(n7638)
         );
  AOI21_X1 U9427 ( .B1(n7639), .B2(n8514), .A(n7638), .ZN(n7640) );
  OAI21_X1 U9428 ( .B1(n7641), .B2(n8518), .A(n7640), .ZN(P2_U3161) );
  XNOR2_X1 U9429 ( .A(n7642), .B(n8237), .ZN(n7783) );
  INV_X1 U9430 ( .A(n7783), .ZN(n7653) );
  INV_X1 U9431 ( .A(n7643), .ZN(n7645) );
  INV_X1 U9432 ( .A(n7682), .ZN(n7644) );
  AOI211_X1 U9433 ( .C1(n7947), .C2(n7645), .A(n9682), .B(n7644), .ZN(n7782)
         );
  NOR2_X1 U9434 ( .A1(n7788), .A2(n9629), .ZN(n7648) );
  OAI22_X1 U9435 ( .A1(n9633), .A2(n7646), .B1(n7945), .B2(n9630), .ZN(n7647)
         );
  AOI211_X1 U9436 ( .C1(n7782), .C2(n9616), .A(n7648), .B(n7647), .ZN(n7652)
         );
  OAI211_X1 U9437 ( .C1(n4433), .C2(n4804), .A(n9640), .B(n7687), .ZN(n7650)
         );
  AOI22_X1 U9438 ( .A1(n7831), .A2(n9644), .B1(n9643), .B2(n7943), .ZN(n7649)
         );
  NAND2_X1 U9439 ( .A1(n7650), .A2(n7649), .ZN(n7781) );
  NAND2_X1 U9440 ( .A1(n7781), .A2(n9633), .ZN(n7651) );
  OAI211_X1 U9441 ( .C1(n7653), .C2(n9650), .A(n7652), .B(n7651), .ZN(P1_U3278) );
  INV_X1 U9442 ( .A(n8568), .ZN(n7659) );
  XNOR2_X1 U9443 ( .A(n7654), .B(n7659), .ZN(n7658) );
  NAND2_X1 U9444 ( .A1(n10132), .A2(n10129), .ZN(n7655) );
  OAI21_X1 U9445 ( .B1(n7656), .B2(n8976), .A(n7655), .ZN(n7657) );
  AOI21_X1 U9446 ( .B1(n7658), .B2(n10134), .A(n7657), .ZN(n10174) );
  XNOR2_X1 U9447 ( .A(n7660), .B(n7659), .ZN(n10171) );
  NOR2_X1 U9448 ( .A1(n10145), .A2(n6037), .ZN(n7664) );
  OAI22_X1 U9449 ( .A1(n8855), .A2(n7662), .B1(n7661), .B2(n8977), .ZN(n7663)
         );
  AOI211_X1 U9450 ( .C1(n10171), .C2(n10142), .A(n7664), .B(n7663), .ZN(n7665)
         );
  OAI21_X1 U9451 ( .B1(n10146), .B2(n10174), .A(n7665), .ZN(P2_U3227) );
  INV_X1 U9452 ( .A(n7666), .ZN(n8357) );
  OAI222_X1 U9453 ( .A1(n9775), .A2(n7668), .B1(n7667), .B2(P1_U3086), .C1(
        n8017), .C2(n8357), .ZN(P1_U3330) );
  NAND2_X1 U9454 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9815) );
  INV_X1 U9455 ( .A(n9815), .ZN(n7669) );
  AOI21_X1 U9456 ( .B1(n9291), .B2(n9250), .A(n7669), .ZN(n7671) );
  NAND2_X1 U9457 ( .A1(n9293), .A2(n9277), .ZN(n7670) );
  OAI211_X1 U9458 ( .C1(n9260), .C2(n7672), .A(n7671), .B(n7670), .ZN(n7678)
         );
  AOI21_X1 U9459 ( .B1(n7675), .B2(n7674), .A(n7673), .ZN(n7676) );
  NOR2_X1 U9460 ( .A1(n7676), .A2(n9267), .ZN(n7677) );
  AOI211_X1 U9461 ( .C1(n7679), .C2(n9265), .A(n7678), .B(n7677), .ZN(n7680)
         );
  INV_X1 U9462 ( .A(n7680), .ZN(P1_U3217) );
  XNOR2_X1 U9463 ( .A(n7681), .B(n7688), .ZN(n9722) );
  AOI211_X1 U9464 ( .C1(n9720), .C2(n7682), .A(n9682), .B(n5884), .ZN(n9719)
         );
  INV_X1 U9465 ( .A(n9720), .ZN(n7684) );
  OAI22_X1 U9466 ( .A1(n7684), .A2(n9629), .B1(n7683), .B2(n9633), .ZN(n7685)
         );
  AOI21_X1 U9467 ( .B1(n9719), .B2(n9616), .A(n7685), .ZN(n7695) );
  NAND2_X1 U9468 ( .A1(n7687), .A2(n7686), .ZN(n7689) );
  INV_X1 U9469 ( .A(n7688), .ZN(n8239) );
  XNOR2_X1 U9470 ( .A(n7689), .B(n8239), .ZN(n7690) );
  OAI222_X1 U9471 ( .A1(n9549), .A2(n9218), .B1(n9551), .B2(n7691), .C1(n9546), 
        .C2(n7690), .ZN(n9718) );
  NOR2_X1 U9472 ( .A1(n9630), .A2(n9216), .ZN(n7693) );
  OAI21_X1 U9473 ( .B1(n9718), .B2(n7693), .A(n7692), .ZN(n7694) );
  OAI211_X1 U9474 ( .C1(n9722), .C2(n9650), .A(n7695), .B(n7694), .ZN(P1_U3277) );
  NAND2_X1 U9475 ( .A1(n7696), .A2(n8632), .ZN(n7697) );
  XNOR2_X1 U9476 ( .A(n7697), .B(n8574), .ZN(n10194) );
  OR2_X1 U9477 ( .A1(n7518), .A2(n7698), .ZN(n7699) );
  AND2_X1 U9478 ( .A1(n7700), .A2(n7699), .ZN(n7705) );
  INV_X1 U9479 ( .A(n8574), .ZN(n7702) );
  NAND3_X1 U9480 ( .A1(n7703), .A2(n7702), .A3(n7701), .ZN(n7704) );
  NAND2_X1 U9481 ( .A1(n7705), .A2(n7704), .ZN(n7706) );
  NAND2_X1 U9482 ( .A1(n7706), .A2(n10134), .ZN(n7708) );
  AOI22_X1 U9483 ( .A1(n10129), .A2(n8779), .B1(n8777), .B2(n10131), .ZN(n7707) );
  NAND2_X1 U9484 ( .A1(n7708), .A2(n7707), .ZN(n7709) );
  AOI21_X1 U9485 ( .B1(n10194), .B2(n7710), .A(n7709), .ZN(n10196) );
  NOR2_X1 U9486 ( .A1(n8855), .A2(n7711), .ZN(n7713) );
  OAI22_X1 U9487 ( .A1(n10145), .A2(n7736), .B1(n7846), .B2(n8977), .ZN(n7712)
         );
  AOI211_X1 U9488 ( .C1(n10194), .C2(n7714), .A(n7713), .B(n7712), .ZN(n7715)
         );
  OAI21_X1 U9489 ( .B1(n10196), .B2(n10146), .A(n7715), .ZN(P2_U3223) );
  XNOR2_X1 U9490 ( .A(n7716), .B(n8575), .ZN(n7718) );
  OAI22_X1 U9491 ( .A1(n7908), .A2(n8974), .B1(n8662), .B2(n8976), .ZN(n7717)
         );
  AOI21_X1 U9492 ( .B1(n7718), .B2(n10134), .A(n7717), .ZN(n10203) );
  XNOR2_X1 U9493 ( .A(n7719), .B(n8575), .ZN(n10199) );
  INV_X1 U9494 ( .A(n10201), .ZN(n7903) );
  NOR2_X1 U9495 ( .A1(n8855), .A2(n7903), .ZN(n7721) );
  INV_X1 U9496 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7882) );
  OAI22_X1 U9497 ( .A1(n10145), .A2(n7882), .B1(n7896), .B2(n8977), .ZN(n7720)
         );
  AOI211_X1 U9498 ( .C1(n10199), .C2(n10142), .A(n7721), .B(n7720), .ZN(n7722)
         );
  OAI21_X1 U9499 ( .B1(n10146), .B2(n10203), .A(n7722), .ZN(P2_U3222) );
  MUX2_X1 U9500 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7524), .S(n10026), .Z(n10028) );
  NAND2_X1 U9501 ( .A1(n10026), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7724) );
  NOR2_X1 U9502 ( .A1(n7725), .A2(n7792), .ZN(n7727) );
  AOI22_X1 U9503 ( .A1(n7875), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7736), .B2(
        n7880), .ZN(n7726) );
  NOR2_X1 U9504 ( .A1(n7727), .A2(n7726), .ZN(n7879) );
  AOI21_X1 U9505 ( .B1(n7727), .B2(n7726), .A(n7879), .ZN(n7761) );
  INV_X1 U9506 ( .A(n7728), .ZN(n7729) );
  MUX2_X1 U9507 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8799), .Z(n7733) );
  XNOR2_X1 U9508 ( .A(n7733), .B(n10026), .ZN(n10037) );
  INV_X1 U9509 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10219) );
  MUX2_X1 U9510 ( .A(n7624), .B(n10219), .S(n8799), .Z(n7734) );
  OR2_X1 U9511 ( .A1(n7734), .A2(n7796), .ZN(n7802) );
  NAND2_X1 U9512 ( .A1(n7734), .A2(n7796), .ZN(n7804) );
  MUX2_X1 U9513 ( .A(n7736), .B(n7735), .S(n8799), .Z(n7737) );
  NAND2_X1 U9514 ( .A1(n7737), .A2(n7875), .ZN(n7869) );
  INV_X1 U9515 ( .A(n7737), .ZN(n7738) );
  NAND2_X1 U9516 ( .A1(n7738), .A2(n7880), .ZN(n7739) );
  NAND2_X1 U9517 ( .A1(n7869), .A2(n7739), .ZN(n7740) );
  AND3_X1 U9518 ( .A1(n7800), .A2(n7804), .A3(n7740), .ZN(n7741) );
  OAI21_X1 U9519 ( .B1(n7871), .B2(n7741), .A(n10115), .ZN(n7760) );
  AOI22_X1 U9520 ( .A1(n7875), .A2(n7735), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7880), .ZN(n7753) );
  NAND2_X1 U9521 ( .A1(n7742), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U9522 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  NAND2_X1 U9523 ( .A1(n7746), .A2(n7745), .ZN(n10022) );
  INV_X1 U9524 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7747) );
  MUX2_X1 U9525 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7747), .S(n10026), .Z(n10023) );
  NAND2_X1 U9526 ( .A1(n10022), .A2(n10023), .ZN(n10021) );
  NAND2_X1 U9527 ( .A1(n10026), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U9528 ( .A1(n7750), .A2(n7749), .ZN(n7751) );
  XNOR2_X1 U9529 ( .A(n7750), .B(n7796), .ZN(n7790) );
  NAND2_X1 U9530 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n7790), .ZN(n7789) );
  OAI21_X1 U9531 ( .B1(n7753), .B2(n7752), .A(n7874), .ZN(n7758) );
  INV_X1 U9532 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7756) );
  NOR2_X1 U9533 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7754), .ZN(n7843) );
  AOI21_X1 U9534 ( .B1(n10107), .B2(n7875), .A(n7843), .ZN(n7755) );
  OAI21_X1 U9535 ( .B1(n10020), .B2(n7756), .A(n7755), .ZN(n7757) );
  AOI21_X1 U9536 ( .B1(n7758), .B2(n10116), .A(n7757), .ZN(n7759) );
  OAI211_X1 U9537 ( .C1(n7761), .C2(n10122), .A(n7760), .B(n7759), .ZN(
        P2_U3192) );
  INV_X1 U9538 ( .A(n7762), .ZN(n7765) );
  OAI222_X1 U9539 ( .A1(n7764), .A2(P2_U3151), .B1(n9175), .B2(n7765), .C1(
        n7763), .C2(n9172), .ZN(P2_U3269) );
  INV_X1 U9540 ( .A(n5779), .ZN(n7766) );
  OAI222_X1 U9541 ( .A1(n9775), .A2(n7767), .B1(n7766), .B2(P1_U3086), .C1(
        n8017), .C2(n7765), .ZN(P1_U3329) );
  OAI21_X1 U9542 ( .B1(n7770), .B2(n7768), .A(n7769), .ZN(n7771) );
  NAND2_X1 U9543 ( .A1(n7771), .A2(n9274), .ZN(n7776) );
  NAND2_X1 U9544 ( .A1(n9289), .A2(n9277), .ZN(n7772) );
  NAND2_X1 U9545 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9896) );
  OAI211_X1 U9546 ( .C1(n9279), .C2(n9218), .A(n7772), .B(n9896), .ZN(n7773)
         );
  AOI21_X1 U9547 ( .B1(n7774), .B2(n9282), .A(n7773), .ZN(n7775) );
  OAI211_X1 U9548 ( .C1(n7777), .C2(n9285), .A(n7776), .B(n7775), .ZN(P1_U3215) );
  INV_X1 U9549 ( .A(n7778), .ZN(n8331) );
  AOI21_X1 U9550 ( .B1(n9169), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7779), .ZN(
        n7780) );
  OAI21_X1 U9551 ( .B1(n8331), .B2(n9175), .A(n7780), .ZN(P2_U3268) );
  AOI211_X1 U9552 ( .C1(n7783), .C2(n9978), .A(n7782), .B(n7781), .ZN(n7786)
         );
  MUX2_X1 U9553 ( .A(n7784), .B(n7786), .S(n9981), .Z(n7785) );
  OAI21_X1 U9554 ( .B1(n7788), .B2(n9770), .A(n7785), .ZN(P1_U3498) );
  MUX2_X1 U9555 ( .A(n9901), .B(n7786), .S(n9988), .Z(n7787) );
  OAI21_X1 U9556 ( .B1(n7788), .B2(n9717), .A(n7787), .ZN(P1_U3537) );
  OAI21_X1 U9557 ( .B1(n7790), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7789), .ZN(
        n7809) );
  INV_X1 U9558 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U9559 ( .A1(n7791), .A2(n7624), .ZN(n7794) );
  INV_X1 U9560 ( .A(n7792), .ZN(n7793) );
  NAND2_X1 U9561 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  NAND2_X1 U9562 ( .A1(n10010), .A2(n7795), .ZN(n7798) );
  NOR2_X1 U9563 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6070), .ZN(n7905) );
  AOI21_X1 U9564 ( .B1(n10107), .B2(n7796), .A(n7905), .ZN(n7797) );
  OAI211_X1 U9565 ( .C1(n10020), .C2(n7799), .A(n7798), .B(n7797), .ZN(n7808)
         );
  INV_X1 U9566 ( .A(n7800), .ZN(n7805) );
  AOI21_X1 U9567 ( .B1(n7802), .B2(n7804), .A(n7801), .ZN(n7803) );
  AOI21_X1 U9568 ( .B1(n7805), .B2(n7804), .A(n7803), .ZN(n7806) );
  NOR2_X1 U9569 ( .A1(n7806), .A2(n10004), .ZN(n7807) );
  AOI211_X1 U9570 ( .C1(n10116), .C2(n7809), .A(n7808), .B(n7807), .ZN(n7810)
         );
  INV_X1 U9571 ( .A(n7810), .ZN(P2_U3191) );
  AOI21_X1 U9572 ( .B1(n8660), .B2(n7811), .A(n4447), .ZN(n7818) );
  NAND2_X1 U9573 ( .A1(n10225), .A2(n10198), .ZN(n9078) );
  INV_X1 U9574 ( .A(n9078), .ZN(n8000) );
  AOI22_X1 U9575 ( .A1(n7818), .A2(n8000), .B1(n9075), .B2(n8663), .ZN(n7817)
         );
  NOR2_X1 U9576 ( .A1(n4440), .A2(n8660), .ZN(n7813) );
  OR3_X1 U9577 ( .A1(n7813), .A2(n7812), .A3(n8972), .ZN(n7815) );
  AOI22_X1 U9578 ( .A1(n10131), .A2(n8775), .B1(n8777), .B2(n10129), .ZN(n7814) );
  NAND2_X1 U9579 ( .A1(n7815), .A2(n7814), .ZN(n7890) );
  INV_X1 U9580 ( .A(n7890), .ZN(n7820) );
  MUX2_X1 U9581 ( .A(n7980), .B(n7820), .S(n10225), .Z(n7816) );
  NAND2_X1 U9582 ( .A1(n7817), .A2(n7816), .ZN(P2_U3471) );
  INV_X1 U9583 ( .A(n7818), .ZN(n7889) );
  INV_X1 U9584 ( .A(n7819), .ZN(n7963) );
  AOI22_X1 U9585 ( .A1(n10138), .A2(n8663), .B1(n10140), .B2(n7963), .ZN(n7822) );
  MUX2_X1 U9586 ( .A(n7820), .B(n7976), .S(n10146), .Z(n7821) );
  OAI211_X1 U9587 ( .C1(n7889), .C2(n9026), .A(n7822), .B(n7821), .ZN(P2_U3221) );
  XOR2_X1 U9588 ( .A(n7823), .B(n7828), .Z(n9714) );
  INV_X1 U9589 ( .A(n9714), .ZN(n7837) );
  AOI211_X1 U9590 ( .C1(n7866), .C2(n7824), .A(n9682), .B(n7930), .ZN(n9713)
         );
  INV_X1 U9591 ( .A(n7866), .ZN(n9771) );
  NOR2_X1 U9592 ( .A1(n9771), .A2(n9629), .ZN(n7826) );
  OAI22_X1 U9593 ( .A1(n9633), .A2(n9427), .B1(n7864), .B2(n9630), .ZN(n7825)
         );
  AOI211_X1 U9594 ( .C1(n9713), .C2(n9616), .A(n7826), .B(n7825), .ZN(n7836)
         );
  NAND2_X1 U9595 ( .A1(n7827), .A2(n9640), .ZN(n7834) );
  INV_X1 U9596 ( .A(n7828), .ZN(n7829) );
  AOI21_X1 U9597 ( .B1(n7830), .B2(n8108), .A(n7829), .ZN(n7833) );
  AOI22_X1 U9598 ( .A1(n7831), .A2(n9643), .B1(n9644), .B2(n9642), .ZN(n7832)
         );
  OAI21_X1 U9599 ( .B1(n7834), .B2(n7833), .A(n7832), .ZN(n9712) );
  NAND2_X1 U9600 ( .A1(n9712), .A2(n9633), .ZN(n7835) );
  OAI211_X1 U9601 ( .C1(n7837), .C2(n9650), .A(n7836), .B(n7835), .ZN(P1_U3276) );
  INV_X1 U9602 ( .A(n7838), .ZN(n7909) );
  NOR2_X1 U9603 ( .A1(n7909), .A2(n7839), .ZN(n7842) );
  XNOR2_X1 U9604 ( .A(n7840), .B(n8778), .ZN(n7841) );
  XNOR2_X1 U9605 ( .A(n7842), .B(n7841), .ZN(n7849) );
  AOI21_X1 U9606 ( .B1(n8527), .B2(n8779), .A(n7843), .ZN(n7845) );
  OR2_X1 U9607 ( .A1(n8523), .A2(n7961), .ZN(n7844) );
  OAI211_X1 U9608 ( .C1(n8524), .C2(n7846), .A(n7845), .B(n7844), .ZN(n7847)
         );
  AOI21_X1 U9609 ( .B1(n6092), .B2(n8478), .A(n7847), .ZN(n7848) );
  OAI21_X1 U9610 ( .B1(n7849), .B2(n8518), .A(n7848), .ZN(P2_U3157) );
  NAND2_X1 U9611 ( .A1(n7854), .A2(n7850), .ZN(n7852) );
  OAI211_X1 U9612 ( .C1(n9172), .C2(n7853), .A(n7852), .B(n7851), .ZN(P2_U3267) );
  INV_X1 U9613 ( .A(n7854), .ZN(n7857) );
  OAI222_X1 U9614 ( .A1(n8017), .A2(n7857), .B1(n7856), .B2(P1_U3086), .C1(
        n7855), .C2(n9775), .ZN(P1_U3327) );
  XNOR2_X1 U9615 ( .A(n7859), .B(n7858), .ZN(n7860) );
  XNOR2_X1 U9616 ( .A(n7861), .B(n7860), .ZN(n7868) );
  NAND2_X1 U9617 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9937) );
  OAI21_X1 U9618 ( .B1(n9252), .B2(n7941), .A(n9937), .ZN(n7862) );
  AOI21_X1 U9619 ( .B1(n9250), .B2(n9642), .A(n7862), .ZN(n7863) );
  OAI21_X1 U9620 ( .B1(n9260), .B2(n7864), .A(n7863), .ZN(n7865) );
  AOI21_X1 U9621 ( .B1(n7866), .B2(n9265), .A(n7865), .ZN(n7867) );
  OAI21_X1 U9622 ( .B1(n7868), .B2(n9267), .A(n7867), .ZN(P1_U3228) );
  INV_X1 U9623 ( .A(n7869), .ZN(n7870) );
  NOR2_X1 U9624 ( .A1(n7871), .A2(n7870), .ZN(n7873) );
  MUX2_X1 U9625 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8799), .Z(n7972) );
  XNOR2_X1 U9626 ( .A(n7972), .B(n7982), .ZN(n7872) );
  NOR2_X1 U9627 ( .A1(n7873), .A2(n7872), .ZN(n7973) );
  AOI21_X1 U9628 ( .B1(n7873), .B2(n7872), .A(n7973), .ZN(n7888) );
  OAI21_X1 U9629 ( .B1(n7875), .B2(n7735), .A(n7874), .ZN(n7981) );
  XOR2_X1 U9630 ( .A(n7981), .B(n7982), .Z(n7876) );
  OAI21_X1 U9631 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7876), .A(n7983), .ZN(
        n7886) );
  INV_X1 U9632 ( .A(n10020), .ZN(n10106) );
  NAND2_X1 U9633 ( .A1(n10106), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7878) );
  OR2_X1 U9634 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7877), .ZN(n7897) );
  OAI211_X1 U9635 ( .C1(n10027), .C2(n7982), .A(n7878), .B(n7897), .ZN(n7885)
         );
  AOI21_X1 U9636 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7880), .A(n7879), .ZN(
        n7967) );
  AOI21_X1 U9637 ( .B1(n7882), .B2(n7881), .A(n7968), .ZN(n7883) );
  NOR2_X1 U9638 ( .A1(n7883), .A2(n10122), .ZN(n7884) );
  AOI211_X1 U9639 ( .C1(n10116), .C2(n7886), .A(n7885), .B(n7884), .ZN(n7887)
         );
  OAI21_X1 U9640 ( .B1(n7888), .B2(n10004), .A(n7887), .ZN(P2_U3193) );
  INV_X1 U9641 ( .A(n8663), .ZN(n7966) );
  OAI22_X1 U9642 ( .A1(n7889), .A2(n9164), .B1(n7966), .B2(n9118), .ZN(n7892)
         );
  MUX2_X1 U9643 ( .A(n7890), .B(P2_REG0_REG_12__SCAN_IN), .S(n10207), .Z(n7891) );
  OR2_X1 U9644 ( .A1(n7892), .A2(n7891), .ZN(P2_U3426) );
  OAI211_X1 U9645 ( .C1(n7895), .C2(n7894), .A(n7893), .B(n8507), .ZN(n7902)
         );
  INV_X1 U9646 ( .A(n7896), .ZN(n7900) );
  NAND2_X1 U9647 ( .A1(n8527), .A2(n8778), .ZN(n7898) );
  OAI211_X1 U9648 ( .C1(n8523), .C2(n8662), .A(n7898), .B(n7897), .ZN(n7899)
         );
  AOI21_X1 U9649 ( .B1(n8514), .B2(n7900), .A(n7899), .ZN(n7901) );
  OAI211_X1 U9650 ( .C1(n7903), .C2(n8530), .A(n7902), .B(n7901), .ZN(P2_U3176) );
  NAND2_X1 U9651 ( .A1(n8478), .A2(n7904), .ZN(n7907) );
  AOI21_X1 U9652 ( .B1(n8527), .B2(n8780), .A(n7905), .ZN(n7906) );
  OAI211_X1 U9653 ( .C1(n7908), .C2(n8523), .A(n7907), .B(n7906), .ZN(n7913)
         );
  AOI211_X1 U9654 ( .C1(n7911), .C2(n7910), .A(n8518), .B(n7909), .ZN(n7912)
         );
  AOI211_X1 U9655 ( .C1(n7914), .C2(n8514), .A(n7913), .B(n7912), .ZN(n7915)
         );
  INV_X1 U9656 ( .A(n7915), .ZN(P2_U3171) );
  INV_X1 U9657 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7919) );
  INV_X1 U9658 ( .A(n8674), .ZN(n7916) );
  OR2_X1 U9659 ( .A1(n8668), .A2(n7916), .ZN(n8577) );
  XOR2_X1 U9660 ( .A(n8577), .B(n7917), .Z(n7918) );
  AOI222_X1 U9661 ( .A1(n10134), .A2(n7918), .B1(n9019), .B2(n10131), .C1(
        n8776), .C2(n10129), .ZN(n7950) );
  MUX2_X1 U9662 ( .A(n7919), .B(n7950), .S(n10205), .Z(n7921) );
  XNOR2_X1 U9663 ( .A(n4442), .B(n8577), .ZN(n7953) );
  INV_X1 U9664 ( .A(n9164), .ZN(n8005) );
  AOI22_X1 U9665 ( .A1(n7953), .A2(n8005), .B1(n9161), .B2(n8479), .ZN(n7920)
         );
  NAND2_X1 U9666 ( .A1(n7921), .A2(n7920), .ZN(P2_U3429) );
  INV_X1 U9667 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7922) );
  MUX2_X1 U9668 ( .A(n7922), .B(n7950), .S(n10225), .Z(n7924) );
  AOI22_X1 U9669 ( .A1(n7953), .A2(n8000), .B1(n9075), .B2(n8479), .ZN(n7923)
         );
  NAND2_X1 U9670 ( .A1(n7924), .A2(n7923), .ZN(P2_U3472) );
  XNOR2_X1 U9671 ( .A(n7925), .B(n7927), .ZN(n9711) );
  OAI211_X1 U9672 ( .C1(n7927), .C2(n7926), .A(n9637), .B(n9640), .ZN(n7929)
         );
  AOI22_X1 U9673 ( .A1(n9610), .A2(n9644), .B1(n9287), .B2(n9643), .ZN(n7928)
         );
  NAND2_X1 U9674 ( .A1(n7929), .A2(n7928), .ZN(n9708) );
  INV_X1 U9675 ( .A(n7930), .ZN(n7931) );
  AOI211_X1 U9676 ( .C1(n9709), .C2(n7931), .A(n9682), .B(n9625), .ZN(n9707)
         );
  NAND2_X1 U9677 ( .A1(n9707), .A2(n9616), .ZN(n7934) );
  INV_X1 U9678 ( .A(n9259), .ZN(n7932) );
  AOI22_X1 U9679 ( .A1(n9469), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n7932), .B2(
        n9617), .ZN(n7933) );
  OAI211_X1 U9680 ( .C1(n7935), .C2(n9629), .A(n7934), .B(n7933), .ZN(n7936)
         );
  AOI21_X1 U9681 ( .B1(n9633), .B2(n9708), .A(n7936), .ZN(n7937) );
  OAI21_X1 U9682 ( .B1(n9711), .B2(n9650), .A(n7937), .ZN(P1_U3275) );
  XNOR2_X1 U9683 ( .A(n7938), .B(n9211), .ZN(n7940) );
  NOR2_X1 U9684 ( .A1(n7940), .A2(n7939), .ZN(n9210) );
  AOI21_X1 U9685 ( .B1(n7940), .B2(n7939), .A(n9210), .ZN(n7949) );
  NAND2_X1 U9686 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9909) );
  OAI21_X1 U9687 ( .B1(n9279), .B2(n7941), .A(n9909), .ZN(n7942) );
  AOI21_X1 U9688 ( .B1(n9277), .B2(n7943), .A(n7942), .ZN(n7944) );
  OAI21_X1 U9689 ( .B1(n9260), .B2(n7945), .A(n7944), .ZN(n7946) );
  AOI21_X1 U9690 ( .B1(n7947), .B2(n9265), .A(n7946), .ZN(n7948) );
  OAI21_X1 U9691 ( .B1(n7949), .B2(n9267), .A(n7948), .ZN(P1_U3241) );
  INV_X1 U9692 ( .A(n7950), .ZN(n7952) );
  OAI22_X1 U9693 ( .A1(n8669), .A2(n8899), .B1(n8471), .B2(n8977), .ZN(n7951)
         );
  OAI21_X1 U9694 ( .B1(n7952), .B2(n7951), .A(n10145), .ZN(n7955) );
  AOI22_X1 U9695 ( .A1(n7953), .A2(n10142), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10146), .ZN(n7954) );
  NAND2_X1 U9696 ( .A1(n7955), .A2(n7954), .ZN(P2_U3220) );
  OAI211_X1 U9697 ( .C1(n7958), .C2(n7957), .A(n7956), .B(n8507), .ZN(n7965)
         );
  INV_X1 U9698 ( .A(n8527), .ZN(n8511) );
  INV_X1 U9699 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7959) );
  NOR2_X1 U9700 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7959), .ZN(n7987) );
  AOI21_X1 U9701 ( .B1(n8468), .B2(n8775), .A(n7987), .ZN(n7960) );
  OAI21_X1 U9702 ( .B1(n7961), .B2(n8511), .A(n7960), .ZN(n7962) );
  AOI21_X1 U9703 ( .B1(n7963), .B2(n8514), .A(n7962), .ZN(n7964) );
  OAI211_X1 U9704 ( .C1(n7966), .C2(n8530), .A(n7965), .B(n7964), .ZN(P2_U3164) );
  NOR2_X1 U9705 ( .A1(n7975), .A2(n7967), .ZN(n7969) );
  NAND2_X1 U9706 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8827), .ZN(n7970) );
  OAI21_X1 U9707 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8827), .A(n7970), .ZN(
        n7971) );
  AOI21_X1 U9708 ( .B1(n4444), .B2(n7971), .A(n8785), .ZN(n7995) );
  INV_X1 U9709 ( .A(n7972), .ZN(n7974) );
  MUX2_X1 U9710 ( .A(n7976), .B(n7980), .S(n8799), .Z(n7977) );
  NOR2_X1 U9711 ( .A1(n7977), .A2(n7988), .ZN(n8800) );
  NOR2_X1 U9712 ( .A1(n8800), .A2(n4449), .ZN(n7979) );
  NAND2_X1 U9713 ( .A1(n4427), .A2(n7979), .ZN(n7978) );
  OAI211_X1 U9714 ( .C1(n4427), .C2(n7979), .A(n10115), .B(n7978), .ZN(n7994)
         );
  AOI22_X1 U9715 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8827), .B1(n7988), .B2(
        n7980), .ZN(n7986) );
  NAND2_X1 U9716 ( .A1(n7982), .A2(n7981), .ZN(n7984) );
  NAND2_X1 U9717 ( .A1(n7986), .A2(n7985), .ZN(n8828) );
  OAI21_X1 U9718 ( .B1(n7986), .B2(n7985), .A(n8828), .ZN(n7992) );
  INV_X1 U9719 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7990) );
  AOI21_X1 U9720 ( .B1(n10107), .B2(n7988), .A(n7987), .ZN(n7989) );
  OAI21_X1 U9721 ( .B1(n10020), .B2(n7990), .A(n7989), .ZN(n7991) );
  AOI21_X1 U9722 ( .B1(n7992), .B2(n10116), .A(n7991), .ZN(n7993) );
  OAI211_X1 U9723 ( .C1(n7995), .C2(n10122), .A(n7994), .B(n7993), .ZN(
        P2_U3194) );
  INV_X1 U9724 ( .A(n7997), .ZN(n8679) );
  OR2_X1 U9725 ( .A1(n8678), .A2(n8679), .ZN(n8561) );
  XNOR2_X1 U9726 ( .A(n7996), .B(n8561), .ZN(n7998) );
  OAI222_X1 U9727 ( .A1(n8976), .A2(n8366), .B1(n8974), .B2(n8670), .C1(n7998), 
        .C2(n8972), .ZN(n8008) );
  INV_X1 U9728 ( .A(n8008), .ZN(n8003) );
  MUX2_X1 U9729 ( .A(n8825), .B(n8003), .S(n10225), .Z(n8002) );
  XNOR2_X1 U9730 ( .A(n7999), .B(n8561), .ZN(n8011) );
  AOI22_X1 U9731 ( .A1(n8011), .A2(n8000), .B1(n9075), .B2(n8372), .ZN(n8001)
         );
  NAND2_X1 U9732 ( .A1(n8002), .A2(n8001), .ZN(P2_U3473) );
  INV_X1 U9733 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8004) );
  MUX2_X1 U9734 ( .A(n8004), .B(n8003), .S(n10205), .Z(n8007) );
  AOI22_X1 U9735 ( .A1(n8011), .A2(n8005), .B1(n9161), .B2(n8372), .ZN(n8006)
         );
  NAND2_X1 U9736 ( .A1(n8007), .A2(n8006), .ZN(P2_U3432) );
  INV_X1 U9737 ( .A(n8899), .ZN(n8909) );
  AOI21_X1 U9738 ( .B1(n8909), .B2(n8372), .A(n8008), .ZN(n8013) );
  OAI22_X1 U9739 ( .A1(n10145), .A2(n8009), .B1(n8370), .B2(n8977), .ZN(n8010)
         );
  AOI21_X1 U9740 ( .B1(n8011), .B2(n10142), .A(n8010), .ZN(n8012) );
  OAI21_X1 U9741 ( .B1(n8013), .B2(n10146), .A(n8012), .ZN(P2_U3219) );
  INV_X1 U9742 ( .A(n8014), .ZN(n9174) );
  OAI222_X1 U9743 ( .A1(n8017), .A2(n9174), .B1(P1_U3086), .B2(n8016), .C1(
        n8015), .C2(n9775), .ZN(P1_U3326) );
  INV_X1 U9744 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8345) );
  INV_X1 U9745 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U9746 ( .A1(n8024), .A2(n7133), .ZN(n8027) );
  INV_X1 U9747 ( .A(n8024), .ZN(n8025) );
  NAND2_X1 U9748 ( .A1(n8025), .A2(SI_30_), .ZN(n8026) );
  NAND2_X1 U9749 ( .A1(n8027), .A2(n8026), .ZN(n8170) );
  XNOR2_X1 U9750 ( .A(n8029), .B(n8028), .ZN(n8030) );
  NAND2_X1 U9751 ( .A1(n9781), .A2(n8172), .ZN(n8033) );
  INV_X1 U9752 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9776) );
  OR2_X1 U9753 ( .A1(n8173), .A2(n9776), .ZN(n8032) );
  INV_X1 U9754 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9653) );
  INV_X1 U9755 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8034) );
  OR2_X1 U9756 ( .A1(n8035), .A2(n8034), .ZN(n8037) );
  INV_X1 U9757 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9732) );
  OR2_X1 U9758 ( .A1(n5907), .A2(n9732), .ZN(n8036) );
  OAI211_X1 U9759 ( .C1(n5095), .C2(n9653), .A(n8037), .B(n8036), .ZN(n9461)
         );
  INV_X1 U9760 ( .A(n9461), .ZN(n8038) );
  NAND2_X1 U9761 ( .A1(n8137), .A2(n8039), .ZN(n8184) );
  NAND2_X1 U9762 ( .A1(n9543), .A2(n8040), .ZN(n8193) );
  MUX2_X1 U9763 ( .A(n8184), .B(n8193), .S(n8176), .Z(n8139) );
  OR2_X1 U9764 ( .A1(n9615), .A2(n8041), .ZN(n8043) );
  AND2_X1 U9765 ( .A1(n8195), .A2(n8043), .ZN(n8057) );
  NAND2_X1 U9766 ( .A1(n8051), .A2(n8129), .ZN(n8216) );
  INV_X1 U9767 ( .A(n8241), .ZN(n8042) );
  AOI21_X1 U9768 ( .B1(n8296), .B2(n8216), .A(n8042), .ZN(n8302) );
  INV_X1 U9769 ( .A(n8176), .ZN(n8179) );
  AOI21_X1 U9770 ( .B1(n8302), .B2(n8058), .A(n8179), .ZN(n8045) );
  AND2_X1 U9771 ( .A1(n8131), .A2(n8058), .ZN(n8194) );
  AOI21_X1 U9772 ( .B1(n8043), .B2(n8242), .A(n8176), .ZN(n8044) );
  AOI22_X1 U9773 ( .A1(n8057), .A2(n8045), .B1(n8194), .B2(n8044), .ZN(n8135)
         );
  NAND2_X1 U9774 ( .A1(n8058), .A2(n8241), .ZN(n8049) );
  AND2_X1 U9775 ( .A1(n9636), .A2(n8046), .ZN(n8295) );
  AND2_X1 U9776 ( .A1(n8051), .A2(n8179), .ZN(n8059) );
  INV_X1 U9777 ( .A(n8059), .ZN(n8047) );
  OR3_X1 U9778 ( .A1(n8049), .A2(n8295), .A3(n8047), .ZN(n8048) );
  NAND2_X1 U9779 ( .A1(n9611), .A2(n8179), .ZN(n8050) );
  NAND2_X1 U9780 ( .A1(n8048), .A2(n8050), .ZN(n8056) );
  INV_X1 U9781 ( .A(n9597), .ZN(n9757) );
  INV_X1 U9782 ( .A(n8049), .ZN(n8055) );
  INV_X1 U9783 ( .A(n8295), .ZN(n8053) );
  INV_X1 U9784 ( .A(n8050), .ZN(n8052) );
  AND3_X1 U9785 ( .A1(n8053), .A2(n8052), .A3(n8051), .ZN(n8054) );
  AOI22_X1 U9786 ( .A1(n8056), .A2(n9757), .B1(n8055), .B2(n8054), .ZN(n8134)
         );
  INV_X1 U9787 ( .A(n8057), .ZN(n8187) );
  NAND3_X1 U9788 ( .A1(n8295), .A2(n8242), .A3(n8176), .ZN(n8061) );
  NAND4_X1 U9789 ( .A1(n8131), .A2(n8059), .A3(n8241), .A4(n8058), .ZN(n8060)
         );
  OAI21_X1 U9790 ( .B1(n8187), .B2(n8061), .A(n8060), .ZN(n8130) );
  INV_X1 U9791 ( .A(n8106), .ZN(n8062) );
  NAND2_X1 U9792 ( .A1(n8063), .A2(n8062), .ZN(n8064) );
  AND2_X1 U9793 ( .A1(n8064), .A2(n8108), .ZN(n8111) );
  NAND2_X1 U9794 ( .A1(n8070), .A2(n8179), .ZN(n8069) );
  NAND2_X1 U9795 ( .A1(n8266), .A2(n8071), .ZN(n8065) );
  NOR2_X1 U9796 ( .A1(n8069), .A2(n8065), .ZN(n8066) );
  NAND2_X1 U9797 ( .A1(n8067), .A2(n8066), .ZN(n8079) );
  NAND2_X1 U9798 ( .A1(n8068), .A2(n8268), .ZN(n8073) );
  INV_X1 U9799 ( .A(n8069), .ZN(n8072) );
  NAND2_X1 U9800 ( .A1(n8071), .A2(n8070), .ZN(n8270) );
  AOI22_X1 U9801 ( .A1(n8073), .A2(n8072), .B1(n8270), .B2(n8176), .ZN(n8078)
         );
  NAND2_X1 U9802 ( .A1(n8074), .A2(n8266), .ZN(n8076) );
  NAND4_X1 U9803 ( .A1(n8076), .A2(n8075), .A3(n8268), .A4(n8176), .ZN(n8077)
         );
  NAND3_X1 U9804 ( .A1(n8079), .A2(n8078), .A3(n8077), .ZN(n8084) );
  INV_X1 U9805 ( .A(n8080), .ZN(n8081) );
  OAI21_X1 U9806 ( .B1(n8084), .B2(n8081), .A(n8086), .ZN(n8083) );
  NAND2_X1 U9807 ( .A1(n8083), .A2(n8082), .ZN(n8088) );
  INV_X1 U9808 ( .A(n8084), .ZN(n8087) );
  NAND2_X1 U9809 ( .A1(n8089), .A2(n8090), .ZN(n8098) );
  NAND2_X1 U9810 ( .A1(n8098), .A2(n8090), .ZN(n8092) );
  NAND2_X1 U9811 ( .A1(n8092), .A2(n8091), .ZN(n8094) );
  NAND2_X1 U9812 ( .A1(n8094), .A2(n8093), .ZN(n8100) );
  INV_X1 U9813 ( .A(n8095), .ZN(n8097) );
  AOI21_X1 U9814 ( .B1(n8098), .B2(n8097), .A(n8096), .ZN(n8099) );
  MUX2_X1 U9815 ( .A(n8100), .B(n8099), .S(n8176), .Z(n8112) );
  NAND2_X1 U9816 ( .A1(n8118), .A2(n8279), .ZN(n8103) );
  NAND2_X1 U9817 ( .A1(n8124), .A2(n8121), .ZN(n8287) );
  AOI21_X1 U9818 ( .B1(n8104), .B2(n8261), .A(n8287), .ZN(n8107) );
  NAND2_X1 U9819 ( .A1(n8106), .A2(n8105), .ZN(n8260) );
  OAI21_X1 U9820 ( .B1(n8107), .B2(n8260), .A(n8291), .ZN(n8109) );
  NAND2_X1 U9821 ( .A1(n8109), .A2(n8108), .ZN(n8110) );
  MUX2_X1 U9822 ( .A(n8111), .B(n8110), .S(n8179), .Z(n8127) );
  INV_X1 U9823 ( .A(n8112), .ZN(n8114) );
  NAND2_X1 U9824 ( .A1(n8114), .A2(n8113), .ZN(n8117) );
  NAND2_X1 U9825 ( .A1(n8116), .A2(n8115), .ZN(n8281) );
  AOI21_X1 U9826 ( .B1(n8117), .B2(n8279), .A(n8281), .ZN(n8120) );
  NAND2_X1 U9827 ( .A1(n8119), .A2(n8118), .ZN(n8285) );
  OAI21_X1 U9828 ( .B1(n8120), .B2(n8285), .A(n8284), .ZN(n8122) );
  NAND2_X1 U9829 ( .A1(n8122), .A2(n8121), .ZN(n8123) );
  NAND3_X1 U9830 ( .A1(n8123), .A2(n8235), .A3(n8261), .ZN(n8125) );
  NAND4_X1 U9831 ( .A1(n8125), .A2(n8291), .A3(n8176), .A4(n8124), .ZN(n8126)
         );
  NAND2_X1 U9832 ( .A1(n8127), .A2(n8126), .ZN(n8128) );
  NAND3_X1 U9833 ( .A1(n8130), .A2(n8129), .A3(n8128), .ZN(n8133) );
  OR2_X1 U9834 ( .A1(n8131), .A2(n8179), .ZN(n8132) );
  NAND4_X1 U9835 ( .A1(n8135), .A2(n8134), .A3(n8133), .A4(n8132), .ZN(n8136)
         );
  MUX2_X1 U9836 ( .A(n9543), .B(n8137), .S(n8176), .Z(n8138) );
  MUX2_X1 U9837 ( .A(n8185), .B(n8198), .S(n8176), .Z(n8140) );
  INV_X1 U9838 ( .A(n8152), .ZN(n8141) );
  AOI21_X1 U9839 ( .B1(n8154), .B2(n8200), .A(n8141), .ZN(n8144) );
  AND3_X1 U9840 ( .A1(n8303), .A2(n8179), .A3(n8153), .ZN(n8142) );
  OAI211_X1 U9841 ( .C1(n4795), .C2(n8144), .A(n8143), .B(n8142), .ZN(n8165)
         );
  NAND3_X1 U9842 ( .A1(n9486), .A2(n9280), .A3(n8179), .ZN(n8145) );
  NAND2_X1 U9843 ( .A1(n9496), .A2(n8179), .ZN(n8146) );
  NAND2_X1 U9844 ( .A1(n8145), .A2(n8146), .ZN(n8150) );
  OAI21_X1 U9845 ( .B1(n9513), .B2(n8146), .A(n9486), .ZN(n8149) );
  OR2_X1 U9846 ( .A1(n9496), .A2(n8179), .ZN(n8159) );
  NOR2_X1 U9847 ( .A1(n8159), .A2(n9280), .ZN(n8147) );
  OR2_X1 U9848 ( .A1(n9486), .A2(n8147), .ZN(n8148) );
  AOI22_X1 U9849 ( .A1(n8151), .A2(n8150), .B1(n8149), .B2(n8148), .ZN(n8164)
         );
  AND2_X1 U9850 ( .A1(n8190), .A2(n8176), .ZN(n8157) );
  AND2_X1 U9851 ( .A1(n8153), .A2(n8152), .ZN(n8203) );
  NAND4_X1 U9852 ( .A1(n8158), .A2(n8157), .A3(n8156), .A4(n8155), .ZN(n8163)
         );
  OR3_X1 U9853 ( .A1(n9486), .A2(n9280), .A3(n8179), .ZN(n8160) );
  NAND2_X1 U9854 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  NAND2_X1 U9855 ( .A1(n8339), .A2(n8161), .ZN(n8162) );
  NAND4_X1 U9856 ( .A1(n8165), .A2(n8164), .A3(n8163), .A4(n8162), .ZN(n8169)
         );
  INV_X1 U9857 ( .A(n8166), .ZN(n8209) );
  INV_X1 U9858 ( .A(n8167), .ZN(n8207) );
  AOI21_X1 U9859 ( .B1(n4797), .B2(n8169), .A(n8168), .ZN(n8178) );
  NAND2_X1 U9860 ( .A1(n8533), .A2(n8172), .ZN(n8175) );
  OR2_X1 U9861 ( .A1(n8173), .A2(n8345), .ZN(n8174) );
  MUX2_X1 U9862 ( .A(n8178), .B(n8176), .S(n9467), .Z(n8177) );
  MUX2_X1 U9863 ( .A(n8179), .B(n8178), .S(n9467), .Z(n8180) );
  INV_X1 U9864 ( .A(n9286), .ZN(n8210) );
  NOR3_X1 U9865 ( .A1(n8180), .A2(n9734), .A3(n8210), .ZN(n8181) );
  NOR3_X1 U9866 ( .A1(n8182), .A2(n8181), .A3(n8212), .ZN(n8255) );
  OAI211_X1 U9867 ( .C1(n8315), .C2(n8317), .A(n8264), .B(n8254), .ZN(n8258)
         );
  INV_X1 U9868 ( .A(n8203), .ZN(n8188) );
  NAND3_X1 U9869 ( .A1(n8198), .A2(n9543), .A3(n8184), .ZN(n8186) );
  NAND2_X1 U9870 ( .A1(n8186), .A2(n8185), .ZN(n8192) );
  NOR3_X1 U9871 ( .A1(n8188), .A2(n8187), .A3(n8192), .ZN(n8299) );
  NAND2_X1 U9872 ( .A1(n8299), .A2(n9608), .ZN(n8191) );
  INV_X1 U9873 ( .A(n8303), .ZN(n8189) );
  AOI21_X1 U9874 ( .B1(n8191), .B2(n8190), .A(n8189), .ZN(n8208) );
  NAND2_X1 U9875 ( .A1(n8192), .A2(n8200), .ZN(n8202) );
  INV_X1 U9876 ( .A(n8193), .ZN(n8199) );
  INV_X1 U9877 ( .A(n8194), .ZN(n8196) );
  NAND2_X1 U9878 ( .A1(n8196), .A2(n8195), .ZN(n8197) );
  NAND4_X1 U9879 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), .ZN(n8201)
         );
  NAND4_X1 U9880 ( .A1(n8303), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n8204)
         );
  NAND2_X1 U9881 ( .A1(n8205), .A2(n8204), .ZN(n8259) );
  NOR2_X1 U9882 ( .A1(n8207), .A2(n8206), .ZN(n8305) );
  OAI21_X1 U9883 ( .B1(n8208), .B2(n8259), .A(n8305), .ZN(n8211) );
  AOI21_X1 U9884 ( .B1(n8210), .B2(n9467), .A(n8209), .ZN(n8309) );
  NOR2_X1 U9885 ( .A1(n9467), .A2(n8210), .ZN(n8310) );
  AOI22_X1 U9886 ( .A1(n8211), .A2(n8309), .B1(n8310), .B2(n9461), .ZN(n8215)
         );
  OAI21_X1 U9887 ( .B1(n9738), .B2(n9461), .A(n8315), .ZN(n8214) );
  OAI211_X1 U9888 ( .C1(n8215), .C2(n8214), .A(n8213), .B(n8312), .ZN(n8253)
         );
  INV_X1 U9889 ( .A(n8216), .ZN(n8240) );
  NOR2_X1 U9890 ( .A1(n8217), .A2(n8264), .ZN(n8224) );
  NOR2_X1 U9891 ( .A1(n8219), .A2(n8218), .ZN(n8223) );
  INV_X1 U9892 ( .A(n8220), .ZN(n8222) );
  NAND4_X1 U9893 ( .A1(n8224), .A2(n8223), .A3(n8222), .A4(n8221), .ZN(n8226)
         );
  NOR2_X1 U9894 ( .A1(n8226), .A2(n8225), .ZN(n8227) );
  NAND4_X1 U9895 ( .A1(n8276), .A2(n8229), .A3(n8228), .A4(n8227), .ZN(n8231)
         );
  NOR3_X1 U9896 ( .A1(n8232), .A2(n8231), .A3(n8230), .ZN(n8233) );
  NAND3_X1 U9897 ( .A1(n8235), .A2(n8234), .A3(n8233), .ZN(n8236) );
  NOR2_X1 U9898 ( .A1(n8237), .A2(n8236), .ZN(n8238) );
  NAND4_X1 U9899 ( .A1(n8295), .A2(n8240), .A3(n8239), .A4(n8238), .ZN(n8243)
         );
  NAND2_X1 U9900 ( .A1(n8242), .A2(n8241), .ZN(n9638) );
  NOR2_X1 U9901 ( .A1(n8243), .A2(n9638), .ZN(n8244) );
  AND4_X1 U9902 ( .A1(n9582), .A2(n9591), .A3(n8244), .A4(n9607), .ZN(n8245)
         );
  NAND3_X1 U9903 ( .A1(n9545), .A2(n9558), .A3(n8245), .ZN(n8246) );
  NOR2_X1 U9904 ( .A1(n9519), .A2(n8246), .ZN(n8247) );
  NAND4_X1 U9905 ( .A1(n8248), .A2(n9493), .A3(n9511), .A4(n8247), .ZN(n8249)
         );
  NOR2_X1 U9906 ( .A1(n8250), .A2(n8249), .ZN(n8252) );
  XNOR2_X1 U9907 ( .A(n9467), .B(n9286), .ZN(n8251) );
  NAND4_X1 U9908 ( .A1(n8315), .A2(n8312), .A3(n8252), .A4(n8251), .ZN(n8256)
         );
  AND2_X1 U9909 ( .A1(n8253), .A2(n8256), .ZN(n8257) );
  INV_X1 U9910 ( .A(n8259), .ZN(n8308) );
  INV_X1 U9911 ( .A(n8260), .ZN(n8294) );
  INV_X1 U9912 ( .A(n8261), .ZN(n8290) );
  INV_X1 U9913 ( .A(n8262), .ZN(n8265) );
  NAND2_X1 U9914 ( .A1(n9300), .A2(n5835), .ZN(n8263) );
  NAND4_X1 U9915 ( .A1(n8266), .A2(n8265), .A3(n8264), .A4(n8263), .ZN(n8267)
         );
  NAND3_X1 U9916 ( .A1(n8269), .A2(n8268), .A3(n8267), .ZN(n8274) );
  INV_X1 U9917 ( .A(n8270), .ZN(n8273) );
  INV_X1 U9918 ( .A(n8271), .ZN(n8272) );
  AOI21_X1 U9919 ( .B1(n8274), .B2(n8273), .A(n8272), .ZN(n8278) );
  INV_X1 U9920 ( .A(n8275), .ZN(n8277) );
  OAI21_X1 U9921 ( .B1(n8278), .B2(n8277), .A(n8276), .ZN(n8283) );
  AND2_X1 U9922 ( .A1(n8280), .A2(n8279), .ZN(n8282) );
  AOI21_X1 U9923 ( .B1(n8283), .B2(n8282), .A(n8281), .ZN(n8286) );
  OAI21_X1 U9924 ( .B1(n8286), .B2(n8285), .A(n8284), .ZN(n8289) );
  INV_X1 U9925 ( .A(n8287), .ZN(n8288) );
  OAI21_X1 U9926 ( .B1(n8290), .B2(n8289), .A(n8288), .ZN(n8293) );
  INV_X1 U9927 ( .A(n8291), .ZN(n8292) );
  AOI21_X1 U9928 ( .B1(n8294), .B2(n8293), .A(n8292), .ZN(n8297) );
  OAI211_X1 U9929 ( .C1(n8298), .C2(n8297), .A(n8296), .B(n8295), .ZN(n8301)
         );
  INV_X1 U9930 ( .A(n8299), .ZN(n8300) );
  AOI21_X1 U9931 ( .B1(n8302), .B2(n8301), .A(n8300), .ZN(n8304) );
  OAI21_X1 U9932 ( .B1(n8304), .B2(n4795), .A(n8303), .ZN(n8307) );
  INV_X1 U9933 ( .A(n8305), .ZN(n8306) );
  AOI21_X1 U9934 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(n8314) );
  INV_X1 U9935 ( .A(n8309), .ZN(n8313) );
  INV_X1 U9936 ( .A(n8310), .ZN(n8311) );
  OAI211_X1 U9937 ( .C1(n8314), .C2(n8313), .A(n8312), .B(n8311), .ZN(n8316)
         );
  NAND2_X1 U9938 ( .A1(n8316), .A2(n8315), .ZN(n8320) );
  NOR2_X1 U9939 ( .A1(n8320), .A2(n8317), .ZN(n8318) );
  NAND2_X1 U9940 ( .A1(n8318), .A2(n5818), .ZN(n8322) );
  NAND2_X1 U9941 ( .A1(n8320), .A2(n8319), .ZN(n8321) );
  NAND2_X1 U9942 ( .A1(n8322), .A2(n8321), .ZN(n8323) );
  NOR4_X1 U9943 ( .A1(n9549), .A2(n8325), .A3(n5796), .A4(n5904), .ZN(n8328)
         );
  OAI21_X1 U9944 ( .B1(n8329), .B2(n8326), .A(P1_B_REG_SCAN_IN), .ZN(n8327) );
  OAI222_X1 U9945 ( .A1(n8017), .A2(n8331), .B1(n5904), .B2(P1_U3086), .C1(
        n8330), .C2(n9775), .ZN(P1_U3328) );
  INV_X1 U9946 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8334) );
  OAI222_X1 U9947 ( .A1(n9775), .A2(n8334), .B1(n8017), .B2(n8333), .C1(
        P1_U3086), .C2(n8317), .ZN(P1_U3336) );
  NAND2_X1 U9948 ( .A1(n8335), .A2(n9616), .ZN(n8338) );
  AOI22_X1 U9949 ( .A1(n8336), .A2(n9617), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9469), .ZN(n8337) );
  OAI211_X1 U9950 ( .C1(n8339), .C2(n9629), .A(n8338), .B(n8337), .ZN(n8340)
         );
  AOI21_X1 U9951 ( .B1(n8341), .B2(n9633), .A(n8340), .ZN(n8342) );
  OAI21_X1 U9952 ( .B1(n8343), .B2(n9650), .A(n8342), .ZN(P1_U3265) );
  INV_X1 U9953 ( .A(n8533), .ZN(n8359) );
  OAI222_X1 U9954 ( .A1(n9775), .A2(n8345), .B1(n8017), .B2(n8359), .C1(
        P1_U3086), .C2(n8344), .ZN(P1_U3325) );
  AND2_X1 U9955 ( .A1(n8347), .A2(n8346), .ZN(n8349) );
  OAI21_X1 U9956 ( .B1(n8349), .B2(n8348), .A(n8507), .ZN(n8355) );
  NAND2_X1 U9957 ( .A1(n8514), .A2(n8876), .ZN(n8351) );
  AOI22_X1 U9958 ( .A1(n8527), .A2(n8895), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8350) );
  OAI211_X1 U9959 ( .C1(n8591), .C2(n8523), .A(n8351), .B(n8350), .ZN(n8352)
         );
  AOI21_X1 U9960 ( .B1(n9095), .B2(n8478), .A(n8352), .ZN(n8353) );
  OAI21_X1 U9961 ( .B1(n8355), .B2(n8354), .A(n8353), .ZN(P2_U3154) );
  OAI222_X1 U9962 ( .A1(n6364), .A2(P2_U3151), .B1(n9175), .B2(n8357), .C1(
        n8356), .C2(n9172), .ZN(P2_U3270) );
  OAI222_X1 U9963 ( .A1(n9172), .A2(n8534), .B1(n9175), .B2(n8359), .C1(n8358), 
        .C2(P2_U3151), .ZN(P2_U3265) );
  OAI222_X1 U9964 ( .A1(n6361), .A2(P2_U3151), .B1(n9175), .B2(n8361), .C1(
        n8360), .C2(n9172), .ZN(P2_U3271) );
  INV_X1 U9965 ( .A(n8362), .ZN(n8363) );
  AOI21_X1 U9966 ( .B1(n8365), .B2(n8364), .A(n8363), .ZN(n8374) );
  NAND2_X1 U9967 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n10071) );
  INV_X1 U9968 ( .A(n10071), .ZN(n8368) );
  NOR2_X1 U9969 ( .A1(n8523), .A2(n8366), .ZN(n8367) );
  AOI211_X1 U9970 ( .C1(n8527), .C2(n8775), .A(n8368), .B(n8367), .ZN(n8369)
         );
  OAI21_X1 U9971 ( .B1(n8370), .B2(n8524), .A(n8369), .ZN(n8371) );
  AOI21_X1 U9972 ( .B1(n8372), .B2(n8478), .A(n8371), .ZN(n8373) );
  OAI21_X1 U9973 ( .B1(n8374), .B2(n8518), .A(n8373), .ZN(P2_U3155) );
  INV_X1 U9974 ( .A(n8376), .ZN(n8448) );
  AOI21_X1 U9975 ( .B1(n8932), .B2(n8375), .A(n8448), .ZN(n8382) );
  NOR2_X1 U9976 ( .A1(n8523), .A2(n8922), .ZN(n8379) );
  OAI22_X1 U9977 ( .A1(n8511), .A2(n8921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8377), .ZN(n8378) );
  AOI211_X1 U9978 ( .C1(n8925), .C2(n8514), .A(n8379), .B(n8378), .ZN(n8381)
         );
  NAND2_X1 U9979 ( .A1(n8926), .A2(n8478), .ZN(n8380) );
  OAI211_X1 U9980 ( .C1(n8382), .C2(n8518), .A(n8381), .B(n8380), .ZN(P2_U3156) );
  NAND2_X1 U9981 ( .A1(n8383), .A2(n8492), .ZN(n8384) );
  NAND2_X1 U9982 ( .A1(n8384), .A2(n8493), .ZN(n8387) );
  INV_X1 U9983 ( .A(n8387), .ZN(n8496) );
  INV_X1 U9984 ( .A(n8386), .ZN(n8385) );
  NOR3_X1 U9985 ( .A1(n8496), .A2(n8385), .A3(n8388), .ZN(n8389) );
  NAND2_X1 U9986 ( .A1(n8387), .A2(n8386), .ZN(n8396) );
  OAI21_X1 U9987 ( .B1(n8389), .B2(n8459), .A(n8507), .ZN(n8393) );
  NAND2_X1 U9988 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8820) );
  OAI21_X1 U9989 ( .B1(n8523), .B2(n8975), .A(n8820), .ZN(n8391) );
  NOR2_X1 U9990 ( .A1(n8524), .A2(n8978), .ZN(n8390) );
  AOI211_X1 U9991 ( .C1(n8527), .C2(n9000), .A(n8391), .B(n8390), .ZN(n8392)
         );
  OAI211_X1 U9992 ( .C1(n8394), .C2(n8530), .A(n8393), .B(n8392), .ZN(P2_U3159) );
  NAND2_X1 U9993 ( .A1(n8396), .A2(n8395), .ZN(n8398) );
  INV_X1 U9994 ( .A(n8399), .ZN(n8401) );
  NOR3_X1 U9995 ( .A1(n4946), .A2(n8401), .A3(n8400), .ZN(n8405) );
  NAND2_X1 U9996 ( .A1(n8383), .A2(n8402), .ZN(n8404) );
  AND2_X1 U9997 ( .A1(n8404), .A2(n8403), .ZN(n8483) );
  OAI21_X1 U9998 ( .B1(n8405), .B2(n8483), .A(n8507), .ZN(n8410) );
  OAI22_X1 U9999 ( .A1(n8523), .A2(n8921), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8406), .ZN(n8408) );
  NOR2_X1 U10000 ( .A1(n8511), .A2(n8975), .ZN(n8407) );
  AOI211_X1 U10001 ( .C1(n8954), .C2(n8514), .A(n8408), .B(n8407), .ZN(n8409)
         );
  OAI211_X1 U10002 ( .C1(n8411), .C2(n8530), .A(n8410), .B(n8409), .ZN(
        P2_U3163) );
  INV_X1 U10003 ( .A(n8412), .ZN(n8449) );
  INV_X1 U10004 ( .A(n8413), .ZN(n8415) );
  NOR3_X1 U10005 ( .A1(n8449), .A2(n8415), .A3(n8414), .ZN(n8418) );
  INV_X1 U10006 ( .A(n8416), .ZN(n8417) );
  OAI21_X1 U10007 ( .B1(n8418), .B2(n8417), .A(n8507), .ZN(n8424) );
  OAI22_X1 U10008 ( .A1(n8523), .A2(n8420), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8419), .ZN(n8422) );
  NOR2_X1 U10009 ( .A1(n8511), .A2(n8922), .ZN(n8421) );
  AOI211_X1 U10010 ( .C1(n8897), .C2(n8514), .A(n8422), .B(n8421), .ZN(n8423)
         );
  OAI211_X1 U10011 ( .C1(n8900), .C2(n8530), .A(n8424), .B(n8423), .ZN(
        P2_U3165) );
  INV_X1 U10012 ( .A(n8425), .ZN(n8439) );
  INV_X1 U10013 ( .A(n8426), .ZN(n8429) );
  INV_X1 U10014 ( .A(n8427), .ZN(n8428) );
  AOI21_X1 U10015 ( .B1(n8521), .B2(n8429), .A(n8428), .ZN(n8430) );
  OAI21_X1 U10016 ( .B1(n8439), .B2(n8430), .A(n8507), .ZN(n8435) );
  NAND2_X1 U10017 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10103)
         );
  OAI21_X1 U10018 ( .B1(n8523), .B2(n8431), .A(n10103), .ZN(n8433) );
  NOR2_X1 U10019 ( .A1(n8524), .A2(n9012), .ZN(n8432) );
  AOI211_X1 U10020 ( .C1(n8527), .C2(n9009), .A(n8433), .B(n8432), .ZN(n8434)
         );
  OAI211_X1 U10021 ( .C1(n8436), .C2(n8530), .A(n8435), .B(n8434), .ZN(
        P2_U3166) );
  INV_X1 U10022 ( .A(n9148), .ZN(n8445) );
  NOR3_X1 U10023 ( .A1(n8439), .A2(n4708), .A3(n8438), .ZN(n8440) );
  INV_X1 U10024 ( .A(n8383), .ZN(n8495) );
  OAI21_X1 U10025 ( .B1(n8440), .B2(n8495), .A(n8507), .ZN(n8444) );
  NAND2_X1 U10026 ( .A1(n8468), .A2(n9000), .ZN(n8441) );
  NAND2_X1 U10027 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n10124)
         );
  OAI211_X1 U10028 ( .C1(n8511), .C2(n8774), .A(n8441), .B(n10124), .ZN(n8442)
         );
  AOI21_X1 U10029 ( .B1(n9002), .B2(n8514), .A(n8442), .ZN(n8443) );
  OAI211_X1 U10030 ( .C1(n8445), .C2(n8530), .A(n8444), .B(n8443), .ZN(
        P2_U3168) );
  NOR3_X1 U10031 ( .A1(n8448), .A2(n8447), .A3(n8446), .ZN(n8450) );
  OAI21_X1 U10032 ( .B1(n8450), .B2(n8449), .A(n8507), .ZN(n8455) );
  OAI22_X1 U10033 ( .A1(n8523), .A2(n8773), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8451), .ZN(n8453) );
  NOR2_X1 U10034 ( .A1(n8511), .A2(n8488), .ZN(n8452) );
  AOI211_X1 U10035 ( .C1(n8908), .C2(n8514), .A(n8453), .B(n8452), .ZN(n8454)
         );
  OAI211_X1 U10036 ( .C1(n8456), .C2(n8530), .A(n8455), .B(n8454), .ZN(
        P2_U3169) );
  NOR3_X1 U10037 ( .A1(n8459), .A2(n4677), .A3(n8458), .ZN(n8460) );
  OAI21_X1 U10038 ( .B1(n8460), .B2(n4946), .A(n8507), .ZN(n8465) );
  INV_X1 U10039 ( .A(n8461), .ZN(n8965) );
  AOI22_X1 U10040 ( .A1(n8468), .A2(n8962), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8462) );
  OAI21_X1 U10041 ( .B1(n8498), .B2(n8511), .A(n8462), .ZN(n8463) );
  AOI21_X1 U10042 ( .B1(n8965), .B2(n8514), .A(n8463), .ZN(n8464) );
  OAI211_X1 U10043 ( .C1(n8466), .C2(n8530), .A(n8465), .B(n8464), .ZN(
        P2_U3173) );
  NAND2_X1 U10044 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10055)
         );
  INV_X1 U10045 ( .A(n10055), .ZN(n8467) );
  AOI21_X1 U10046 ( .B1(n8468), .B2(n9019), .A(n8467), .ZN(n8470) );
  NAND2_X1 U10047 ( .A1(n8527), .A2(n8776), .ZN(n8469) );
  OAI211_X1 U10048 ( .C1(n8524), .C2(n8471), .A(n8470), .B(n8469), .ZN(n8477)
         );
  XNOR2_X1 U10049 ( .A(n8472), .B(n8775), .ZN(n8473) );
  XNOR2_X1 U10050 ( .A(n8474), .B(n8473), .ZN(n8475) );
  NOR2_X1 U10051 ( .A1(n8475), .A2(n8518), .ZN(n8476) );
  AOI211_X1 U10052 ( .C1(n8479), .C2(n8478), .A(n8477), .B(n8476), .ZN(n8480)
         );
  INV_X1 U10053 ( .A(n8480), .ZN(P2_U3174) );
  NOR3_X1 U10054 ( .A1(n8483), .A2(n8482), .A3(n8481), .ZN(n8486) );
  INV_X1 U10055 ( .A(n8484), .ZN(n8485) );
  OAI21_X1 U10056 ( .B1(n8486), .B2(n8485), .A(n8507), .ZN(n8491) );
  AOI22_X1 U10057 ( .A1(n8527), .A2(n8962), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8487) );
  OAI21_X1 U10058 ( .B1(n8488), .B2(n8523), .A(n8487), .ZN(n8489) );
  AOI21_X1 U10059 ( .B1(n8934), .B2(n8514), .A(n8489), .ZN(n8490) );
  OAI211_X1 U10060 ( .C1(n9054), .C2(n8530), .A(n8491), .B(n8490), .ZN(
        P2_U3175) );
  INV_X1 U10061 ( .A(n8492), .ZN(n8494) );
  NOR3_X1 U10062 ( .A1(n8495), .A2(n8494), .A3(n8493), .ZN(n8497) );
  OAI21_X1 U10063 ( .B1(n8497), .B2(n8496), .A(n8507), .ZN(n8502) );
  NAND2_X1 U10064 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9792) );
  OAI21_X1 U10065 ( .B1(n8523), .B2(n8498), .A(n9792), .ZN(n8500) );
  NOR2_X1 U10066 ( .A1(n8524), .A2(n8993), .ZN(n8499) );
  AOI211_X1 U10067 ( .C1(n8527), .C2(n9008), .A(n8500), .B(n8499), .ZN(n8501)
         );
  OAI211_X1 U10068 ( .C1(n8503), .C2(n8530), .A(n8502), .B(n8501), .ZN(
        P2_U3178) );
  XNOR2_X1 U10069 ( .A(n8505), .B(n8895), .ZN(n8506) );
  XNOR2_X1 U10070 ( .A(n8504), .B(n8506), .ZN(n8508) );
  NAND2_X1 U10071 ( .A1(n8508), .A2(n8507), .ZN(n8516) );
  NOR2_X1 U10072 ( .A1(n8523), .A2(n8509), .ZN(n8513) );
  OAI22_X1 U10073 ( .A1(n8511), .A2(n8773), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8510), .ZN(n8512) );
  AOI211_X1 U10074 ( .C1(n8886), .C2(n8514), .A(n8513), .B(n8512), .ZN(n8515)
         );
  OAI211_X1 U10075 ( .C1(n8517), .C2(n8530), .A(n8516), .B(n8515), .ZN(
        P2_U3180) );
  AOI21_X1 U10076 ( .B1(n8520), .B2(n8519), .A(n8518), .ZN(n8522) );
  NAND2_X1 U10077 ( .A1(n8522), .A2(n8521), .ZN(n8529) );
  NAND2_X1 U10078 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10087)
         );
  OAI21_X1 U10079 ( .B1(n8523), .B2(n8774), .A(n10087), .ZN(n8526) );
  NOR2_X1 U10080 ( .A1(n8524), .A2(n9022), .ZN(n8525) );
  AOI211_X1 U10081 ( .C1(n8527), .C2(n9019), .A(n8526), .B(n8525), .ZN(n8528)
         );
  OAI211_X1 U10082 ( .C1(n8560), .C2(n8530), .A(n8529), .B(n8528), .ZN(
        P2_U3181) );
  INV_X1 U10083 ( .A(n8746), .ZN(n8531) );
  NAND2_X1 U10084 ( .A1(n8533), .A2(n8544), .ZN(n8536) );
  OR2_X1 U10085 ( .A1(n6008), .A2(n8534), .ZN(n8535) );
  NOR2_X1 U10086 ( .A1(n9086), .A2(n8771), .ZN(n8586) );
  INV_X1 U10087 ( .A(n8537), .ZN(n8538) );
  NOR2_X1 U10088 ( .A1(n8586), .A2(n8538), .ZN(n8741) );
  NAND2_X1 U10089 ( .A1(n6012), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U10090 ( .A1(n4958), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U10091 ( .A1(n8539), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8540) );
  NAND4_X1 U10092 ( .A1(n8543), .A2(n8542), .A3(n8541), .A4(n8540), .ZN(n8848)
         );
  NAND2_X1 U10093 ( .A1(n9781), .A2(n8544), .ZN(n8547) );
  INV_X1 U10094 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8545) );
  OR2_X1 U10095 ( .A1(n6008), .A2(n8545), .ZN(n8546) );
  OAI21_X1 U10096 ( .B1(n9029), .B2(n8848), .A(n8852), .ZN(n8548) );
  INV_X1 U10097 ( .A(n8771), .ZN(n8589) );
  INV_X1 U10098 ( .A(n8550), .ZN(n8551) );
  OAI21_X1 U10099 ( .B1(n8748), .B2(n8852), .A(n8551), .ZN(n8552) );
  INV_X1 U10100 ( .A(n8738), .ZN(n8739) );
  INV_X1 U10101 ( .A(n8555), .ZN(n8732) );
  INV_X1 U10102 ( .A(n8556), .ZN(n8730) );
  INV_X1 U10103 ( .A(n8557), .ZN(n8558) );
  NOR2_X1 U10104 ( .A1(n8718), .A2(n8558), .ZN(n8914) );
  NAND2_X1 U10105 ( .A1(n8719), .A2(n8912), .ZN(n8919) );
  INV_X1 U10106 ( .A(n8960), .ZN(n8957) );
  AND2_X1 U10107 ( .A1(n8986), .A2(n8559), .ZN(n8693) );
  INV_X1 U10108 ( .A(n8693), .ZN(n8580) );
  XNOR2_X1 U10109 ( .A(n8560), .B(n9009), .ZN(n9017) );
  INV_X1 U10110 ( .A(n8561), .ZN(n8676) );
  NOR2_X1 U10111 ( .A1(n8562), .A2(n7463), .ZN(n8567) );
  NOR2_X1 U10112 ( .A1(n8563), .A2(n8592), .ZN(n8564) );
  NAND4_X1 U10113 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n8569)
         );
  INV_X1 U10114 ( .A(n10136), .ZN(n10127) );
  NOR3_X1 U10115 ( .A1(n8569), .A2(n10127), .A3(n8568), .ZN(n8573) );
  INV_X1 U10116 ( .A(n8571), .ZN(n8572) );
  NAND4_X1 U10117 ( .A1(n8573), .A2(n8635), .A3(n6081), .A4(n8572), .ZN(n8576)
         );
  NOR4_X1 U10118 ( .A1(n8576), .A2(n8660), .A3(n8575), .A4(n8574), .ZN(n8578)
         );
  NAND4_X1 U10119 ( .A1(n9007), .A2(n8676), .A3(n8578), .A4(n8577), .ZN(n8579)
         );
  NOR4_X1 U10120 ( .A1(n8690), .A2(n8580), .A3(n9017), .A4(n8579), .ZN(n8581)
         );
  NAND3_X1 U10121 ( .A1(n8957), .A2(n8970), .A3(n8581), .ZN(n8582) );
  NOR4_X1 U10122 ( .A1(n8919), .A2(n8931), .A3(n8945), .A4(n8582), .ZN(n8583)
         );
  NAND4_X1 U10123 ( .A1(n8879), .A2(n8725), .A3(n8914), .A4(n8583), .ZN(n8584)
         );
  NOR4_X1 U10124 ( .A1(n8739), .A2(n8585), .A3(n8871), .A4(n8584), .ZN(n8588)
         );
  INV_X1 U10125 ( .A(n8586), .ZN(n8587) );
  NAND2_X1 U10126 ( .A1(n8852), .A2(n8848), .ZN(n8743) );
  NAND4_X1 U10127 ( .A1(n8588), .A2(n8587), .A3(n8748), .A4(n8743), .ZN(n8757)
         );
  OAI21_X1 U10128 ( .B1(n8589), .B2(n4354), .A(n9029), .ZN(n8590) );
  OAI211_X1 U10129 ( .C1(n8747), .C2(n8771), .A(n8743), .B(n8590), .ZN(n8754)
         );
  MUX2_X1 U10130 ( .A(n8591), .B(n8752), .S(n4354), .Z(n8740) );
  NAND2_X1 U10131 ( .A1(n8593), .A2(n8592), .ZN(n8598) );
  NAND3_X1 U10132 ( .A1(n8598), .A2(n8595), .A3(n8594), .ZN(n8596) );
  MUX2_X1 U10133 ( .A(n8596), .B(n8595), .S(n8747), .Z(n8603) );
  NOR2_X1 U10134 ( .A1(n8598), .A2(n8597), .ZN(n8600) );
  MUX2_X1 U10135 ( .A(n4354), .B(n8600), .S(n8599), .Z(n8601) );
  INV_X1 U10136 ( .A(n8601), .ZN(n8602) );
  NAND3_X1 U10137 ( .A1(n8603), .A2(n7238), .A3(n8602), .ZN(n8610) );
  NAND2_X1 U10138 ( .A1(n8617), .A2(n8604), .ZN(n8607) );
  NAND2_X1 U10139 ( .A1(n8612), .A2(n8605), .ZN(n8606) );
  MUX2_X1 U10140 ( .A(n8607), .B(n8606), .S(n8747), .Z(n8608) );
  INV_X1 U10141 ( .A(n8608), .ZN(n8609) );
  NAND2_X1 U10142 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  NAND2_X1 U10143 ( .A1(n8611), .A2(n10136), .ZN(n8622) );
  INV_X1 U10144 ( .A(n8612), .ZN(n8614) );
  OAI211_X1 U10145 ( .C1(n8622), .C2(n8614), .A(n8623), .B(n8613), .ZN(n8616)
         );
  AND2_X1 U10146 ( .A1(n8625), .A2(n8619), .ZN(n8615) );
  AOI21_X1 U10147 ( .B1(n8616), .B2(n8615), .A(n6047), .ZN(n8630) );
  INV_X1 U10148 ( .A(n8617), .ZN(n8621) );
  NAND2_X1 U10149 ( .A1(n8618), .A2(n10162), .ZN(n8620) );
  OAI211_X1 U10150 ( .C1(n8622), .C2(n8621), .A(n8620), .B(n8619), .ZN(n8628)
         );
  AND2_X1 U10151 ( .A1(n8624), .A2(n8623), .ZN(n8627) );
  INV_X1 U10152 ( .A(n8625), .ZN(n8626) );
  AOI21_X1 U10153 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(n8629) );
  MUX2_X1 U10154 ( .A(n8630), .B(n8629), .S(n8747), .Z(n8638) );
  NAND2_X1 U10155 ( .A1(n8640), .A2(n8641), .ZN(n8634) );
  NAND2_X1 U10156 ( .A1(n8632), .A2(n8631), .ZN(n8633) );
  INV_X1 U10157 ( .A(n8635), .ZN(n8636) );
  NOR2_X1 U10158 ( .A1(n8645), .A2(n8636), .ZN(n8637) );
  NAND2_X1 U10159 ( .A1(n8638), .A2(n8637), .ZN(n8650) );
  AND2_X1 U10160 ( .A1(n8640), .A2(n8639), .ZN(n8642) );
  OAI211_X1 U10161 ( .C1(n8645), .C2(n8642), .A(n8651), .B(n8641), .ZN(n8647)
         );
  OAI21_X1 U10162 ( .B1(n8645), .B2(n8644), .A(n8643), .ZN(n8646) );
  MUX2_X1 U10163 ( .A(n8647), .B(n8646), .S(n4354), .Z(n8648) );
  INV_X1 U10164 ( .A(n8648), .ZN(n8649) );
  NAND2_X1 U10165 ( .A1(n8650), .A2(n8649), .ZN(n8659) );
  AND2_X1 U10166 ( .A1(n8656), .A2(n8651), .ZN(n8653) );
  INV_X1 U10167 ( .A(n8655), .ZN(n8652) );
  AND2_X1 U10168 ( .A1(n8655), .A2(n8654), .ZN(n8658) );
  INV_X1 U10169 ( .A(n8656), .ZN(n8657) );
  INV_X1 U10170 ( .A(n8660), .ZN(n8661) );
  AND2_X1 U10171 ( .A1(n8663), .A2(n8662), .ZN(n8665) );
  MUX2_X1 U10172 ( .A(n8665), .B(n8664), .S(n8747), .Z(n8666) );
  INV_X1 U10173 ( .A(n8666), .ZN(n8667) );
  INV_X1 U10174 ( .A(n8672), .ZN(n8675) );
  MUX2_X1 U10175 ( .A(n8670), .B(n8669), .S(n8747), .Z(n8671) );
  OAI21_X1 U10176 ( .B1(n8675), .B2(n8674), .A(n8673), .ZN(n8677) );
  NAND2_X1 U10177 ( .A1(n8677), .A2(n8676), .ZN(n8687) );
  MUX2_X1 U10178 ( .A(n8679), .B(n8678), .S(n8747), .Z(n8680) );
  NOR2_X1 U10179 ( .A1(n9017), .A2(n8680), .ZN(n8686) );
  INV_X1 U10180 ( .A(n8681), .ZN(n8682) );
  MUX2_X1 U10181 ( .A(n8683), .B(n8682), .S(n8747), .Z(n8684) );
  NAND2_X1 U10182 ( .A1(n9007), .A2(n8684), .ZN(n8685) );
  AOI21_X1 U10183 ( .B1(n8687), .B2(n8686), .A(n8685), .ZN(n8689) );
  INV_X1 U10184 ( .A(n8690), .ZN(n8691) );
  NAND2_X1 U10185 ( .A1(n8695), .A2(n8691), .ZN(n8692) );
  NAND2_X1 U10186 ( .A1(n8692), .A2(n8986), .ZN(n8696) );
  OAI211_X1 U10187 ( .C1(n8709), .C2(n8698), .A(n8710), .B(n8697), .ZN(n8699)
         );
  NAND3_X1 U10188 ( .A1(n8699), .A2(n8713), .A3(n8708), .ZN(n8700) );
  NAND2_X1 U10189 ( .A1(n8700), .A2(n8711), .ZN(n8701) );
  NOR2_X1 U10190 ( .A1(n8702), .A2(n8747), .ZN(n8703) );
  NAND2_X1 U10191 ( .A1(n8721), .A2(n8703), .ZN(n8705) );
  NAND4_X1 U10192 ( .A1(n8719), .A2(n8747), .A3(n8921), .A4(n8938), .ZN(n8704)
         );
  OAI211_X1 U10193 ( .C1(n8721), .C2(n4354), .A(n8705), .B(n8704), .ZN(n8706)
         );
  INV_X1 U10194 ( .A(n8706), .ZN(n8717) );
  NAND3_X1 U10195 ( .A1(n8709), .A2(n8708), .A3(n8707), .ZN(n8712) );
  NAND3_X1 U10196 ( .A1(n8712), .A2(n8711), .A3(n8710), .ZN(n8714) );
  NAND2_X1 U10197 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  NAND4_X1 U10198 ( .A1(n8715), .A2(n8747), .A3(n8939), .A4(n8719), .ZN(n8716)
         );
  INV_X1 U10199 ( .A(n8718), .ZN(n8724) );
  INV_X1 U10200 ( .A(n8719), .ZN(n8720) );
  NAND2_X1 U10201 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  AOI21_X1 U10202 ( .B1(n8722), .B2(n8724), .A(n8747), .ZN(n8723) );
  MUX2_X1 U10203 ( .A(n8727), .B(n8726), .S(n8747), .Z(n8728) );
  MUX2_X1 U10204 ( .A(n8730), .B(n8729), .S(n8747), .Z(n8731) );
  NOR2_X1 U10205 ( .A1(n8871), .A2(n8731), .ZN(n8735) );
  MUX2_X1 U10206 ( .A(n8733), .B(n8732), .S(n4354), .Z(n8734) );
  AOI21_X1 U10207 ( .B1(n8736), .B2(n8735), .A(n8734), .ZN(n8737) );
  INV_X1 U10208 ( .A(n8751), .ZN(n8745) );
  INV_X1 U10209 ( .A(n8741), .ZN(n8742) );
  NOR2_X1 U10210 ( .A1(n8749), .A2(n8742), .ZN(n8744) );
  OAI211_X1 U10211 ( .C1(n8745), .C2(n8873), .A(n8744), .B(n8743), .ZN(n8753)
         );
  NAND3_X1 U10212 ( .A1(n8748), .A2(n8747), .A3(n8746), .ZN(n8750) );
  INV_X1 U10213 ( .A(n8848), .ZN(n8758) );
  XNOR2_X1 U10214 ( .A(n8763), .B(n8762), .ZN(n8770) );
  NAND3_X1 U10215 ( .A1(n8765), .A2(n8764), .A3(n8806), .ZN(n8766) );
  OAI211_X1 U10216 ( .C1(n8767), .C2(n8769), .A(n8766), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8768) );
  OAI21_X1 U10217 ( .B1(n8770), .B2(n8769), .A(n8768), .ZN(P2_U3296) );
  MUX2_X1 U10218 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8848), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10219 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8771), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10220 ( .A(n8772), .ZN(n8860) );
  MUX2_X1 U10221 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8860), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10222 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8873), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10223 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8883), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10224 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8895), .S(P2_U3893), .Z(
        P2_U3517) );
  INV_X1 U10225 ( .A(n8773), .ZN(n8906) );
  MUX2_X1 U10226 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8906), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10227 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8894), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10228 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8932), .S(P2_U3893), .Z(
        P2_U3514) );
  INV_X1 U10229 ( .A(n8921), .ZN(n8950) );
  MUX2_X1 U10230 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8950), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10231 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8962), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10232 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8951), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10233 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8991), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10234 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9000), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10235 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9008), .S(P2_U3893), .Z(
        P2_U3508) );
  INV_X1 U10236 ( .A(n8774), .ZN(n9020) );
  MUX2_X1 U10237 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9020), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10238 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9009), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10239 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9019), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10240 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8775), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10241 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8776), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10242 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8777), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10243 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8778), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10244 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8779), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10245 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8780), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10246 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8781), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10247 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n10130), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10248 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8782), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10249 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8783), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10250 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8784), .S(P2_U3893), .Z(
        P2_U3491) );
  NOR2_X1 U10251 ( .A1(n10042), .A2(n8786), .ZN(n8787) );
  INV_X1 U10252 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U10253 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8826), .ZN(n8788) );
  OAI21_X1 U10254 ( .B1(n8826), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8788), .ZN(
        n10068) );
  NOR2_X1 U10255 ( .A1(n10074), .A2(n8789), .ZN(n8790) );
  NAND2_X1 U10256 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8824), .ZN(n8791) );
  OAI21_X1 U10257 ( .B1(n8824), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8791), .ZN(
        n10100) );
  NOR2_X1 U10258 ( .A1(n10108), .A2(n8792), .ZN(n8793) );
  INV_X1 U10259 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8794) );
  AOI22_X1 U10260 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n9805), .B1(n9803), .B2(
        n8794), .ZN(n9795) );
  AOI21_X1 U10261 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n9803), .A(n9794), .ZN(
        n8795) );
  MUX2_X1 U10262 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8979), .S(n4353), .Z(n8816) );
  NOR2_X1 U10263 ( .A1(n8795), .A2(n8816), .ZN(n8846) );
  INV_X1 U10264 ( .A(n8816), .ZN(n8812) );
  OAI21_X1 U10265 ( .B1(n9794), .B2(n8812), .A(n10010), .ZN(n8845) );
  MUX2_X1 U10266 ( .A(n10119), .B(n9068), .S(n8799), .Z(n8805) );
  XNOR2_X1 U10267 ( .A(n8836), .B(n8805), .ZN(n10113) );
  MUX2_X1 U10268 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8799), .Z(n8796) );
  OR2_X1 U10269 ( .A1(n8796), .A2(n8824), .ZN(n8804) );
  XNOR2_X1 U10270 ( .A(n8796), .B(n10090), .ZN(n10096) );
  MUX2_X1 U10271 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8799), .Z(n8797) );
  OR2_X1 U10272 ( .A1(n8797), .A2(n4730), .ZN(n8803) );
  XNOR2_X1 U10273 ( .A(n8797), .B(n10074), .ZN(n10079) );
  MUX2_X1 U10274 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8799), .Z(n8798) );
  OR2_X1 U10275 ( .A1(n8798), .A2(n8826), .ZN(n8802) );
  XNOR2_X1 U10276 ( .A(n8798), .B(n10058), .ZN(n10064) );
  MUX2_X1 U10277 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8799), .Z(n8801) );
  XNOR2_X1 U10278 ( .A(n8801), .B(n10042), .ZN(n10047) );
  NAND2_X1 U10279 ( .A1(n10064), .A2(n10063), .ZN(n10062) );
  NAND2_X1 U10280 ( .A1(n8804), .A2(n10094), .ZN(n10112) );
  MUX2_X1 U10281 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8806), .Z(n8809) );
  INV_X1 U10282 ( .A(n8809), .ZN(n8807) );
  NAND2_X1 U10283 ( .A1(n8808), .A2(n8807), .ZN(n9784) );
  AND2_X1 U10284 ( .A1(n8810), .A2(n8809), .ZN(n9786) );
  AOI21_X1 U10285 ( .B1(n9803), .B2(n9784), .A(n9786), .ZN(n8813) );
  XNOR2_X1 U10286 ( .A(n4353), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8839) );
  MUX2_X1 U10287 ( .A(n8839), .B(n8812), .S(n8811), .Z(n8817) );
  INV_X1 U10288 ( .A(n9786), .ZN(n8814) );
  NAND3_X1 U10289 ( .A1(n10115), .A2(n8817), .A3(n9784), .ZN(n8819) );
  INV_X1 U10290 ( .A(n8839), .ZN(n8843) );
  NAND3_X1 U10291 ( .A1(n10116), .A2(P2_REG1_REG_18__SCAN_IN), .A3(n8843), 
        .ZN(n8818) );
  NAND2_X1 U10292 ( .A1(n10106), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8821) );
  OAI211_X1 U10293 ( .C1(n10027), .C2(n4353), .A(n8821), .B(n8820), .ZN(n8823)
         );
  AOI22_X1 U10294 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n9803), .B1(n9805), .B2(
        n9065), .ZN(n9791) );
  AOI22_X1 U10295 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8824), .B1(n10090), 
        .B2(n9071), .ZN(n10093) );
  NAND2_X1 U10296 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8826), .ZN(n8833) );
  AOI22_X1 U10297 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8826), .B1(n10058), 
        .B2(n8825), .ZN(n10061) );
  NAND2_X1 U10298 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8827), .ZN(n8829) );
  NAND2_X1 U10299 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  NAND2_X1 U10300 ( .A1(n8830), .A2(n8831), .ZN(n8832) );
  XOR2_X1 U10301 ( .A(n8831), .B(n8830), .Z(n10044) );
  NAND2_X1 U10302 ( .A1(n10061), .A2(n10060), .ZN(n10059) );
  NAND2_X1 U10303 ( .A1(n4730), .A2(n8834), .ZN(n8835) );
  XNOR2_X1 U10304 ( .A(n10074), .B(n8834), .ZN(n10076) );
  NAND2_X1 U10305 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10076), .ZN(n10075) );
  NAND2_X1 U10306 ( .A1(n8835), .A2(n10075), .ZN(n10092) );
  NAND2_X1 U10307 ( .A1(n10093), .A2(n10092), .ZN(n10091) );
  NAND2_X1 U10308 ( .A1(n8836), .A2(n8837), .ZN(n8838) );
  XNOR2_X1 U10309 ( .A(n10108), .B(n8837), .ZN(n10110) );
  NAND2_X1 U10310 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n10110), .ZN(n10109) );
  OAI21_X1 U10311 ( .B1(n9805), .B2(n9065), .A(n8839), .ZN(n8841) );
  AOI21_X1 U10312 ( .B1(n9789), .B2(n8841), .A(n8840), .ZN(n8842) );
  OAI21_X1 U10313 ( .B1(n9789), .B2(n8843), .A(n8842), .ZN(n8844) );
  NAND2_X1 U10314 ( .A1(n10146), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8851) );
  AND2_X1 U10315 ( .A1(n8848), .A2(n8847), .ZN(n9081) );
  AND2_X1 U10316 ( .A1(n8849), .A2(n10140), .ZN(n8850) );
  OAI21_X1 U10317 ( .B1(n9081), .B2(n8850), .A(n10145), .ZN(n8853) );
  OAI211_X1 U10318 ( .C1(n8852), .C2(n8855), .A(n8851), .B(n8853), .ZN(
        P2_U3202) );
  NAND2_X1 U10319 ( .A1(n10146), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8854) );
  OAI211_X1 U10320 ( .C1(n9086), .C2(n8855), .A(n8854), .B(n8853), .ZN(
        P2_U3203) );
  XNOR2_X1 U10321 ( .A(n8859), .B(n8858), .ZN(n8864) );
  AOI21_X1 U10322 ( .B1(n8864), .B2(n10134), .A(n8863), .ZN(n9087) );
  MUX2_X1 U10323 ( .A(n8865), .B(n9087), .S(n10145), .Z(n8869) );
  INV_X1 U10324 ( .A(n8866), .ZN(n8867) );
  AOI22_X1 U10325 ( .A1(n9089), .A2(n10138), .B1(n10140), .B2(n8867), .ZN(
        n8868) );
  OAI211_X1 U10326 ( .C1(n9092), .C2(n9026), .A(n8869), .B(n8868), .ZN(
        P2_U3205) );
  XNOR2_X1 U10327 ( .A(n8870), .B(n8871), .ZN(n9098) );
  INV_X1 U10328 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8875) );
  XNOR2_X1 U10329 ( .A(n8872), .B(n8871), .ZN(n8874) );
  AOI222_X1 U10330 ( .A1(n10134), .A2(n8874), .B1(n8895), .B2(n10129), .C1(
        n8873), .C2(n10131), .ZN(n9093) );
  MUX2_X1 U10331 ( .A(n8875), .B(n9093), .S(n10145), .Z(n8878) );
  AOI22_X1 U10332 ( .A1(n9095), .A2(n10138), .B1(n10140), .B2(n8876), .ZN(
        n8877) );
  OAI211_X1 U10333 ( .C1(n9098), .C2(n9026), .A(n8878), .B(n8877), .ZN(
        P2_U3206) );
  XNOR2_X1 U10334 ( .A(n8880), .B(n8879), .ZN(n9104) );
  INV_X1 U10335 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8885) );
  XNOR2_X1 U10336 ( .A(n8882), .B(n8881), .ZN(n8884) );
  AOI222_X1 U10337 ( .A1(n10134), .A2(n8884), .B1(n8883), .B2(n10131), .C1(
        n8906), .C2(n10129), .ZN(n9099) );
  MUX2_X1 U10338 ( .A(n8885), .B(n9099), .S(n10145), .Z(n8888) );
  AOI22_X1 U10339 ( .A1(n9101), .A2(n10138), .B1(n10140), .B2(n8886), .ZN(
        n8887) );
  OAI211_X1 U10340 ( .C1(n9104), .C2(n9026), .A(n8888), .B(n8887), .ZN(
        P2_U3207) );
  XNOR2_X1 U10341 ( .A(n8889), .B(n8892), .ZN(n9110) );
  INV_X1 U10342 ( .A(n8890), .ZN(n8893) );
  OAI21_X1 U10343 ( .B1(n8893), .B2(n8892), .A(n8891), .ZN(n8896) );
  AOI222_X1 U10344 ( .A1(n10134), .A2(n8896), .B1(n8895), .B2(n10131), .C1(
        n8894), .C2(n10129), .ZN(n9105) );
  INV_X1 U10345 ( .A(n9105), .ZN(n8902) );
  INV_X1 U10346 ( .A(n8897), .ZN(n8898) );
  OAI22_X1 U10347 ( .A1(n8900), .A2(n8899), .B1(n8898), .B2(n8977), .ZN(n8901)
         );
  OAI21_X1 U10348 ( .B1(n8902), .B2(n8901), .A(n10145), .ZN(n8904) );
  NAND2_X1 U10349 ( .A1(n10146), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8903) );
  OAI211_X1 U10350 ( .C1(n9110), .C2(n9026), .A(n8904), .B(n8903), .ZN(
        P2_U3208) );
  XOR2_X1 U10351 ( .A(n8914), .B(n8905), .Z(n8907) );
  AOI222_X1 U10352 ( .A1(n10134), .A2(n8907), .B1(n8906), .B2(n10131), .C1(
        n8932), .C2(n10129), .ZN(n9111) );
  AOI22_X1 U10353 ( .A1(n9113), .A2(n8909), .B1(n10140), .B2(n8908), .ZN(n8910) );
  AOI21_X1 U10354 ( .B1(n9111), .B2(n8910), .A(n10146), .ZN(n8917) );
  NAND2_X1 U10355 ( .A1(n8911), .A2(n8912), .ZN(n8913) );
  XOR2_X1 U10356 ( .A(n8914), .B(n8913), .Z(n9116) );
  OAI22_X1 U10357 ( .A1(n9116), .A2(n9026), .B1(n8915), .B2(n10145), .ZN(n8916) );
  OR2_X1 U10358 ( .A1(n8917), .A2(n8916), .ZN(P2_U3209) );
  XNOR2_X1 U10359 ( .A(n4405), .B(n8919), .ZN(n9120) );
  INV_X1 U10360 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8924) );
  XOR2_X1 U10361 ( .A(n8919), .B(n8918), .Z(n8920) );
  OAI222_X1 U10362 ( .A1(n8976), .A2(n8922), .B1(n8974), .B2(n8921), .C1(n8972), .C2(n8920), .ZN(n9117) );
  INV_X1 U10363 ( .A(n9117), .ZN(n8923) );
  MUX2_X1 U10364 ( .A(n8924), .B(n8923), .S(n10145), .Z(n8928) );
  AOI22_X1 U10365 ( .A1(n8926), .A2(n10138), .B1(n10140), .B2(n8925), .ZN(
        n8927) );
  OAI211_X1 U10366 ( .C1(n9120), .C2(n9026), .A(n8928), .B(n8927), .ZN(
        P2_U3210) );
  OAI21_X1 U10367 ( .B1(n8931), .B2(n8930), .A(n8929), .ZN(n8933) );
  AOI222_X1 U10368 ( .A1(n10134), .A2(n8933), .B1(n8932), .B2(n10131), .C1(
        n8962), .C2(n10129), .ZN(n9053) );
  INV_X1 U10369 ( .A(n8934), .ZN(n8935) );
  OAI22_X1 U10370 ( .A1(n10145), .A2(n8936), .B1(n8935), .B2(n8977), .ZN(n8937) );
  AOI21_X1 U10371 ( .B1(n8938), .B2(n10138), .A(n8937), .ZN(n8943) );
  OR2_X1 U10372 ( .A1(n8940), .A2(n8939), .ZN(n9051) );
  NAND3_X1 U10373 ( .A1(n9051), .A2(n8941), .A3(n10142), .ZN(n8942) );
  OAI211_X1 U10374 ( .C1(n9053), .C2(n10146), .A(n8943), .B(n8942), .ZN(
        P2_U3211) );
  XNOR2_X1 U10375 ( .A(n8944), .B(n8945), .ZN(n9129) );
  INV_X1 U10376 ( .A(n8945), .ZN(n8947) );
  NAND3_X1 U10377 ( .A1(n8959), .A2(n8947), .A3(n8946), .ZN(n8948) );
  NAND2_X1 U10378 ( .A1(n8949), .A2(n8948), .ZN(n8952) );
  AOI222_X1 U10379 ( .A1(n10134), .A2(n8952), .B1(n8951), .B2(n10129), .C1(
        n8950), .C2(n10131), .ZN(n9124) );
  MUX2_X1 U10380 ( .A(n8953), .B(n9124), .S(n10145), .Z(n8956) );
  AOI22_X1 U10381 ( .A1(n9126), .A2(n10138), .B1(n10140), .B2(n8954), .ZN(
        n8955) );
  OAI211_X1 U10382 ( .C1(n9129), .C2(n9026), .A(n8956), .B(n8955), .ZN(
        P2_U3212) );
  XNOR2_X1 U10383 ( .A(n8958), .B(n8957), .ZN(n9135) );
  OAI21_X1 U10384 ( .B1(n8961), .B2(n8960), .A(n8959), .ZN(n8963) );
  AOI222_X1 U10385 ( .A1(n10134), .A2(n8963), .B1(n8962), .B2(n10131), .C1(
        n8991), .C2(n10129), .ZN(n9130) );
  MUX2_X1 U10386 ( .A(n8964), .B(n9130), .S(n10145), .Z(n8967) );
  AOI22_X1 U10387 ( .A1(n9132), .A2(n10138), .B1(n10140), .B2(n8965), .ZN(
        n8966) );
  OAI211_X1 U10388 ( .C1(n9135), .C2(n9026), .A(n8967), .B(n8966), .ZN(
        P2_U3213) );
  XOR2_X1 U10389 ( .A(n8970), .B(n8968), .Z(n9139) );
  XOR2_X1 U10390 ( .A(n8970), .B(n8969), .Z(n8971) );
  OAI222_X1 U10391 ( .A1(n8976), .A2(n8975), .B1(n8974), .B2(n8973), .C1(n8972), .C2(n8971), .ZN(n9061) );
  NAND2_X1 U10392 ( .A1(n9061), .A2(n10145), .ZN(n8982) );
  OAI22_X1 U10393 ( .A1(n10145), .A2(n8979), .B1(n8978), .B2(n8977), .ZN(n8980) );
  AOI21_X1 U10394 ( .B1(n9062), .B2(n10138), .A(n8980), .ZN(n8981) );
  OAI211_X1 U10395 ( .C1(n9139), .C2(n9026), .A(n8982), .B(n8981), .ZN(
        P2_U3214) );
  INV_X1 U10396 ( .A(n8983), .ZN(n8984) );
  NOR2_X1 U10397 ( .A1(n8985), .A2(n8984), .ZN(n8988) );
  NAND2_X1 U10398 ( .A1(n8987), .A2(n8986), .ZN(n8989) );
  XNOR2_X1 U10399 ( .A(n8988), .B(n8989), .ZN(n9145) );
  XNOR2_X1 U10400 ( .A(n8990), .B(n8989), .ZN(n8992) );
  AOI222_X1 U10401 ( .A1(n10134), .A2(n8992), .B1(n8991), .B2(n10131), .C1(
        n9008), .C2(n10129), .ZN(n9140) );
  MUX2_X1 U10402 ( .A(n8794), .B(n9140), .S(n10145), .Z(n8996) );
  INV_X1 U10403 ( .A(n8993), .ZN(n8994) );
  AOI22_X1 U10404 ( .A1(n9142), .A2(n10138), .B1(n10140), .B2(n8994), .ZN(
        n8995) );
  OAI211_X1 U10405 ( .C1(n9145), .C2(n9026), .A(n8996), .B(n8995), .ZN(
        P2_U3215) );
  XNOR2_X1 U10406 ( .A(n8997), .B(n8999), .ZN(n9151) );
  XOR2_X1 U10407 ( .A(n8999), .B(n8998), .Z(n9001) );
  AOI222_X1 U10408 ( .A1(n10134), .A2(n9001), .B1(n9000), .B2(n10131), .C1(
        n9020), .C2(n10129), .ZN(n9146) );
  MUX2_X1 U10409 ( .A(n10119), .B(n9146), .S(n10145), .Z(n9004) );
  AOI22_X1 U10410 ( .A1(n9148), .A2(n10138), .B1(n10140), .B2(n9002), .ZN(
        n9003) );
  OAI211_X1 U10411 ( .C1(n9151), .C2(n9026), .A(n9004), .B(n9003), .ZN(
        P2_U3216) );
  XNOR2_X1 U10412 ( .A(n9005), .B(n9007), .ZN(n9157) );
  XOR2_X1 U10413 ( .A(n9007), .B(n9006), .Z(n9010) );
  AOI222_X1 U10414 ( .A1(n10134), .A2(n9010), .B1(n9009), .B2(n10129), .C1(
        n9008), .C2(n10131), .ZN(n9152) );
  MUX2_X1 U10415 ( .A(n9011), .B(n9152), .S(n10145), .Z(n9015) );
  INV_X1 U10416 ( .A(n9012), .ZN(n9013) );
  AOI22_X1 U10417 ( .A1(n9154), .A2(n10138), .B1(n10140), .B2(n9013), .ZN(
        n9014) );
  OAI211_X1 U10418 ( .C1(n9157), .C2(n9026), .A(n9015), .B(n9014), .ZN(
        P2_U3217) );
  XNOR2_X1 U10419 ( .A(n9016), .B(n9017), .ZN(n9165) );
  XNOR2_X1 U10420 ( .A(n9018), .B(n9017), .ZN(n9021) );
  AOI222_X1 U10421 ( .A1(n10134), .A2(n9021), .B1(n9020), .B2(n10131), .C1(
        n9019), .C2(n10129), .ZN(n9158) );
  MUX2_X1 U10422 ( .A(n10083), .B(n9158), .S(n10145), .Z(n9025) );
  INV_X1 U10423 ( .A(n9022), .ZN(n9023) );
  AOI22_X1 U10424 ( .A1(n9160), .A2(n10138), .B1(n10140), .B2(n9023), .ZN(
        n9024) );
  OAI211_X1 U10425 ( .C1(n9165), .C2(n9026), .A(n9025), .B(n9024), .ZN(
        P2_U3218) );
  INV_X1 U10426 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U10427 ( .A1(n9080), .A2(n9075), .ZN(n9027) );
  NAND2_X1 U10428 ( .A1(n10225), .A2(n9081), .ZN(n9030) );
  OAI211_X1 U10429 ( .C1(n10225), .C2(n9028), .A(n9027), .B(n9030), .ZN(
        P2_U3490) );
  INV_X1 U10430 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U10431 ( .A1(n9029), .A2(n9075), .ZN(n9031) );
  OAI211_X1 U10432 ( .C1(n10225), .C2(n9032), .A(n9031), .B(n9030), .ZN(
        P2_U3489) );
  INV_X1 U10433 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9033) );
  MUX2_X1 U10434 ( .A(n9033), .B(n9087), .S(n10225), .Z(n9035) );
  NAND2_X1 U10435 ( .A1(n9089), .A2(n9075), .ZN(n9034) );
  OAI211_X1 U10436 ( .C1(n9092), .C2(n9078), .A(n9035), .B(n9034), .ZN(
        P2_U3487) );
  MUX2_X1 U10437 ( .A(n9036), .B(n9093), .S(n10225), .Z(n9038) );
  NAND2_X1 U10438 ( .A1(n9095), .A2(n9075), .ZN(n9037) );
  OAI211_X1 U10439 ( .C1(n9078), .C2(n9098), .A(n9038), .B(n9037), .ZN(
        P2_U3486) );
  MUX2_X1 U10440 ( .A(n9039), .B(n9099), .S(n10225), .Z(n9041) );
  NAND2_X1 U10441 ( .A1(n9101), .A2(n9075), .ZN(n9040) );
  OAI211_X1 U10442 ( .C1(n9104), .C2(n9078), .A(n9041), .B(n9040), .ZN(
        P2_U3485) );
  INV_X1 U10443 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9042) );
  MUX2_X1 U10444 ( .A(n9042), .B(n9105), .S(n10225), .Z(n9044) );
  NAND2_X1 U10445 ( .A1(n9107), .A2(n9075), .ZN(n9043) );
  OAI211_X1 U10446 ( .C1(n9110), .C2(n9078), .A(n9044), .B(n9043), .ZN(
        P2_U3484) );
  INV_X1 U10447 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9045) );
  MUX2_X1 U10448 ( .A(n9045), .B(n9111), .S(n10225), .Z(n9047) );
  NAND2_X1 U10449 ( .A1(n9113), .A2(n9075), .ZN(n9046) );
  OAI211_X1 U10450 ( .C1(n9078), .C2(n9116), .A(n9047), .B(n9046), .ZN(
        P2_U3483) );
  MUX2_X1 U10451 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9117), .S(n10225), .Z(
        n9050) );
  OAI22_X1 U10452 ( .A1(n9120), .A2(n9078), .B1(n9119), .B2(n9048), .ZN(n9049)
         );
  OR2_X1 U10453 ( .A1(n9050), .A2(n9049), .ZN(P2_U3482) );
  NAND3_X1 U10454 ( .A1(n9051), .A2(n8941), .A3(n10198), .ZN(n9052) );
  OAI211_X1 U10455 ( .C1(n9054), .C2(n10186), .A(n9053), .B(n9052), .ZN(n9123)
         );
  MUX2_X1 U10456 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9123), .S(n10225), .Z(
        P2_U3481) );
  MUX2_X1 U10457 ( .A(n9055), .B(n9124), .S(n10225), .Z(n9057) );
  NAND2_X1 U10458 ( .A1(n9126), .A2(n9075), .ZN(n9056) );
  OAI211_X1 U10459 ( .C1(n9078), .C2(n9129), .A(n9057), .B(n9056), .ZN(
        P2_U3480) );
  INV_X1 U10460 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9058) );
  MUX2_X1 U10461 ( .A(n9058), .B(n9130), .S(n10225), .Z(n9060) );
  NAND2_X1 U10462 ( .A1(n9132), .A2(n9075), .ZN(n9059) );
  OAI211_X1 U10463 ( .C1(n9078), .C2(n9135), .A(n9060), .B(n9059), .ZN(
        P2_U3479) );
  AOI21_X1 U10464 ( .B1(n10200), .B2(n9062), .A(n9061), .ZN(n9136) );
  MUX2_X1 U10465 ( .A(n9063), .B(n9136), .S(n10225), .Z(n9064) );
  OAI21_X1 U10466 ( .B1(n9078), .B2(n9139), .A(n9064), .ZN(P2_U3478) );
  MUX2_X1 U10467 ( .A(n9065), .B(n9140), .S(n10225), .Z(n9067) );
  NAND2_X1 U10468 ( .A1(n9142), .A2(n9075), .ZN(n9066) );
  OAI211_X1 U10469 ( .C1(n9145), .C2(n9078), .A(n9067), .B(n9066), .ZN(
        P2_U3477) );
  MUX2_X1 U10470 ( .A(n9068), .B(n9146), .S(n10225), .Z(n9070) );
  NAND2_X1 U10471 ( .A1(n9148), .A2(n9075), .ZN(n9069) );
  OAI211_X1 U10472 ( .C1(n9151), .C2(n9078), .A(n9070), .B(n9069), .ZN(
        P2_U3476) );
  MUX2_X1 U10473 ( .A(n9071), .B(n9152), .S(n10225), .Z(n9073) );
  NAND2_X1 U10474 ( .A1(n9154), .A2(n9075), .ZN(n9072) );
  OAI211_X1 U10475 ( .C1(n9157), .C2(n9078), .A(n9073), .B(n9072), .ZN(
        P2_U3475) );
  MUX2_X1 U10476 ( .A(n9074), .B(n9158), .S(n10225), .Z(n9077) );
  NAND2_X1 U10477 ( .A1(n9160), .A2(n9075), .ZN(n9076) );
  OAI211_X1 U10478 ( .C1(n9165), .C2(n9078), .A(n9077), .B(n9076), .ZN(
        P2_U3474) );
  MUX2_X1 U10479 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9079), .S(n10225), .Z(
        P2_U3459) );
  INV_X1 U10480 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U10481 ( .A1(n9080), .A2(n9161), .ZN(n9082) );
  NAND2_X1 U10482 ( .A1(n10205), .A2(n9081), .ZN(n9084) );
  OAI211_X1 U10483 ( .C1(n9083), .C2(n10205), .A(n9082), .B(n9084), .ZN(
        P2_U3458) );
  NAND2_X1 U10484 ( .A1(n10207), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9085) );
  OAI211_X1 U10485 ( .C1(n9086), .C2(n9118), .A(n9085), .B(n9084), .ZN(
        P2_U3457) );
  MUX2_X1 U10486 ( .A(n9088), .B(n9087), .S(n10205), .Z(n9091) );
  NAND2_X1 U10487 ( .A1(n9089), .A2(n9161), .ZN(n9090) );
  OAI211_X1 U10488 ( .C1(n9092), .C2(n9164), .A(n9091), .B(n9090), .ZN(
        P2_U3455) );
  INV_X1 U10489 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9094) );
  MUX2_X1 U10490 ( .A(n9094), .B(n9093), .S(n10205), .Z(n9097) );
  NAND2_X1 U10491 ( .A1(n9095), .A2(n9161), .ZN(n9096) );
  OAI211_X1 U10492 ( .C1(n9098), .C2(n9164), .A(n9097), .B(n9096), .ZN(
        P2_U3454) );
  INV_X1 U10493 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9100) );
  MUX2_X1 U10494 ( .A(n9100), .B(n9099), .S(n10205), .Z(n9103) );
  NAND2_X1 U10495 ( .A1(n9101), .A2(n9161), .ZN(n9102) );
  OAI211_X1 U10496 ( .C1(n9104), .C2(n9164), .A(n9103), .B(n9102), .ZN(
        P2_U3453) );
  INV_X1 U10497 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9106) );
  MUX2_X1 U10498 ( .A(n9106), .B(n9105), .S(n10205), .Z(n9109) );
  NAND2_X1 U10499 ( .A1(n9107), .A2(n9161), .ZN(n9108) );
  OAI211_X1 U10500 ( .C1(n9110), .C2(n9164), .A(n9109), .B(n9108), .ZN(
        P2_U3452) );
  INV_X1 U10501 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9112) );
  MUX2_X1 U10502 ( .A(n9112), .B(n9111), .S(n10205), .Z(n9115) );
  NAND2_X1 U10503 ( .A1(n9113), .A2(n9161), .ZN(n9114) );
  OAI211_X1 U10504 ( .C1(n9116), .C2(n9164), .A(n9115), .B(n9114), .ZN(
        P2_U3451) );
  MUX2_X1 U10505 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9117), .S(n10205), .Z(
        n9122) );
  OAI22_X1 U10506 ( .A1(n9120), .A2(n9164), .B1(n9119), .B2(n9118), .ZN(n9121)
         );
  OR2_X1 U10507 ( .A1(n9122), .A2(n9121), .ZN(P2_U3450) );
  MUX2_X1 U10508 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9123), .S(n10205), .Z(
        P2_U3449) );
  MUX2_X1 U10509 ( .A(n9125), .B(n9124), .S(n10205), .Z(n9128) );
  NAND2_X1 U10510 ( .A1(n9126), .A2(n9161), .ZN(n9127) );
  OAI211_X1 U10511 ( .C1(n9129), .C2(n9164), .A(n9128), .B(n9127), .ZN(
        P2_U3448) );
  MUX2_X1 U10512 ( .A(n9131), .B(n9130), .S(n10205), .Z(n9134) );
  NAND2_X1 U10513 ( .A1(n9132), .A2(n9161), .ZN(n9133) );
  OAI211_X1 U10514 ( .C1(n9135), .C2(n9164), .A(n9134), .B(n9133), .ZN(
        P2_U3447) );
  INV_X1 U10515 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9137) );
  MUX2_X1 U10516 ( .A(n9137), .B(n9136), .S(n10205), .Z(n9138) );
  OAI21_X1 U10517 ( .B1(n9139), .B2(n9164), .A(n9138), .ZN(P2_U3446) );
  INV_X1 U10518 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U10519 ( .A(n9141), .B(n9140), .S(n10205), .Z(n9144) );
  NAND2_X1 U10520 ( .A1(n9142), .A2(n9161), .ZN(n9143) );
  OAI211_X1 U10521 ( .C1(n9145), .C2(n9164), .A(n9144), .B(n9143), .ZN(
        P2_U3444) );
  INV_X1 U10522 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9147) );
  MUX2_X1 U10523 ( .A(n9147), .B(n9146), .S(n10205), .Z(n9150) );
  NAND2_X1 U10524 ( .A1(n9148), .A2(n9161), .ZN(n9149) );
  OAI211_X1 U10525 ( .C1(n9151), .C2(n9164), .A(n9150), .B(n9149), .ZN(
        P2_U3441) );
  INV_X1 U10526 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9153) );
  MUX2_X1 U10527 ( .A(n9153), .B(n9152), .S(n10205), .Z(n9156) );
  NAND2_X1 U10528 ( .A1(n9154), .A2(n9161), .ZN(n9155) );
  OAI211_X1 U10529 ( .C1(n9157), .C2(n9164), .A(n9156), .B(n9155), .ZN(
        P2_U3438) );
  INV_X1 U10530 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9159) );
  MUX2_X1 U10531 ( .A(n9159), .B(n9158), .S(n10205), .Z(n9163) );
  NAND2_X1 U10532 ( .A1(n9161), .A2(n9160), .ZN(n9162) );
  OAI211_X1 U10533 ( .C1(n9165), .C2(n9164), .A(n9163), .B(n9162), .ZN(
        P2_U3435) );
  INV_X1 U10534 ( .A(n9781), .ZN(n9171) );
  NOR4_X1 U10535 ( .A1(n9167), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9166), .ZN(n9168) );
  AOI21_X1 U10536 ( .B1(n9169), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9168), .ZN(
        n9170) );
  OAI21_X1 U10537 ( .B1(n9171), .B2(n9175), .A(n9170), .ZN(P2_U3264) );
  OAI222_X1 U10538 ( .A1(P2_U3151), .A2(n9176), .B1(n9175), .B2(n9174), .C1(
        n9173), .C2(n9172), .ZN(P2_U3266) );
  MUX2_X1 U10539 ( .A(n9178), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10540 ( .A(n9562), .ZN(n9752) );
  INV_X1 U10541 ( .A(n9225), .ZN(n9181) );
  NOR3_X1 U10542 ( .A1(n9242), .A2(n9246), .A3(n9179), .ZN(n9180) );
  OAI21_X1 U10543 ( .B1(n9181), .B2(n9180), .A(n9274), .ZN(n9186) );
  AOI22_X1 U10544 ( .A1(n9560), .A2(n9250), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9182) );
  OAI21_X1 U10545 ( .B1(n9183), .B2(n9252), .A(n9182), .ZN(n9184) );
  AOI21_X1 U10546 ( .B1(n9555), .B2(n9282), .A(n9184), .ZN(n9185) );
  OAI211_X1 U10547 ( .C1(n9752), .C2(n9285), .A(n9186), .B(n9185), .ZN(
        P1_U3216) );
  NAND2_X1 U10548 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  XNOR2_X1 U10549 ( .A(n9187), .B(n9190), .ZN(n9195) );
  AND2_X1 U10550 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9455) );
  AOI21_X1 U10551 ( .B1(n9645), .B2(n9250), .A(n9455), .ZN(n9192) );
  NAND2_X1 U10552 ( .A1(n9277), .A2(n9642), .ZN(n9191) );
  OAI211_X1 U10553 ( .C1(n9260), .C2(n9631), .A(n9192), .B(n9191), .ZN(n9193)
         );
  AOI21_X1 U10554 ( .B1(n9628), .B2(n9265), .A(n9193), .ZN(n9194) );
  OAI21_X1 U10555 ( .B1(n9195), .B2(n9267), .A(n9194), .ZN(P1_U3219) );
  XOR2_X1 U10556 ( .A(n9197), .B(n9196), .Z(n9202) );
  AOI22_X1 U10557 ( .A1(n9593), .A2(n9250), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9199) );
  NAND2_X1 U10558 ( .A1(n9645), .A2(n9277), .ZN(n9198) );
  OAI211_X1 U10559 ( .C1(n9260), .C2(n9598), .A(n9199), .B(n9198), .ZN(n9200)
         );
  AOI21_X1 U10560 ( .B1(n9597), .B2(n9265), .A(n9200), .ZN(n9201) );
  OAI21_X1 U10561 ( .B1(n9202), .B2(n9267), .A(n9201), .ZN(P1_U3223) );
  AOI21_X1 U10562 ( .B1(n4396), .B2(n9203), .A(n9272), .ZN(n9209) );
  AOI22_X1 U10563 ( .A1(n9524), .A2(n9250), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9205) );
  NAND2_X1 U10564 ( .A1(n9530), .A2(n9282), .ZN(n9204) );
  OAI211_X1 U10565 ( .C1(n9206), .C2(n9252), .A(n9205), .B(n9204), .ZN(n9207)
         );
  AOI21_X1 U10566 ( .B1(n9529), .B2(n9265), .A(n9207), .ZN(n9208) );
  OAI21_X1 U10567 ( .B1(n9209), .B2(n9267), .A(n9208), .ZN(P1_U3225) );
  AOI21_X1 U10568 ( .B1(n9211), .B2(n7938), .A(n9210), .ZN(n9215) );
  XNOR2_X1 U10569 ( .A(n9213), .B(n9212), .ZN(n9214) );
  XNOR2_X1 U10570 ( .A(n9215), .B(n9214), .ZN(n9222) );
  NOR2_X1 U10571 ( .A1(n9260), .A2(n9216), .ZN(n9220) );
  NAND2_X1 U10572 ( .A1(n9250), .A2(n9287), .ZN(n9217) );
  NAND2_X1 U10573 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9923) );
  OAI211_X1 U10574 ( .C1(n9252), .C2(n9218), .A(n9217), .B(n9923), .ZN(n9219)
         );
  AOI211_X1 U10575 ( .C1(n9720), .C2(n9265), .A(n9220), .B(n9219), .ZN(n9221)
         );
  OAI21_X1 U10576 ( .B1(n9222), .B2(n9267), .A(n9221), .ZN(P1_U3226) );
  INV_X1 U10577 ( .A(n9676), .ZN(n9538) );
  AND3_X1 U10578 ( .A1(n9225), .A2(n9224), .A3(n9223), .ZN(n9226) );
  OAI21_X1 U10579 ( .B1(n9227), .B2(n9226), .A(n9274), .ZN(n9232) );
  NOR2_X1 U10580 ( .A1(n9260), .A2(n9540), .ZN(n9230) );
  OAI22_X1 U10581 ( .A1(n9550), .A2(n9279), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9228), .ZN(n9229) );
  AOI211_X1 U10582 ( .C1(n9277), .C2(n9583), .A(n9230), .B(n9229), .ZN(n9231)
         );
  OAI211_X1 U10583 ( .C1(n9538), .C2(n9285), .A(n9232), .B(n9231), .ZN(
        P1_U3229) );
  XNOR2_X1 U10584 ( .A(n9235), .B(n9234), .ZN(n9236) );
  XNOR2_X1 U10585 ( .A(n9233), .B(n9236), .ZN(n9241) );
  NAND2_X1 U10586 ( .A1(n9282), .A2(n9618), .ZN(n9238) );
  AOI22_X1 U10587 ( .A1(n9611), .A2(n9250), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9237) );
  OAI211_X1 U10588 ( .C1(n9262), .C2(n9252), .A(n9238), .B(n9237), .ZN(n9239)
         );
  AOI21_X1 U10589 ( .B1(n9615), .B2(n9265), .A(n9239), .ZN(n9240) );
  OAI21_X1 U10590 ( .B1(n9241), .B2(n9267), .A(n9240), .ZN(P1_U3233) );
  INV_X1 U10591 ( .A(n9242), .ZN(n9247) );
  OAI21_X1 U10592 ( .B1(n9244), .B2(n9246), .A(n9243), .ZN(n9245) );
  OAI21_X1 U10593 ( .B1(n9247), .B2(n9246), .A(n9245), .ZN(n9248) );
  NAND2_X1 U10594 ( .A1(n9248), .A2(n9274), .ZN(n9256) );
  INV_X1 U10595 ( .A(n9249), .ZN(n9577) );
  AOI22_X1 U10596 ( .A1(n9583), .A2(n9250), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9251) );
  OAI21_X1 U10597 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n9254) );
  AOI21_X1 U10598 ( .B1(n9577), .B2(n9282), .A(n9254), .ZN(n9255) );
  OAI211_X1 U10599 ( .C1(n9579), .C2(n9285), .A(n9256), .B(n9255), .ZN(
        P1_U3235) );
  AOI21_X1 U10600 ( .B1(n9258), .B2(n9257), .A(n4439), .ZN(n9268) );
  NOR2_X1 U10601 ( .A1(n9260), .A2(n9259), .ZN(n9264) );
  NAND2_X1 U10602 ( .A1(n9277), .A2(n9287), .ZN(n9261) );
  NAND2_X1 U10603 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9954) );
  OAI211_X1 U10604 ( .C1(n9279), .C2(n9262), .A(n9261), .B(n9954), .ZN(n9263)
         );
  AOI211_X1 U10605 ( .C1(n9709), .C2(n9265), .A(n9264), .B(n9263), .ZN(n9266)
         );
  OAI21_X1 U10606 ( .B1(n9268), .B2(n9267), .A(n9266), .ZN(P1_U3238) );
  INV_X1 U10607 ( .A(n9269), .ZN(n9275) );
  OAI21_X1 U10608 ( .B1(n9272), .B2(n9271), .A(n9270), .ZN(n9273) );
  NAND3_X1 U10609 ( .A1(n9275), .A2(n9274), .A3(n9273), .ZN(n9284) );
  INV_X1 U10610 ( .A(n9276), .ZN(n9506) );
  AOI22_X1 U10611 ( .A1(n9512), .A2(n9277), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9278) );
  OAI21_X1 U10612 ( .B1(n9280), .B2(n9279), .A(n9278), .ZN(n9281) );
  AOI21_X1 U10613 ( .B1(n9506), .B2(n9282), .A(n9281), .ZN(n9283) );
  OAI211_X1 U10614 ( .C1(n9508), .C2(n9285), .A(n9284), .B(n9283), .ZN(
        P1_U3240) );
  MUX2_X1 U10615 ( .A(n9461), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9301), .Z(
        P1_U3585) );
  MUX2_X1 U10616 ( .A(n9286), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9301), .Z(
        P1_U3584) );
  MUX2_X1 U10617 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n4837), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10618 ( .A(n9524), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9301), .Z(
        P1_U3580) );
  MUX2_X1 U10619 ( .A(n9512), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9301), .Z(
        P1_U3579) );
  MUX2_X1 U10620 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9560), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10621 ( .A(n9593), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9301), .Z(
        P1_U3576) );
  MUX2_X1 U10622 ( .A(n9611), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9301), .Z(
        P1_U3575) );
  MUX2_X1 U10623 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9645), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10624 ( .A(n9610), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9301), .Z(
        P1_U3573) );
  MUX2_X1 U10625 ( .A(n9642), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9301), .Z(
        P1_U3572) );
  MUX2_X1 U10626 ( .A(n9287), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9301), .Z(
        P1_U3571) );
  MUX2_X1 U10627 ( .A(n9288), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9301), .Z(
        P1_U3569) );
  MUX2_X1 U10628 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9289), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10629 ( .A(n9290), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9301), .Z(
        P1_U3566) );
  MUX2_X1 U10630 ( .A(n9291), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9301), .Z(
        P1_U3565) );
  MUX2_X1 U10631 ( .A(n9292), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9301), .Z(
        P1_U3564) );
  MUX2_X1 U10632 ( .A(n9293), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9301), .Z(
        P1_U3563) );
  MUX2_X1 U10633 ( .A(n9294), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9301), .Z(
        P1_U3562) );
  MUX2_X1 U10634 ( .A(n9295), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9301), .Z(
        P1_U3561) );
  MUX2_X1 U10635 ( .A(n9296), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9301), .Z(
        P1_U3560) );
  MUX2_X1 U10636 ( .A(n9297), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9301), .Z(
        P1_U3559) );
  MUX2_X1 U10637 ( .A(n9298), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9301), .Z(
        P1_U3557) );
  MUX2_X1 U10638 ( .A(n9299), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9301), .Z(
        P1_U3556) );
  MUX2_X1 U10639 ( .A(n9300), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9301), .Z(
        P1_U3555) );
  MUX2_X1 U10640 ( .A(n9302), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9301), .Z(
        P1_U3554) );
  INV_X1 U10641 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9304) );
  OAI22_X1 U10642 ( .A1(n9956), .A2(n9304), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9303), .ZN(n9305) );
  AOI21_X1 U10643 ( .B1(n9306), .B2(n9908), .A(n9305), .ZN(n9315) );
  OAI211_X1 U10644 ( .C1(n9309), .C2(n9308), .A(n9946), .B(n9307), .ZN(n9314)
         );
  OAI211_X1 U10645 ( .C1(n9312), .C2(n9311), .A(n9942), .B(n9310), .ZN(n9313)
         );
  NAND3_X1 U10646 ( .A1(n9315), .A2(n9314), .A3(n9313), .ZN(P1_U3244) );
  NOR2_X1 U10647 ( .A1(n9952), .A2(n9316), .ZN(n9320) );
  INV_X1 U10648 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9318) );
  OAI22_X1 U10649 ( .A1(n9956), .A2(n9318), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9317), .ZN(n9319) );
  NOR2_X1 U10650 ( .A1(n9320), .A2(n9319), .ZN(n9329) );
  OAI211_X1 U10651 ( .C1(n9323), .C2(n9322), .A(n9942), .B(n9321), .ZN(n9328)
         );
  OAI211_X1 U10652 ( .C1(n9326), .C2(n9325), .A(n9946), .B(n9324), .ZN(n9327)
         );
  NAND4_X1 U10653 ( .A1(n9330), .A2(n9329), .A3(n9328), .A4(n9327), .ZN(
        P1_U3245) );
  INV_X1 U10654 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9332) );
  OAI21_X1 U10655 ( .B1(n9956), .B2(n9332), .A(n9331), .ZN(n9333) );
  AOI21_X1 U10656 ( .B1(n9334), .B2(n9908), .A(n9333), .ZN(n9343) );
  OAI211_X1 U10657 ( .C1(n9337), .C2(n9336), .A(n9942), .B(n9335), .ZN(n9342)
         );
  OAI211_X1 U10658 ( .C1(n9340), .C2(n9339), .A(n9946), .B(n9338), .ZN(n9341)
         );
  NAND3_X1 U10659 ( .A1(n9343), .A2(n9342), .A3(n9341), .ZN(P1_U3246) );
  INV_X1 U10660 ( .A(n9370), .ZN(n9347) );
  INV_X1 U10661 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9345) );
  OAI21_X1 U10662 ( .B1(n9956), .B2(n9345), .A(n9344), .ZN(n9346) );
  AOI21_X1 U10663 ( .B1(n9347), .B2(n9908), .A(n9346), .ZN(n9359) );
  MUX2_X1 U10664 ( .A(n9363), .B(P1_REG2_REG_5__SCAN_IN), .S(n9370), .Z(n9351)
         );
  NAND2_X1 U10665 ( .A1(n9352), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U10666 ( .A1(n9349), .A2(n9348), .ZN(n9350) );
  NAND2_X1 U10667 ( .A1(n9350), .A2(n9351), .ZN(n9365) );
  OAI211_X1 U10668 ( .C1(n9351), .C2(n9350), .A(n9942), .B(n9365), .ZN(n9358)
         );
  MUX2_X1 U10669 ( .A(n9369), .B(P1_REG1_REG_5__SCAN_IN), .S(n9370), .Z(n9356)
         );
  NAND2_X1 U10670 ( .A1(n9352), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U10671 ( .A1(n9354), .A2(n9353), .ZN(n9355) );
  NAND2_X1 U10672 ( .A1(n9355), .A2(n9356), .ZN(n9372) );
  OAI211_X1 U10673 ( .C1(n9356), .C2(n9355), .A(n9946), .B(n9372), .ZN(n9357)
         );
  NAND3_X1 U10674 ( .A1(n9359), .A2(n9358), .A3(n9357), .ZN(P1_U3248) );
  INV_X1 U10675 ( .A(n9368), .ZN(n9386) );
  INV_X1 U10676 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9361) );
  OAI21_X1 U10677 ( .B1(n9956), .B2(n9361), .A(n9360), .ZN(n9362) );
  AOI21_X1 U10678 ( .B1(n9386), .B2(n9908), .A(n9362), .ZN(n9377) );
  XNOR2_X1 U10679 ( .A(n9368), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9367) );
  OR2_X1 U10680 ( .A1(n9370), .A2(n9363), .ZN(n9364) );
  NAND2_X1 U10681 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  NAND2_X1 U10682 ( .A1(n9366), .A2(n9367), .ZN(n9388) );
  OAI211_X1 U10683 ( .C1(n9367), .C2(n9366), .A(n9942), .B(n9388), .ZN(n9376)
         );
  XNOR2_X1 U10684 ( .A(n9368), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9374) );
  OR2_X1 U10685 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  NAND2_X1 U10686 ( .A1(n9372), .A2(n9371), .ZN(n9373) );
  NAND2_X1 U10687 ( .A1(n9373), .A2(n9374), .ZN(n9383) );
  OAI211_X1 U10688 ( .C1(n9374), .C2(n9373), .A(n9946), .B(n9383), .ZN(n9375)
         );
  NAND3_X1 U10689 ( .A1(n9377), .A2(n9376), .A3(n9375), .ZN(P1_U3249) );
  INV_X1 U10690 ( .A(n9405), .ZN(n9381) );
  INV_X1 U10691 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9379) );
  OAI21_X1 U10692 ( .B1(n9956), .B2(n9379), .A(n9378), .ZN(n9380) );
  AOI21_X1 U10693 ( .B1(n9381), .B2(n9908), .A(n9380), .ZN(n9393) );
  MUX2_X1 U10694 ( .A(n9398), .B(P1_REG1_REG_7__SCAN_IN), .S(n9405), .Z(n9385)
         );
  NAND2_X1 U10695 ( .A1(n9386), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U10696 ( .A1(n9383), .A2(n9382), .ZN(n9384) );
  NAND2_X1 U10697 ( .A1(n9384), .A2(n9385), .ZN(n9400) );
  OAI211_X1 U10698 ( .C1(n9385), .C2(n9384), .A(n9946), .B(n9400), .ZN(n9392)
         );
  MUX2_X1 U10699 ( .A(n9404), .B(P1_REG2_REG_7__SCAN_IN), .S(n9405), .Z(n9390)
         );
  NAND2_X1 U10700 ( .A1(n9386), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U10701 ( .A1(n9388), .A2(n9387), .ZN(n9389) );
  NAND2_X1 U10702 ( .A1(n9389), .A2(n9390), .ZN(n9407) );
  OAI211_X1 U10703 ( .C1(n9390), .C2(n9389), .A(n9942), .B(n9407), .ZN(n9391)
         );
  NAND3_X1 U10704 ( .A1(n9393), .A2(n9392), .A3(n9391), .ZN(P1_U3250) );
  INV_X1 U10705 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9395) );
  OAI21_X1 U10706 ( .B1(n9956), .B2(n9395), .A(n9394), .ZN(n9396) );
  AOI21_X1 U10707 ( .B1(n9430), .B2(n9908), .A(n9396), .ZN(n9412) );
  XNOR2_X1 U10708 ( .A(n9430), .B(n9397), .ZN(n9402) );
  OR2_X1 U10709 ( .A1(n9405), .A2(n9398), .ZN(n9399) );
  NAND2_X1 U10710 ( .A1(n9400), .A2(n9399), .ZN(n9401) );
  NAND2_X1 U10711 ( .A1(n9401), .A2(n9402), .ZN(n9416) );
  OAI211_X1 U10712 ( .C1(n9402), .C2(n9401), .A(n9946), .B(n9416), .ZN(n9411)
         );
  XNOR2_X1 U10713 ( .A(n9430), .B(n9403), .ZN(n9409) );
  OR2_X1 U10714 ( .A1(n9405), .A2(n9404), .ZN(n9406) );
  NAND2_X1 U10715 ( .A1(n9407), .A2(n9406), .ZN(n9408) );
  NAND2_X1 U10716 ( .A1(n9408), .A2(n9409), .ZN(n9432) );
  OAI211_X1 U10717 ( .C1(n9409), .C2(n9408), .A(n9942), .B(n9432), .ZN(n9410)
         );
  NAND3_X1 U10718 ( .A1(n9412), .A2(n9411), .A3(n9410), .ZN(P1_U3251) );
  XNOR2_X1 U10719 ( .A(n9926), .B(n9715), .ZN(n9931) );
  OR2_X1 U10720 ( .A1(n9443), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9422) );
  XNOR2_X1 U10721 ( .A(n9443), .B(n9413), .ZN(n9913) );
  XNOR2_X1 U10722 ( .A(n9437), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U10723 ( .A1(n9814), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9414) );
  OAI21_X1 U10724 ( .B1(n9814), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9414), .ZN(
        n9807) );
  NAND2_X1 U10725 ( .A1(n9430), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U10726 ( .A1(n9416), .A2(n9415), .ZN(n9824) );
  NAND2_X1 U10727 ( .A1(n9435), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9418) );
  OR2_X1 U10728 ( .A1(n9435), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U10729 ( .A1(n9418), .A2(n9417), .ZN(n9823) );
  OAI21_X1 U10730 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9435), .A(n9826), .ZN(
        n9808) );
  NOR2_X1 U10731 ( .A1(n9807), .A2(n9808), .ZN(n9806) );
  AOI21_X1 U10732 ( .B1(n9814), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9806), .ZN(
        n9843) );
  XNOR2_X1 U10733 ( .A(n9836), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n9842) );
  NOR2_X1 U10734 ( .A1(n9843), .A2(n9842), .ZN(n9841) );
  AOI21_X1 U10735 ( .B1(n9836), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9841), .ZN(
        n9858) );
  XNOR2_X1 U10736 ( .A(n9852), .B(n9419), .ZN(n9859) );
  NAND2_X1 U10737 ( .A1(n9858), .A2(n9859), .ZN(n9857) );
  OAI21_X1 U10738 ( .B1(n9852), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9857), .ZN(
        n9873) );
  NOR2_X1 U10739 ( .A1(n9874), .A2(n9873), .ZN(n9872) );
  AOI21_X1 U10740 ( .B1(n9437), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9872), .ZN(
        n9886) );
  XNOR2_X1 U10741 ( .A(n9883), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9885) );
  NOR2_X1 U10742 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  AOI21_X1 U10743 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9883), .A(n9884), .ZN(
        n9420) );
  NOR2_X1 U10744 ( .A1(n9420), .A2(n9440), .ZN(n9421) );
  XNOR2_X1 U10745 ( .A(n9440), .B(n9420), .ZN(n9902) );
  NOR2_X1 U10746 ( .A1(n9901), .A2(n9902), .ZN(n9900) );
  NOR2_X1 U10747 ( .A1(n9421), .A2(n9900), .ZN(n9914) );
  NAND2_X1 U10748 ( .A1(n9913), .A2(n9914), .ZN(n9912) );
  NAND2_X1 U10749 ( .A1(n9422), .A2(n9912), .ZN(n9930) );
  NOR2_X1 U10750 ( .A1(n9926), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9423) );
  AOI21_X1 U10751 ( .B1(n9931), .B2(n9930), .A(n9423), .ZN(n9948) );
  OR2_X1 U10752 ( .A1(n9940), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U10753 ( .A1(n9940), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9425) );
  AND2_X1 U10754 ( .A1(n9424), .A2(n9425), .ZN(n9947) );
  NAND2_X1 U10755 ( .A1(n9948), .A2(n9947), .ZN(n9945) );
  NAND2_X1 U10756 ( .A1(n9945), .A2(n9425), .ZN(n9426) );
  XNOR2_X1 U10757 ( .A(n9426), .B(n9705), .ZN(n9449) );
  XNOR2_X1 U10758 ( .A(n9926), .B(n9427), .ZN(n9928) );
  AOI22_X1 U10759 ( .A1(n9437), .A2(n7387), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n9878), .ZN(n9870) );
  NOR2_X1 U10760 ( .A1(n9852), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9428) );
  AOI21_X1 U10761 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9852), .A(n9428), .ZN(
        n9855) );
  NAND2_X1 U10762 ( .A1(n9814), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9429) );
  OAI21_X1 U10763 ( .B1(n9814), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9429), .ZN(
        n9810) );
  NAND2_X1 U10764 ( .A1(n9430), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U10765 ( .A1(n9432), .A2(n9431), .ZN(n9819) );
  NAND2_X1 U10766 ( .A1(n9435), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9434) );
  OR2_X1 U10767 ( .A1(n9435), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U10768 ( .A1(n9434), .A2(n9433), .ZN(n9818) );
  OAI21_X1 U10769 ( .B1(n9435), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9821), .ZN(
        n9811) );
  NOR2_X1 U10770 ( .A1(n9810), .A2(n9811), .ZN(n9809) );
  AOI21_X1 U10771 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9814), .A(n9809), .ZN(
        n9838) );
  NAND2_X1 U10772 ( .A1(n9836), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9436) );
  OAI21_X1 U10773 ( .B1(n9836), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9436), .ZN(
        n9839) );
  NOR2_X1 U10774 ( .A1(n9838), .A2(n9839), .ZN(n9837) );
  AOI21_X1 U10775 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9836), .A(n9837), .ZN(
        n9854) );
  NAND2_X1 U10776 ( .A1(n9855), .A2(n9854), .ZN(n9853) );
  OAI21_X1 U10777 ( .B1(n9852), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9853), .ZN(
        n9869) );
  NOR2_X1 U10778 ( .A1(n9870), .A2(n9869), .ZN(n9868) );
  AOI21_X1 U10779 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9437), .A(n9868), .ZN(
        n9889) );
  NAND2_X1 U10780 ( .A1(n9883), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9438) );
  OAI21_X1 U10781 ( .B1(n9883), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9438), .ZN(
        n9890) );
  NOR2_X1 U10782 ( .A1(n9889), .A2(n9890), .ZN(n9888) );
  AOI21_X1 U10783 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9883), .A(n9888), .ZN(
        n9439) );
  NOR2_X1 U10784 ( .A1(n9439), .A2(n9440), .ZN(n9441) );
  XNOR2_X1 U10785 ( .A(n9440), .B(n9439), .ZN(n9904) );
  NOR2_X1 U10786 ( .A1(n7646), .A2(n9904), .ZN(n9903) );
  NOR2_X1 U10787 ( .A1(n9441), .A2(n9903), .ZN(n9919) );
  NAND2_X1 U10788 ( .A1(n9443), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9442) );
  OAI21_X1 U10789 ( .B1(n9443), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9442), .ZN(
        n9918) );
  NOR2_X1 U10790 ( .A1(n9919), .A2(n9918), .ZN(n9917) );
  AOI21_X1 U10791 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9443), .A(n9917), .ZN(
        n9927) );
  NOR2_X1 U10792 ( .A1(n9926), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9444) );
  AOI21_X1 U10793 ( .B1(n9928), .B2(n9927), .A(n9444), .ZN(n9943) );
  OR2_X1 U10794 ( .A1(n9940), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U10795 ( .A1(n9940), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9446) );
  AND2_X1 U10796 ( .A1(n9445), .A2(n9446), .ZN(n9944) );
  NAND2_X1 U10797 ( .A1(n9943), .A2(n9944), .ZN(n9941) );
  NAND2_X1 U10798 ( .A1(n9941), .A2(n9446), .ZN(n9447) );
  XNOR2_X1 U10799 ( .A(n9447), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9451) );
  AOI21_X1 U10800 ( .B1(n9942), .B2(n9451), .A(n9908), .ZN(n9448) );
  OAI21_X1 U10801 ( .B1(n9899), .B2(n9449), .A(n9448), .ZN(n9453) );
  INV_X1 U10802 ( .A(n9449), .ZN(n9450) );
  OAI22_X1 U10803 ( .A1(n9451), .A2(n9916), .B1(n9899), .B2(n9450), .ZN(n9452)
         );
  MUX2_X1 U10804 ( .A(n9453), .B(n9452), .S(n8317), .Z(n9454) );
  AOI211_X1 U10805 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n9456), .A(n9455), .B(
        n9454), .ZN(n9457) );
  INV_X1 U10806 ( .A(n9457), .ZN(P1_U3262) );
  NAND2_X1 U10807 ( .A1(n9652), .A2(n9616), .ZN(n9464) );
  AND2_X1 U10808 ( .A1(n9461), .A2(n9460), .ZN(n9655) );
  INV_X1 U10809 ( .A(n9655), .ZN(n9462) );
  NOR2_X1 U10810 ( .A1(n9462), .A2(n9469), .ZN(n9468) );
  AOI21_X1 U10811 ( .B1(n9469), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9468), .ZN(
        n9463) );
  OAI211_X1 U10812 ( .C1(n9734), .C2(n9629), .A(n9464), .B(n9463), .ZN(
        P1_U3263) );
  INV_X1 U10813 ( .A(n9465), .ZN(n9466) );
  AOI211_X1 U10814 ( .C1(n9467), .C2(n9466), .A(n9682), .B(n4392), .ZN(n9656)
         );
  NAND2_X1 U10815 ( .A1(n9656), .A2(n9616), .ZN(n9471) );
  AOI21_X1 U10816 ( .B1(n9469), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9468), .ZN(
        n9470) );
  OAI211_X1 U10817 ( .C1(n9738), .C2(n9629), .A(n9471), .B(n9470), .ZN(
        P1_U3264) );
  INV_X1 U10818 ( .A(n9472), .ZN(n9483) );
  NAND2_X1 U10819 ( .A1(n9473), .A2(n9616), .ZN(n9478) );
  NOR3_X1 U10820 ( .A1(n9475), .A2(n9474), .A3(n9630), .ZN(n9476) );
  AOI21_X1 U10821 ( .B1(n9469), .B2(P1_REG2_REG_29__SCAN_IN), .A(n9476), .ZN(
        n9477) );
  OAI211_X1 U10822 ( .C1(n9479), .C2(n9629), .A(n9478), .B(n9477), .ZN(n9480)
         );
  AOI21_X1 U10823 ( .B1(n9481), .B2(n9633), .A(n9480), .ZN(n9482) );
  OAI21_X1 U10824 ( .B1(n9483), .B2(n9650), .A(n9482), .ZN(P1_U3356) );
  XNOR2_X1 U10825 ( .A(n9484), .B(n9493), .ZN(n9661) );
  INV_X1 U10826 ( .A(n9661), .ZN(n9502) );
  AOI211_X1 U10827 ( .C1(n9486), .C2(n9504), .A(n9682), .B(n5885), .ZN(n9660)
         );
  NOR2_X1 U10828 ( .A1(n9742), .A2(n9629), .ZN(n9490) );
  OAI22_X1 U10829 ( .A1(n9488), .A2(n9630), .B1(n9487), .B2(n7692), .ZN(n9489)
         );
  AOI211_X1 U10830 ( .C1(n9660), .C2(n9616), .A(n9490), .B(n9489), .ZN(n9501)
         );
  OAI21_X1 U10831 ( .B1(n9493), .B2(n9492), .A(n9491), .ZN(n9494) );
  NAND2_X1 U10832 ( .A1(n9494), .A2(n9640), .ZN(n9499) );
  OAI22_X1 U10833 ( .A1(n9496), .A2(n9551), .B1(n9495), .B2(n9549), .ZN(n9497)
         );
  INV_X1 U10834 ( .A(n9497), .ZN(n9498) );
  NAND2_X1 U10835 ( .A1(n9499), .A2(n9498), .ZN(n9659) );
  NAND2_X1 U10836 ( .A1(n9659), .A2(n9633), .ZN(n9500) );
  OAI211_X1 U10837 ( .C1(n9502), .C2(n9650), .A(n9501), .B(n9500), .ZN(
        P1_U3266) );
  XNOR2_X1 U10838 ( .A(n9503), .B(n9511), .ZN(n9668) );
  INV_X1 U10839 ( .A(n9527), .ZN(n9505) );
  AOI211_X1 U10840 ( .C1(n9665), .C2(n9505), .A(n9682), .B(n4754), .ZN(n9664)
         );
  AOI22_X1 U10841 ( .A1(n9506), .A2(n9617), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9469), .ZN(n9507) );
  OAI21_X1 U10842 ( .B1(n9508), .B2(n9629), .A(n9507), .ZN(n9516) );
  OAI21_X1 U10843 ( .B1(n9511), .B2(n9510), .A(n9509), .ZN(n9514) );
  AOI222_X1 U10844 ( .A1(n9640), .A2(n9514), .B1(n9513), .B2(n9644), .C1(n9512), .C2(n9643), .ZN(n9667) );
  NOR2_X1 U10845 ( .A1(n9667), .A2(n9469), .ZN(n9515) );
  AOI211_X1 U10846 ( .C1(n9664), .C2(n9616), .A(n9516), .B(n9515), .ZN(n9517)
         );
  OAI21_X1 U10847 ( .B1(n9668), .B2(n9650), .A(n9517), .ZN(P1_U3267) );
  XOR2_X1 U10848 ( .A(n9519), .B(n9518), .Z(n9671) );
  INV_X1 U10849 ( .A(n9671), .ZN(n9535) );
  NAND2_X1 U10850 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  NAND2_X1 U10851 ( .A1(n9522), .A2(n9521), .ZN(n9523) );
  NAND2_X1 U10852 ( .A1(n9523), .A2(n9640), .ZN(n9526) );
  AOI22_X1 U10853 ( .A1(n9524), .A2(n9644), .B1(n9643), .B2(n9560), .ZN(n9525)
         );
  NAND2_X1 U10854 ( .A1(n9526), .A2(n9525), .ZN(n9669) );
  INV_X1 U10855 ( .A(n9537), .ZN(n9528) );
  AOI211_X1 U10856 ( .C1(n9529), .C2(n9528), .A(n9682), .B(n9527), .ZN(n9670)
         );
  NAND2_X1 U10857 ( .A1(n9670), .A2(n9616), .ZN(n9532) );
  AOI22_X1 U10858 ( .A1(n9530), .A2(n9617), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9469), .ZN(n9531) );
  OAI211_X1 U10859 ( .C1(n9747), .C2(n9629), .A(n9532), .B(n9531), .ZN(n9533)
         );
  AOI21_X1 U10860 ( .B1(n9633), .B2(n9669), .A(n9533), .ZN(n9534) );
  OAI21_X1 U10861 ( .B1(n9535), .B2(n9650), .A(n9534), .ZN(P1_U3268) );
  XOR2_X1 U10862 ( .A(n9536), .B(n9545), .Z(n9678) );
  AOI211_X1 U10863 ( .C1(n9676), .C2(n4944), .A(n9682), .B(n9537), .ZN(n9675)
         );
  NOR2_X1 U10864 ( .A1(n9538), .A2(n9629), .ZN(n9542) );
  OAI22_X1 U10865 ( .A1(n9540), .A2(n9630), .B1(n9539), .B2(n9633), .ZN(n9541)
         );
  AOI211_X1 U10866 ( .C1(n9675), .C2(n9616), .A(n9542), .B(n9541), .ZN(n9553)
         );
  NAND2_X1 U10867 ( .A1(n9556), .A2(n9543), .ZN(n9544) );
  XOR2_X1 U10868 ( .A(n9545), .B(n9544), .Z(n9547) );
  OAI222_X1 U10869 ( .A1(n9551), .A2(n9550), .B1(n9549), .B2(n9548), .C1(n9547), .C2(n9546), .ZN(n9674) );
  NAND2_X1 U10870 ( .A1(n9674), .A2(n7692), .ZN(n9552) );
  OAI211_X1 U10871 ( .C1(n9678), .C2(n9650), .A(n9553), .B(n9552), .ZN(
        P1_U3269) );
  XOR2_X1 U10872 ( .A(n9558), .B(n9554), .Z(n9684) );
  INV_X1 U10873 ( .A(n9684), .ZN(n9569) );
  INV_X1 U10874 ( .A(n9555), .ZN(n9561) );
  OAI21_X1 U10875 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9559) );
  NAND2_X1 U10876 ( .A1(n9559), .A2(n9640), .ZN(n9680) );
  AOI22_X1 U10877 ( .A1(n9560), .A2(n9644), .B1(n9643), .B2(n9593), .ZN(n9679)
         );
  OAI211_X1 U10878 ( .C1(n9630), .C2(n9561), .A(n9680), .B(n9679), .ZN(n9567)
         );
  XNOR2_X1 U10879 ( .A(n9562), .B(n9574), .ZN(n9681) );
  NOR2_X1 U10880 ( .A1(n9681), .A2(n9563), .ZN(n9566) );
  OAI22_X1 U10881 ( .A1(n9752), .A2(n9629), .B1(n9564), .B2(n9633), .ZN(n9565)
         );
  AOI211_X1 U10882 ( .C1(n9567), .C2(n9633), .A(n9566), .B(n9565), .ZN(n9568)
         );
  OAI21_X1 U10883 ( .B1(n9569), .B2(n9650), .A(n9568), .ZN(P1_U3270) );
  OR2_X1 U10884 ( .A1(n9588), .A2(n9570), .ZN(n9572) );
  NAND2_X1 U10885 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  XNOR2_X1 U10886 ( .A(n9573), .B(n9582), .ZN(n9691) );
  INV_X1 U10887 ( .A(n9596), .ZN(n9576) );
  INV_X1 U10888 ( .A(n9574), .ZN(n9575) );
  AOI211_X1 U10889 ( .C1(n9688), .C2(n9576), .A(n9682), .B(n9575), .ZN(n9687)
         );
  AOI22_X1 U10890 ( .A1(n9577), .A2(n9617), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9469), .ZN(n9578) );
  OAI21_X1 U10891 ( .B1(n9579), .B2(n9629), .A(n9578), .ZN(n9586) );
  OAI21_X1 U10892 ( .B1(n9582), .B2(n9581), .A(n9580), .ZN(n9584) );
  AOI222_X1 U10893 ( .A1(n9640), .A2(n9584), .B1(n9611), .B2(n9643), .C1(n9583), .C2(n9644), .ZN(n9690) );
  NOR2_X1 U10894 ( .A1(n9690), .A2(n9469), .ZN(n9585) );
  AOI211_X1 U10895 ( .C1(n9687), .C2(n9616), .A(n9586), .B(n9585), .ZN(n9587)
         );
  OAI21_X1 U10896 ( .B1(n9691), .B2(n9650), .A(n9587), .ZN(P1_U3271) );
  XNOR2_X1 U10897 ( .A(n9588), .B(n9591), .ZN(n9694) );
  INV_X1 U10898 ( .A(n9694), .ZN(n9604) );
  OAI21_X1 U10899 ( .B1(n9591), .B2(n9590), .A(n9589), .ZN(n9592) );
  NAND2_X1 U10900 ( .A1(n9592), .A2(n9640), .ZN(n9595) );
  AOI22_X1 U10901 ( .A1(n9593), .A2(n9644), .B1(n9643), .B2(n9645), .ZN(n9594)
         );
  NAND2_X1 U10902 ( .A1(n9595), .A2(n9594), .ZN(n9692) );
  AOI211_X1 U10903 ( .C1(n9597), .C2(n9614), .A(n9682), .B(n9596), .ZN(n9693)
         );
  NAND2_X1 U10904 ( .A1(n9693), .A2(n9616), .ZN(n9601) );
  INV_X1 U10905 ( .A(n9598), .ZN(n9599) );
  AOI22_X1 U10906 ( .A1(n9599), .A2(n9617), .B1(n9469), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9600) );
  OAI211_X1 U10907 ( .C1(n9757), .C2(n9629), .A(n9601), .B(n9600), .ZN(n9602)
         );
  AOI21_X1 U10908 ( .B1(n9633), .B2(n9692), .A(n9602), .ZN(n9603) );
  OAI21_X1 U10909 ( .B1(n9604), .B2(n9650), .A(n9603), .ZN(P1_U3272) );
  XOR2_X1 U10910 ( .A(n9607), .B(n9605), .Z(n9699) );
  INV_X1 U10911 ( .A(n9699), .ZN(n9623) );
  OAI21_X1 U10912 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9609) );
  NAND2_X1 U10913 ( .A1(n9609), .A2(n9640), .ZN(n9613) );
  AOI22_X1 U10914 ( .A1(n9611), .A2(n9644), .B1(n9643), .B2(n9610), .ZN(n9612)
         );
  NAND2_X1 U10915 ( .A1(n9613), .A2(n9612), .ZN(n9697) );
  INV_X1 U10916 ( .A(n9615), .ZN(n9761) );
  AOI211_X1 U10917 ( .C1(n9615), .C2(n9626), .A(n9682), .B(n4758), .ZN(n9698)
         );
  NAND2_X1 U10918 ( .A1(n9698), .A2(n9616), .ZN(n9620) );
  AOI22_X1 U10919 ( .A1(n9469), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9618), .B2(
        n9617), .ZN(n9619) );
  OAI211_X1 U10920 ( .C1(n9761), .C2(n9629), .A(n9620), .B(n9619), .ZN(n9621)
         );
  AOI21_X1 U10921 ( .B1(n9633), .B2(n9697), .A(n9621), .ZN(n9622) );
  OAI21_X1 U10922 ( .B1(n9623), .B2(n9650), .A(n9622), .ZN(P1_U3273) );
  XOR2_X1 U10923 ( .A(n9638), .B(n9624), .Z(n9704) );
  INV_X1 U10924 ( .A(n9704), .ZN(n9651) );
  INV_X1 U10925 ( .A(n9625), .ZN(n9627) );
  AOI211_X1 U10926 ( .C1(n9628), .C2(n9627), .A(n9682), .B(n4759), .ZN(n9703)
         );
  NOR2_X1 U10927 ( .A1(n9765), .A2(n9629), .ZN(n9635) );
  OAI22_X1 U10928 ( .A1(n9633), .A2(n9632), .B1(n9631), .B2(n9630), .ZN(n9634)
         );
  AOI211_X1 U10929 ( .C1(n9703), .C2(n9616), .A(n9635), .B(n9634), .ZN(n9649)
         );
  NAND2_X1 U10930 ( .A1(n9637), .A2(n9636), .ZN(n9639) );
  XNOR2_X1 U10931 ( .A(n9639), .B(n9638), .ZN(n9641) );
  NAND2_X1 U10932 ( .A1(n9641), .A2(n9640), .ZN(n9647) );
  AOI22_X1 U10933 ( .A1(n9645), .A2(n9644), .B1(n9643), .B2(n9642), .ZN(n9646)
         );
  NAND2_X1 U10934 ( .A1(n9647), .A2(n9646), .ZN(n9702) );
  NAND2_X1 U10935 ( .A1(n9702), .A2(n7692), .ZN(n9648) );
  OAI211_X1 U10936 ( .C1(n9651), .C2(n9650), .A(n9649), .B(n9648), .ZN(
        P1_U3274) );
  NOR2_X1 U10937 ( .A1(n9652), .A2(n9655), .ZN(n9731) );
  MUX2_X1 U10938 ( .A(n9653), .B(n9731), .S(n9988), .Z(n9654) );
  OAI21_X1 U10939 ( .B1(n9734), .B2(n9717), .A(n9654), .ZN(P1_U3553) );
  NOR2_X1 U10940 ( .A1(n9656), .A2(n9655), .ZN(n9735) );
  MUX2_X1 U10941 ( .A(n9657), .B(n9735), .S(n9988), .Z(n9658) );
  OAI21_X1 U10942 ( .B1(n9738), .B2(n9717), .A(n9658), .ZN(P1_U3552) );
  AOI211_X1 U10943 ( .C1(n9661), .C2(n9978), .A(n9660), .B(n9659), .ZN(n9739)
         );
  MUX2_X1 U10944 ( .A(n9662), .B(n9739), .S(n9988), .Z(n9663) );
  OAI21_X1 U10945 ( .B1(n9742), .B2(n9717), .A(n9663), .ZN(P1_U3549) );
  AOI21_X1 U10946 ( .B1(n9726), .B2(n9665), .A(n9664), .ZN(n9666) );
  OAI211_X1 U10947 ( .C1(n9668), .C2(n9728), .A(n9667), .B(n9666), .ZN(n9743)
         );
  MUX2_X1 U10948 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9743), .S(n9988), .Z(
        P1_U3548) );
  AOI211_X1 U10949 ( .C1(n9671), .C2(n9978), .A(n9670), .B(n9669), .ZN(n9744)
         );
  MUX2_X1 U10950 ( .A(n9672), .B(n9744), .S(n9988), .Z(n9673) );
  OAI21_X1 U10951 ( .B1(n9747), .B2(n9717), .A(n9673), .ZN(P1_U3547) );
  AOI211_X1 U10952 ( .C1(n9726), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9677)
         );
  OAI21_X1 U10953 ( .B1(n9678), .B2(n9728), .A(n9677), .ZN(n9748) );
  MUX2_X1 U10954 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9748), .S(n9988), .Z(
        P1_U3546) );
  OAI211_X1 U10955 ( .C1(n9682), .C2(n9681), .A(n9680), .B(n9679), .ZN(n9683)
         );
  AOI21_X1 U10956 ( .B1(n9684), .B2(n9978), .A(n9683), .ZN(n9749) );
  MUX2_X1 U10957 ( .A(n9685), .B(n9749), .S(n9988), .Z(n9686) );
  OAI21_X1 U10958 ( .B1(n9752), .B2(n9717), .A(n9686), .ZN(P1_U3545) );
  AOI21_X1 U10959 ( .B1(n9726), .B2(n9688), .A(n9687), .ZN(n9689) );
  OAI211_X1 U10960 ( .C1(n9691), .C2(n9728), .A(n9690), .B(n9689), .ZN(n9753)
         );
  MUX2_X1 U10961 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9753), .S(n9988), .Z(
        P1_U3544) );
  INV_X1 U10962 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9695) );
  AOI211_X1 U10963 ( .C1(n9694), .C2(n9978), .A(n9693), .B(n9692), .ZN(n9754)
         );
  MUX2_X1 U10964 ( .A(n9695), .B(n9754), .S(n9988), .Z(n9696) );
  OAI21_X1 U10965 ( .B1(n9757), .B2(n9717), .A(n9696), .ZN(P1_U3543) );
  AOI211_X1 U10966 ( .C1(n9699), .C2(n9978), .A(n9698), .B(n9697), .ZN(n9758)
         );
  MUX2_X1 U10967 ( .A(n9700), .B(n9758), .S(n9988), .Z(n9701) );
  OAI21_X1 U10968 ( .B1(n9761), .B2(n9717), .A(n9701), .ZN(P1_U3542) );
  AOI211_X1 U10969 ( .C1(n9704), .C2(n9978), .A(n9703), .B(n9702), .ZN(n9762)
         );
  MUX2_X1 U10970 ( .A(n9705), .B(n9762), .S(n9988), .Z(n9706) );
  OAI21_X1 U10971 ( .B1(n9765), .B2(n9717), .A(n9706), .ZN(P1_U3541) );
  AOI211_X1 U10972 ( .C1(n9726), .C2(n9709), .A(n9708), .B(n9707), .ZN(n9710)
         );
  OAI21_X1 U10973 ( .B1(n9711), .B2(n9728), .A(n9710), .ZN(n9766) );
  MUX2_X1 U10974 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9766), .S(n9988), .Z(
        P1_U3540) );
  AOI211_X1 U10975 ( .C1(n9714), .C2(n9978), .A(n9713), .B(n9712), .ZN(n9767)
         );
  MUX2_X1 U10976 ( .A(n9715), .B(n9767), .S(n9988), .Z(n9716) );
  OAI21_X1 U10977 ( .B1(n9771), .B2(n9717), .A(n9716), .ZN(P1_U3539) );
  AOI211_X1 U10978 ( .C1(n9726), .C2(n9720), .A(n9719), .B(n9718), .ZN(n9721)
         );
  OAI21_X1 U10979 ( .B1(n9722), .B2(n9728), .A(n9721), .ZN(n9772) );
  MUX2_X1 U10980 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9772), .S(n9988), .Z(
        P1_U3538) );
  AOI211_X1 U10981 ( .C1(n9726), .C2(n9725), .A(n9724), .B(n9723), .ZN(n9727)
         );
  OAI21_X1 U10982 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9773) );
  MUX2_X1 U10983 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9773), .S(n9988), .Z(
        P1_U3536) );
  MUX2_X1 U10984 ( .A(n9730), .B(P1_REG1_REG_0__SCAN_IN), .S(n9986), .Z(
        P1_U3522) );
  MUX2_X1 U10985 ( .A(n9732), .B(n9731), .S(n9981), .Z(n9733) );
  OAI21_X1 U10986 ( .B1(n9734), .B2(n9770), .A(n9733), .ZN(P1_U3521) );
  MUX2_X1 U10987 ( .A(n9736), .B(n9735), .S(n9981), .Z(n9737) );
  OAI21_X1 U10988 ( .B1(n9738), .B2(n9770), .A(n9737), .ZN(P1_U3520) );
  MUX2_X1 U10989 ( .A(n9740), .B(n9739), .S(n9981), .Z(n9741) );
  OAI21_X1 U10990 ( .B1(n9742), .B2(n9770), .A(n9741), .ZN(P1_U3517) );
  MUX2_X1 U10991 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9743), .S(n9981), .Z(
        P1_U3516) );
  MUX2_X1 U10992 ( .A(n9745), .B(n9744), .S(n9981), .Z(n9746) );
  OAI21_X1 U10993 ( .B1(n9747), .B2(n9770), .A(n9746), .ZN(P1_U3515) );
  MUX2_X1 U10994 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9748), .S(n9981), .Z(
        P1_U3514) );
  MUX2_X1 U10995 ( .A(n9750), .B(n9749), .S(n9981), .Z(n9751) );
  OAI21_X1 U10996 ( .B1(n9752), .B2(n9770), .A(n9751), .ZN(P1_U3513) );
  MUX2_X1 U10997 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9753), .S(n9981), .Z(
        P1_U3512) );
  MUX2_X1 U10998 ( .A(n9755), .B(n9754), .S(n9981), .Z(n9756) );
  OAI21_X1 U10999 ( .B1(n9757), .B2(n9770), .A(n9756), .ZN(P1_U3511) );
  MUX2_X1 U11000 ( .A(n9759), .B(n9758), .S(n9981), .Z(n9760) );
  OAI21_X1 U11001 ( .B1(n9761), .B2(n9770), .A(n9760), .ZN(P1_U3510) );
  MUX2_X1 U11002 ( .A(n9763), .B(n9762), .S(n9981), .Z(n9764) );
  OAI21_X1 U11003 ( .B1(n9765), .B2(n9770), .A(n9764), .ZN(P1_U3509) );
  MUX2_X1 U11004 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9766), .S(n9981), .Z(
        P1_U3507) );
  MUX2_X1 U11005 ( .A(n9768), .B(n9767), .S(n9981), .Z(n9769) );
  OAI21_X1 U11006 ( .B1(n9771), .B2(n9770), .A(n9769), .ZN(P1_U3504) );
  MUX2_X1 U11007 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9772), .S(n9981), .Z(
        P1_U3501) );
  MUX2_X1 U11008 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9773), .S(n9981), .Z(
        P1_U3495) );
  MUX2_X1 U11009 ( .A(n9774), .B(P1_D_REG_1__SCAN_IN), .S(n9957), .Z(P1_U3440)
         );
  NAND2_X1 U11010 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .ZN(n9777) );
  OAI22_X1 U11011 ( .A1(n9778), .A2(n9777), .B1(n9776), .B2(n9775), .ZN(n9779)
         );
  AOI21_X1 U11012 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9782) );
  INV_X1 U11013 ( .A(n9782), .ZN(P1_U3324) );
  MUX2_X1 U11014 ( .A(n9783), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11015 ( .A(n9784), .ZN(n9785) );
  NAND2_X1 U11016 ( .A1(n10115), .A2(n9787), .ZN(n9804) );
  INV_X1 U11017 ( .A(n9787), .ZN(n9788) );
  AOI21_X1 U11018 ( .B1(P2_U3893), .B2(n9788), .A(n10107), .ZN(n9802) );
  OAI21_X1 U11019 ( .B1(n9791), .B2(n9790), .A(n9789), .ZN(n9800) );
  INV_X1 U11020 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9793) );
  OAI21_X1 U11021 ( .B1(n10020), .B2(n9793), .A(n9792), .ZN(n9799) );
  AOI211_X1 U11022 ( .C1(n10116), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9801)
         );
  OAI221_X1 U11023 ( .B1(n9805), .B2(n9804), .C1(n9803), .C2(n9802), .A(n9801), 
        .ZN(P2_U3200) );
  INV_X1 U11024 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9817) );
  AOI211_X1 U11025 ( .C1(n9808), .C2(n9807), .A(n9806), .B(n9899), .ZN(n9813)
         );
  AOI211_X1 U11026 ( .C1(n9811), .C2(n9810), .A(n9809), .B(n9916), .ZN(n9812)
         );
  AOI211_X1 U11027 ( .C1(n9908), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9816)
         );
  OAI211_X1 U11028 ( .C1(n9956), .C2(n9817), .A(n9816), .B(n9815), .ZN(
        P1_U3253) );
  INV_X1 U11029 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U11030 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  NAND2_X1 U11031 ( .A1(n9821), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U11032 ( .A1(n9942), .A2(n9822), .ZN(n9829) );
  NAND2_X1 U11033 ( .A1(n9824), .A2(n9823), .ZN(n9825) );
  NAND2_X1 U11034 ( .A1(n9826), .A2(n9825), .ZN(n9827) );
  NAND2_X1 U11035 ( .A1(n9946), .A2(n9827), .ZN(n9828) );
  OAI211_X1 U11036 ( .C1(n9952), .C2(n9830), .A(n9829), .B(n9828), .ZN(n9831)
         );
  INV_X1 U11037 ( .A(n9831), .ZN(n9833) );
  OAI211_X1 U11038 ( .C1(n9956), .C2(n9834), .A(n9833), .B(n9832), .ZN(
        P1_U3252) );
  XOR2_X1 U11039 ( .A(n9835), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XOR2_X1 U11040 ( .A(n5006), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  INV_X1 U11041 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9851) );
  INV_X1 U11042 ( .A(n9836), .ZN(n9847) );
  AOI21_X1 U11043 ( .B1(n9839), .B2(n9838), .A(n9837), .ZN(n9840) );
  NAND2_X1 U11044 ( .A1(n9942), .A2(n9840), .ZN(n9846) );
  AOI21_X1 U11045 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9844) );
  NAND2_X1 U11046 ( .A1(n9946), .A2(n9844), .ZN(n9845) );
  OAI211_X1 U11047 ( .C1(n9952), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9848)
         );
  INV_X1 U11048 ( .A(n9848), .ZN(n9850) );
  OAI211_X1 U11049 ( .C1(n9956), .C2(n9851), .A(n9850), .B(n9849), .ZN(
        P1_U3254) );
  INV_X1 U11050 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9867) );
  INV_X1 U11051 ( .A(n9852), .ZN(n9863) );
  OAI21_X1 U11052 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(n9856) );
  NAND2_X1 U11053 ( .A1(n9942), .A2(n9856), .ZN(n9862) );
  OAI21_X1 U11054 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9860) );
  NAND2_X1 U11055 ( .A1(n9946), .A2(n9860), .ZN(n9861) );
  OAI211_X1 U11056 ( .C1(n9952), .C2(n9863), .A(n9862), .B(n9861), .ZN(n9864)
         );
  INV_X1 U11057 ( .A(n9864), .ZN(n9866) );
  OAI211_X1 U11058 ( .C1(n9956), .C2(n9867), .A(n9866), .B(n9865), .ZN(
        P1_U3255) );
  INV_X1 U11059 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9882) );
  AOI21_X1 U11060 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9871) );
  NAND2_X1 U11061 ( .A1(n9942), .A2(n9871), .ZN(n9877) );
  AOI21_X1 U11062 ( .B1(n9874), .B2(n9873), .A(n9872), .ZN(n9875) );
  NAND2_X1 U11063 ( .A1(n9946), .A2(n9875), .ZN(n9876) );
  OAI211_X1 U11064 ( .C1(n9952), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9879)
         );
  INV_X1 U11065 ( .A(n9879), .ZN(n9881) );
  OAI211_X1 U11066 ( .C1(n9956), .C2(n9882), .A(n9881), .B(n9880), .ZN(
        P1_U3256) );
  INV_X1 U11067 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9898) );
  INV_X1 U11068 ( .A(n9883), .ZN(n9894) );
  AOI21_X1 U11069 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9887) );
  NAND2_X1 U11070 ( .A1(n9946), .A2(n9887), .ZN(n9893) );
  AOI21_X1 U11071 ( .B1(n9890), .B2(n9889), .A(n9888), .ZN(n9891) );
  NAND2_X1 U11072 ( .A1(n9942), .A2(n9891), .ZN(n9892) );
  OAI211_X1 U11073 ( .C1(n9952), .C2(n9894), .A(n9893), .B(n9892), .ZN(n9895)
         );
  INV_X1 U11074 ( .A(n9895), .ZN(n9897) );
  OAI211_X1 U11075 ( .C1(n9956), .C2(n9898), .A(n9897), .B(n9896), .ZN(
        P1_U3257) );
  INV_X1 U11076 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9911) );
  AOI211_X1 U11077 ( .C1(n9902), .C2(n9901), .A(n9900), .B(n9899), .ZN(n9906)
         );
  AOI211_X1 U11078 ( .C1(n9904), .C2(n7646), .A(n9903), .B(n9916), .ZN(n9905)
         );
  AOI211_X1 U11079 ( .C1(n9908), .C2(n9907), .A(n9906), .B(n9905), .ZN(n9910)
         );
  OAI211_X1 U11080 ( .C1(n9956), .C2(n9911), .A(n9910), .B(n9909), .ZN(
        P1_U3258) );
  INV_X1 U11081 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9925) );
  OAI21_X1 U11082 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(n9922) );
  NOR2_X1 U11083 ( .A1(n9952), .A2(n9915), .ZN(n9921) );
  AOI211_X1 U11084 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9920)
         );
  AOI211_X1 U11085 ( .C1(n9946), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9924)
         );
  OAI211_X1 U11086 ( .C1(n9956), .C2(n9925), .A(n9924), .B(n9923), .ZN(
        P1_U3259) );
  INV_X1 U11087 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9939) );
  INV_X1 U11088 ( .A(n9926), .ZN(n9935) );
  XNOR2_X1 U11089 ( .A(n9928), .B(n9927), .ZN(n9929) );
  NAND2_X1 U11090 ( .A1(n9942), .A2(n9929), .ZN(n9934) );
  XNOR2_X1 U11091 ( .A(n9931), .B(n9930), .ZN(n9932) );
  NAND2_X1 U11092 ( .A1(n9946), .A2(n9932), .ZN(n9933) );
  OAI211_X1 U11093 ( .C1(n9952), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9936)
         );
  INV_X1 U11094 ( .A(n9936), .ZN(n9938) );
  OAI211_X1 U11095 ( .C1(n9956), .C2(n9939), .A(n9938), .B(n9937), .ZN(
        P1_U3260) );
  INV_X1 U11096 ( .A(n9940), .ZN(n9951) );
  OAI211_X1 U11097 ( .C1(n9944), .C2(n9943), .A(n9942), .B(n9941), .ZN(n9950)
         );
  OAI211_X1 U11098 ( .C1(n9948), .C2(n9947), .A(n9946), .B(n9945), .ZN(n9949)
         );
  OAI211_X1 U11099 ( .C1(n9952), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9953)
         );
  INV_X1 U11100 ( .A(n9953), .ZN(n9955) );
  OAI211_X1 U11101 ( .C1(n9956), .C2(n10232), .A(n9955), .B(n9954), .ZN(
        P1_U3261) );
  AND2_X1 U11102 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9957), .ZN(P1_U3294) );
  AND2_X1 U11103 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9957), .ZN(P1_U3295) );
  AND2_X1 U11104 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9957), .ZN(P1_U3296) );
  AND2_X1 U11105 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9957), .ZN(P1_U3297) );
  AND2_X1 U11106 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9957), .ZN(P1_U3298) );
  AND2_X1 U11107 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9957), .ZN(P1_U3299) );
  AND2_X1 U11108 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9957), .ZN(P1_U3300) );
  AND2_X1 U11109 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9957), .ZN(P1_U3301) );
  AND2_X1 U11110 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9957), .ZN(P1_U3302) );
  AND2_X1 U11111 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9957), .ZN(P1_U3303) );
  AND2_X1 U11112 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9957), .ZN(P1_U3304) );
  AND2_X1 U11113 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9957), .ZN(P1_U3305) );
  AND2_X1 U11114 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9957), .ZN(P1_U3306) );
  AND2_X1 U11115 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9957), .ZN(P1_U3307) );
  AND2_X1 U11116 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9957), .ZN(P1_U3308) );
  AND2_X1 U11117 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9957), .ZN(P1_U3309) );
  AND2_X1 U11118 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9957), .ZN(P1_U3310) );
  AND2_X1 U11119 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9957), .ZN(P1_U3311) );
  AND2_X1 U11120 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9957), .ZN(P1_U3312) );
  AND2_X1 U11121 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9957), .ZN(P1_U3313) );
  AND2_X1 U11122 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9957), .ZN(P1_U3314) );
  AND2_X1 U11123 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9957), .ZN(P1_U3315) );
  AND2_X1 U11124 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9957), .ZN(P1_U3316) );
  AND2_X1 U11125 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9957), .ZN(P1_U3317) );
  AND2_X1 U11126 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9957), .ZN(P1_U3318) );
  AND2_X1 U11127 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9957), .ZN(P1_U3319) );
  AND2_X1 U11128 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9957), .ZN(P1_U3320) );
  AND2_X1 U11129 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9957), .ZN(P1_U3321) );
  AND2_X1 U11130 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9957), .ZN(P1_U3322) );
  AND2_X1 U11131 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9957), .ZN(P1_U3323) );
  OAI21_X1 U11132 ( .B1(n9959), .B2(n9975), .A(n9958), .ZN(n9961) );
  AOI211_X1 U11133 ( .C1(n9978), .C2(n9962), .A(n9961), .B(n9960), .ZN(n9982)
         );
  AOI22_X1 U11134 ( .A1(n9981), .A2(n9982), .B1(n5115), .B2(n9980), .ZN(
        P1_U3465) );
  OAI21_X1 U11135 ( .B1(n9964), .B2(n9975), .A(n9963), .ZN(n9966) );
  AOI211_X1 U11136 ( .C1(n9978), .C2(n9967), .A(n9966), .B(n9965), .ZN(n9984)
         );
  AOI22_X1 U11137 ( .A1(n9981), .A2(n9984), .B1(n5170), .B2(n9980), .ZN(
        P1_U3471) );
  OAI211_X1 U11138 ( .C1(n4763), .C2(n9975), .A(n9970), .B(n9969), .ZN(n9971)
         );
  AOI21_X1 U11139 ( .B1(n9978), .B2(n9972), .A(n9971), .ZN(n9985) );
  AOI22_X1 U11140 ( .A1(n9981), .A2(n9985), .B1(n5245), .B2(n9980), .ZN(
        P1_U3480) );
  OAI211_X1 U11141 ( .C1(n9976), .C2(n9975), .A(n9974), .B(n9973), .ZN(n9977)
         );
  AOI21_X1 U11142 ( .B1(n9979), .B2(n9978), .A(n9977), .ZN(n9987) );
  AOI22_X1 U11143 ( .A1(n9981), .A2(n9987), .B1(n5328), .B2(n9980), .ZN(
        P1_U3483) );
  AOI22_X1 U11144 ( .A1(n9988), .A2(n9982), .B1(n5114), .B2(n9986), .ZN(
        P1_U3526) );
  INV_X1 U11145 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U11146 ( .A1(n9988), .A2(n9984), .B1(n9983), .B2(n9986), .ZN(
        P1_U3528) );
  AOI22_X1 U11147 ( .A1(n9988), .A2(n9985), .B1(n5244), .B2(n9986), .ZN(
        P1_U3531) );
  AOI22_X1 U11148 ( .A1(n9988), .A2(n9987), .B1(n5327), .B2(n9986), .ZN(
        P1_U3532) );
  XNOR2_X1 U11149 ( .A(n9989), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n9993) );
  OAI21_X1 U11150 ( .B1(n9991), .B2(P2_REG2_REG_3__SCAN_IN), .A(n9990), .ZN(
        n9992) );
  AOI22_X1 U11151 ( .A1(n10116), .A2(n9993), .B1(n10010), .B2(n9992), .ZN(
        n9994) );
  INV_X1 U11152 ( .A(n9994), .ZN(n9995) );
  AOI211_X1 U11153 ( .C1(n4734), .C2(n10107), .A(n9996), .B(n9995), .ZN(n10002) );
  OAI21_X1 U11154 ( .B1(n9999), .B2(n9998), .A(n9997), .ZN(n10000) );
  AOI22_X1 U11155 ( .A1(n10000), .A2(n10115), .B1(n10106), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U11156 ( .A1(n10002), .A2(n10001), .ZN(P2_U3185) );
  INV_X1 U11157 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10019) );
  AOI211_X1 U11158 ( .C1(n10006), .C2(n10005), .A(n10004), .B(n10003), .ZN(
        n10017) );
  XNOR2_X1 U11159 ( .A(n10007), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n10011) );
  OAI21_X1 U11160 ( .B1(n4448), .B2(P2_REG2_REG_5__SCAN_IN), .A(n10008), .ZN(
        n10009) );
  AOI22_X1 U11161 ( .A1(n10116), .A2(n10011), .B1(n10010), .B2(n10009), .ZN(
        n10014) );
  INV_X1 U11162 ( .A(n10012), .ZN(n10013) );
  OAI211_X1 U11163 ( .C1(n10027), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10016) );
  NOR2_X1 U11164 ( .A1(n10017), .A2(n10016), .ZN(n10018) );
  OAI21_X1 U11165 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(P2_U3187) );
  OAI21_X1 U11166 ( .B1(n10023), .B2(n10022), .A(n10021), .ZN(n10036) );
  INV_X1 U11167 ( .A(n10024), .ZN(n10025) );
  OAI21_X1 U11168 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(n10035) );
  INV_X1 U11169 ( .A(n10028), .ZN(n10030) );
  NAND3_X1 U11170 ( .A1(n10031), .A2(n10030), .A3(n10029), .ZN(n10032) );
  AOI21_X1 U11171 ( .B1(n10033), .B2(n10032), .A(n10122), .ZN(n10034) );
  AOI211_X1 U11172 ( .C1(n10116), .C2(n10036), .A(n10035), .B(n10034), .ZN(
        n10041) );
  XNOR2_X1 U11173 ( .A(n10038), .B(n10037), .ZN(n10039) );
  AOI22_X1 U11174 ( .A1(n10039), .A2(n10115), .B1(n10106), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U11175 ( .A1(n10041), .A2(n10040), .ZN(P2_U3190) );
  AOI22_X1 U11176 ( .A1(n10042), .A2(n10107), .B1(n10106), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10057) );
  OAI21_X1 U11177 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10044), .A(n10043), 
        .ZN(n10049) );
  OAI21_X1 U11178 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(n10048) );
  AOI22_X1 U11179 ( .A1(n10049), .A2(n10116), .B1(n10115), .B2(n10048), .ZN(
        n10056) );
  AOI21_X1 U11180 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(n10053) );
  OR2_X1 U11181 ( .A1(n10053), .A2(n10122), .ZN(n10054) );
  NAND4_X1 U11182 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        P2_U3195) );
  AOI22_X1 U11183 ( .A1(n10058), .A2(n10107), .B1(n10106), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10073) );
  OAI21_X1 U11184 ( .B1(n10061), .B2(n10060), .A(n10059), .ZN(n10066) );
  OAI21_X1 U11185 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(n10065) );
  AOI22_X1 U11186 ( .A1(n10066), .A2(n10116), .B1(n10115), .B2(n10065), .ZN(
        n10072) );
  AOI21_X1 U11187 ( .B1(n4432), .B2(n10068), .A(n10067), .ZN(n10069) );
  OR2_X1 U11188 ( .A1(n10069), .A2(n10122), .ZN(n10070) );
  NAND4_X1 U11189 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        P2_U3196) );
  AOI22_X1 U11190 ( .A1(n10074), .A2(n10107), .B1(n10106), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n10089) );
  OAI21_X1 U11191 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10076), .A(n10075), 
        .ZN(n10081) );
  OAI21_X1 U11192 ( .B1(n10079), .B2(n10078), .A(n10077), .ZN(n10080) );
  AOI22_X1 U11193 ( .A1(n10081), .A2(n10116), .B1(n10115), .B2(n10080), .ZN(
        n10088) );
  AOI21_X1 U11194 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(n10085) );
  OR2_X1 U11195 ( .A1(n10122), .A2(n10085), .ZN(n10086) );
  NAND4_X1 U11196 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        P2_U3197) );
  AOI22_X1 U11197 ( .A1(n10090), .A2(n10107), .B1(n10106), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10105) );
  OAI21_X1 U11198 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(n10098) );
  OAI21_X1 U11199 ( .B1(n10096), .B2(n10095), .A(n10094), .ZN(n10097) );
  AOI22_X1 U11200 ( .A1(n10098), .A2(n10116), .B1(n10115), .B2(n10097), .ZN(
        n10104) );
  AOI21_X1 U11201 ( .B1(n4430), .B2(n10100), .A(n10099), .ZN(n10101) );
  OR2_X1 U11202 ( .A1(n10101), .A2(n10122), .ZN(n10102) );
  NAND4_X1 U11203 ( .A1(n10105), .A2(n10104), .A3(n10103), .A4(n10102), .ZN(
        P2_U3198) );
  AOI22_X1 U11204 ( .A1(n10108), .A2(n10107), .B1(n10106), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10126) );
  OAI21_X1 U11205 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10110), .A(n10109), 
        .ZN(n10117) );
  OAI21_X1 U11206 ( .B1(n10113), .B2(n10112), .A(n10111), .ZN(n10114) );
  AOI22_X1 U11207 ( .A1(n10117), .A2(n10116), .B1(n10115), .B2(n10114), .ZN(
        n10125) );
  AOI21_X1 U11208 ( .B1(n10120), .B2(n10119), .A(n10118), .ZN(n10121) );
  OR2_X1 U11209 ( .A1(n10122), .A2(n10121), .ZN(n10123) );
  NAND4_X1 U11210 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        P2_U3199) );
  XNOR2_X1 U11211 ( .A(n10128), .B(n10127), .ZN(n10133) );
  AOI222_X1 U11212 ( .A1(n10134), .A2(n10133), .B1(n10132), .B2(n10131), .C1(
        n10130), .C2(n10129), .ZN(n10161) );
  INV_X1 U11213 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10144) );
  XNOR2_X1 U11214 ( .A(n10135), .B(n10136), .ZN(n10164) );
  INV_X1 U11215 ( .A(n10137), .ZN(n10141) );
  AOI222_X1 U11216 ( .A1(n10164), .A2(n10142), .B1(n10141), .B2(n10140), .C1(
        n10139), .C2(n10138), .ZN(n10143) );
  OAI221_X1 U11217 ( .B1(n10146), .B2(n10161), .C1(n10145), .C2(n10144), .A(
        n10143), .ZN(P2_U3229) );
  INV_X1 U11218 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10151) );
  OAI22_X1 U11219 ( .A1(n10148), .A2(n10192), .B1(n10147), .B2(n10186), .ZN(
        n10149) );
  NOR2_X1 U11220 ( .A1(n10150), .A2(n10149), .ZN(n10209) );
  AOI22_X1 U11221 ( .A1(n10207), .A2(n10151), .B1(n10209), .B2(n10205), .ZN(
        P2_U3393) );
  INV_X1 U11222 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10155) );
  OAI22_X1 U11223 ( .A1(n10152), .A2(n10192), .B1(n6402), .B2(n10186), .ZN(
        n10153) );
  NOR2_X1 U11224 ( .A1(n10154), .A2(n10153), .ZN(n10210) );
  AOI22_X1 U11225 ( .A1(n10207), .A2(n10155), .B1(n10210), .B2(n10205), .ZN(
        P2_U3396) );
  INV_X1 U11226 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U11227 ( .A1(n10157), .A2(n10198), .B1(n10200), .B2(n10156), .ZN(
        n10158) );
  AND2_X1 U11228 ( .A1(n10159), .A2(n10158), .ZN(n10211) );
  AOI22_X1 U11229 ( .A1(n10207), .A2(n10160), .B1(n10211), .B2(n10205), .ZN(
        P2_U3399) );
  INV_X1 U11230 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10165) );
  OAI21_X1 U11231 ( .B1(n10162), .B2(n10186), .A(n10161), .ZN(n10163) );
  AOI21_X1 U11232 ( .B1(n10198), .B2(n10164), .A(n10163), .ZN(n10212) );
  AOI22_X1 U11233 ( .A1(n10207), .A2(n10165), .B1(n10212), .B2(n10205), .ZN(
        P2_U3402) );
  INV_X1 U11234 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10170) );
  NOR2_X1 U11235 ( .A1(n10166), .A2(n10186), .ZN(n10168) );
  AOI211_X1 U11236 ( .C1(n10198), .C2(n10169), .A(n10168), .B(n10167), .ZN(
        n10214) );
  AOI22_X1 U11237 ( .A1(n10207), .A2(n10170), .B1(n10214), .B2(n10205), .ZN(
        P2_U3405) );
  INV_X1 U11238 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U11239 ( .A1(n10171), .A2(n10198), .ZN(n10175) );
  NAND2_X1 U11240 ( .A1(n10172), .A2(n10200), .ZN(n10173) );
  AND3_X1 U11241 ( .A1(n10175), .A2(n10174), .A3(n10173), .ZN(n10215) );
  AOI22_X1 U11242 ( .A1(n10207), .A2(n10176), .B1(n10215), .B2(n10205), .ZN(
        P2_U3408) );
  INV_X1 U11243 ( .A(n10177), .ZN(n10179) );
  OAI22_X1 U11244 ( .A1(n10179), .A2(n10192), .B1(n10178), .B2(n10186), .ZN(
        n10180) );
  NOR2_X1 U11245 ( .A1(n10181), .A2(n10180), .ZN(n10217) );
  AOI22_X1 U11246 ( .A1(n10207), .A2(n6048), .B1(n10217), .B2(n10205), .ZN(
        P2_U3411) );
  NOR2_X1 U11247 ( .A1(n10182), .A2(n10186), .ZN(n10184) );
  AOI211_X1 U11248 ( .C1(n10198), .C2(n10185), .A(n10184), .B(n10183), .ZN(
        n10218) );
  AOI22_X1 U11249 ( .A1(n10207), .A2(n6060), .B1(n10218), .B2(n10205), .ZN(
        P2_U3414) );
  INV_X1 U11250 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10191) );
  OAI22_X1 U11251 ( .A1(n10188), .A2(n10192), .B1(n10187), .B2(n10186), .ZN(
        n10189) );
  NOR2_X1 U11252 ( .A1(n10190), .A2(n10189), .ZN(n10220) );
  AOI22_X1 U11253 ( .A1(n10207), .A2(n10191), .B1(n10220), .B2(n10205), .ZN(
        P2_U3417) );
  INV_X1 U11254 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10197) );
  INV_X1 U11255 ( .A(n10192), .ZN(n10193) );
  AOI22_X1 U11256 ( .A1(n10194), .A2(n10193), .B1(n10200), .B2(n6092), .ZN(
        n10195) );
  AND2_X1 U11257 ( .A1(n10196), .A2(n10195), .ZN(n10221) );
  AOI22_X1 U11258 ( .A1(n10207), .A2(n10197), .B1(n10221), .B2(n10205), .ZN(
        P2_U3420) );
  INV_X1 U11259 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10206) );
  NAND2_X1 U11260 ( .A1(n10199), .A2(n10198), .ZN(n10204) );
  NAND2_X1 U11261 ( .A1(n10201), .A2(n10200), .ZN(n10202) );
  AND3_X1 U11262 ( .A1(n10204), .A2(n10203), .A3(n10202), .ZN(n10224) );
  AOI22_X1 U11263 ( .A1(n10207), .A2(n10206), .B1(n10224), .B2(n10205), .ZN(
        P2_U3423) );
  INV_X1 U11264 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U11265 ( .A1(n10225), .A2(n10209), .B1(n10208), .B2(n10222), .ZN(
        P2_U3460) );
  AOI22_X1 U11266 ( .A1(n10225), .A2(n10210), .B1(n7331), .B2(n10222), .ZN(
        P2_U3461) );
  AOI22_X1 U11267 ( .A1(n10225), .A2(n10211), .B1(n6002), .B2(n10222), .ZN(
        P2_U3462) );
  AOI22_X1 U11268 ( .A1(n10225), .A2(n10212), .B1(n7330), .B2(n10222), .ZN(
        P2_U3463) );
  INV_X1 U11269 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U11270 ( .A1(n10225), .A2(n10214), .B1(n10213), .B2(n10222), .ZN(
        P2_U3464) );
  AOI22_X1 U11271 ( .A1(n10225), .A2(n10215), .B1(n7412), .B2(n10222), .ZN(
        P2_U3465) );
  INV_X1 U11272 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U11273 ( .A1(n10225), .A2(n10217), .B1(n10216), .B2(n10222), .ZN(
        P2_U3466) );
  AOI22_X1 U11274 ( .A1(n10225), .A2(n10218), .B1(n7747), .B2(n10222), .ZN(
        P2_U3467) );
  AOI22_X1 U11275 ( .A1(n10225), .A2(n10220), .B1(n10219), .B2(n10222), .ZN(
        P2_U3468) );
  AOI22_X1 U11276 ( .A1(n10225), .A2(n10221), .B1(n7735), .B2(n10222), .ZN(
        P2_U3469) );
  INV_X1 U11277 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U11278 ( .A1(n10225), .A2(n10224), .B1(n10223), .B2(n10222), .ZN(
        P2_U3470) );
  OAI222_X1 U11279 ( .A1(n10230), .A2(n10229), .B1(n10230), .B2(n10228), .C1(
        n10227), .C2(n10226), .ZN(ADD_1068_U5) );
  XOR2_X1 U11280 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11281 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(n10234) );
  XOR2_X1 U11282 ( .A(n10234), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11283 ( .B1(n10237), .B2(n10236), .A(n10235), .ZN(ADD_1068_U56) );
  OAI21_X1 U11284 ( .B1(n10240), .B2(n10239), .A(n10238), .ZN(ADD_1068_U57) );
  OAI21_X1 U11285 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(ADD_1068_U58) );
  OAI21_X1 U11286 ( .B1(n10246), .B2(n10245), .A(n10244), .ZN(ADD_1068_U59) );
  OAI21_X1 U11287 ( .B1(n10249), .B2(n10248), .A(n10247), .ZN(ADD_1068_U60) );
  OAI21_X1 U11288 ( .B1(n10252), .B2(n10251), .A(n10250), .ZN(ADD_1068_U61) );
  OAI21_X1 U11289 ( .B1(n10255), .B2(n10254), .A(n10253), .ZN(ADD_1068_U62) );
  OAI21_X1 U11290 ( .B1(n10258), .B2(n10257), .A(n10256), .ZN(ADD_1068_U63) );
  AOI21_X1 U11291 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(ADD_1068_U54) );
  OAI21_X1 U11292 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(ADD_1068_U47) );
  OAI21_X1 U11293 ( .B1(n10267), .B2(n10266), .A(n10265), .ZN(ADD_1068_U48) );
  OAI21_X1 U11294 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(ADD_1068_U49) );
  OAI21_X1 U11295 ( .B1(n10273), .B2(n10272), .A(n10271), .ZN(ADD_1068_U50) );
  OAI21_X1 U11296 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(ADD_1068_U51) );
  AOI21_X1 U11297 ( .B1(n10279), .B2(n10278), .A(n10277), .ZN(ADD_1068_U53) );
  OAI21_X1 U11298 ( .B1(n10282), .B2(n10281), .A(n10280), .ZN(ADD_1068_U52) );
  NAND2_X1 U4931 ( .A1(n6431), .A2(n6430), .ZN(n8362) );
  CLKBUF_X1 U4978 ( .A(n5052), .Z(n6611) );
  CLKBUF_X1 U5082 ( .A(n8822), .Z(n4353) );
endmodule

