

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108;

  AND2_X1 U5175 ( .A1(n5491), .A2(n5489), .ZN(n7241) );
  OAI21_X1 U5176 ( .B1(n7088), .B2(n7087), .A(n6981), .ZN(n6984) );
  XNOR2_X1 U5177 ( .A(n6218), .B(n6217), .ZN(n10085) );
  XNOR2_X1 U5178 ( .A(n6230), .B(n6231), .ZN(n10081) );
  AND2_X1 U5179 ( .A1(n5221), .A2(n5219), .ZN(n9060) );
  CLKBUF_X2 U5181 ( .A(n6327), .Z(n9756) );
  CLKBUF_X2 U5182 ( .A(n5889), .Z(n9251) );
  NAND2_X1 U5183 ( .A1(n5308), .A2(n5307), .ZN(n9326) );
  AND4_X1 U5185 ( .A1(n6512), .A2(n6511), .A3(n6510), .A4(n6509), .ZN(n7011)
         );
  NAND2_X1 U5186 ( .A1(n6407), .A2(n6410), .ZN(n10795) );
  NAND2_X1 U5187 ( .A1(n6406), .A2(n6405), .ZN(n6959) );
  AOI22_X1 U5188 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n9175), .B1(n9174), .B2(
        n9173), .ZN(n9667) );
  AND2_X1 U5189 ( .A1(n6321), .A2(n5630), .ZN(n5282) );
  NOR2_X1 U5190 ( .A1(n5621), .A2(n7860), .ZN(n5307) );
  AOI21_X1 U5191 ( .B1(n10186), .B2(n5655), .A(n5657), .ZN(n5653) );
  XNOR2_X1 U5192 ( .A(n10257), .B(n7009), .ZN(n7620) );
  NAND2_X1 U5193 ( .A1(n8953), .A2(n10980), .ZN(n9173) );
  NOR2_X1 U5194 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  NAND2_X1 U5195 ( .A1(n7082), .A2(n7081), .ZN(n10620) );
  NAND2_X1 U5196 ( .A1(n6050), .A2(n5531), .ZN(n5528) );
  AND2_X1 U5197 ( .A1(n6400), .A2(n8479), .ZN(n5674) );
  OR2_X1 U5198 ( .A1(n9497), .A2(n9496), .ZN(n9575) );
  INV_X1 U5200 ( .A(n6250), .ZN(n9249) );
  BUF_X1 U5201 ( .A(n5854), .Z(n7449) );
  INV_X1 U5202 ( .A(n7257), .ZN(n6485) );
  INV_X1 U5203 ( .A(n6946), .ZN(n6444) );
  INV_X1 U5204 ( .A(n8701), .ZN(n8110) );
  AND3_X1 U5205 ( .A1(n6532), .A2(n6531), .A3(n6530), .ZN(n7919) );
  MUX2_X1 U5206 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6404), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n6406) );
  OAI21_X1 U5207 ( .B1(n6425), .B2(n6424), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6426) );
  INV_X1 U5208 ( .A(n5851), .ZN(n9266) );
  OAI211_X1 U5209 ( .C1(n6872), .C2(n7295), .A(n6508), .B(n6507), .ZN(n10198)
         );
  MUX2_X1 U5210 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6409), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n6410) );
  NAND2_X1 U5212 ( .A1(n7257), .A2(n6885), .ZN(n6497) );
  INV_X2 U5213 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8479) );
  OR2_X1 U5214 ( .A1(n9861), .A2(n6312), .ZN(n6314) );
  NAND4_X1 U5215 ( .A1(n6495), .A2(n6494), .A3(n6492), .A4(n6493), .ZN(n10257)
         );
  NAND2_X2 U5216 ( .A1(n5855), .A2(n7342), .ZN(n7441) );
  NOR2_X1 U5217 ( .A1(n7582), .A2(n7581), .ZN(n7681) );
  NAND2_X2 U5218 ( .A1(n6824), .A2(n6823), .ZN(n10545) );
  OAI21_X2 U5219 ( .B1(n7643), .B2(n6277), .A(n6276), .ZN(n7787) );
  NAND2_X2 U5220 ( .A1(n6275), .A2(n6274), .ZN(n7643) );
  INV_X1 U5221 ( .A(n6497), .ZN(n5112) );
  INV_X1 U5222 ( .A(n5112), .ZN(n5113) );
  AOI21_X2 U5223 ( .B1(n6190), .B2(n6189), .A(n5784), .ZN(n6204) );
  AOI21_X2 U5224 ( .B1(n5282), .B2(n5280), .A(n9436), .ZN(n5279) );
  OAI21_X2 U5225 ( .B1(n8910), .B2(n9644), .A(n5687), .ZN(n8965) );
  XNOR2_X2 U5226 ( .A(n8909), .B(n8908), .ZN(n8910) );
  XNOR2_X2 U5228 ( .A(n7088), .B(n7087), .ZN(n9244) );
  OAI21_X2 U5229 ( .B1(n7827), .B2(n6280), .A(n6279), .ZN(n8011) );
  OAI22_X2 U5230 ( .A1(n7787), .A2(n6278), .B1(n7559), .B2(n7644), .ZN(n7827)
         );
  AND2_X1 U5231 ( .A1(n7217), .A2(n7159), .ZN(n9073) );
  OR2_X1 U5232 ( .A1(n8827), .A2(n5222), .ZN(n5221) );
  INV_X2 U5233 ( .A(n8717), .ZN(n10253) );
  AND4_X1 U5234 ( .A1(n6563), .A2(n6562), .A3(n6561), .A4(n6560), .ZN(n8717)
         );
  NAND4_X2 U5235 ( .A1(n6523), .A2(n6522), .A3(n6521), .A4(n6520), .ZN(n10255)
         );
  INV_X1 U5236 ( .A(n6271), .ZN(n5573) );
  NAND2_X1 U5237 ( .A1(n6995), .A2(n6518), .ZN(n6522) );
  INV_X1 U5238 ( .A(n8634), .ZN(n10254) );
  CLKBUF_X2 U5239 ( .A(n6525), .Z(n5115) );
  INV_X1 U5240 ( .A(n7644), .ZN(n7828) );
  INV_X2 U5241 ( .A(n6273), .ZN(n5427) );
  NAND2_X1 U5242 ( .A1(n6942), .A2(n6431), .ZN(n6483) );
  CLKBUF_X2 U5243 ( .A(n5899), .Z(n6250) );
  AND2_X1 U5244 ( .A1(n5640), .A2(n5805), .ZN(n5299) );
  INV_X1 U5245 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5689) );
  OAI21_X1 U5246 ( .B1(n6337), .B2(n11105), .A(n5678), .ZN(n5199) );
  AOI21_X1 U5247 ( .B1(n9791), .B2(n6325), .A(n9790), .ZN(n9968) );
  XNOR2_X1 U5248 ( .A(n9264), .B(n6254), .ZN(n9775) );
  OR2_X1 U5249 ( .A1(n10379), .A2(n7102), .ZN(n7245) );
  NAND2_X1 U5250 ( .A1(n10520), .A2(n10417), .ZN(n10504) );
  NAND2_X1 U5251 ( .A1(n6987), .A2(n6986), .ZN(n10379) );
  AND2_X1 U5252 ( .A1(n9269), .A2(n9268), .ZN(n5683) );
  OAI21_X1 U5253 ( .B1(n9440), .B2(n9439), .A(n9438), .ZN(n9444) );
  NAND2_X1 U5254 ( .A1(n10550), .A2(n10555), .ZN(n10549) );
  NAND2_X1 U5255 ( .A1(n6234), .A2(n6233), .ZN(n6268) );
  NAND2_X1 U5256 ( .A1(n6888), .A2(n6887), .ZN(n10487) );
  NAND2_X1 U5257 ( .A1(n6221), .A2(n6220), .ZN(n9630) );
  NAND2_X1 U5258 ( .A1(n6874), .A2(n6873), .ZN(n10647) );
  CLKBUF_X1 U5259 ( .A(n7070), .Z(n10529) );
  NAND2_X1 U5260 ( .A1(n5575), .A2(n5574), .ZN(n9566) );
  OAI21_X1 U5261 ( .B1(n6177), .B2(n6176), .A(n5781), .ZN(n6190) );
  AOI21_X1 U5262 ( .B1(n5434), .B2(n5433), .A(n5430), .ZN(n9398) );
  OR2_X1 U5263 ( .A1(n9717), .A2(n9716), .ZN(n5475) );
  OR2_X1 U5264 ( .A1(n5776), .A2(n5775), .ZN(n5777) );
  NOR2_X1 U5265 ( .A1(n9053), .A2(n5386), .ZN(n5384) );
  NAND2_X1 U5266 ( .A1(n8664), .A2(n8122), .ZN(n8124) );
  NAND2_X1 U5267 ( .A1(n8770), .A2(n5670), .ZN(n8827) );
  INV_X1 U5268 ( .A(n9805), .ZN(n9636) );
  OAI21_X1 U5269 ( .B1(n8628), .B2(n8631), .A(n8629), .ZN(n8608) );
  INV_X1 U5270 ( .A(n8681), .ZN(n9064) );
  NAND2_X1 U5271 ( .A1(n5248), .A2(n6632), .ZN(n8681) );
  INV_X1 U5272 ( .A(n9092), .ZN(n8646) );
  NOR3_X2 U5273 ( .A1(n7681), .A2(n7680), .A3(n7679), .ZN(n7965) );
  AND2_X1 U5274 ( .A1(n5953), .A2(n5952), .ZN(n8548) );
  NAND2_X1 U5275 ( .A1(n6596), .A2(n6595), .ZN(n8701) );
  AND2_X1 U5276 ( .A1(n5972), .A2(n5971), .ZN(n8803) );
  NAND2_X1 U5277 ( .A1(n7592), .A2(n7591), .ZN(n7921) );
  NAND2_X1 U5278 ( .A1(n7760), .A2(n7761), .ZN(n7878) );
  INV_X1 U5279 ( .A(n7919), .ZN(n8748) );
  INV_X1 U5280 ( .A(n9280), .ZN(n6269) );
  NAND2_X1 U5281 ( .A1(n7701), .A2(n7702), .ZN(n7756) );
  AND3_X1 U5282 ( .A1(n5885), .A2(n5884), .A3(n5883), .ZN(n7648) );
  NAND2_X2 U5283 ( .A1(n6489), .A2(n6483), .ZN(n6885) );
  NAND2_X1 U5284 ( .A1(n5876), .A2(n5875), .ZN(n5878) );
  NAND4_X1 U5285 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n10258)
         );
  NAND2_X1 U5286 ( .A1(n5485), .A2(n5484), .ZN(n7699) );
  OR2_X1 U5287 ( .A1(n5851), .A2(n7288), .ZN(n5437) );
  INV_X1 U5288 ( .A(n5817), .ZN(n9267) );
  NAND2_X1 U5289 ( .A1(n7697), .A2(n7698), .ZN(n10926) );
  NAND2_X1 U5290 ( .A1(n6443), .A2(n6944), .ZN(n6946) );
  CLKBUF_X1 U5291 ( .A(n6959), .Z(n10271) );
  INV_X2 U5292 ( .A(n5845), .ZN(n5817) );
  INV_X1 U5293 ( .A(n9026), .ZN(n7734) );
  NOR2_X1 U5294 ( .A1(n6430), .A2(n6429), .ZN(n10797) );
  OR2_X1 U5295 ( .A1(n9458), .A2(n9762), .ZN(n9026) );
  NAND2_X2 U5296 ( .A1(n5832), .A2(n5829), .ZN(n6237) );
  OR2_X1 U5297 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  OR2_X1 U5298 ( .A1(n6448), .A2(n8518), .ZN(n5207) );
  OAI21_X1 U5299 ( .B1(n7453), .B2(n7811), .A(n10899), .ZN(n7695) );
  NAND2_X2 U5300 ( .A1(n7359), .A2(n6327), .ZN(n5852) );
  NAND2_X1 U5301 ( .A1(n6434), .A2(n6433), .ZN(n8920) );
  NAND2_X1 U5302 ( .A1(n6753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6438) );
  XNOR2_X1 U5303 ( .A(n5821), .B(n10069), .ZN(n5828) );
  NAND2_X1 U5304 ( .A1(n6349), .A2(n6348), .ZN(n10088) );
  XNOR2_X1 U5305 ( .A(n5825), .B(n5824), .ZN(n5826) );
  AND2_X1 U5306 ( .A1(n6343), .A2(n5146), .ZN(n6369) );
  NAND2_X1 U5307 ( .A1(n5727), .A2(SI_7_), .ZN(n5730) );
  XNOR2_X1 U5308 ( .A(n6255), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U5309 ( .A1(n10068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  OR2_X1 U5310 ( .A1(n5823), .A2(n5822), .ZN(n5825) );
  MUX2_X1 U5311 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5813), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5815) );
  NOR2_X1 U5312 ( .A1(n5700), .A2(n6475), .ZN(n5846) );
  XNOR2_X1 U5313 ( .A(n5911), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10934) );
  OR2_X1 U5314 ( .A1(n7345), .A2(n7344), .ZN(n7451) );
  NAND2_X1 U5315 ( .A1(n5814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5812) );
  AND3_X2 U5316 ( .A1(n5867), .A2(n5487), .A3(n5378), .ZN(n7453) );
  NOR2_X1 U5317 ( .A1(n5209), .A2(n5314), .ZN(n5679) );
  OR2_X1 U5318 ( .A1(n7449), .A2(n5379), .ZN(n5378) );
  AND2_X1 U5319 ( .A1(n5809), .A2(n5810), .ZN(n5640) );
  AND3_X1 U5320 ( .A1(n6261), .A2(n6260), .A3(n6259), .ZN(n6338) );
  AND4_X1 U5321 ( .A1(n5808), .A2(n5807), .A3(n5806), .A4(n6260), .ZN(n5809)
         );
  OAI21_X2 U5322 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n5689), .ZN(n5693) );
  AND2_X1 U5323 ( .A1(n6420), .A2(n6419), .ZN(n5313) );
  AND2_X1 U5324 ( .A1(n8311), .A2(n5312), .ZN(n5311) );
  INV_X1 U5325 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6260) );
  NOR2_X1 U5326 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5801) );
  NOR2_X1 U5327 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5802) );
  NOR2_X1 U5328 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5797) );
  NOR2_X1 U5329 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5798) );
  NOR2_X1 U5330 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5799) );
  INV_X1 U5331 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5690) );
  INV_X4 U5332 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X2 U5333 ( .B1(n5931), .B2(n5129), .A(n5244), .ZN(n5243) );
  AND2_X1 U5334 ( .A1(n5828), .A2(n5826), .ZN(n5899) );
  NAND2_X1 U5335 ( .A1(n5828), .A2(n5829), .ZN(n6181) );
  AOI21_X1 U5336 ( .B1(n5402), .B2(n5400), .A(n5398), .ZN(n9433) );
  AOI22_X2 U5337 ( .A1(n9060), .A2(n6645), .B1(n6644), .B2(n9057), .ZN(n9186)
         );
  OAI222_X1 U5338 ( .A1(n8895), .A2(P1_U3086), .B1(n9234), .B2(n8693), .C1(
        n8692), .C2(n10792), .ZN(P1_U3336) );
  NAND2_X1 U5339 ( .A1(n6444), .A2(n8895), .ZN(n7594) );
  INV_X1 U5341 ( .A(n6872), .ZN(n6525) );
  NOR2_X1 U5342 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6396) );
  INV_X1 U5343 ( .A(n5828), .ZN(n5832) );
  INV_X1 U5344 ( .A(n5826), .ZN(n5829) );
  OR2_X1 U5345 ( .A1(n9996), .A2(n9863), .ZN(n9414) );
  OR2_X1 U5346 ( .A1(n10620), .A2(n10626), .ZN(n7172) );
  NAND2_X1 U5347 ( .A1(n6033), .A2(n5749), .ZN(n6050) );
  INV_X1 U5348 ( .A(n5594), .ZN(n9144) );
  NAND2_X1 U5349 ( .A1(n5601), .A2(n9142), .ZN(n5598) );
  INV_X1 U5350 ( .A(n5596), .ZN(n5595) );
  AND2_X1 U5351 ( .A1(n9545), .A2(n5176), .ZN(n5579) );
  CLKBUF_X1 U5352 ( .A(n6181), .Z(n9247) );
  INV_X1 U5353 ( .A(n6181), .ZN(n6330) );
  NAND2_X1 U5354 ( .A1(n5832), .A2(n5826), .ZN(n5889) );
  INV_X1 U5355 ( .A(n9243), .ZN(n6942) );
  INV_X1 U5356 ( .A(n10421), .ZN(n5549) );
  NAND2_X1 U5357 ( .A1(n6271), .A2(n7860), .ZN(n9321) );
  NOR2_X1 U5358 ( .A1(n9358), .A2(n5414), .ZN(n9360) );
  NAND2_X1 U5359 ( .A1(n5416), .A2(n5415), .ZN(n5414) );
  NOR2_X1 U5360 ( .A1(n9355), .A2(n9356), .ZN(n5415) );
  OR2_X1 U5361 ( .A1(n10009), .A2(n9906), .ZN(n9394) );
  NAND2_X1 U5362 ( .A1(n6268), .A2(n9786), .ZN(n5469) );
  NOR2_X1 U5363 ( .A1(n5645), .A2(n5644), .ZN(n5643) );
  INV_X1 U5364 ( .A(n10206), .ZN(n5644) );
  NOR2_X1 U5365 ( .A1(n5646), .A2(n5647), .ZN(n5645) );
  XNOR2_X1 U5366 ( .A(n6500), .B(n6867), .ZN(n6503) );
  NAND2_X1 U5367 ( .A1(n7180), .A2(n7095), .ZN(n7098) );
  NOR2_X1 U5368 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6506) );
  INV_X1 U5369 ( .A(n8678), .ZN(n5544) );
  XNOR2_X1 U5370 ( .A(n5759), .B(n8165), .ZN(n6098) );
  NAND2_X1 U5371 ( .A1(n5758), .A2(n5757), .ZN(n6099) );
  NOR2_X1 U5372 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6397) );
  NOR2_X1 U5373 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6395) );
  AOI21_X1 U5374 ( .B1(n5497), .B2(n5245), .A(n5168), .ZN(n5495) );
  XNOR2_X1 U5375 ( .A(n5731), .B(SI_8_), .ZN(n5946) );
  OR2_X1 U5376 ( .A1(n7965), .A2(n5617), .ZN(n8018) );
  OR2_X1 U5377 ( .A1(n6237), .A2(n9260), .ZN(n9255) );
  XNOR2_X1 U5378 ( .A(n7699), .B(n10944), .ZN(n10943) );
  OR2_X1 U5379 ( .A1(n9673), .A2(n9672), .ZN(n5477) );
  AOI21_X1 U5380 ( .B1(n5279), .B2(n5281), .A(n5276), .ZN(n5275) );
  AND2_X1 U5381 ( .A1(n5820), .A2(n5819), .ZN(n9441) );
  NAND2_X1 U5382 ( .A1(n5158), .A2(n6228), .ZN(n5630) );
  AND4_X1 U5383 ( .A1(n6199), .A2(n6198), .A3(n6197), .A4(n6196), .ZN(n9830)
         );
  AND4_X1 U5384 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n9841)
         );
  AND4_X1 U5385 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .ZN(n9863)
         );
  INV_X1 U5386 ( .A(n5451), .ZN(n5450) );
  OAI21_X1 U5387 ( .B1(n6304), .B2(n5452), .A(n6306), .ZN(n5451) );
  AND4_X1 U5388 ( .A1(n6109), .A2(n6108), .A3(n6107), .A4(n6106), .ZN(n9955)
         );
  INV_X1 U5389 ( .A(n5446), .ZN(n5445) );
  OAI21_X1 U5390 ( .B1(n5133), .B2(n6291), .A(n6292), .ZN(n5446) );
  AOI21_X1 U5391 ( .B1(n5305), .B2(n5117), .A(n9287), .ZN(n5302) );
  AND4_X1 U5392 ( .A1(n5929), .A2(n5928), .A3(n5927), .A4(n5926), .ZN(n8001)
         );
  INV_X1 U5393 ( .A(n9934), .ZN(n9954) );
  NAND2_X1 U5394 ( .A1(n5852), .A2(n7287), .ZN(n5845) );
  INV_X1 U5395 ( .A(n5852), .ZN(n5879) );
  NAND2_X1 U5396 ( .A1(n7429), .A2(n5422), .ZN(n9956) );
  CLKBUF_X1 U5397 ( .A(n6378), .Z(n7726) );
  OR2_X1 U5398 ( .A1(n9323), .A2(n9465), .ZN(n10027) );
  INV_X1 U5399 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6261) );
  AOI22_X1 U5400 ( .A1(n5643), .A2(n5646), .B1(n5652), .B2(n5649), .ZN(n5641)
         );
  NOR2_X1 U5401 ( .A1(n5224), .A2(n5226), .ZN(n5222) );
  INV_X1 U5402 ( .A(n6771), .ZN(n5652) );
  NAND2_X1 U5403 ( .A1(n6445), .A2(n7594), .ZN(n6446) );
  INV_X1 U5404 ( .A(n6543), .ZN(n6463) );
  NAND2_X1 U5405 ( .A1(n6519), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6492) );
  AND2_X1 U5406 ( .A1(n10620), .A2(n10427), .ZN(n10428) );
  NAND2_X1 U5407 ( .A1(n6992), .A2(n6991), .ZN(n10618) );
  NAND2_X1 U5408 ( .A1(n7171), .A2(n10402), .ZN(n5563) );
  INV_X1 U5409 ( .A(n5563), .ZN(n10471) );
  NAND2_X1 U5410 ( .A1(n10504), .A2(n10418), .ZN(n10420) );
  NAND2_X1 U5411 ( .A1(n10569), .A2(n10378), .ZN(n10570) );
  NAND2_X1 U5412 ( .A1(n10411), .A2(n10410), .ZN(n10568) );
  AOI21_X1 U5413 ( .B1(n9159), .B2(n5538), .A(n5150), .ZN(n5537) );
  INV_X1 U5414 ( .A(n9153), .ZN(n5538) );
  NAND2_X1 U5415 ( .A1(n8853), .A2(n5685), .ZN(n5553) );
  CLKBUF_X3 U5416 ( .A(n6600), .Z(n7090) );
  AND2_X1 U5417 ( .A1(n9473), .A2(n10791), .ZN(n6600) );
  NAND2_X1 U5418 ( .A1(n8895), .A2(n8920), .ZN(n7593) );
  NOR2_X1 U5419 ( .A1(n10627), .A2(n10628), .ZN(n5345) );
  OR2_X1 U5420 ( .A1(n7652), .A2(n6872), .ZN(n6705) );
  INV_X1 U5421 ( .A(n11020), .ZN(n10725) );
  INV_X1 U5422 ( .A(n6450), .ZN(n5206) );
  AND2_X1 U5423 ( .A1(n5679), .A2(n5565), .ZN(n5564) );
  INV_X1 U5424 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U5425 ( .A1(n5528), .A2(n5529), .ZN(n6079) );
  XNOR2_X1 U5426 ( .A(n5573), .B(n7860), .ZN(n5572) );
  AOI21_X1 U5427 ( .B1(n5122), .B2(n5577), .A(n5164), .ZN(n5574) );
  INV_X1 U5428 ( .A(n6113), .ZN(n6126) );
  NAND2_X1 U5429 ( .A1(n8772), .A2(n8771), .ZN(n8770) );
  AOI21_X1 U5430 ( .B1(n10448), .B2(n10447), .A(n10404), .ZN(n10405) );
  NAND2_X1 U5431 ( .A1(n5429), .A2(n5426), .ZN(n5425) );
  NAND2_X1 U5432 ( .A1(n9327), .A2(n9326), .ZN(n5429) );
  NAND2_X1 U5433 ( .A1(n5418), .A2(n5417), .ZN(n9358) );
  OR2_X1 U5434 ( .A1(n9349), .A2(n9449), .ZN(n5417) );
  NAND2_X1 U5435 ( .A1(n5432), .A2(n5431), .ZN(n5430) );
  NOR2_X1 U5436 ( .A1(n9388), .A2(n9389), .ZN(n5433) );
  NAND2_X1 U5437 ( .A1(n5436), .A2(n5435), .ZN(n5434) );
  NAND2_X1 U5438 ( .A1(n5259), .A2(n7221), .ZN(n5258) );
  NAND2_X1 U5439 ( .A1(n5264), .A2(n5147), .ZN(n5259) );
  NAND2_X1 U5440 ( .A1(n5263), .A2(n7190), .ZN(n5262) );
  NAND2_X1 U5441 ( .A1(n5264), .A2(n7217), .ZN(n5263) );
  NOR2_X1 U5442 ( .A1(n7054), .A2(n7096), .ZN(n5261) );
  NAND2_X1 U5443 ( .A1(n5406), .A2(n9421), .ZN(n5405) );
  AND2_X1 U5444 ( .A1(n9855), .A2(n5404), .ZN(n5403) );
  INV_X1 U5445 ( .A(n9420), .ZN(n5404) );
  INV_X1 U5446 ( .A(n9428), .ZN(n5399) );
  INV_X1 U5447 ( .A(n9845), .ZN(n5401) );
  INV_X1 U5448 ( .A(n10092), .ZN(n5669) );
  INV_X1 U5449 ( .A(n10399), .ZN(n5250) );
  NAND2_X1 U5450 ( .A1(n5170), .A2(n5252), .ZN(n5251) );
  AND2_X1 U5451 ( .A1(n7073), .A2(n7069), .ZN(n5255) );
  INV_X1 U5452 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8311) );
  INV_X1 U5453 ( .A(n5683), .ZN(n9305) );
  AND2_X1 U5454 ( .A1(n10021), .A2(n9568), .ZN(n9389) );
  NAND2_X1 U5455 ( .A1(n5444), .A2(n9377), .ZN(n5443) );
  NAND2_X1 U5456 ( .A1(n5445), .A2(n5133), .ZN(n5444) );
  OR2_X1 U5457 ( .A1(n10647), .A2(n10634), .ZN(n7105) );
  NAND2_X1 U5458 ( .A1(n6247), .A2(n6246), .ZN(n6973) );
  AND2_X1 U5459 ( .A1(n6203), .A2(n5791), .ZN(n5520) );
  OAI21_X1 U5460 ( .B1(n5599), .B2(n5597), .A(n5165), .ZN(n5596) );
  INV_X1 U5461 ( .A(n9142), .ZN(n5597) );
  AOI21_X1 U5462 ( .B1(n5412), .B2(n9455), .A(n9272), .ZN(n5411) );
  NAND2_X1 U5463 ( .A1(n5347), .A2(n5144), .ZN(n10921) );
  NAND2_X1 U5464 ( .A1(n7756), .A2(n5483), .ZN(n7758) );
  OR2_X1 U5465 ( .A1(n7757), .A2(n5925), .ZN(n5483) );
  NAND2_X1 U5466 ( .A1(n7878), .A2(n7879), .ZN(n8946) );
  NAND2_X1 U5467 ( .A1(n9855), .A2(n9419), .ZN(n5632) );
  NAND2_X1 U5468 ( .A1(n5843), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5441) );
  OR2_X1 U5469 ( .A1(n6237), .A2(n7859), .ZN(n5440) );
  NOR2_X1 U5470 ( .A1(n9800), .A2(n5468), .ZN(n5467) );
  INV_X1 U5471 ( .A(n6319), .ZN(n5468) );
  NOR2_X1 U5472 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5638) );
  INV_X1 U5473 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U5474 ( .A1(n6482), .A2(n5672), .ZN(n6490) );
  AND2_X1 U5475 ( .A1(n6481), .A2(n6489), .ZN(n5672) );
  NOR2_X1 U5476 ( .A1(n5658), .A2(n5656), .ZN(n5655) );
  INV_X1 U5477 ( .A(n10188), .ZN(n5656) );
  AND2_X1 U5478 ( .A1(n6858), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6875) );
  INV_X1 U5479 ( .A(n5680), .ZN(n5229) );
  AND2_X1 U5480 ( .A1(n8030), .A2(n6558), .ZN(n6572) );
  OAI21_X1 U5481 ( .B1(n9186), .B2(n5119), .A(n5237), .ZN(n6714) );
  INV_X1 U5482 ( .A(n5238), .ZN(n5237) );
  OAI21_X1 U5483 ( .B1(n5119), .B2(n9187), .A(n5660), .ZN(n5238) );
  AND2_X1 U5484 ( .A1(n5662), .A2(n5661), .ZN(n5660) );
  NAND2_X1 U5485 ( .A1(n7241), .A2(n10383), .ZN(n7180) );
  OR2_X1 U5486 ( .A1(n10618), .A2(n10450), .ZN(n7177) );
  AND2_X1 U5487 ( .A1(n5330), .A2(n5327), .ZN(n5326) );
  NAND2_X1 U5488 ( .A1(n10392), .A2(n7230), .ZN(n5327) );
  NAND2_X1 U5489 ( .A1(n9053), .A2(n10138), .ZN(n7159) );
  NOR2_X1 U5490 ( .A1(n5161), .A2(n5552), .ZN(n5551) );
  NOR2_X1 U5491 ( .A1(n8854), .A2(n9006), .ZN(n5388) );
  AND2_X1 U5492 ( .A1(n7108), .A2(n7151), .ZN(n8123) );
  AND2_X1 U5493 ( .A1(n6947), .A2(n8920), .ZN(n6470) );
  NAND2_X1 U5494 ( .A1(n8716), .A2(n8748), .ZN(n7200) );
  NAND2_X1 U5495 ( .A1(n10560), .A2(n10768), .ZN(n10541) );
  INV_X1 U5496 ( .A(n7620), .ZN(n7618) );
  INV_X1 U5497 ( .A(n8920), .ZN(n7603) );
  INV_X1 U5498 ( .A(n5338), .ZN(n5336) );
  NOR2_X1 U5499 ( .A1(n6217), .A2(n5526), .ZN(n5525) );
  INV_X1 U5500 ( .A(n5788), .ZN(n5526) );
  NAND2_X1 U5501 ( .A1(n6433), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6439) );
  AND2_X1 U5502 ( .A1(n5688), .A2(n6419), .ZN(n5676) );
  NAND2_X1 U5503 ( .A1(n5503), .A2(n5499), .ZN(n6137) );
  INV_X1 U5504 ( .A(n5500), .ZN(n5499) );
  OAI21_X1 U5505 ( .B1(n5505), .B2(n5501), .A(n5767), .ZN(n5500) );
  AOI21_X1 U5506 ( .B1(n5510), .B2(n5508), .A(n5507), .ZN(n5506) );
  INV_X1 U5507 ( .A(n5764), .ZN(n5507) );
  INV_X1 U5508 ( .A(n6098), .ZN(n5508) );
  INV_X1 U5509 ( .A(n5510), .ZN(n5509) );
  NOR2_X1 U5510 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6436) );
  NAND2_X1 U5511 ( .A1(n5753), .A2(SI_15_), .ZN(n5754) );
  INV_X1 U5512 ( .A(SI_14_), .ZN(n8160) );
  INV_X1 U5513 ( .A(SI_13_), .ZN(n8164) );
  INV_X1 U5514 ( .A(n5962), .ZN(n5494) );
  INV_X1 U5515 ( .A(n5730), .ZN(n5498) );
  NAND2_X1 U5516 ( .A1(n5729), .A2(n5730), .ZN(n5245) );
  NAND2_X1 U5517 ( .A1(n5816), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U5518 ( .A1(n9498), .A2(n9862), .ZN(n5583) );
  AOI21_X1 U5519 ( .B1(n9522), .B2(n5593), .A(n9512), .ZN(n5592) );
  INV_X1 U5520 ( .A(n9620), .ZN(n5593) );
  INV_X1 U5521 ( .A(n5592), .ZN(n5590) );
  NAND2_X1 U5522 ( .A1(n6021), .A2(n6020), .ZN(n9367) );
  OR2_X1 U5523 ( .A1(n9210), .A2(n9953), .ZN(n9211) );
  NOR2_X1 U5524 ( .A1(n5609), .A2(n7580), .ZN(n5608) );
  INV_X1 U5525 ( .A(n5613), .ZN(n5609) );
  AND2_X1 U5526 ( .A1(n7540), .A2(n7538), .ZN(n5613) );
  NOR2_X1 U5527 ( .A1(n7553), .A2(n5611), .ZN(n5610) );
  INV_X1 U5528 ( .A(n5612), .ZN(n5611) );
  OR2_X1 U5529 ( .A1(n5618), .A2(n5619), .ZN(n5617) );
  NAND2_X1 U5530 ( .A1(n5581), .A2(n9489), .ZN(n9587) );
  INV_X1 U5531 ( .A(n9589), .ZN(n5581) );
  NAND2_X1 U5532 ( .A1(n9557), .A2(n5568), .ZN(n5567) );
  INV_X1 U5533 ( .A(n9503), .ZN(n5568) );
  AOI21_X1 U5534 ( .B1(n5411), .B2(n5413), .A(n9458), .ZN(n5409) );
  INV_X1 U5535 ( .A(n5411), .ZN(n5410) );
  AND2_X1 U5536 ( .A1(n9307), .A2(n5624), .ZN(n5627) );
  AND2_X1 U5537 ( .A1(n9306), .A2(n5125), .ZN(n9307) );
  AND2_X1 U5538 ( .A1(n9451), .A2(n9323), .ZN(n5626) );
  NAND2_X1 U5539 ( .A1(n9276), .A2(n5629), .ZN(n5628) );
  AND2_X1 U5540 ( .A1(n9275), .A2(n9323), .ZN(n5629) );
  NAND2_X1 U5541 ( .A1(n5844), .A2(n5439), .ZN(n5621) );
  OR2_X1 U5542 ( .A1(n5889), .A2(n7344), .ZN(n5439) );
  OR2_X1 U5543 ( .A1(n6237), .A2(n10898), .ZN(n5840) );
  XNOR2_X1 U5544 ( .A(n7691), .B(n10944), .ZN(n10947) );
  OR2_X1 U5545 ( .A1(n10934), .A2(n5890), .ZN(n5484) );
  INV_X1 U5546 ( .A(n10927), .ZN(n5486) );
  XNOR2_X1 U5547 ( .A(n7758), .B(n7766), .ZN(n7838) );
  NOR2_X1 U5548 ( .A1(n7757), .A2(n7749), .ZN(n7750) );
  XNOR2_X1 U5549 ( .A(n8946), .B(n8927), .ZN(n7880) );
  AOI21_X1 U5550 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7877), .A(n7875), .ZN(
        n8926) );
  OAI21_X1 U5551 ( .B1(n7876), .B2(n5374), .A(n5373), .ZN(n10968) );
  NAND2_X1 U5552 ( .A1(n5377), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U5553 ( .A1(n8929), .A2(n5377), .ZN(n5373) );
  INV_X1 U5554 ( .A(n10969), .ZN(n5377) );
  INV_X1 U5555 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6035) );
  OR2_X1 U5556 ( .A1(n10986), .A2(n5367), .ZN(n5366) );
  OR2_X1 U5557 ( .A1(n8933), .A2(n6005), .ZN(n5367) );
  NAND2_X1 U5558 ( .A1(n8932), .A2(n5365), .ZN(n5364) );
  INV_X1 U5559 ( .A(n8933), .ZN(n5365) );
  INV_X1 U5560 ( .A(n5214), .ZN(n9710) );
  OR2_X1 U5561 ( .A1(n9682), .A2(n5361), .ZN(n5358) );
  OR2_X1 U5562 ( .A1(n9702), .A2(n6071), .ZN(n5361) );
  NAND2_X1 U5563 ( .A1(n9701), .A2(n5360), .ZN(n5359) );
  INV_X1 U5564 ( .A(n9702), .ZN(n5360) );
  NOR2_X1 U5565 ( .A1(n11007), .A2(n11006), .ZN(n11005) );
  OR2_X1 U5566 ( .A1(n9725), .A2(n5195), .ZN(n5348) );
  NAND2_X1 U5567 ( .A1(n9746), .A2(n5350), .ZN(n5349) );
  INV_X1 U5568 ( .A(n11010), .ZN(n5350) );
  INV_X1 U5569 ( .A(n5282), .ZN(n5281) );
  INV_X1 U5570 ( .A(n5137), .ZN(n5280) );
  AND2_X1 U5571 ( .A1(n5470), .A2(n5469), .ZN(n9785) );
  INV_X1 U5572 ( .A(n9796), .ZN(n5276) );
  AND2_X1 U5573 ( .A1(n6193), .A2(n9581), .ZN(n6209) );
  NAND2_X1 U5574 ( .A1(n6209), .A2(n9559), .ZN(n6222) );
  NAND2_X1 U5575 ( .A1(n6202), .A2(n6201), .ZN(n9835) );
  NAND2_X1 U5576 ( .A1(n6215), .A2(n9429), .ZN(n9834) );
  NAND2_X1 U5577 ( .A1(n5460), .A2(n5459), .ZN(n9828) );
  AOI21_X1 U5578 ( .B1(n5123), .B2(n5116), .A(n5155), .ZN(n5459) );
  AND4_X1 U5579 ( .A1(n6227), .A2(n6226), .A3(n6225), .A4(n6224), .ZN(n9831)
         );
  NAND2_X1 U5580 ( .A1(n9885), .A2(n9414), .ZN(n9869) );
  NAND2_X1 U5581 ( .A1(n9869), .A2(n9868), .ZN(n9871) );
  AND2_X1 U5582 ( .A1(n6309), .A2(n9886), .ZN(n6310) );
  AND2_X1 U5583 ( .A1(n6308), .A2(n9412), .ZN(n9900) );
  AND4_X1 U5584 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n9907)
         );
  NAND2_X1 U5585 ( .A1(n5292), .A2(n5291), .ZN(n9119) );
  AOI21_X1 U5586 ( .B1(n5294), .B2(n9376), .A(n9382), .ZN(n5291) );
  NAND2_X1 U5587 ( .A1(n6053), .A2(n6052), .ZN(n9138) );
  NOR2_X1 U5588 ( .A1(n6048), .A2(n9368), .ZN(n5296) );
  NOR2_X1 U5589 ( .A1(n5295), .A2(n9377), .ZN(n5294) );
  NOR2_X1 U5590 ( .A1(n5296), .A2(n9376), .ZN(n5295) );
  OR2_X1 U5591 ( .A1(n8983), .A2(n9376), .ZN(n5290) );
  AND4_X1 U5592 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n9197)
         );
  NAND2_X1 U5593 ( .A1(n5454), .A2(n5453), .ZN(n8792) );
  AOI21_X1 U5594 ( .B1(n5121), .B2(n5458), .A(n5154), .ZN(n5453) );
  INV_X1 U5595 ( .A(n5306), .ZN(n5305) );
  OAI21_X1 U5596 ( .B1(n5140), .B2(n5117), .A(n5997), .ZN(n5306) );
  NAND2_X1 U5597 ( .A1(n5961), .A2(n9354), .ZN(n5635) );
  AND2_X1 U5598 ( .A1(n9348), .A2(n9345), .ZN(n5637) );
  NAND2_X1 U5599 ( .A1(n5285), .A2(n5284), .ZN(n8009) );
  AOI21_X1 U5600 ( .B1(n5286), .B2(n5289), .A(n5167), .ZN(n5284) );
  NAND2_X1 U5601 ( .A1(n7785), .A2(n5286), .ZN(n5285) );
  AOI21_X1 U5602 ( .B1(n9281), .B2(n5288), .A(n5287), .ZN(n5286) );
  OR2_X1 U5603 ( .A1(n9651), .A2(n7747), .ZN(n7436) );
  INV_X1 U5604 ( .A(n9956), .ZN(n9936) );
  AOI21_X1 U5605 ( .B1(n9775), .B2(n8840), .A(n5310), .ZN(n5473) );
  INV_X1 U5606 ( .A(n6336), .ZN(n5310) );
  NAND2_X1 U5607 ( .A1(n6208), .A2(n6207), .ZN(n9554) );
  OR2_X1 U5608 ( .A1(n9242), .A2(n5851), .ZN(n6208) );
  NAND2_X1 U5609 ( .A1(n6369), .A2(n6368), .ZN(n7405) );
  XNOR2_X1 U5610 ( .A(n6372), .B(n6371), .ZN(n7404) );
  INV_X1 U5611 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6371) );
  AND2_X1 U5612 ( .A1(n5471), .A2(n5811), .ZN(n5298) );
  NAND2_X1 U5613 ( .A1(n6256), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6265) );
  OR2_X1 U5614 ( .A1(n6700), .A2(n6699), .ZN(n5668) );
  AND2_X1 U5615 ( .A1(n5665), .A2(n6699), .ZN(n5664) );
  OR2_X1 U5616 ( .A1(n6680), .A2(n6700), .ZN(n5665) );
  XNOR2_X1 U5617 ( .A(n6513), .B(n6489), .ZN(n6514) );
  OAI22_X1 U5618 ( .A1(n5112), .A2(n8103), .B1(n7011), .B2(n7262), .ZN(n6513)
         );
  AND2_X1 U5619 ( .A1(n6919), .A2(n6918), .ZN(n7268) );
  NAND2_X1 U5620 ( .A1(n5392), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U5621 ( .A1(n10165), .A2(n10166), .ZN(n5673) );
  AOI21_X1 U5622 ( .B1(n5136), .B2(n5641), .A(n5235), .ZN(n5234) );
  INV_X1 U5623 ( .A(n10110), .ZN(n5235) );
  AND2_X1 U5624 ( .A1(n10174), .A2(n10175), .ZN(n6680) );
  OR2_X1 U5625 ( .A1(n6667), .A2(n6666), .ZN(n6690) );
  AOI21_X1 U5626 ( .B1(n5227), .B2(n5229), .A(n5225), .ZN(n5224) );
  INV_X1 U5627 ( .A(n9090), .ZN(n5225) );
  AND2_X1 U5628 ( .A1(n5230), .A2(n5680), .ZN(n5226) );
  AND2_X1 U5629 ( .A1(n5651), .A2(n5650), .ZN(n5649) );
  NOR2_X1 U5630 ( .A1(n6770), .A2(n6766), .ZN(n5651) );
  OR2_X1 U5631 ( .A1(n5652), .A2(n10134), .ZN(n5650) );
  NOR2_X1 U5632 ( .A1(n5132), .A2(n5648), .ZN(n5647) );
  INV_X1 U5633 ( .A(n10134), .ZN(n5648) );
  NOR2_X1 U5634 ( .A1(n5132), .A2(n6769), .ZN(n5646) );
  NAND2_X1 U5635 ( .A1(n6718), .A2(n10230), .ZN(n10133) );
  NAND2_X1 U5636 ( .A1(n10125), .A2(n10126), .ZN(n10218) );
  AND2_X1 U5637 ( .A1(n6943), .A2(n10784), .ZN(n6951) );
  AND2_X1 U5638 ( .A1(n5271), .A2(n5172), .ZN(n5270) );
  NAND2_X1 U5639 ( .A1(n7243), .A2(n5274), .ZN(n5271) );
  NAND2_X1 U5640 ( .A1(n7099), .A2(n7245), .ZN(n5274) );
  NOR2_X1 U5641 ( .A1(n10447), .A2(n5561), .ZN(n5560) );
  INV_X1 U5642 ( .A(n10426), .ZN(n5561) );
  AND2_X1 U5643 ( .A1(n7172), .A2(n10403), .ZN(n10447) );
  AND2_X1 U5644 ( .A1(n6994), .A2(n6909), .ZN(n10465) );
  NAND2_X1 U5645 ( .A1(n10495), .A2(n10758), .ZN(n10484) );
  AND2_X1 U5646 ( .A1(n10514), .A2(n10397), .ZN(n10491) );
  NAND2_X1 U5647 ( .A1(n10532), .A2(n5152), .ZN(n10520) );
  INV_X1 U5648 ( .A(n10394), .ZN(n10535) );
  AND4_X1 U5649 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n9219)
         );
  AND2_X1 U5650 ( .A1(n9047), .A2(n7159), .ZN(n9081) );
  OR2_X1 U5651 ( .A1(n10729), .A2(n10179), .ZN(n9045) );
  NAND3_X1 U5652 ( .A1(n9046), .A2(n9073), .A3(n9045), .ZN(n9047) );
  NAND2_X1 U5653 ( .A1(n7152), .A2(n5333), .ZN(n8722) );
  INV_X1 U5654 ( .A(n5334), .ZN(n5333) );
  AOI21_X1 U5655 ( .B1(n5542), .B2(n5544), .A(n5157), .ZN(n5540) );
  INV_X1 U5656 ( .A(n8123), .ZN(n8125) );
  NAND2_X1 U5657 ( .A1(n8124), .A2(n8125), .ZN(n8679) );
  NAND2_X1 U5658 ( .A1(n8714), .A2(n7197), .ZN(n7927) );
  NAND2_X1 U5659 ( .A1(n7631), .A2(n7590), .ZN(n7592) );
  NAND2_X1 U5660 ( .A1(n7815), .A2(n5383), .ZN(n7635) );
  NOR2_X1 U5661 ( .A1(n10198), .A2(n7657), .ZN(n5383) );
  NAND2_X1 U5662 ( .A1(n10803), .A2(n6962), .ZN(n10435) );
  OR2_X1 U5663 ( .A1(n6948), .A2(n8043), .ZN(n11088) );
  INV_X1 U5664 ( .A(n10667), .ZN(n10731) );
  INV_X1 U5665 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8323) );
  INV_X1 U5666 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U5667 ( .A1(n6165), .A2(n5778), .ZN(n6177) );
  XNOR2_X1 U5668 ( .A(n6945), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7328) );
  OR2_X1 U5669 ( .A1(n6163), .A2(n8349), .ZN(n6165) );
  INV_X1 U5670 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6441) );
  NOR2_X1 U5671 ( .A1(n5760), .A2(n6110), .ZN(n5510) );
  AND2_X1 U5672 ( .A1(n5532), .A2(n5752), .ZN(n5531) );
  INV_X1 U5673 ( .A(n6063), .ZN(n5532) );
  AND3_X1 U5674 ( .A1(n5674), .A2(n5312), .A3(n8495), .ZN(n5239) );
  AND2_X1 U5675 ( .A1(n5517), .A2(n5743), .ZN(n5516) );
  INV_X1 U5676 ( .A(n6014), .ZN(n5517) );
  INV_X1 U5677 ( .A(n5998), .ZN(n5202) );
  NAND2_X1 U5678 ( .A1(n5933), .A2(n5730), .ZN(n5947) );
  NAND2_X1 U5679 ( .A1(n5918), .A2(n5726), .ZN(n5931) );
  INV_X1 U5680 ( .A(n5245), .ZN(n5930) );
  NAND2_X1 U5681 ( .A1(n6129), .A2(n6128), .ZN(n9910) );
  AND4_X1 U5682 ( .A1(n6047), .A2(n6046), .A3(n6045), .A4(n6044), .ZN(n9139)
         );
  INV_X1 U5683 ( .A(n9613), .ZN(n9624) );
  AND2_X1 U5684 ( .A1(n5914), .A2(n5913), .ZN(n7826) );
  OR2_X1 U5685 ( .A1(n7551), .A2(n7789), .ZN(n5612) );
  NAND2_X1 U5686 ( .A1(n7539), .A2(n5613), .ZN(n7550) );
  NAND2_X1 U5687 ( .A1(n6040), .A2(n6039), .ZN(n9022) );
  XNOR2_X1 U5688 ( .A(n9513), .B(n7860), .ZN(n5571) );
  OR2_X1 U5689 ( .A1(n9481), .A2(n9955), .ZN(n5682) );
  AND2_X1 U5690 ( .A1(n7426), .A2(n7733), .ZN(n9629) );
  XNOR2_X1 U5691 ( .A(n6264), .B(P2_IR_REG_22__SCAN_IN), .ZN(n9465) );
  OR2_X1 U5692 ( .A1(n7836), .A2(n7764), .ZN(n5356) );
  OR2_X1 U5693 ( .A1(n7876), .A2(n5973), .ZN(n5376) );
  XNOR2_X1 U5694 ( .A(n8926), .B(n8927), .ZN(n7876) );
  NAND2_X1 U5695 ( .A1(n5461), .A2(n6315), .ZN(n9839) );
  OR2_X1 U5696 ( .A1(n9849), .A2(n5116), .ZN(n5461) );
  NAND2_X1 U5697 ( .A1(n6116), .A2(n6115), .ZN(n10009) );
  OR2_X1 U5698 ( .A1(n8054), .A2(n5851), .ZN(n6116) );
  AND2_X1 U5699 ( .A1(n6070), .A2(n6069), .ZN(n10028) );
  AND2_X1 U5700 ( .A1(n5898), .A2(n5897), .ZN(n7852) );
  NAND2_X1 U5701 ( .A1(n7732), .A2(n7731), .ZN(n7742) );
  INV_X1 U5702 ( .A(n5463), .ZN(n5462) );
  AND2_X1 U5703 ( .A1(n5473), .A2(n5309), .ZN(n5472) );
  NAND2_X1 U5704 ( .A1(n9775), .A2(n7833), .ZN(n5309) );
  AND2_X1 U5705 ( .A1(n7404), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7305) );
  AND2_X1 U5706 ( .A1(n6929), .A2(n10797), .ZN(n6431) );
  INV_X1 U5707 ( .A(n7328), .ZN(n7325) );
  NAND2_X1 U5708 ( .A1(n6776), .A2(n6775), .ZN(n10593) );
  INV_X1 U5709 ( .A(n7267), .ZN(n7277) );
  AND2_X1 U5710 ( .A1(n7269), .A2(n10223), .ZN(n7276) );
  AND2_X1 U5711 ( .A1(n6721), .A2(n6720), .ZN(n10714) );
  OR2_X1 U5712 ( .A1(n6872), .A2(n7300), .ZN(n6568) );
  NAND2_X1 U5713 ( .A1(n6737), .A2(n6736), .ZN(n10706) );
  NAND2_X1 U5714 ( .A1(n6857), .A2(n6856), .ZN(n10654) );
  NAND2_X1 U5715 ( .A1(n6608), .A2(n6609), .ZN(n5670) );
  AND4_X1 U5716 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n9063)
         );
  AND2_X1 U5717 ( .A1(n6908), .A2(n6892), .ZN(n10481) );
  OR2_X1 U5718 ( .A1(n7188), .A2(n5684), .ZN(n7251) );
  INV_X1 U5719 ( .A(n10643), .ZN(n10464) );
  INV_X1 U5720 ( .A(n9063), .ZN(n10246) );
  NAND2_X1 U5721 ( .A1(n6543), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U5722 ( .A1(n6635), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U5723 ( .A1(n6757), .A2(n6756), .ZN(n10406) );
  NAND2_X1 U5724 ( .A1(n5343), .A2(n5346), .ZN(n10750) );
  NAND2_X1 U5725 ( .A1(n10629), .A2(n10725), .ZN(n5346) );
  NAND2_X1 U5726 ( .A1(n10752), .A2(n10631), .ZN(n5342) );
  NOR2_X1 U5727 ( .A1(n10616), .A2(n5197), .ZN(n5196) );
  NAND2_X1 U5728 ( .A1(n10750), .A2(n11079), .ZN(n5201) );
  INV_X1 U5729 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5200) );
  AND2_X1 U5730 ( .A1(n6417), .A2(n6416), .ZN(n9092) );
  NOR2_X1 U5731 ( .A1(n5338), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5337) );
  INV_X1 U5732 ( .A(n9357), .ZN(n5416) );
  OR2_X1 U5733 ( .A1(n9343), .A2(n5422), .ZN(n5421) );
  OR2_X1 U5734 ( .A1(n9344), .A2(n9449), .ZN(n5423) );
  NOR2_X1 U5735 ( .A1(n9352), .A2(n5420), .ZN(n5419) );
  NAND2_X1 U5736 ( .A1(n9348), .A2(n9347), .ZN(n5420) );
  OR2_X1 U5737 ( .A1(n9379), .A2(n5162), .ZN(n5436) );
  NOR2_X1 U5738 ( .A1(n9383), .A2(n9384), .ZN(n5435) );
  NAND2_X1 U5739 ( .A1(n9391), .A2(n5422), .ZN(n5431) );
  NAND2_X1 U5740 ( .A1(n5266), .A2(n5265), .ZN(n5264) );
  NAND2_X1 U5741 ( .A1(n7052), .A2(n7096), .ZN(n5265) );
  NAND2_X1 U5742 ( .A1(n7053), .A2(n7095), .ZN(n5266) );
  NAND2_X1 U5743 ( .A1(n5260), .A2(n5257), .ZN(n7055) );
  NAND2_X1 U5744 ( .A1(n5262), .A2(n5261), .ZN(n5260) );
  NAND2_X1 U5745 ( .A1(n5258), .A2(n7096), .ZN(n5257) );
  INV_X1 U5746 ( .A(SI_19_), .ZN(n8155) );
  NOR2_X1 U5747 ( .A1(n9425), .A2(n5401), .ZN(n5400) );
  NAND2_X1 U5748 ( .A1(n6216), .A2(n5399), .ZN(n5398) );
  NAND2_X1 U5749 ( .A1(n5405), .A2(n5403), .ZN(n5402) );
  AOI21_X1 U5750 ( .B1(n8618), .B2(n5457), .A(n5160), .ZN(n5456) );
  INV_X1 U5751 ( .A(n6284), .ZN(n5457) );
  NOR2_X2 U5752 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5964) );
  INV_X1 U5753 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U5754 ( .A1(n5666), .A2(n5668), .ZN(n5661) );
  NAND2_X1 U5755 ( .A1(n5664), .A2(n6700), .ZN(n5662) );
  INV_X1 U5756 ( .A(n5664), .ZN(n5663) );
  OAI21_X1 U5757 ( .B1(n5254), .B2(n5253), .A(n5249), .ZN(n7074) );
  INV_X1 U5758 ( .A(n7068), .ZN(n5254) );
  AOI21_X1 U5759 ( .B1(n5151), .B2(n5251), .A(n5250), .ZN(n5249) );
  AOI21_X1 U5760 ( .B1(n7068), .B2(n5255), .A(n5251), .ZN(n7076) );
  INV_X1 U5761 ( .A(n8855), .ZN(n5552) );
  INV_X1 U5762 ( .A(n5523), .ZN(n5522) );
  OAI21_X1 U5763 ( .B1(n5525), .B2(n5524), .A(n6231), .ZN(n5523) );
  INV_X1 U5764 ( .A(n5506), .ZN(n5505) );
  NAND2_X1 U5765 ( .A1(n5509), .A2(n5502), .ZN(n5501) );
  INV_X1 U5766 ( .A(n6124), .ZN(n5502) );
  NOR2_X1 U5767 ( .A1(n5505), .A2(n6124), .ZN(n5504) );
  INV_X1 U5768 ( .A(SI_20_), .ZN(n8354) );
  INV_X1 U5769 ( .A(SI_17_), .ZN(n8165) );
  INV_X1 U5770 ( .A(n6078), .ZN(n5527) );
  OAI21_X1 U5771 ( .B1(n7287), .B2(n5247), .A(n5246), .ZN(n5731) );
  NAND2_X1 U5772 ( .A1(n7287), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n5246) );
  AND2_X1 U5773 ( .A1(n5130), .A2(n9323), .ZN(n5625) );
  AND2_X1 U5774 ( .A1(n9274), .A2(n9273), .ZN(n9275) );
  NOR2_X1 U5775 ( .A1(n9455), .A2(n9272), .ZN(n9273) );
  NAND2_X1 U5776 ( .A1(n10900), .A2(n10901), .ZN(n10899) );
  AOI21_X1 U5777 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n10912), .A(n10907), .ZN(
        n7456) );
  OR2_X1 U5778 ( .A1(n7458), .A2(n7446), .ZN(n5347) );
  INV_X1 U5779 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5965) );
  INV_X1 U5780 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8401) );
  AOI21_X1 U5781 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n8945), .A(n10968), .ZN(
        n8931) );
  NAND2_X1 U5782 ( .A1(n5477), .A2(n5476), .ZN(n5214) );
  NAND2_X1 U5783 ( .A1(n9689), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5476) );
  AND2_X1 U5784 ( .A1(n5475), .A2(n5474), .ZN(n9763) );
  NAND2_X1 U5785 ( .A1(n9736), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5474) );
  INV_X1 U5786 ( .A(n9389), .ZN(n9396) );
  AOI21_X1 U5787 ( .B1(n8977), .B2(n5445), .A(n5443), .ZN(n5442) );
  INV_X1 U5788 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8419) );
  AND2_X1 U5789 ( .A1(n5939), .A2(n8401), .ZN(n5954) );
  INV_X1 U5790 ( .A(n9337), .ZN(n5288) );
  INV_X1 U5791 ( .A(n9338), .ZN(n5287) );
  NAND2_X1 U5792 ( .A1(n5455), .A2(n5456), .ZN(n8839) );
  OR2_X1 U5793 ( .A1(n6285), .A2(n5458), .ZN(n5455) );
  INV_X1 U5794 ( .A(P2_B_REG_SCAN_IN), .ZN(n8430) );
  AND2_X1 U5795 ( .A1(n6840), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6858) );
  AND2_X1 U5796 ( .A1(n6825), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6840) );
  AND2_X1 U5797 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n6794), .ZN(n6809) );
  AND2_X1 U5798 ( .A1(n6809), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6825) );
  NOR2_X1 U5799 ( .A1(n10245), .A2(n5490), .ZN(n5489) );
  INV_X1 U5800 ( .A(n7089), .ZN(n5490) );
  AND2_X1 U5801 ( .A1(n6889), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6906) );
  AOI21_X1 U5802 ( .B1(n7221), .B2(n5320), .A(n9159), .ZN(n5319) );
  AND2_X1 U5803 ( .A1(n7221), .A2(n7190), .ZN(n9078) );
  INV_X1 U5804 ( .A(n8863), .ZN(n5332) );
  OR2_X1 U5805 ( .A1(n7154), .A2(n5335), .ZN(n5334) );
  INV_X1 U5806 ( .A(n7151), .ZN(n5335) );
  OR2_X1 U5807 ( .A1(n8854), .A2(n9063), .ZN(n7107) );
  INV_X1 U5808 ( .A(n5543), .ZN(n5542) );
  OAI21_X1 U5809 ( .B1(n8125), .B2(n5544), .A(n8725), .ZN(n5543) );
  AND2_X1 U5810 ( .A1(n7149), .A2(n7148), .ZN(n7208) );
  OR2_X1 U5811 ( .A1(n7147), .A2(n7146), .ZN(n7148) );
  AND2_X1 U5812 ( .A1(n7143), .A2(n7110), .ZN(n7203) );
  INV_X1 U5813 ( .A(n7920), .ZN(n5557) );
  NAND2_X1 U5814 ( .A1(n6977), .A2(n6976), .ZN(n7088) );
  XNOR2_X1 U5815 ( .A(n6973), .B(n6974), .ZN(n6972) );
  INV_X1 U5816 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U5817 ( .A1(n6401), .A2(n6402), .ZN(n5314) );
  INV_X1 U5818 ( .A(SI_21_), .ZN(n8347) );
  INV_X1 U5819 ( .A(SI_18_), .ZN(n8159) );
  AOI21_X1 U5820 ( .B1(n5531), .B2(n6049), .A(n5530), .ZN(n5529) );
  INV_X1 U5821 ( .A(n5754), .ZN(n5530) );
  INV_X1 U5822 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8480) );
  OAI21_X1 U5823 ( .B1(n7287), .B2(n5709), .A(n5708), .ZN(n5711) );
  INV_X1 U5824 ( .A(n5816), .ZN(n5703) );
  NAND2_X1 U5825 ( .A1(n8965), .A2(n8964), .ZN(n5603) );
  OR2_X1 U5826 ( .A1(n9200), .A2(n5577), .ZN(n5576) );
  INV_X1 U5827 ( .A(n9211), .ZN(n5577) );
  AOI21_X1 U5828 ( .B1(n5601), .B2(n5600), .A(n5148), .ZN(n5599) );
  INV_X1 U5829 ( .A(n8964), .ZN(n5600) );
  NOR2_X1 U5830 ( .A1(n6006), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6022) );
  OR2_X1 U5831 ( .A1(n9564), .A2(n9918), .ZN(n9480) );
  NAND2_X1 U5832 ( .A1(n6258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U5833 ( .A1(n6113), .A2(n5604), .ZN(n6258) );
  OR2_X1 U5834 ( .A1(n6237), .A2(n10902), .ZN(n5860) );
  AND2_X1 U5835 ( .A1(n10906), .A2(n10905), .ZN(n10907) );
  INV_X1 U5836 ( .A(n5881), .ZN(n5969) );
  AND2_X1 U5837 ( .A1(n10925), .A2(n7690), .ZN(n7691) );
  NAND2_X1 U5838 ( .A1(n7837), .A2(n7759), .ZN(n7760) );
  AND3_X1 U5839 ( .A1(n5366), .A2(n5364), .A3(n5188), .ZN(n9652) );
  XNOR2_X1 U5840 ( .A(n5214), .B(n5213), .ZN(n9690) );
  NOR2_X1 U5841 ( .A1(n9681), .A2(n9680), .ZN(n9699) );
  XNOR2_X1 U5842 ( .A(n9763), .B(n9764), .ZN(n9737) );
  NOR2_X1 U5843 ( .A1(n9940), .A2(n9737), .ZN(n9765) );
  AND3_X1 U5844 ( .A1(n5359), .A2(n5358), .A3(n5192), .ZN(n9744) );
  AND4_X1 U5845 ( .A1(n5836), .A2(n5835), .A3(n5834), .A4(n5833), .ZN(n9805)
         );
  AND4_X1 U5846 ( .A1(n6241), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n9819)
         );
  OAI21_X1 U5847 ( .B1(n9885), .B2(n5139), .A(n5300), .ZN(n9846) );
  NOR2_X1 U5848 ( .A1(n5139), .A2(n9414), .ZN(n5301) );
  OR2_X1 U5849 ( .A1(n6168), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6182) );
  AOI21_X1 U5850 ( .B1(n6148), .B2(n9407), .A(n9409), .ZN(n5634) );
  INV_X1 U5851 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U5852 ( .A1(n6156), .A2(n9547), .ZN(n6168) );
  AND2_X1 U5853 ( .A1(n9414), .A2(n9413), .ZN(n9886) );
  AND2_X1 U5854 ( .A1(n6130), .A2(n9537), .ZN(n6142) );
  INV_X1 U5855 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U5856 ( .A1(n5450), .A2(n5118), .ZN(n5449) );
  AOI21_X1 U5857 ( .B1(n5450), .B2(n5126), .A(n5156), .ZN(n5448) );
  INV_X1 U5858 ( .A(n6104), .ZN(n6118) );
  NAND2_X1 U5859 ( .A1(n9942), .A2(n5432), .ZN(n5636) );
  NOR2_X1 U5860 ( .A1(n6105), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U5861 ( .A1(n9213), .A2(n6089), .ZN(n6105) );
  INV_X1 U5862 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9147) );
  NOR2_X1 U5863 ( .A1(n6042), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6056) );
  AND4_X1 U5864 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n8975)
         );
  NAND2_X1 U5865 ( .A1(n8615), .A2(n5981), .ZN(n8837) );
  OR2_X1 U5866 ( .A1(n5991), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U5867 ( .A1(n11065), .A2(n8620), .ZN(n9312) );
  NAND2_X1 U5868 ( .A1(n5635), .A2(n5140), .ZN(n8615) );
  OR2_X1 U5869 ( .A1(n5923), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U5870 ( .A1(n7785), .A2(n9337), .ZN(n7824) );
  NAND2_X1 U5871 ( .A1(n7824), .A2(n9281), .ZN(n8007) );
  INV_X1 U5872 ( .A(n9649), .ZN(n8013) );
  AND2_X1 U5873 ( .A1(n9337), .A2(n9333), .ZN(n9331) );
  AND2_X1 U5874 ( .A1(n5424), .A2(n9336), .ZN(n9279) );
  INV_X1 U5875 ( .A(n7436), .ZN(n9324) );
  NAND2_X1 U5876 ( .A1(n9324), .A2(n9280), .ZN(n7566) );
  AND2_X1 U5877 ( .A1(n9449), .A2(n6383), .ZN(n6385) );
  AND2_X1 U5878 ( .A1(n6382), .A2(n6381), .ZN(n7731) );
  OAI22_X1 U5879 ( .A1(n6322), .A2(n5469), .B1(n9441), .B2(n9805), .ZN(n5463)
         );
  AND2_X1 U5880 ( .A1(n5467), .A2(n5466), .ZN(n5465) );
  INV_X1 U5881 ( .A(n6322), .ZN(n5466) );
  NAND2_X1 U5882 ( .A1(n6192), .A2(n6191), .ZN(n9574) );
  INV_X1 U5883 ( .A(n10025), .ZN(n10017) );
  INV_X1 U5884 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6066) );
  INV_X1 U5885 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6689) );
  NOR2_X1 U5886 ( .A1(n6836), .A2(n5654), .ZN(n10102) );
  INV_X1 U5887 ( .A(n10185), .ZN(n6836) );
  AND2_X1 U5888 ( .A1(n10186), .A2(n10188), .ZN(n5654) );
  OR2_X1 U5889 ( .A1(n8827), .A2(n5229), .ZN(n5223) );
  OAI21_X1 U5890 ( .B1(n8608), .B2(n5686), .A(n6591), .ZN(n6592) );
  INV_X1 U5891 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6653) );
  NOR2_X1 U5892 ( .A1(n10185), .A2(n5658), .ZN(n5217) );
  INV_X1 U5893 ( .A(n5653), .ZN(n5218) );
  INV_X1 U5894 ( .A(n8032), .ZN(n6555) );
  NAND2_X1 U5895 ( .A1(n8590), .A2(n8591), .ZN(n5675) );
  OR2_X1 U5896 ( .A1(n6599), .A2(n6464), .ZN(n6614) );
  INV_X1 U5897 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6613) );
  NOR2_X1 U5898 ( .A1(n6614), .A2(n6613), .ZN(n6616) );
  AND2_X1 U5899 ( .A1(n6481), .A2(n6484), .ZN(n5671) );
  AND2_X1 U5900 ( .A1(n6616), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6633) );
  AND2_X1 U5901 ( .A1(n6758), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6777) );
  NOR2_X1 U5902 ( .A1(n6572), .A2(n6571), .ZN(n8628) );
  INV_X1 U5903 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6573) );
  OR2_X1 U5904 ( .A1(n6963), .A2(n7254), .ZN(n6961) );
  NAND2_X1 U5905 ( .A1(n7243), .A2(n5273), .ZN(n5272) );
  INV_X1 U5906 ( .A(n7101), .ZN(n5273) );
  OR2_X1 U5907 ( .A1(n7130), .A2(n5268), .ZN(n5267) );
  NOR2_X1 U5908 ( .A1(n5270), .A2(n8824), .ZN(n5268) );
  NOR3_X1 U5909 ( .A1(n7100), .A2(n8824), .A3(n5272), .ZN(n5269) );
  AND4_X1 U5910 ( .A1(n6620), .A2(n6619), .A3(n6618), .A4(n6617), .ZN(n8121)
         );
  OR2_X1 U5911 ( .A1(n6581), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6593) );
  NOR2_X1 U5912 ( .A1(n10618), .A2(n10454), .ZN(n10431) );
  NAND2_X1 U5913 ( .A1(n5114), .A2(n5396), .ZN(n10454) );
  NAND2_X1 U5914 ( .A1(n10400), .A2(n7170), .ZN(n10476) );
  NOR2_X1 U5915 ( .A1(n10493), .A2(n5546), .ZN(n5550) );
  INV_X1 U5916 ( .A(n10419), .ZN(n5546) );
  INV_X1 U5917 ( .A(n10512), .ZN(n5215) );
  INV_X1 U5918 ( .A(n10393), .ZN(n5324) );
  INV_X1 U5919 ( .A(n5326), .ZN(n5325) );
  NAND2_X1 U5920 ( .A1(n5329), .A2(n5328), .ZN(n10391) );
  INV_X1 U5921 ( .A(n7230), .ZN(n5328) );
  NAND2_X1 U5922 ( .A1(n5545), .A2(n10414), .ZN(n10532) );
  OAI21_X1 U5923 ( .B1(n9223), .B2(n9222), .A(n7162), .ZN(n10584) );
  NAND2_X1 U5924 ( .A1(n5317), .A2(n5315), .ZN(n9223) );
  AOI21_X1 U5925 ( .B1(n5319), .B2(n7054), .A(n5316), .ZN(n5315) );
  NAND2_X1 U5926 ( .A1(n9081), .A2(n5319), .ZN(n5317) );
  INV_X1 U5927 ( .A(n7161), .ZN(n5316) );
  AOI21_X1 U5928 ( .B1(n5537), .B2(n7160), .A(n5535), .ZN(n5534) );
  INV_X1 U5929 ( .A(n9222), .ZN(n5535) );
  OR2_X1 U5930 ( .A1(n9018), .A2(n9017), .ZN(n9046) );
  NAND2_X1 U5931 ( .A1(n8729), .A2(n5388), .ZN(n9012) );
  NAND2_X1 U5932 ( .A1(n8729), .A2(n11089), .ZN(n8857) );
  NAND2_X1 U5933 ( .A1(n5395), .A2(n5394), .ZN(n8680) );
  NOR2_X1 U5934 ( .A1(n8646), .A2(n8673), .ZN(n5394) );
  INV_X1 U5935 ( .A(n8667), .ZN(n5395) );
  AND2_X1 U5936 ( .A1(n8660), .A2(n7111), .ZN(n8560) );
  NAND2_X1 U5937 ( .A1(n8555), .A2(n8781), .ZN(n8667) );
  AND2_X1 U5938 ( .A1(n7985), .A2(n8110), .ZN(n8555) );
  AND2_X1 U5939 ( .A1(n7146), .A2(n7980), .ZN(n7951) );
  OAI21_X1 U5940 ( .B1(n7927), .B2(n7141), .A(n7202), .ZN(n7982) );
  NOR2_X1 U5941 ( .A1(n7953), .A2(n8651), .ZN(n7985) );
  OR2_X1 U5942 ( .A1(n8708), .A2(n11046), .ZN(n7953) );
  NAND2_X1 U5943 ( .A1(n7140), .A2(n7200), .ZN(n8714) );
  INV_X1 U5944 ( .A(n7922), .ZN(n8713) );
  NAND2_X1 U5945 ( .A1(n7921), .A2(n7920), .ZN(n8707) );
  NOR2_X1 U5946 ( .A1(n8748), .A2(n7635), .ZN(n8709) );
  INV_X1 U5947 ( .A(n7591), .ZN(n7601) );
  NAND2_X1 U5948 ( .A1(n7815), .A2(n8042), .ZN(n7634) );
  OR2_X1 U5949 ( .A1(n8043), .A2(n7603), .ZN(n10591) );
  NAND2_X1 U5950 ( .A1(n6946), .A2(n8824), .ZN(n8043) );
  INV_X1 U5951 ( .A(n5382), .ZN(n5197) );
  AOI21_X1 U5952 ( .B1(n10618), .B2(n10707), .A(n10617), .ZN(n5382) );
  AND4_X1 U5953 ( .A1(n6882), .A2(n6881), .A3(n6880), .A4(n6879), .ZN(n10634)
         );
  OR2_X1 U5954 ( .A1(n9242), .A2(n6872), .ZN(n6874) );
  AND4_X1 U5955 ( .A1(n6816), .A2(n6815), .A3(n6814), .A4(n6813), .ZN(n10669)
         );
  NAND2_X1 U5956 ( .A1(n6808), .A2(n6807), .ZN(n10561) );
  OR2_X1 U5957 ( .A1(n8823), .A2(n6872), .ZN(n6808) );
  NAND2_X1 U5958 ( .A1(n6665), .A2(n6664), .ZN(n9006) );
  NAND2_X1 U5959 ( .A1(n7337), .A2(n5115), .ZN(n5248) );
  NAND2_X1 U5960 ( .A1(n7599), .A2(n10271), .ZN(n10667) );
  AND2_X1 U5961 ( .A1(n8040), .A2(n7613), .ZN(n7793) );
  AND2_X1 U5962 ( .A1(n7605), .A2(n7604), .ZN(n11020) );
  INV_X1 U5963 ( .A(n11091), .ZN(n11021) );
  NAND2_X1 U5964 ( .A1(n8316), .A2(n5339), .ZN(n5338) );
  INV_X1 U5965 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5339) );
  XNOR2_X1 U5966 ( .A(n6243), .B(n6242), .ZN(n9471) );
  NAND2_X1 U5967 ( .A1(n5521), .A2(n5791), .ZN(n6230) );
  NAND2_X1 U5968 ( .A1(n6205), .A2(n5525), .ZN(n5521) );
  AND2_X1 U5969 ( .A1(n5788), .A2(n5787), .ZN(n6203) );
  INV_X1 U5970 ( .A(SI_22_), .ZN(n8349) );
  NAND2_X1 U5971 ( .A1(n6440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6442) );
  OAI21_X1 U5972 ( .B1(n6099), .B2(n5509), .A(n5506), .ZN(n6125) );
  NAND2_X1 U5973 ( .A1(n6735), .A2(n6436), .ZN(n6753) );
  OR2_X1 U5974 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6752) );
  AOI21_X1 U5975 ( .B1(n5516), .B2(n5998), .A(n5514), .ZN(n5513) );
  INV_X1 U5976 ( .A(n5745), .ZN(n5514) );
  AND2_X1 U5977 ( .A1(n5749), .A2(n5748), .ZN(n6030) );
  AND2_X1 U5978 ( .A1(n6549), .A2(n5674), .ZN(n5539) );
  OAI21_X1 U5979 ( .B1(n5495), .B2(n5494), .A(n5166), .ZN(n5493) );
  OAI21_X1 U5980 ( .B1(n5931), .B2(n5496), .A(n5495), .ZN(n5963) );
  AND2_X1 U5981 ( .A1(n5726), .A2(n5725), .ZN(n5915) );
  INV_X1 U5982 ( .A(n5697), .ZN(n5696) );
  NOR2_X1 U5983 ( .A1(n7965), .A2(n5619), .ZN(n7967) );
  INV_X1 U5984 ( .A(n5583), .ZN(n5582) );
  NAND2_X1 U5985 ( .A1(n9575), .A2(n9498), .ZN(n9529) );
  NOR2_X1 U5986 ( .A1(n9514), .A2(n5590), .ZN(n5585) );
  NAND2_X1 U5987 ( .A1(n5588), .A2(n5587), .ZN(n5586) );
  OAI21_X1 U5988 ( .B1(n9514), .B2(n9522), .A(n5592), .ZN(n5587) );
  NAND2_X1 U5989 ( .A1(n5590), .A2(n5589), .ZN(n5588) );
  INV_X1 U5990 ( .A(n9514), .ZN(n5589) );
  NAND2_X1 U5991 ( .A1(n9514), .A2(n9522), .ZN(n5591) );
  NAND2_X1 U5992 ( .A1(n8018), .A2(n8017), .ZN(n8084) );
  NAND2_X1 U5993 ( .A1(n9587), .A2(n9490), .ZN(n9544) );
  AND2_X1 U5994 ( .A1(n5603), .A2(n5141), .ZN(n8967) );
  NAND2_X1 U5995 ( .A1(n5603), .A2(n5601), .ZN(n8995) );
  NAND2_X1 U5996 ( .A1(n9556), .A2(n9557), .ZN(n9555) );
  NAND2_X1 U5997 ( .A1(n9578), .A2(n9503), .ZN(n9556) );
  NAND2_X1 U5998 ( .A1(n7539), .A2(n5608), .ZN(n5607) );
  INV_X1 U5999 ( .A(n5610), .ZN(n5606) );
  OR2_X1 U6000 ( .A1(n7431), .A2(n7428), .ZN(n9613) );
  AOI21_X1 U6001 ( .B1(n5617), .B2(n5120), .A(n5615), .ZN(n5614) );
  INV_X1 U6002 ( .A(n8083), .ZN(n5615) );
  OR2_X1 U6003 ( .A1(n9536), .A2(n6307), .ZN(n9486) );
  OAI21_X1 U6004 ( .B1(n8965), .B2(n5602), .A(n5599), .ZN(n9143) );
  AND2_X1 U6005 ( .A1(n9601), .A2(n9597), .ZN(n9493) );
  AND4_X1 U6006 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n8021)
         );
  INV_X1 U6007 ( .A(n9557), .ZN(n5569) );
  AND2_X1 U6008 ( .A1(n5567), .A2(n9506), .ZN(n5566) );
  AND4_X1 U6009 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n9568)
         );
  NAND2_X1 U6010 ( .A1(n9201), .A2(n9200), .ZN(n9212) );
  INV_X1 U6011 ( .A(n9632), .ZN(n9600) );
  AND2_X1 U6012 ( .A1(n7425), .A2(n7741), .ZN(n9463) );
  NAND2_X1 U6013 ( .A1(n5628), .A2(n5627), .ZN(n9460) );
  NAND2_X1 U6014 ( .A1(n5409), .A2(n5410), .ZN(n5408) );
  INV_X1 U6015 ( .A(n9831), .ZN(n9637) );
  INV_X1 U6016 ( .A(n9830), .ZN(n9850) );
  INV_X1 U6017 ( .A(n9548), .ZN(n9881) );
  INV_X1 U6018 ( .A(n8001), .ZN(n9648) );
  INV_X1 U6019 ( .A(n5621), .ZN(n5623) );
  NAND4_X1 U6020 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n9651)
         );
  OR2_X1 U6021 ( .A1(n7405), .A2(n7281), .ZN(n11001) );
  NAND2_X1 U6022 ( .A1(n10942), .A2(n7700), .ZN(n7701) );
  INV_X1 U6023 ( .A(n7753), .ZN(n5355) );
  OAI21_X1 U6024 ( .B1(n7836), .B2(n5354), .A(n5353), .ZN(n7875) );
  NAND2_X1 U6025 ( .A1(n5357), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6026 ( .A1(n7753), .A2(n5357), .ZN(n5353) );
  INV_X1 U6027 ( .A(n7755), .ZN(n5357) );
  INV_X1 U6028 ( .A(n8929), .ZN(n5375) );
  AND2_X1 U6029 ( .A1(n6018), .A2(n6002), .ZN(n10975) );
  OR2_X1 U6030 ( .A1(n10986), .A2(n6005), .ZN(n5369) );
  NAND2_X1 U6031 ( .A1(n5366), .A2(n5364), .ZN(n9166) );
  NOR2_X1 U6032 ( .A1(n9167), .A2(n6043), .ZN(n9653) );
  INV_X1 U6033 ( .A(n5477), .ZN(n9688) );
  OAI21_X1 U6034 ( .B1(n9167), .B2(n5371), .A(n5370), .ZN(n9681) );
  NAND2_X1 U6035 ( .A1(n5372), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6036 ( .A1(n9654), .A2(n5372), .ZN(n5370) );
  INV_X1 U6037 ( .A(n9656), .ZN(n5372) );
  OR2_X1 U6038 ( .A1(n9682), .A2(n6071), .ZN(n5363) );
  INV_X1 U6039 ( .A(n5475), .ZN(n9735) );
  NAND2_X1 U6040 ( .A1(n5359), .A2(n5358), .ZN(n9724) );
  NAND2_X1 U6041 ( .A1(n5349), .A2(n5348), .ZN(n11013) );
  NAND2_X1 U6042 ( .A1(n9771), .A2(n10996), .ZN(n5480) );
  INV_X1 U6043 ( .A(n9770), .ZN(n5479) );
  XNOR2_X1 U6044 ( .A(n5482), .B(n9769), .ZN(n5481) );
  NOR2_X1 U6045 ( .A1(n11005), .A2(n9768), .ZN(n5482) );
  NOR2_X1 U6046 ( .A1(n9772), .A2(n11011), .ZN(n5211) );
  AND3_X1 U6047 ( .A1(n5349), .A2(n9747), .A3(n5348), .ZN(n9748) );
  INV_X1 U6048 ( .A(n6323), .ZN(n6254) );
  AND2_X1 U6049 ( .A1(n9260), .A2(n5831), .ZN(n9792) );
  NAND2_X1 U6050 ( .A1(n5278), .A2(n5279), .ZN(n9797) );
  OR2_X1 U6051 ( .A1(n9835), .A2(n5281), .ZN(n5278) );
  INV_X1 U6052 ( .A(n9441), .ZN(n9966) );
  NAND2_X1 U6053 ( .A1(n9789), .A2(n9788), .ZN(n9790) );
  NAND2_X1 U6054 ( .A1(n5630), .A2(n5283), .ZN(n9813) );
  NAND2_X1 U6055 ( .A1(n9835), .A2(n5137), .ZN(n5283) );
  AND2_X1 U6056 ( .A1(n6236), .A2(n6223), .ZN(n9822) );
  NAND2_X1 U6057 ( .A1(n5631), .A2(n6215), .ZN(n9821) );
  NAND2_X1 U6058 ( .A1(n9835), .A2(n6216), .ZN(n5631) );
  NAND2_X1 U6059 ( .A1(n9856), .A2(n9855), .ZN(n9854) );
  NAND2_X1 U6060 ( .A1(n9871), .A2(n6175), .ZN(n9856) );
  NAND2_X1 U6061 ( .A1(n6179), .A2(n6178), .ZN(n9987) );
  NAND2_X1 U6062 ( .A1(n6167), .A2(n6166), .ZN(n9874) );
  NAND2_X1 U6063 ( .A1(n6155), .A2(n6154), .ZN(n9996) );
  OR2_X1 U6064 ( .A1(n8823), .A2(n5851), .ZN(n6155) );
  OR2_X1 U6065 ( .A1(n9909), .A2(n9407), .ZN(n9899) );
  NAND2_X1 U6066 ( .A1(n6140), .A2(n6139), .ZN(n10000) );
  OAI21_X1 U6067 ( .B1(n6305), .B2(n5452), .A(n5450), .ZN(n9904) );
  NAND2_X1 U6068 ( .A1(n6305), .A2(n6304), .ZN(n9917) );
  NAND2_X1 U6069 ( .A1(n6103), .A2(n6102), .ZN(n10013) );
  NAND2_X1 U6070 ( .A1(n6087), .A2(n6086), .ZN(n10021) );
  OR2_X1 U6071 ( .A1(n10027), .A2(n7734), .ZN(n9843) );
  NAND2_X1 U6072 ( .A1(n5293), .A2(n9375), .ZN(n9109) );
  NAND2_X1 U6073 ( .A1(n5290), .A2(n5294), .ZN(n9108) );
  OAI21_X1 U6074 ( .B1(n8977), .B2(n5133), .A(n5445), .ZN(n9106) );
  NAND2_X1 U6075 ( .A1(n8977), .A2(n6291), .ZN(n9024) );
  NAND2_X1 U6076 ( .A1(n8983), .A2(n6029), .ZN(n9027) );
  NAND2_X1 U6077 ( .A1(n5304), .A2(n5305), .ZN(n8796) );
  OR2_X1 U6078 ( .A1(n5635), .A2(n5117), .ZN(n5304) );
  NAND2_X1 U6079 ( .A1(n5990), .A2(n5989), .ZN(n8906) );
  INV_X1 U6080 ( .A(n8548), .ZN(n11065) );
  NAND2_X1 U6081 ( .A1(n8009), .A2(n9345), .ZN(n7997) );
  INV_X1 U6082 ( .A(n11064), .ZN(n9913) );
  INV_X2 U6083 ( .A(n10023), .ZN(n10033) );
  INV_X1 U6084 ( .A(n6268), .ZN(n10040) );
  INV_X1 U6085 ( .A(n9630), .ZN(n10044) );
  INV_X1 U6086 ( .A(n9554), .ZN(n10048) );
  INV_X1 U6087 ( .A(n9574), .ZN(n10052) );
  INV_X1 U6088 ( .A(n9874), .ZN(n10057) );
  OR3_X1 U6089 ( .A1(n10031), .A2(n10030), .A3(n10029), .ZN(n11102) );
  NAND2_X1 U6090 ( .A1(n6353), .A2(n6352), .ZN(n7728) );
  OR2_X1 U6091 ( .A1(n7302), .A2(n7301), .ZN(n9238) );
  INV_X1 U6092 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n10069) );
  AND2_X1 U6093 ( .A1(n5299), .A2(n5824), .ZN(n5297) );
  NAND2_X1 U6094 ( .A1(n6257), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5570) );
  INV_X1 U6095 ( .A(n10957), .ZN(n8945) );
  INV_X1 U6096 ( .A(n7772), .ZN(n7877) );
  INV_X1 U6097 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U6098 ( .A1(n5659), .A2(n5664), .ZN(n10091) );
  OR2_X1 U6099 ( .A1(n9185), .A2(n6700), .ZN(n5659) );
  OR2_X1 U6100 ( .A1(n10230), .A2(n5136), .ZN(n5232) );
  OR2_X1 U6101 ( .A1(n6718), .A2(n5136), .ZN(n5233) );
  NAND2_X1 U6102 ( .A1(n10222), .A2(n6926), .ZN(n7267) );
  NAND2_X1 U6103 ( .A1(n5216), .A2(n8694), .ZN(n8772) );
  NAND2_X1 U6104 ( .A1(n6592), .A2(n5189), .ZN(n5216) );
  NAND2_X1 U6105 ( .A1(n7326), .A2(n5390), .ZN(n5389) );
  OAI21_X1 U6106 ( .B1(n7288), .B2(n5392), .A(n5391), .ZN(n5390) );
  AND4_X1 U6107 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n9191)
         );
  INV_X1 U6108 ( .A(n10647), .ZN(n10496) );
  AND2_X1 U6109 ( .A1(n6891), .A2(n6878), .ZN(n10497) );
  NAND2_X1 U6110 ( .A1(n10101), .A2(n6855), .ZN(n10159) );
  INV_X1 U6111 ( .A(n8711), .ZN(n11036) );
  NAND2_X1 U6112 ( .A1(n8827), .A2(n8826), .ZN(n8825) );
  INV_X1 U6113 ( .A(n10233), .ZN(n10169) );
  OR2_X1 U6114 ( .A1(n6787), .A2(n6786), .ZN(n6788) );
  NAND2_X1 U6115 ( .A1(n6791), .A2(n6790), .ZN(n10684) );
  AND4_X1 U6116 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n10179)
         );
  AND2_X1 U6117 ( .A1(n9185), .A2(n6680), .ZN(n10173) );
  AOI22_X1 U6118 ( .A1(n5224), .A2(n5228), .B1(n5226), .B2(n5220), .ZN(n5219)
         );
  INV_X1 U6119 ( .A(n8826), .ZN(n5220) );
  INV_X1 U6120 ( .A(n10236), .ZN(n10200) );
  INV_X1 U6121 ( .A(n5642), .ZN(n10205) );
  AOI21_X1 U6122 ( .B1(n10133), .B2(n5647), .A(n5646), .ZN(n5642) );
  NAND2_X1 U6123 ( .A1(n6953), .A2(n10435), .ZN(n10215) );
  AND2_X1 U6124 ( .A1(n6951), .A2(n6949), .ZN(n10223) );
  AND2_X1 U6125 ( .A1(n6966), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10241) );
  INV_X1 U6126 ( .A(n10223), .ZN(n10243) );
  INV_X1 U6127 ( .A(n10634), .ZN(n10480) );
  INV_X1 U6128 ( .A(n10669), .ZN(n10577) );
  INV_X1 U6129 ( .A(n10209), .ZN(n10694) );
  INV_X1 U6130 ( .A(n9191), .ZN(n10733) );
  OR2_X1 U6131 ( .A1(n7329), .A2(n7331), .ZN(n10367) );
  AOI21_X1 U6132 ( .B1(n10461), .B2(n5560), .A(n5208), .ZN(n10430) );
  AOI21_X1 U6133 ( .B1(n10471), .B2(n5560), .A(n10428), .ZN(n5559) );
  AND2_X1 U6134 ( .A1(n5562), .A2(n5560), .ZN(n10444) );
  NAND2_X1 U6135 ( .A1(n5562), .A2(n10426), .ZN(n10445) );
  XNOR2_X1 U6136 ( .A(n10461), .B(n5563), .ZN(n10630) );
  AND4_X1 U6137 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(n10633)
         );
  AND4_X1 U6138 ( .A1(n6896), .A2(n6895), .A3(n6894), .A4(n6893), .ZN(n10643)
         );
  NAND2_X1 U6139 ( .A1(n10420), .A2(n5550), .ZN(n10649) );
  NAND2_X1 U6140 ( .A1(n10420), .A2(n10419), .ZN(n10494) );
  AND4_X1 U6141 ( .A1(n6865), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(n10644)
         );
  AND4_X1 U6142 ( .A1(n6847), .A2(n6846), .A3(n6845), .A4(n6844), .ZN(n10668)
         );
  NAND2_X1 U6143 ( .A1(n5318), .A2(n7221), .ZN(n9160) );
  NAND2_X1 U6144 ( .A1(n9081), .A2(n7190), .ZN(n5318) );
  NAND2_X1 U6145 ( .A1(n9155), .A2(n9159), .ZN(n9220) );
  NAND2_X1 U6146 ( .A1(n9154), .A2(n9153), .ZN(n9155) );
  NAND2_X1 U6147 ( .A1(n8722), .A2(n7155), .ZN(n8864) );
  NAND2_X1 U6148 ( .A1(n5553), .A2(n8855), .ZN(n9005) );
  NAND2_X1 U6149 ( .A1(n7152), .A2(n7151), .ZN(n8686) );
  NAND2_X1 U6150 ( .A1(n8679), .A2(n8678), .ZN(n8726) );
  INV_X1 U6151 ( .A(n10599), .ZN(n11047) );
  AND4_X1 U6152 ( .A1(n6580), .A2(n6579), .A3(n6578), .A4(n6577), .ZN(n8698)
         );
  AND4_X1 U6153 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n8697)
         );
  OR2_X1 U6154 ( .A1(n10596), .A2(n11020), .ZN(n10548) );
  INV_X1 U6155 ( .A(n10603), .ZN(n11053) );
  INV_X1 U6156 ( .A(n10440), .ZN(n10536) );
  OR2_X1 U6157 ( .A1(n10596), .A2(n6773), .ZN(n11050) );
  NAND2_X1 U6158 ( .A1(n6462), .A2(n6461), .ZN(n8564) );
  NAND2_X1 U6159 ( .A1(n6774), .A2(n10283), .ZN(n6507) );
  INV_X1 U6160 ( .A(n10379), .ZN(n10743) );
  INV_X1 U6161 ( .A(n7124), .ZN(n10747) );
  INV_X1 U6162 ( .A(n10529), .ZN(n10764) );
  INV_X1 U6163 ( .A(n10561), .ZN(n10772) );
  INV_X1 U6164 ( .A(n9006), .ZN(n10184) );
  INV_X1 U6165 ( .A(n7009), .ZN(n7815) );
  AND3_X1 U6166 ( .A1(n6483), .A2(P1_STATE_REG_SCAN_IN), .A3(n7325), .ZN(
        n10803) );
  NAND2_X1 U6167 ( .A1(n6450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6451) );
  NOR2_X1 U6168 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5205) );
  INV_X1 U6169 ( .A(n6428), .ZN(n6430) );
  XNOR2_X1 U6170 ( .A(n6177), .B(n6176), .ZN(n9134) );
  MUX2_X1 U6171 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6432), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6434) );
  NAND2_X1 U6172 ( .A1(n5511), .A2(n5510), .ZN(n6112) );
  NAND2_X1 U6173 ( .A1(n5533), .A2(n5531), .ZN(n6062) );
  NAND2_X1 U6174 ( .A1(n5533), .A2(n5752), .ZN(n6064) );
  NAND2_X1 U6175 ( .A1(n5518), .A2(n5516), .ZN(n6016) );
  AND2_X1 U6176 ( .A1(n6630), .A2(n6415), .ZN(n7531) );
  OR2_X1 U6177 ( .A1(n5931), .A2(n5930), .ZN(n5932) );
  NAND2_X1 U6178 ( .A1(n5910), .A2(n5909), .ZN(n7300) );
  NAND2_X1 U6179 ( .A1(n7550), .A2(n5612), .ZN(n7554) );
  INV_X1 U6180 ( .A(n5356), .ZN(n7835) );
  INV_X1 U6181 ( .A(n5376), .ZN(n8928) );
  NAND2_X1 U6182 ( .A1(n5212), .A2(n5210), .ZN(P2_U3201) );
  NOR2_X1 U6183 ( .A1(n5211), .A2(n5478), .ZN(n5210) );
  NAND2_X1 U6184 ( .A1(n5481), .A2(n10983), .ZN(n5212) );
  NAND2_X1 U6185 ( .A1(n5480), .A2(n5479), .ZN(n5478) );
  OAI21_X1 U6186 ( .B1(n5472), .B2(n11105), .A(n5198), .ZN(P2_U3456) );
  INV_X1 U6187 ( .A(n5199), .ZN(n5198) );
  NAND2_X1 U6188 ( .A1(n11093), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6189 ( .A1(n10748), .A2(n11094), .ZN(n5381) );
  AOI21_X1 U6190 ( .B1(n10750), .B2(n11094), .A(n5340), .ZN(n10632) );
  NAND2_X1 U6191 ( .A1(n5342), .A2(n5341), .ZN(n5340) );
  NAND2_X1 U6192 ( .A1(n11093), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6193 ( .A1(n5201), .A2(n5186), .ZN(n10751) );
  AND2_X1 U6194 ( .A1(n9987), .A2(n9639), .ZN(n5116) );
  INV_X1 U6195 ( .A(n8618), .ZN(n5458) );
  OR2_X1 U6196 ( .A1(n9355), .A2(n9356), .ZN(n5117) );
  NAND2_X1 U6197 ( .A1(n9910), .A2(n9919), .ZN(n5118) );
  AND2_X1 U6198 ( .A1(n5663), .A2(n5667), .ZN(n5119) );
  INV_X1 U6199 ( .A(n9281), .ZN(n5289) );
  AND2_X1 U6200 ( .A1(n8017), .A2(n5193), .ZN(n5120) );
  AND2_X1 U6201 ( .A1(n5456), .A2(n5149), .ZN(n5121) );
  AND2_X1 U6202 ( .A1(n5576), .A2(n9476), .ZN(n5122) );
  AND2_X1 U6203 ( .A1(n5169), .A2(n6315), .ZN(n5123) );
  OR3_X1 U6204 ( .A1(n10044), .A2(n5422), .A3(n9637), .ZN(n5124) );
  INV_X1 U6205 ( .A(n10511), .ZN(n5252) );
  AND2_X1 U6206 ( .A1(n9454), .A2(n9458), .ZN(n5125) );
  AND2_X1 U6207 ( .A1(n5452), .A2(n5118), .ZN(n5126) );
  NAND2_X1 U6208 ( .A1(n5571), .A2(n5573), .ZN(n5127) );
  INV_X1 U6209 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U6210 ( .A1(n5511), .A2(n5512), .ZN(n5128) );
  INV_X1 U6211 ( .A(n5386), .ZN(n5385) );
  NAND2_X1 U6212 ( .A1(n5388), .A2(n5387), .ZN(n5386) );
  NAND2_X1 U6213 ( .A1(n5497), .A2(n5962), .ZN(n5129) );
  NOR2_X1 U6214 ( .A1(n9650), .A2(n7648), .ZN(n9334) );
  INV_X1 U6215 ( .A(n9334), .ZN(n5424) );
  AND2_X1 U6216 ( .A1(n9452), .A2(n9305), .ZN(n5130) );
  AND2_X1 U6217 ( .A1(n5223), .A2(n5227), .ZN(n5131) );
  NAND2_X1 U6218 ( .A1(n8966), .A2(n5141), .ZN(n5602) );
  NAND2_X1 U6219 ( .A1(n5675), .A2(n6541), .ZN(n8029) );
  NOR2_X1 U6220 ( .A1(n6772), .A2(n10145), .ZN(n5132) );
  INV_X1 U6221 ( .A(n6635), .ZN(n6990) );
  INV_X1 U6222 ( .A(n6505), .ZN(n6569) );
  INV_X1 U6223 ( .A(n7287), .ZN(n5392) );
  AND2_X1 U6224 ( .A1(n6549), .A2(n8479), .ZN(n6411) );
  NOR2_X1 U6225 ( .A1(n9022), .A2(n9642), .ZN(n5133) );
  INV_X1 U6226 ( .A(n7757), .ZN(n7748) );
  AND2_X1 U6227 ( .A1(n9575), .A2(n5582), .ZN(n5134) );
  OR2_X1 U6228 ( .A1(n9508), .A2(n9637), .ZN(n5135) );
  NOR2_X1 U6229 ( .A1(n5643), .A2(n5649), .ZN(n5136) );
  AND2_X1 U6230 ( .A1(n6216), .A2(n6228), .ZN(n5137) );
  AND2_X1 U6231 ( .A1(n6818), .A2(n6806), .ZN(n5138) );
  NAND2_X1 U6232 ( .A1(n9855), .A2(n9868), .ZN(n5139) );
  AND2_X1 U6233 ( .A1(n5458), .A2(n9312), .ZN(n5140) );
  NAND2_X1 U6234 ( .A1(n8963), .A2(n8975), .ZN(n5141) );
  NAND2_X1 U6235 ( .A1(n10649), .A2(n10421), .ZN(n10478) );
  AND2_X1 U6236 ( .A1(n10391), .A2(n10392), .ZN(n5142) );
  NAND2_X1 U6237 ( .A1(n7177), .A2(n7178), .ZN(n10429) );
  AND2_X1 U6238 ( .A1(n5464), .A2(n5462), .ZN(n5143) );
  NAND2_X1 U6239 ( .A1(n5389), .A2(n5393), .ZN(n7009) );
  INV_X1 U6240 ( .A(n10620), .ZN(n5396) );
  INV_X1 U6241 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6437) );
  AND2_X1 U6242 ( .A1(n6506), .A2(n6394), .ZN(n6549) );
  INV_X1 U6243 ( .A(n9390), .ZN(n5432) );
  NAND2_X1 U6244 ( .A1(n10102), .A2(n10103), .ZN(n10101) );
  OAI21_X1 U6245 ( .B1(n10133), .B2(n5652), .A(n5649), .ZN(n10204) );
  OR2_X1 U6246 ( .A1(n7456), .A2(n7708), .ZN(n5144) );
  NAND2_X1 U6247 ( .A1(n5673), .A2(n5138), .ZN(n10119) );
  NAND2_X1 U6248 ( .A1(n10218), .A2(n6903), .ZN(n10222) );
  XOR2_X1 U6249 ( .A(n5572), .B(n9513), .Z(n5145) );
  NAND2_X1 U6250 ( .A1(n9319), .A2(n9328), .ZN(n9325) );
  INV_X1 U6251 ( .A(n9325), .ZN(n5426) );
  OAI21_X1 U6252 ( .B1(n5218), .B2(n5217), .A(n10156), .ZN(n10125) );
  NAND2_X1 U6253 ( .A1(n6113), .A2(n5809), .ZN(n5146) );
  INV_X1 U6254 ( .A(n7054), .ZN(n7221) );
  AND2_X1 U6255 ( .A1(n7159), .A2(n7190), .ZN(n5147) );
  AND2_X1 U6256 ( .A1(n8993), .A2(n8994), .ZN(n5148) );
  INV_X1 U6257 ( .A(n5228), .ZN(n5227) );
  OAI21_X1 U6258 ( .B1(n8826), .B2(n5229), .A(n6629), .ZN(n5228) );
  OR2_X1 U6259 ( .A1(n8906), .A2(n9644), .ZN(n5149) );
  INV_X1 U6260 ( .A(n8854), .ZN(n11089) );
  NAND2_X1 U6261 ( .A1(n6652), .A2(n6651), .ZN(n8854) );
  INV_X1 U6262 ( .A(n9348), .ZN(n7998) );
  AND2_X1 U6263 ( .A1(n9353), .A2(n9311), .ZN(n9348) );
  INV_X1 U6264 ( .A(n5114), .ZN(n10462) );
  NOR2_X1 U6265 ( .A1(n10484), .A2(n10752), .ZN(n5397) );
  AND2_X1 U6266 ( .A1(n10706), .A2(n10711), .ZN(n5150) );
  AND2_X1 U6267 ( .A1(n7105), .A2(n10397), .ZN(n5151) );
  AND2_X1 U6268 ( .A1(n10521), .A2(n10415), .ZN(n5152) );
  INV_X1 U6269 ( .A(n5667), .ZN(n5666) );
  OAI21_X1 U6270 ( .B1(n6680), .B2(n5668), .A(n5669), .ZN(n5667) );
  NAND2_X1 U6271 ( .A1(n9630), .A2(n9637), .ZN(n5153) );
  NAND2_X1 U6272 ( .A1(n9394), .A2(n9399), .ZN(n9927) );
  INV_X1 U6273 ( .A(n9927), .ZN(n5452) );
  AND2_X1 U6274 ( .A1(n8906), .A2(n9644), .ZN(n5154) );
  INV_X1 U6275 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8507) );
  INV_X1 U6276 ( .A(n6629), .ZN(n5230) );
  AND2_X1 U6277 ( .A1(n9574), .A2(n9850), .ZN(n5155) );
  NOR2_X1 U6278 ( .A1(n9910), .A2(n9919), .ZN(n5156) );
  AND2_X1 U6279 ( .A1(n9064), .A2(n8727), .ZN(n5157) );
  OR2_X1 U6280 ( .A1(n6229), .A2(n9430), .ZN(n5158) );
  NAND2_X1 U6281 ( .A1(n10521), .A2(n7071), .ZN(n5159) );
  AND2_X1 U6282 ( .A1(n8803), .A2(n8783), .ZN(n5160) );
  AND2_X1 U6283 ( .A1(n9006), .A2(n10733), .ZN(n5161) );
  OR2_X1 U6284 ( .A1(n9378), .A2(n9377), .ZN(n5162) );
  INV_X1 U6285 ( .A(n5243), .ZN(n5982) );
  NAND2_X1 U6286 ( .A1(n6435), .A2(n5688), .ZN(n5163) );
  NOR2_X1 U6287 ( .A1(n9479), .A2(n9568), .ZN(n5164) );
  NAND2_X1 U6288 ( .A1(n9141), .A2(n9642), .ZN(n5165) );
  INV_X1 U6289 ( .A(n6855), .ZN(n5658) );
  OR2_X1 U6290 ( .A1(n5734), .A2(SI_9_), .ZN(n5166) );
  NAND2_X1 U6291 ( .A1(n9346), .A2(n9345), .ZN(n5167) );
  INV_X1 U6292 ( .A(n5497), .ZN(n5496) );
  NOR2_X1 U6293 ( .A1(n5498), .A2(n5946), .ZN(n5497) );
  AND2_X1 U6294 ( .A1(n5733), .A2(n5732), .ZN(n5168) );
  AND2_X1 U6295 ( .A1(n6013), .A2(n9361), .ZN(n8795) );
  OR2_X1 U6296 ( .A1(n9574), .A2(n9850), .ZN(n5169) );
  OAI21_X1 U6297 ( .B1(n10103), .B2(n5658), .A(n10157), .ZN(n5657) );
  NAND2_X1 U6298 ( .A1(n5440), .A2(n5441), .ZN(n5622) );
  INV_X1 U6299 ( .A(n5622), .ZN(n5308) );
  AND3_X1 U6300 ( .A1(n5870), .A2(n5869), .A3(n5868), .ZN(n7805) );
  INV_X1 U6301 ( .A(n7805), .ZN(n5428) );
  INV_X1 U6302 ( .A(n5602), .ZN(n5601) );
  AND2_X1 U6303 ( .A1(n6705), .A2(n6704), .ZN(n10723) );
  INV_X1 U6304 ( .A(n10723), .ZN(n9053) );
  OR2_X1 U6305 ( .A1(n5159), .A2(n5256), .ZN(n5170) );
  INV_X1 U6306 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8495) );
  AND2_X1 U6307 ( .A1(n5529), .A2(n5527), .ZN(n5171) );
  OR2_X1 U6308 ( .A1(n7243), .A2(n7096), .ZN(n5172) );
  AND2_X1 U6309 ( .A1(n5452), .A2(n9392), .ZN(n5173) );
  INV_X1 U6310 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5604) );
  AND2_X1 U6311 ( .A1(n10619), .A2(n5196), .ZN(n5174) );
  AND2_X1 U6312 ( .A1(n10532), .A2(n10415), .ZN(n5175) );
  OR2_X1 U6313 ( .A1(n9489), .A2(n5580), .ZN(n5176) );
  NAND2_X1 U6314 ( .A1(n7072), .A2(n10395), .ZN(n10521) );
  INV_X1 U6315 ( .A(n7923), .ZN(n5558) );
  AND2_X1 U6316 ( .A1(n5363), .A2(n5362), .ZN(n5177) );
  INV_X1 U6317 ( .A(n7073), .ZN(n5256) );
  AND2_X1 U6318 ( .A1(n5676), .A2(n8507), .ZN(n5178) );
  INV_X1 U6319 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U6320 ( .A1(n5632), .A2(n6188), .ZN(n5179) );
  INV_X1 U6321 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U6322 ( .A1(n5428), .A2(n5427), .ZN(n9328) );
  INV_X1 U6323 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8518) );
  INV_X1 U6324 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5488) );
  INV_X1 U6325 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5312) );
  AND2_X1 U6326 ( .A1(n5352), .A2(n5351), .ZN(n5180) );
  INV_X1 U6327 ( .A(n9449), .ZN(n5422) );
  NAND2_X1 U6328 ( .A1(n9186), .A2(n9187), .ZN(n9185) );
  NAND2_X1 U6329 ( .A1(n6946), .A2(n6773), .ZN(n7096) );
  INV_X1 U6330 ( .A(n7190), .ZN(n5320) );
  NAND2_X1 U6331 ( .A1(n6411), .A2(n6399), .ZN(n6646) );
  NAND2_X1 U6332 ( .A1(n6399), .A2(n5539), .ZN(n6661) );
  NAND2_X1 U6333 ( .A1(n9212), .A2(n9211), .ZN(n9477) );
  NAND2_X1 U6334 ( .A1(n6285), .A2(n6284), .ZN(n8617) );
  OR2_X1 U6335 ( .A1(n6435), .A2(n6447), .ZN(n6735) );
  OR2_X1 U6336 ( .A1(n10173), .A2(n5668), .ZN(n5181) );
  NOR2_X1 U6337 ( .A1(n9653), .A2(n9654), .ZN(n5182) );
  INV_X1 U6338 ( .A(n9490), .ZN(n5580) );
  OR2_X1 U6339 ( .A1(n9412), .A2(n5422), .ZN(n5183) );
  AND2_X1 U6340 ( .A1(n8825), .A2(n5226), .ZN(n5184) );
  AND2_X1 U6341 ( .A1(n5369), .A2(n5368), .ZN(n5185) );
  NAND2_X1 U6342 ( .A1(n6442), .A2(n6441), .ZN(n6944) );
  INV_X1 U6343 ( .A(n5760), .ZN(n5512) );
  INV_X1 U6344 ( .A(n9711), .ZN(n5213) );
  NAND2_X1 U6345 ( .A1(n5303), .A2(n5302), .ZN(n8794) );
  OR2_X1 U6346 ( .A1(n11079), .A2(n5200), .ZN(n5186) );
  AND2_X1 U6347 ( .A1(n8729), .A2(n5385), .ZN(n5187) );
  NAND2_X1 U6348 ( .A1(n6688), .A2(n6687), .ZN(n10729) );
  INV_X1 U6349 ( .A(n10729), .ZN(n5387) );
  OR2_X1 U6350 ( .A1(n8954), .A2(n9165), .ZN(n5188) );
  NAND2_X1 U6351 ( .A1(n5635), .A2(n9312), .ZN(n8614) );
  INV_X1 U6352 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8303) );
  OR2_X1 U6353 ( .A1(n6607), .A2(n6606), .ZN(n5189) );
  AND2_X1 U6354 ( .A1(n5356), .A2(n5355), .ZN(n5190) );
  AND2_X1 U6355 ( .A1(n5376), .A2(n5375), .ZN(n5191) );
  INV_X1 U6356 ( .A(n5791), .ZN(n5524) );
  NAND2_X1 U6357 ( .A1(n9736), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5192) );
  AND2_X2 U6358 ( .A1(n7793), .A2(n10785), .ZN(n11094) );
  NAND2_X1 U6359 ( .A1(n5308), .A2(n5623), .ZN(n6271) );
  INV_X1 U6360 ( .A(n9302), .ZN(n9323) );
  XNOR2_X1 U6361 ( .A(n5570), .B(n6259), .ZN(n9302) );
  OR2_X1 U6362 ( .A1(n8019), .A2(n9646), .ZN(n5193) );
  OR2_X1 U6363 ( .A1(n6504), .A2(n6503), .ZN(n7939) );
  AND2_X1 U6364 ( .A1(n7550), .A2(n5610), .ZN(n5194) );
  OR2_X1 U6365 ( .A1(n11010), .A2(n9726), .ZN(n5195) );
  XNOR2_X1 U6366 ( .A(n6439), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6947) );
  XNOR2_X1 U6367 ( .A(n6265), .B(P2_IR_REG_20__SCAN_IN), .ZN(n9458) );
  XNOR2_X1 U6368 ( .A(n6451), .B(n8323), .ZN(n9473) );
  NAND2_X1 U6369 ( .A1(n5297), .A2(n5298), .ZN(n10068) );
  INV_X1 U6370 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7916) );
  INV_X1 U6371 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5247) );
  INV_X1 U6372 ( .A(n10198), .ZN(n8103) );
  INV_X1 U6373 ( .A(n6429), .ZN(n6408) );
  NAND2_X1 U6374 ( .A1(n5982), .A2(n5739), .ZN(n5985) );
  NAND2_X1 U6375 ( .A1(n5777), .A2(n5778), .ZN(n6163) );
  NOR2_X1 U6376 ( .A1(n5301), .A2(n5179), .ZN(n5300) );
  INV_X1 U6377 ( .A(n10398), .ZN(n10493) );
  INV_X1 U6378 ( .A(n5550), .ZN(n5548) );
  NAND2_X1 U6379 ( .A1(n5548), .A2(n10421), .ZN(n5547) );
  NAND2_X1 U6380 ( .A1(n5578), .A2(n5579), .ZN(n9598) );
  NAND2_X1 U6381 ( .A1(n9523), .A2(n9522), .ZN(n9521) );
  NAND2_X1 U6382 ( .A1(n8786), .A2(n8785), .ZN(n8909) );
  INV_X1 U6383 ( .A(n7968), .ZN(n5618) );
  INV_X1 U6384 ( .A(n9622), .ZN(n9507) );
  NAND2_X1 U6385 ( .A1(n5616), .A2(n5614), .ZN(n8086) );
  NAND3_X1 U6386 ( .A1(n9460), .A2(n5408), .A3(n5407), .ZN(n9461) );
  NAND2_X2 U6387 ( .A1(n6062), .A2(n6065), .ZN(n7652) );
  OR2_X2 U6388 ( .A1(n6050), .A2(n6049), .ZN(n5533) );
  NAND2_X1 U6389 ( .A1(n5277), .A2(n5275), .ZN(n9795) );
  NAND2_X1 U6390 ( .A1(n5215), .A2(n5252), .ZN(n10514) );
  INV_X1 U6391 ( .A(n5559), .ZN(n5208) );
  NAND2_X1 U6392 ( .A1(n5381), .A2(n5380), .ZN(P1_U3551) );
  NAND2_X1 U6393 ( .A1(n5518), .A2(n5743), .ZN(n6015) );
  NAND2_X1 U6394 ( .A1(n5203), .A2(n5202), .ZN(n5518) );
  INV_X1 U6395 ( .A(n5999), .ZN(n5203) );
  OAI21_X1 U6396 ( .B1(n7152), .B2(n7212), .A(n5331), .ZN(n7157) );
  OAI21_X1 U6397 ( .B1(n10625), .B2(n11021), .A(n10624), .ZN(n10749) );
  INV_X1 U6398 ( .A(n5344), .ZN(n5343) );
  INV_X1 U6399 ( .A(n11046), .ZN(n7946) );
  NAND3_X1 U6400 ( .A1(n5240), .A2(n6399), .A3(n6549), .ZN(n6685) );
  AND4_X2 U6401 ( .A1(n6398), .A2(n6397), .A3(n6395), .A4(n6396), .ZN(n6399)
         );
  NOR2_X1 U6402 ( .A1(n5206), .A2(n5205), .ZN(n5204) );
  OAI21_X1 U6403 ( .B1(n10630), .B2(n11021), .A(n5345), .ZN(n5344) );
  NAND2_X2 U6404 ( .A1(n5207), .A2(n5204), .ZN(n10791) );
  NAND2_X1 U6405 ( .A1(n5541), .A2(n5540), .ZN(n8852) );
  NAND4_X1 U6406 ( .A1(n6436), .A2(n5311), .A3(n5313), .A4(n6437), .ZN(n5209)
         );
  OAI211_X1 U6407 ( .C1(n10420), .C2(n5549), .A(n5547), .B(n10422), .ZN(n10424) );
  NAND2_X1 U6408 ( .A1(n10926), .A2(n5486), .ZN(n5485) );
  NOR2_X1 U6409 ( .A1(n9669), .A2(n9670), .ZN(n9673) );
  NOR2_X1 U6410 ( .A1(n9712), .A2(n9713), .ZN(n9717) );
  NAND2_X1 U6411 ( .A1(n5528), .A2(n5171), .ZN(n5758) );
  INV_X4 U6412 ( .A(n5816), .ZN(n7287) );
  NAND2_X2 U6413 ( .A1(n5692), .A2(n5693), .ZN(n5816) );
  NAND2_X1 U6414 ( .A1(n5515), .A2(n5513), .ZN(n6031) );
  NAND2_X1 U6415 ( .A1(n6031), .A2(n6030), .ZN(n6033) );
  INV_X1 U6416 ( .A(n10394), .ZN(n5330) );
  INV_X2 U6417 ( .A(n10545), .ZN(n10768) );
  AOI21_X1 U6418 ( .B1(n5323), .B2(n5325), .A(n10521), .ZN(n5321) );
  OAI21_X1 U6419 ( .B1(n10614), .B2(n11020), .A(n5174), .ZN(n10748) );
  NAND2_X1 U6420 ( .A1(n7278), .A2(n7279), .ZN(P1_U3220) );
  NAND2_X1 U6421 ( .A1(n5231), .A2(n5234), .ZN(n6789) );
  NAND3_X1 U6422 ( .A1(n6718), .A2(n10230), .A3(n5641), .ZN(n5231) );
  NAND3_X1 U6423 ( .A1(n5233), .A2(n5641), .A3(n5232), .ZN(n10109) );
  AND2_X1 U6424 ( .A1(n5236), .A2(n7940), .ZN(n10195) );
  NAND2_X1 U6425 ( .A1(n7939), .A2(n7941), .ZN(n5236) );
  INV_X1 U6426 ( .A(n6714), .ZN(n6717) );
  NAND3_X1 U6427 ( .A1(n6555), .A2(n5675), .A3(n6541), .ZN(n8030) );
  NAND3_X1 U6428 ( .A1(n6399), .A2(n6549), .A3(n5239), .ZN(n6701) );
  AND2_X1 U6429 ( .A1(n5674), .A2(n8495), .ZN(n5240) );
  NAND2_X1 U6430 ( .A1(n5241), .A2(n7095), .ZN(n7063) );
  NAND2_X1 U6431 ( .A1(n5242), .A2(n7162), .ZN(n5241) );
  OR2_X1 U6432 ( .A1(n7058), .A2(n7120), .ZN(n5242) );
  INV_X1 U6433 ( .A(n5493), .ZN(n5244) );
  XNOR2_X1 U6434 ( .A(n5999), .B(n5998), .ZN(n7337) );
  NAND2_X1 U6435 ( .A1(n5151), .A2(n5255), .ZN(n5253) );
  OAI21_X1 U6436 ( .B1(n7100), .B2(n5272), .A(n5270), .ZN(n7129) );
  NOR2_X1 U6437 ( .A1(n5269), .A2(n5267), .ZN(n7188) );
  NAND2_X1 U6438 ( .A1(n9835), .A2(n5279), .ZN(n5277) );
  NAND2_X1 U6439 ( .A1(n8983), .A2(n5294), .ZN(n5292) );
  NAND2_X1 U6440 ( .A1(n8983), .A2(n5296), .ZN(n5293) );
  AND2_X1 U6441 ( .A1(n5298), .A2(n5299), .ZN(n5823) );
  NAND2_X1 U6442 ( .A1(n5299), .A2(n5471), .ZN(n5814) );
  NAND2_X1 U6443 ( .A1(n9846), .A2(n6200), .ZN(n6202) );
  NAND2_X1 U6444 ( .A1(n5635), .A2(n5305), .ZN(n5303) );
  AND2_X2 U6445 ( .A1(n5620), .A2(n9326), .ZN(n9280) );
  NAND2_X1 U6446 ( .A1(n7621), .A2(n7620), .ZN(n7619) );
  OAI21_X1 U6447 ( .B1(n10553), .B2(n5325), .A(n5323), .ZN(n10519) );
  NAND2_X1 U6448 ( .A1(n5322), .A2(n5321), .ZN(n10396) );
  NAND2_X1 U6449 ( .A1(n10553), .A2(n5323), .ZN(n5322) );
  AOI21_X2 U6450 ( .B1(n5326), .B2(n10390), .A(n5324), .ZN(n5323) );
  INV_X1 U6451 ( .A(n10553), .ZN(n5329) );
  AOI21_X1 U6452 ( .B1(n7155), .B2(n5334), .A(n5332), .ZN(n5331) );
  AND2_X1 U6453 ( .A1(n6429), .A2(n5336), .ZN(n6449) );
  NAND2_X1 U6454 ( .A1(n6429), .A2(n8316), .ZN(n6407) );
  NAND2_X1 U6455 ( .A1(n6429), .A2(n5337), .ZN(n6450) );
  INV_X1 U6456 ( .A(n5347), .ZN(n7688) );
  NAND2_X1 U6457 ( .A1(n10921), .A2(n10920), .ZN(n10925) );
  NAND2_X1 U6458 ( .A1(n5144), .A2(n7457), .ZN(n7458) );
  OR2_X1 U6459 ( .A1(n9725), .A2(n9726), .ZN(n5352) );
  INV_X1 U6460 ( .A(n5352), .ZN(n9745) );
  INV_X1 U6461 ( .A(n9746), .ZN(n5351) );
  XNOR2_X1 U6462 ( .A(n7752), .B(n7766), .ZN(n7836) );
  INV_X1 U6463 ( .A(n5363), .ZN(n9700) );
  INV_X1 U6464 ( .A(n9701), .ZN(n5362) );
  INV_X1 U6465 ( .A(n5369), .ZN(n10985) );
  INV_X1 U6466 ( .A(n8932), .ZN(n5368) );
  MUX2_X1 U6467 ( .A(n5857), .B(P2_REG1_REG_2__SCAN_IN), .S(n7453), .Z(n10906)
         );
  NAND2_X1 U6468 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5379) );
  NOR2_X2 U6469 ( .A1(n10541), .A2(n10529), .ZN(n10505) );
  NOR2_X2 U6470 ( .A1(n10570), .A2(n10561), .ZN(n10560) );
  AND2_X2 U6471 ( .A1(n8729), .A2(n5384), .ZN(n9082) );
  NAND2_X2 U6472 ( .A1(n7326), .A2(n7287), .ZN(n6872) );
  AND2_X2 U6473 ( .A1(n7326), .A2(n5392), .ZN(n6505) );
  NAND2_X2 U6474 ( .A1(n6959), .A2(n10795), .ZN(n7326) );
  NAND3_X1 U6475 ( .A1(n6959), .A2(n10795), .A3(n10266), .ZN(n5393) );
  INV_X2 U6476 ( .A(n7326), .ZN(n6774) );
  NOR2_X2 U6477 ( .A1(n10506), .A2(n10647), .ZN(n10495) );
  AND2_X2 U6478 ( .A1(n5564), .A2(n6403), .ZN(n6429) );
  NAND3_X1 U6479 ( .A1(n9411), .A2(n9886), .A3(n5183), .ZN(n5406) );
  NAND2_X1 U6480 ( .A1(n9456), .A2(n5409), .ZN(n5407) );
  INV_X1 U6481 ( .A(n5413), .ZN(n5412) );
  NAND2_X1 U6482 ( .A1(n9454), .A2(n9453), .ZN(n5413) );
  NAND3_X1 U6483 ( .A1(n5423), .A2(n5421), .A3(n5419), .ZN(n5418) );
  NAND3_X1 U6484 ( .A1(n9328), .A2(n5425), .A3(n5424), .ZN(n9329) );
  NAND3_X1 U6485 ( .A1(n6113), .A2(n5639), .A3(n5640), .ZN(n6348) );
  AND2_X2 U6486 ( .A1(n5805), .A2(n5881), .ZN(n6113) );
  AND3_X4 U6487 ( .A1(n5437), .A2(n5438), .A3(n5856), .ZN(n7860) );
  OR2_X1 U6488 ( .A1(n5845), .A2(n7289), .ZN(n5438) );
  INV_X1 U6489 ( .A(n5442), .ZN(n6294) );
  INV_X1 U6490 ( .A(n6305), .ZN(n5447) );
  OAI21_X1 U6491 ( .B1(n5447), .B2(n5449), .A(n5448), .ZN(n9892) );
  NAND2_X1 U6492 ( .A1(n6285), .A2(n5121), .ZN(n5454) );
  NAND2_X1 U6493 ( .A1(n9849), .A2(n5123), .ZN(n5460) );
  NAND2_X1 U6494 ( .A1(n6320), .A2(n5465), .ZN(n5464) );
  NAND2_X1 U6495 ( .A1(n6320), .A2(n5467), .ZN(n5470) );
  NAND2_X1 U6496 ( .A1(n6320), .A2(n6319), .ZN(n9801) );
  INV_X1 U6497 ( .A(n5470), .ZN(n9803) );
  AND2_X1 U6498 ( .A1(n5881), .A2(n5638), .ZN(n5471) );
  AND2_X1 U6499 ( .A1(n6337), .A2(n5472), .ZN(n6393) );
  NAND2_X1 U6500 ( .A1(n6337), .A2(n5473), .ZN(n9776) );
  NAND2_X1 U6501 ( .A1(n7570), .A2(n6272), .ZN(n7806) );
  AOI21_X1 U6502 ( .B1(n9877), .B2(n6311), .A(n6310), .ZN(n9861) );
  NAND2_X1 U6503 ( .A1(n6290), .A2(n8981), .ZN(n8977) );
  OAI22_X1 U6504 ( .A1(n8011), .A2(n6281), .B1(n9648), .B2(n8010), .ZN(n7999)
         );
  NAND2_X1 U6505 ( .A1(n10491), .A2(n10493), .ZN(n10490) );
  NAND2_X1 U6506 ( .A1(n7630), .A2(n7629), .ZN(n7139) );
  NAND2_X1 U6507 ( .A1(n10472), .A2(n10471), .ZN(n10470) );
  NOR2_X1 U6508 ( .A1(n10584), .A2(n7163), .ZN(n10553) );
  MUX2_X1 U6509 ( .A(n9365), .B(n9364), .S(n9449), .Z(n9373) );
  MUX2_X1 U6510 ( .A(n9330), .B(n9329), .S(n9449), .Z(n9332) );
  AOI211_X1 U6511 ( .C1(n9373), .C2(n9372), .A(n9371), .B(n9370), .ZN(n9379)
         );
  OAI21_X2 U6512 ( .B1(n5704), .B2(SI_2_), .A(n5706), .ZN(n5863) );
  NOR3_X1 U6513 ( .A1(n9398), .A2(n9393), .A3(n9927), .ZN(n9395) );
  OAI21_X2 U6514 ( .B1(n5714), .B2(SI_4_), .A(n5716), .ZN(n5895) );
  OR2_X1 U6515 ( .A1(n5845), .A2(n7296), .ZN(n5870) );
  MUX2_X1 U6516 ( .A(n7811), .B(P2_REG2_REG_2__SCAN_IN), .S(n7453), .Z(n10901)
         );
  NAND2_X1 U6517 ( .A1(n5822), .A2(n5488), .ZN(n5487) );
  NAND2_X1 U6518 ( .A1(n5491), .A2(n7089), .ZN(n7124) );
  NAND3_X1 U6519 ( .A1(n5693), .A2(n5692), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n5492) );
  NAND2_X1 U6520 ( .A1(n5694), .A2(n5492), .ZN(n5697) );
  NAND2_X1 U6521 ( .A1(n5931), .A2(n5930), .ZN(n5933) );
  NAND2_X1 U6522 ( .A1(n6099), .A2(n5504), .ZN(n5503) );
  NAND2_X1 U6523 ( .A1(n6099), .A2(n6098), .ZN(n5511) );
  NAND2_X1 U6524 ( .A1(n5999), .A2(n5516), .ZN(n5515) );
  NAND2_X1 U6525 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  NAND2_X1 U6526 ( .A1(n5519), .A2(n5522), .ZN(n5796) );
  NAND2_X1 U6527 ( .A1(n6204), .A2(n5520), .ZN(n5519) );
  NAND2_X1 U6528 ( .A1(n6205), .A2(n5788), .ZN(n6218) );
  OAI21_X1 U6529 ( .B1(n9154), .B2(n7160), .A(n5537), .ZN(n9221) );
  NAND2_X1 U6530 ( .A1(n5536), .A2(n5534), .ZN(n10408) );
  NAND2_X1 U6531 ( .A1(n9154), .A2(n5537), .ZN(n5536) );
  NAND2_X1 U6532 ( .A1(n8124), .A2(n5542), .ZN(n5541) );
  INV_X1 U6533 ( .A(n10534), .ZN(n5545) );
  NAND2_X1 U6534 ( .A1(n5553), .A2(n5551), .ZN(n9008) );
  NAND2_X1 U6535 ( .A1(n7922), .A2(n7923), .ZN(n5555) );
  NAND2_X1 U6536 ( .A1(n7921), .A2(n5554), .ZN(n5556) );
  NOR2_X1 U6537 ( .A1(n5557), .A2(n5558), .ZN(n5554) );
  NAND3_X1 U6538 ( .A1(n5556), .A2(n7924), .A3(n5555), .ZN(n7948) );
  NAND2_X1 U6539 ( .A1(n8706), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U6540 ( .A1(n8707), .A2(n8713), .ZN(n8706) );
  OAI21_X2 U6541 ( .B1(n10568), .B2(n10576), .A(n10412), .ZN(n10550) );
  OR2_X1 U6542 ( .A1(n10461), .A2(n10471), .ZN(n5562) );
  NAND2_X1 U6543 ( .A1(n6403), .A2(n5679), .ZN(n6418) );
  OAI21_X2 U6544 ( .B1(n9578), .B2(n5569), .A(n5566), .ZN(n9622) );
  NAND2_X1 U6545 ( .A1(n5145), .A2(n7416), .ZN(n7469) );
  NAND2_X1 U6546 ( .A1(n9201), .A2(n5122), .ZN(n5575) );
  NAND2_X1 U6547 ( .A1(n9589), .A2(n9490), .ZN(n5578) );
  NAND2_X1 U6548 ( .A1(n5583), .A2(n9575), .ZN(n9502) );
  NAND2_X1 U6549 ( .A1(n9509), .A2(n5585), .ZN(n5584) );
  OAI211_X1 U6550 ( .C1(n9509), .C2(n5591), .A(n5586), .B(n5584), .ZN(n9520)
         );
  NAND2_X1 U6551 ( .A1(n9509), .A2(n9620), .ZN(n9523) );
  OAI21_X1 U6552 ( .B1(n8965), .B2(n5598), .A(n5595), .ZN(n5594) );
  NAND2_X1 U6553 ( .A1(n5607), .A2(n5605), .ZN(n7582) );
  NAND2_X1 U6554 ( .A1(n7579), .A2(n5606), .ZN(n5605) );
  NAND2_X1 U6555 ( .A1(n7965), .A2(n5120), .ZN(n5616) );
  AND2_X1 U6556 ( .A1(n7966), .A2(n9648), .ZN(n5619) );
  NOR2_X2 U6557 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5854) );
  NAND2_X1 U6558 ( .A1(n5854), .A2(n5488), .ZN(n5867) );
  OAI21_X1 U6559 ( .B1(n5621), .B2(n5622), .A(n7860), .ZN(n5620) );
  AOI21_X1 U6560 ( .B1(n9275), .B2(n5626), .A(n5625), .ZN(n5624) );
  NAND2_X1 U6561 ( .A1(n5633), .A2(n5634), .ZN(n9887) );
  NAND2_X1 U6562 ( .A1(n9909), .A2(n6148), .ZN(n5633) );
  NAND2_X1 U6563 ( .A1(n5636), .A2(n5173), .ZN(n9925) );
  NAND2_X1 U6564 ( .A1(n5636), .A2(n9392), .ZN(n9924) );
  NAND2_X1 U6565 ( .A1(n8009), .A2(n5637), .ZN(n7995) );
  NAND2_X1 U6566 ( .A1(n6113), .A2(n5640), .ZN(n6345) );
  NAND2_X1 U6567 ( .A1(n10133), .A2(n10134), .ZN(n10132) );
  INV_X1 U6568 ( .A(n6592), .ZN(n8696) );
  NAND2_X1 U6569 ( .A1(n6482), .A2(n5671), .ZN(n7653) );
  NAND2_X1 U6570 ( .A1(n5673), .A2(n6806), .ZN(n10117) );
  NAND2_X1 U6571 ( .A1(n6435), .A2(n5676), .ZN(n6433) );
  NAND2_X1 U6572 ( .A1(n6435), .A2(n5178), .ZN(n6425) );
  NAND2_X1 U6573 ( .A1(n6113), .A2(n6341), .ZN(n6370) );
  AND2_X1 U6574 ( .A1(P2_U3893), .A2(n7359), .ZN(n10996) );
  NAND2_X1 U6575 ( .A1(n7182), .A2(n7096), .ZN(n7097) );
  NAND2_X1 U6576 ( .A1(n6269), .A2(n6270), .ZN(n7570) );
  OAI21_X1 U6577 ( .B1(n10221), .B2(n10220), .A(n10219), .ZN(n10224) );
  NOR2_X1 U6578 ( .A1(n7597), .A2(n6947), .ZN(n6962) );
  INV_X1 U6579 ( .A(n6947), .ZN(n8824) );
  AND2_X1 U6580 ( .A1(n6444), .A2(n6947), .ZN(n7599) );
  AND2_X4 U6581 ( .A1(n7594), .A2(n6471), .ZN(n6489) );
  OR3_X1 U6582 ( .A1(n9630), .A2(n9831), .A3(n9449), .ZN(n5677) );
  AND2_X1 U6583 ( .A1(n6377), .A2(n6376), .ZN(n5678) );
  AND2_X2 U6584 ( .A1(n6373), .A2(n7425), .ZN(n11108) );
  INV_X1 U6585 ( .A(n10063), .ZN(n6374) );
  AND4_X1 U6586 ( .A1(n6123), .A2(n6122), .A3(n6121), .A4(n6120), .ZN(n9906)
         );
  AOI21_X1 U6587 ( .B1(n10075), .B2(n9266), .A(n6249), .ZN(n6390) );
  AND4_X1 U6588 ( .A1(n6136), .A2(n6135), .A3(n6134), .A4(n6133), .ZN(n6307)
         );
  OR2_X1 U6589 ( .A1(n6627), .A2(n6626), .ZN(n5680) );
  NOR2_X1 U6590 ( .A1(n6633), .A2(n6453), .ZN(n5681) );
  INV_X1 U6591 ( .A(n9458), .ZN(n9459) );
  AND2_X1 U6592 ( .A1(n6324), .A2(n6365), .ZN(n9951) );
  OR2_X1 U6593 ( .A1(n7187), .A2(n8920), .ZN(n5684) );
  INV_X1 U6594 ( .A(n9862), .ZN(n9639) );
  AND4_X1 U6595 ( .A1(n6187), .A2(n6186), .A3(n6185), .A4(n6184), .ZN(n9862)
         );
  INV_X1 U6596 ( .A(n8954), .ZN(n9175) );
  OR2_X1 U6597 ( .A1(n8854), .A2(n10246), .ZN(n5685) );
  AND2_X1 U6598 ( .A1(n8606), .A2(n8605), .ZN(n5686) );
  AND4_X1 U6599 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n9366)
         );
  INV_X1 U6600 ( .A(n9366), .ZN(n8994) );
  OR2_X1 U6601 ( .A1(n8909), .A2(n8908), .ZN(n5687) );
  NAND2_X1 U6602 ( .A1(n8041), .A2(n10435), .ZN(n10601) );
  INV_X2 U6603 ( .A(n10601), .ZN(n10596) );
  AND2_X1 U6604 ( .A1(n6436), .A2(n6437), .ZN(n5688) );
  INV_X1 U6605 ( .A(n7197), .ZN(n7014) );
  AND2_X1 U6606 ( .A1(n10403), .A2(n10402), .ZN(n7175) );
  INV_X1 U6607 ( .A(n9437), .ZN(n9438) );
  INV_X1 U6608 ( .A(n7096), .ZN(n7095) );
  INV_X1 U6609 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U6610 ( .A1(n9303), .A2(n9302), .ZN(n9306) );
  INV_X1 U6611 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U6612 ( .A1(n7098), .A2(n7097), .ZN(n7099) );
  INV_X1 U6613 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6400) );
  INV_X1 U6614 ( .A(n10921), .ZN(n10922) );
  INV_X1 U6615 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7749) );
  INV_X1 U6616 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9165) );
  INV_X1 U6617 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9537) );
  INV_X1 U6618 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8943) );
  AND2_X1 U6619 ( .A1(n6340), .A2(n5604), .ZN(n6341) );
  INV_X1 U6620 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5986) );
  INV_X1 U6621 ( .A(n10535), .ZN(n10414) );
  INV_X1 U6622 ( .A(n10684), .ZN(n10378) );
  INV_X1 U6623 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6420) );
  INV_X1 U6624 ( .A(SI_16_), .ZN(n8361) );
  INV_X1 U6625 ( .A(SI_11_), .ZN(n8172) );
  INV_X1 U6626 ( .A(n9513), .ZN(n9510) );
  INV_X1 U6627 ( .A(n9590), .ZN(n9489) );
  INV_X1 U6628 ( .A(n9626), .ZN(n9615) );
  NOR2_X1 U6629 ( .A1(n6072), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6089) );
  NOR2_X1 U6630 ( .A1(n6236), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6235) );
  OR2_X1 U6631 ( .A1(n6222), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6236) );
  NOR2_X1 U6632 ( .A1(n6182), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6193) );
  AND2_X1 U6633 ( .A1(n6142), .A2(n9591), .ZN(n6156) );
  NOR2_X1 U6634 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n6118), .ZN(n6130) );
  NAND2_X1 U6635 ( .A1(n6022), .A2(n8943), .ZN(n6042) );
  AND2_X1 U6636 ( .A1(n9338), .A2(n9341), .ZN(n9281) );
  OR2_X1 U6637 ( .A1(n6000), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6037) );
  INV_X1 U6638 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6464) );
  AND2_X1 U6639 ( .A1(n6875), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6889) );
  INV_X1 U6640 ( .A(n6951), .ZN(n6963) );
  INV_X1 U6641 ( .A(n10791), .ZN(n6452) );
  AND2_X1 U6642 ( .A1(n6877), .A2(n6861), .ZN(n10508) );
  NOR2_X1 U6643 ( .A1(n10804), .A2(n6941), .ZN(n7610) );
  INV_X1 U6644 ( .A(SI_9_), .ZN(n8176) );
  NOR2_X1 U6645 ( .A1(n5940), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5939) );
  OR2_X1 U6646 ( .A1(n8016), .A2(n9647), .ZN(n8017) );
  AND2_X1 U6647 ( .A1(n9503), .A2(n9501), .ZN(n9576) );
  OR3_X1 U6648 ( .A1(n9323), .A2(n9459), .A3(n6365), .ZN(n7418) );
  OR2_X1 U6649 ( .A1(n7431), .A2(n7430), .ZN(n9626) );
  OR2_X1 U6650 ( .A1(n6237), .A2(n9822), .ZN(n6225) );
  INV_X1 U6651 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8211) );
  NOR2_X1 U6652 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  NAND2_X1 U6653 ( .A1(n5815), .A2(n5814), .ZN(n6327) );
  NAND2_X1 U6654 ( .A1(n9787), .A2(n9936), .ZN(n9788) );
  INV_X1 U6655 ( .A(n9900), .ZN(n9891) );
  NAND2_X2 U6656 ( .A1(n9323), .A2(n9465), .ZN(n9449) );
  NAND2_X1 U6657 ( .A1(n9147), .A2(n6056), .ZN(n6072) );
  AND2_X1 U6658 ( .A1(n7425), .A2(n10022), .ZN(n7733) );
  AND2_X1 U6659 ( .A1(n5422), .A2(n6384), .ZN(n7741) );
  OR2_X1 U6660 ( .A1(n7726), .A2(n7728), .ZN(n6382) );
  OR2_X1 U6661 ( .A1(n9304), .A2(n9257), .ZN(n9262) );
  INV_X1 U6662 ( .A(n9640), .ZN(n9953) );
  NOR2_X1 U6663 ( .A1(n7741), .A2(n6267), .ZN(n8840) );
  OR2_X1 U6664 ( .A1(n6037), .A2(n6036), .ZN(n6051) );
  NAND2_X1 U6665 ( .A1(n6944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6945) );
  NOR2_X1 U6666 ( .A1(n6690), .A2(n6689), .ZN(n6706) );
  OR2_X1 U6667 ( .A1(n6654), .A2(n6653), .ZN(n6667) );
  OR2_X1 U6668 ( .A1(n6723), .A2(n6722), .ZN(n6739) );
  NOR2_X1 U6669 ( .A1(n6739), .A2(n6738), .ZN(n6758) );
  NAND2_X1 U6670 ( .A1(n10195), .A2(n10196), .ZN(n10194) );
  NAND2_X1 U6671 ( .A1(n6960), .A2(n10271), .ZN(n10236) );
  OR2_X1 U6672 ( .A1(n7528), .A2(n7497), .ZN(n7514) );
  INV_X1 U6673 ( .A(n8073), .ZN(n8065) );
  OR2_X1 U6674 ( .A1(n7331), .A2(n7330), .ZN(n7396) );
  INV_X1 U6675 ( .A(n10476), .ZN(n10479) );
  INV_X1 U6676 ( .A(n10658), .ZN(n10559) );
  INV_X1 U6677 ( .A(n10719), .ZN(n10703) );
  INV_X1 U6678 ( .A(n10247), .ZN(n8727) );
  OR2_X1 U6679 ( .A1(n10596), .A2(n10667), .ZN(n10540) );
  NAND2_X1 U6680 ( .A1(n7013), .A2(n7194), .ZN(n7632) );
  NAND2_X1 U6681 ( .A1(n6838), .A2(n6837), .ZN(n7070) );
  NAND2_X1 U6682 ( .A1(n7599), .A2(n7598), .ZN(n10702) );
  OR2_X1 U6683 ( .A1(n7096), .A2(n7603), .ZN(n7597) );
  NOR2_X1 U6684 ( .A1(n7610), .A2(n7609), .ZN(n8040) );
  INV_X1 U6685 ( .A(n5862), .ZN(n5864) );
  INV_X1 U6686 ( .A(n9623), .ZN(n9606) );
  AND4_X1 U6687 ( .A1(n9255), .A2(n9254), .A3(n9253), .A4(n9252), .ZN(n9304)
         );
  AND4_X1 U6688 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(n9548)
         );
  AND4_X1 U6689 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n8836)
         );
  NAND4_X2 U6690 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n6273)
         );
  INV_X1 U6691 ( .A(n11008), .ZN(n10983) );
  XNOR2_X1 U6692 ( .A(n9699), .B(n9711), .ZN(n9682) );
  XNOR2_X1 U6693 ( .A(n9744), .B(n9764), .ZN(n9725) );
  INV_X1 U6694 ( .A(n10940), .ZN(n10999) );
  NAND2_X1 U6695 ( .A1(n7733), .A2(n7734), .ZN(n9957) );
  AND2_X1 U6696 ( .A1(n11071), .A2(n11059), .ZN(n9943) );
  INV_X1 U6697 ( .A(n9957), .ZN(n11066) );
  AND2_X1 U6698 ( .A1(n7730), .A2(n6386), .ZN(n6387) );
  NOR2_X1 U6699 ( .A1(n9026), .A2(n9465), .ZN(n7833) );
  OR2_X1 U6700 ( .A1(n8840), .A2(n7833), .ZN(n10025) );
  INV_X1 U6701 ( .A(n10027), .ZN(n10022) );
  AND2_X1 U6702 ( .A1(n6100), .A2(n6085), .ZN(n9714) );
  AND2_X1 U6703 ( .A1(n6860), .A2(n6843), .ZN(n10522) );
  AND2_X1 U6704 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6559) );
  INV_X1 U6705 ( .A(n7249), .ZN(n7250) );
  AND4_X1 U6706 ( .A1(n6957), .A2(n6956), .A3(n6955), .A4(n6954), .ZN(n10626)
         );
  AND3_X1 U6707 ( .A1(n6781), .A2(n6780), .A3(n6779), .ZN(n10209) );
  AND2_X1 U6708 ( .A1(n7514), .A2(n7513), .ZN(n7516) );
  INV_X1 U6709 ( .A(n10591), .ZN(n10542) );
  AND2_X1 U6710 ( .A1(n7106), .A2(n10554), .ZN(n10576) );
  INV_X1 U6711 ( .A(n9078), .ZN(n9080) );
  INV_X1 U6712 ( .A(n10548), .ZN(n10473) );
  INV_X1 U6713 ( .A(n7978), .ZN(n7984) );
  INV_X1 U6714 ( .A(n10702), .ZN(n10732) );
  INV_X1 U6715 ( .A(n11050), .ZN(n10594) );
  INV_X1 U6716 ( .A(n11088), .ZN(n10707) );
  NAND2_X1 U6717 ( .A1(n8094), .A2(n7597), .ZN(n11091) );
  NAND2_X1 U6718 ( .A1(n6931), .A2(n10797), .ZN(n10804) );
  INV_X1 U6719 ( .A(n10792), .ZN(n10796) );
  AND2_X1 U6720 ( .A1(n7412), .A2(n7411), .ZN(n9623) );
  NAND2_X1 U6721 ( .A1(n7422), .A2(n7421), .ZN(n9632) );
  INV_X1 U6722 ( .A(n9819), .ZN(n9786) );
  INV_X1 U6723 ( .A(n6307), .ZN(n9919) );
  OR2_X1 U6724 ( .A1(P2_U3150), .A2(n7352), .ZN(n10940) );
  NAND2_X1 U6725 ( .A1(n10895), .A2(n9756), .ZN(n11011) );
  INV_X1 U6726 ( .A(n9946), .ZN(n11069) );
  INV_X1 U6727 ( .A(n11071), .ZN(n9946) );
  NAND2_X1 U6728 ( .A1(n7742), .A2(n9957), .ZN(n11071) );
  INV_X1 U6729 ( .A(n9943), .ZN(n9963) );
  NAND2_X1 U6730 ( .A1(n10033), .A2(n10022), .ZN(n10008) );
  NAND2_X1 U6731 ( .A1(n9969), .A2(n9968), .ZN(n10036) );
  NAND2_X1 U6732 ( .A1(n11108), .A2(n10022), .ZN(n10063) );
  INV_X1 U6733 ( .A(n11108), .ZN(n11105) );
  AND2_X1 U6734 ( .A1(n7405), .A2(n7305), .ZN(n7425) );
  INV_X1 U6735 ( .A(n9754), .ZN(n9762) );
  INV_X1 U6736 ( .A(n9714), .ZN(n9736) );
  INV_X1 U6737 ( .A(n9133), .ZN(n10077) );
  INV_X1 U6738 ( .A(n10367), .ZN(n10265) );
  INV_X1 U6739 ( .A(n8564), .ZN(n8781) );
  OR3_X1 U6740 ( .A1(n10173), .A2(n10176), .A3(n10243), .ZN(n10183) );
  INV_X1 U6741 ( .A(n10215), .ZN(n10237) );
  AND4_X1 U6742 ( .A1(n6999), .A2(n6998), .A3(n6997), .A4(n6996), .ZN(n10450)
         );
  INV_X1 U6743 ( .A(n10644), .ZN(n10659) );
  INV_X1 U6744 ( .A(n10179), .ZN(n10720) );
  INV_X1 U6745 ( .A(n8121), .ZN(n10249) );
  OR2_X1 U6746 ( .A1(n10596), .A2(n8100), .ZN(n10599) );
  OR2_X1 U6747 ( .A1(n10596), .A2(n8096), .ZN(n10603) );
  NAND2_X1 U6748 ( .A1(n11094), .A2(n10707), .ZN(n10693) );
  INV_X1 U6749 ( .A(n11094), .ZN(n11093) );
  INV_X1 U6750 ( .A(n10487), .ZN(n10758) );
  NAND2_X1 U6751 ( .A1(n11079), .A2(n10707), .ZN(n10777) );
  NAND2_X1 U6752 ( .A1(n7793), .A2(n8039), .ZN(n11095) );
  AND2_X2 U6753 ( .A1(n10804), .A2(n10803), .ZN(n10835) );
  CLKBUF_X1 U6754 ( .A(n9234), .Z(n10799) );
  INV_X2 U6755 ( .A(n11001), .ZN(P2_U3893) );
  AND2_X2 U6756 ( .A1(n7280), .A2(n7325), .ZN(P1_U3973) );
  NAND2_X1 U6757 ( .A1(n5690), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5691) );
  NAND2_X2 U6758 ( .A1(n5691), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5692) );
  INV_X1 U6759 ( .A(SI_1_), .ZN(n5695) );
  NAND2_X1 U6760 ( .A1(n5696), .A2(n5695), .ZN(n5698) );
  NAND2_X1 U6761 ( .A1(n5697), .A2(SI_1_), .ZN(n5702) );
  NAND2_X1 U6762 ( .A1(n5698), .A2(n5702), .ZN(n5848) );
  INV_X1 U6763 ( .A(n5848), .ZN(n5701) );
  INV_X1 U6764 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5699) );
  INV_X1 U6765 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5841) );
  MUX2_X1 U6766 ( .A(n5699), .B(n5841), .S(n5816), .Z(n5700) );
  INV_X1 U6767 ( .A(SI_0_), .ZN(n6475) );
  NAND2_X1 U6768 ( .A1(n5701), .A2(n5846), .ZN(n5850) );
  NAND2_X1 U6769 ( .A1(n5850), .A2(n5702), .ZN(n5862) );
  MUX2_X1 U6770 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5703), .Z(n5704) );
  NAND2_X1 U6771 ( .A1(n5704), .A2(SI_2_), .ZN(n5706) );
  INV_X1 U6772 ( .A(n5863), .ZN(n5705) );
  NAND2_X1 U6773 ( .A1(n5862), .A2(n5705), .ZN(n5865) );
  NAND2_X1 U6774 ( .A1(n5865), .A2(n5706), .ZN(n5876) );
  INV_X1 U6775 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5707) );
  OR2_X1 U6776 ( .A1(n5816), .A2(n5707), .ZN(n5708) );
  INV_X1 U6777 ( .A(n5711), .ZN(n5710) );
  INV_X1 U6778 ( .A(SI_3_), .ZN(n8379) );
  NAND2_X1 U6779 ( .A1(n5710), .A2(n8379), .ZN(n5712) );
  NAND2_X1 U6780 ( .A1(n5711), .A2(SI_3_), .ZN(n5713) );
  AND2_X2 U6781 ( .A1(n5712), .A2(n5713), .ZN(n5875) );
  NAND2_X1 U6782 ( .A1(n5878), .A2(n5713), .ZN(n5896) );
  MUX2_X1 U6783 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7287), .Z(n5714) );
  NAND2_X1 U6784 ( .A1(n5714), .A2(SI_4_), .ZN(n5716) );
  INV_X1 U6785 ( .A(n5895), .ZN(n5715) );
  NAND2_X1 U6786 ( .A1(n5896), .A2(n5715), .ZN(n5717) );
  NAND2_X1 U6787 ( .A1(n5717), .A2(n5716), .ZN(n5908) );
  MUX2_X1 U6788 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7287), .Z(n5718) );
  NAND2_X1 U6789 ( .A1(n5718), .A2(SI_5_), .ZN(n5721) );
  INV_X1 U6790 ( .A(n5718), .ZN(n5719) );
  INV_X1 U6791 ( .A(SI_5_), .ZN(n8378) );
  NAND2_X1 U6792 ( .A1(n5719), .A2(n8378), .ZN(n5720) );
  AND2_X1 U6793 ( .A1(n5721), .A2(n5720), .ZN(n5907) );
  NAND2_X1 U6794 ( .A1(n5908), .A2(n5907), .ZN(n5910) );
  NAND2_X1 U6795 ( .A1(n5910), .A2(n5721), .ZN(n5916) );
  MUX2_X1 U6796 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7287), .Z(n5722) );
  NAND2_X1 U6797 ( .A1(n5722), .A2(SI_6_), .ZN(n5726) );
  INV_X1 U6798 ( .A(n5722), .ZN(n5724) );
  INV_X1 U6799 ( .A(SI_6_), .ZN(n5723) );
  NAND2_X1 U6800 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  NAND2_X1 U6801 ( .A1(n5916), .A2(n5915), .ZN(n5918) );
  MUX2_X1 U6802 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7287), .Z(n5727) );
  INV_X1 U6803 ( .A(n5727), .ZN(n5728) );
  INV_X1 U6804 ( .A(SI_7_), .ZN(n8374) );
  NAND2_X1 U6805 ( .A1(n5728), .A2(n8374), .ZN(n5729) );
  INV_X1 U6806 ( .A(n5731), .ZN(n5733) );
  INV_X1 U6807 ( .A(SI_8_), .ZN(n5732) );
  MUX2_X1 U6808 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n7287), .Z(n5734) );
  XNOR2_X1 U6809 ( .A(n5734), .B(n8176), .ZN(n5962) );
  MUX2_X1 U6810 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7287), .Z(n5735) );
  NAND2_X1 U6811 ( .A1(n5735), .A2(SI_10_), .ZN(n5740) );
  INV_X1 U6812 ( .A(n5735), .ZN(n5737) );
  INV_X1 U6813 ( .A(SI_10_), .ZN(n5736) );
  NAND2_X1 U6814 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  NAND2_X1 U6815 ( .A1(n5740), .A2(n5738), .ZN(n5983) );
  INV_X1 U6816 ( .A(n5983), .ZN(n5739) );
  NAND2_X1 U6817 ( .A1(n5985), .A2(n5740), .ZN(n5999) );
  MUX2_X1 U6818 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7287), .Z(n5741) );
  XNOR2_X1 U6819 ( .A(n5741), .B(SI_11_), .ZN(n5998) );
  INV_X1 U6820 ( .A(n5741), .ZN(n5742) );
  NAND2_X1 U6821 ( .A1(n5742), .A2(n8172), .ZN(n5743) );
  MUX2_X1 U6822 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7287), .Z(n5744) );
  NAND2_X1 U6823 ( .A1(n5744), .A2(SI_12_), .ZN(n5745) );
  OAI21_X1 U6824 ( .B1(n5744), .B2(SI_12_), .A(n5745), .ZN(n6014) );
  MUX2_X1 U6825 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7287), .Z(n5746) );
  NAND2_X1 U6826 ( .A1(n5746), .A2(SI_13_), .ZN(n5749) );
  INV_X1 U6827 ( .A(n5746), .ZN(n5747) );
  NAND2_X1 U6828 ( .A1(n5747), .A2(n8164), .ZN(n5748) );
  MUX2_X1 U6829 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7287), .Z(n5750) );
  XNOR2_X1 U6830 ( .A(n5750), .B(SI_14_), .ZN(n6049) );
  INV_X1 U6831 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U6832 ( .A1(n5751), .A2(n8160), .ZN(n5752) );
  MUX2_X1 U6833 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7287), .Z(n5753) );
  OAI21_X1 U6834 ( .B1(n5753), .B2(SI_15_), .A(n5754), .ZN(n6063) );
  MUX2_X1 U6835 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7287), .Z(n5755) );
  XNOR2_X1 U6836 ( .A(n5755), .B(SI_16_), .ZN(n6078) );
  INV_X1 U6837 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U6838 ( .A1(n5756), .A2(n8361), .ZN(n5757) );
  MUX2_X1 U6839 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n7287), .Z(n5759) );
  NOR2_X1 U6840 ( .A1(n5759), .A2(SI_17_), .ZN(n5760) );
  MUX2_X1 U6841 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7287), .Z(n5761) );
  NAND2_X1 U6842 ( .A1(n5761), .A2(SI_18_), .ZN(n5764) );
  INV_X1 U6843 ( .A(n5761), .ZN(n5762) );
  NAND2_X1 U6844 ( .A1(n5762), .A2(n8159), .ZN(n5763) );
  NAND2_X1 U6845 ( .A1(n5764), .A2(n5763), .ZN(n6110) );
  MUX2_X1 U6846 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7287), .Z(n5765) );
  XNOR2_X1 U6847 ( .A(n5765), .B(SI_19_), .ZN(n6124) );
  INV_X1 U6848 ( .A(n5765), .ZN(n5766) );
  NAND2_X1 U6849 ( .A1(n5766), .A2(n8155), .ZN(n5767) );
  MUX2_X1 U6850 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7287), .Z(n5768) );
  XNOR2_X1 U6851 ( .A(n5768), .B(n8354), .ZN(n6138) );
  NOR2_X1 U6852 ( .A1(n5768), .A2(SI_20_), .ZN(n5769) );
  AOI21_X2 U6853 ( .B1(n6137), .B2(n6138), .A(n5769), .ZN(n6149) );
  MUX2_X1 U6854 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7287), .Z(n5770) );
  NAND2_X1 U6855 ( .A1(n5770), .A2(SI_21_), .ZN(n5774) );
  INV_X1 U6856 ( .A(n5770), .ZN(n5771) );
  NAND2_X1 U6857 ( .A1(n5771), .A2(n8347), .ZN(n5772) );
  NAND2_X1 U6858 ( .A1(n5774), .A2(n5772), .ZN(n6150) );
  INV_X1 U6859 ( .A(n6150), .ZN(n5773) );
  NAND2_X1 U6860 ( .A1(n6149), .A2(n5773), .ZN(n6153) );
  NAND2_X1 U6861 ( .A1(n6153), .A2(n5774), .ZN(n5776) );
  MUX2_X1 U6862 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7287), .Z(n5775) );
  NAND2_X1 U6863 ( .A1(n5776), .A2(n5775), .ZN(n5778) );
  MUX2_X1 U6864 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n7287), .Z(n5779) );
  XNOR2_X1 U6865 ( .A(n5779), .B(SI_23_), .ZN(n6176) );
  INV_X1 U6866 ( .A(n5779), .ZN(n5780) );
  INV_X1 U6867 ( .A(SI_23_), .ZN(n8348) );
  NAND2_X1 U6868 ( .A1(n5780), .A2(n8348), .ZN(n5781) );
  MUX2_X1 U6869 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7287), .Z(n5783) );
  INV_X1 U6870 ( .A(SI_24_), .ZN(n5782) );
  XNOR2_X1 U6871 ( .A(n5783), .B(n5782), .ZN(n6189) );
  NOR2_X1 U6872 ( .A1(n5783), .A2(SI_24_), .ZN(n5784) );
  MUX2_X1 U6873 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n7287), .Z(n5785) );
  NAND2_X1 U6874 ( .A1(n5785), .A2(SI_25_), .ZN(n5788) );
  INV_X1 U6875 ( .A(n5785), .ZN(n5786) );
  INV_X1 U6876 ( .A(SI_25_), .ZN(n8147) );
  NAND2_X1 U6877 ( .A1(n5786), .A2(n8147), .ZN(n5787) );
  MUX2_X1 U6878 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n7287), .Z(n5789) );
  XNOR2_X1 U6879 ( .A(n5789), .B(SI_26_), .ZN(n6217) );
  INV_X1 U6880 ( .A(n5789), .ZN(n5790) );
  INV_X1 U6881 ( .A(SI_26_), .ZN(n8143) );
  NAND2_X1 U6882 ( .A1(n5790), .A2(n8143), .ZN(n5791) );
  MUX2_X1 U6883 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7287), .Z(n5792) );
  INV_X1 U6884 ( .A(SI_27_), .ZN(n5793) );
  XNOR2_X1 U6885 ( .A(n5792), .B(n5793), .ZN(n6231) );
  INV_X1 U6886 ( .A(n5792), .ZN(n5794) );
  NAND2_X1 U6887 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  NAND2_X1 U6888 ( .A1(n5796), .A2(n5795), .ZN(n6243) );
  MUX2_X1 U6889 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7287), .Z(n6244) );
  INV_X1 U6890 ( .A(SI_28_), .ZN(n8138) );
  XNOR2_X1 U6891 ( .A(n6244), .B(n8138), .ZN(n6242) );
  NOR2_X1 U6892 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5800) );
  NAND4_X1 U6893 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .ZN(n5804)
         );
  NAND3_X1 U6894 ( .A1(n5964), .A2(n5802), .A3(n5801), .ZN(n5803) );
  NOR2_X2 U6895 ( .A1(n5867), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5881) );
  NOR2_X1 U6896 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5808) );
  NOR2_X1 U6897 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5807) );
  NOR2_X1 U6898 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5806) );
  XNOR2_X2 U6899 ( .A(n5812), .B(n5811), .ZN(n7359) );
  NAND2_X1 U6900 ( .A1(n6348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5813) );
  NAND2_X2 U6901 ( .A1(n5852), .A2(n5392), .ZN(n5851) );
  NAND2_X1 U6902 ( .A1(n9471), .A2(n9266), .ZN(n5820) );
  INV_X1 U6903 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5818) );
  OR2_X1 U6904 ( .A1(n9267), .A2(n5818), .ZN(n5819) );
  INV_X1 U6905 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U6906 ( .A1(n6330), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5836) );
  INV_X1 U6907 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5827) );
  OR2_X1 U6908 ( .A1(n9249), .A2(n5827), .ZN(n5835) );
  INV_X1 U6909 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8204) );
  INV_X1 U6910 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9213) );
  NOR2_X1 U6911 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5887) );
  NAND2_X1 U6912 ( .A1(n5887), .A2(n8211), .ZN(n5923) );
  NAND2_X1 U6913 ( .A1(n5954), .A2(n8419), .ZN(n5991) );
  INV_X1 U6914 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9581) );
  INV_X1 U6915 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U6916 ( .A1(n8204), .A2(n6235), .ZN(n9260) );
  INV_X1 U6917 ( .A(n6235), .ZN(n5830) );
  NAND2_X1 U6918 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n5830), .ZN(n5831) );
  OR2_X1 U6919 ( .A1(n6237), .A2(n9792), .ZN(n5834) );
  INV_X1 U6920 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9793) );
  OR2_X1 U6921 ( .A1(n9251), .A2(n9793), .ZN(n5833) );
  INV_X1 U6922 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U6923 ( .A1(n5899), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5839) );
  INV_X1 U6924 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7358) );
  OR2_X1 U6925 ( .A1(n5889), .A2(n7358), .ZN(n5838) );
  INV_X1 U6926 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7357) );
  OR2_X1 U6927 ( .A1(n6181), .A2(n7357), .ZN(n5837) );
  INV_X1 U6928 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U6929 ( .A1(n5392), .A2(SI_0_), .ZN(n5842) );
  XNOR2_X1 U6930 ( .A(n5842), .B(n5841), .ZN(n10089) );
  MUX2_X1 U6931 ( .A(n7347), .B(n10089), .S(n5852), .Z(n7747) );
  INV_X1 U6932 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7859) );
  INV_X1 U6933 ( .A(n6181), .ZN(n5843) );
  INV_X1 U6934 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7344) );
  NAND2_X1 U6935 ( .A1(n5899), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5844) );
  INV_X1 U6936 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7289) );
  INV_X1 U6937 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U6938 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  NAND2_X1 U6939 ( .A1(n5850), .A2(n5849), .ZN(n7288) );
  NAND2_X1 U6940 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5853) );
  MUX2_X1 U6941 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5853), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5855) );
  INV_X1 U6942 ( .A(n7449), .ZN(n7342) );
  INV_X1 U6943 ( .A(n7441), .ZN(n7356) );
  NAND2_X1 U6944 ( .A1(n5879), .A2(n7356), .ZN(n5856) );
  NAND2_X1 U6945 ( .A1(n7566), .A2(n9326), .ZN(n7803) );
  NAND2_X1 U6946 ( .A1(n5899), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5861) );
  INV_X1 U6947 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10902) );
  INV_X1 U6948 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7811) );
  OR2_X1 U6949 ( .A1(n5889), .A2(n7811), .ZN(n5859) );
  INV_X1 U6950 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5857) );
  OR2_X1 U6951 ( .A1(n6181), .A2(n5857), .ZN(n5858) );
  INV_X1 U6952 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7296) );
  NAND2_X1 U6953 ( .A1(n5864), .A2(n5863), .ZN(n5866) );
  NAND2_X1 U6954 ( .A1(n5866), .A2(n5865), .ZN(n7295) );
  OR2_X1 U6955 ( .A1(n5851), .A2(n7295), .ZN(n5869) );
  NAND2_X1 U6956 ( .A1(n5879), .A2(n7453), .ZN(n5868) );
  NAND2_X1 U6957 ( .A1(n6273), .A2(n7805), .ZN(n9319) );
  NAND2_X1 U6958 ( .A1(n7803), .A2(n5426), .ZN(n7802) );
  NAND2_X1 U6959 ( .A1(n7802), .A2(n9328), .ZN(n7642) );
  NAND2_X1 U6960 ( .A1(n6250), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5874) );
  OR2_X1 U6961 ( .A1(n6237), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5873) );
  INV_X1 U6962 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7736) );
  OR2_X1 U6963 ( .A1(n5889), .A2(n7736), .ZN(n5872) );
  INV_X1 U6964 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7446) );
  OR2_X1 U6965 ( .A1(n6181), .A2(n7446), .ZN(n5871) );
  NAND4_X1 U6966 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n9650)
         );
  OR2_X1 U6967 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  NAND2_X1 U6968 ( .A1(n5878), .A2(n5877), .ZN(n7298) );
  OR2_X1 U6969 ( .A1(n7298), .A2(n5851), .ZN(n5885) );
  OR2_X1 U6970 ( .A1(n9267), .A2(n5709), .ZN(n5884) );
  NAND2_X1 U6971 ( .A1(n5867), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5880) );
  MUX2_X1 U6972 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5880), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5882) );
  AND2_X1 U6973 ( .A1(n5882), .A2(n5969), .ZN(n7708) );
  NAND2_X1 U6974 ( .A1(n6127), .A2(n7708), .ZN(n5883) );
  NAND2_X1 U6975 ( .A1(n9650), .A2(n7648), .ZN(n9336) );
  NAND2_X1 U6976 ( .A1(n7642), .A2(n9279), .ZN(n7641) );
  NAND2_X1 U6977 ( .A1(n7641), .A2(n5424), .ZN(n7786) );
  NAND2_X1 U6978 ( .A1(n6330), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5894) );
  INV_X1 U6979 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5886) );
  OR2_X1 U6980 ( .A1(n9249), .A2(n5886), .ZN(n5893) );
  INV_X1 U6981 ( .A(n5887), .ZN(n5901) );
  NAND2_X1 U6982 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5888) );
  AND2_X1 U6983 ( .A1(n5901), .A2(n5888), .ZN(n7851) );
  OR2_X1 U6984 ( .A1(n6237), .A2(n7851), .ZN(n5892) );
  INV_X1 U6985 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5890) );
  OR2_X1 U6986 ( .A1(n9251), .A2(n5890), .ZN(n5891) );
  NAND4_X1 U6987 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n7644)
         );
  NAND2_X1 U6988 ( .A1(n5969), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5911) );
  AOI22_X1 U6989 ( .A1(n5817), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6127), .B2(
        n10934), .ZN(n5898) );
  XNOR2_X1 U6990 ( .A(n5896), .B(n5895), .ZN(n6548) );
  NAND2_X1 U6991 ( .A1(n6548), .A2(n9266), .ZN(n5897) );
  OR2_X1 U6992 ( .A1(n7644), .A2(n7852), .ZN(n9337) );
  NAND2_X1 U6993 ( .A1(n7644), .A2(n7852), .ZN(n9333) );
  NAND2_X1 U6994 ( .A1(n7786), .A2(n9331), .ZN(n7785) );
  NAND2_X1 U6995 ( .A1(n6250), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5906) );
  INV_X1 U6996 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5900) );
  OR2_X1 U6997 ( .A1(n6181), .A2(n5900), .ZN(n5905) );
  NAND2_X1 U6998 ( .A1(n5901), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5902) );
  AND2_X1 U6999 ( .A1(n5923), .A2(n5902), .ZN(n7583) );
  OR2_X1 U7000 ( .A1(n6237), .A2(n7583), .ZN(n5904) );
  INV_X1 U7001 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7869) );
  OR2_X1 U7002 ( .A1(n9251), .A2(n7869), .ZN(n5903) );
  NAND4_X1 U7003 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n9649)
         );
  OR2_X1 U7004 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  OR2_X1 U7005 ( .A1(n7300), .A2(n5851), .ZN(n5914) );
  NAND2_X1 U7006 ( .A1(n5911), .A2(n5965), .ZN(n5912) );
  NAND2_X1 U7007 ( .A1(n5912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5919) );
  XNOR2_X1 U7008 ( .A(n5919), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U7009 ( .A1(n5817), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6127), .B2(
        n10944), .ZN(n5913) );
  INV_X1 U7010 ( .A(n7826), .ZN(n7871) );
  NAND2_X1 U7011 ( .A1(n8013), .A2(n7871), .ZN(n9338) );
  NAND2_X1 U7012 ( .A1(n7826), .A2(n9649), .ZN(n9341) );
  OR2_X1 U7013 ( .A1(n5916), .A2(n5915), .ZN(n5917) );
  NAND2_X1 U7014 ( .A1(n5918), .A2(n5917), .ZN(n7309) );
  OR2_X1 U7015 ( .A1(n7309), .A2(n5851), .ZN(n5922) );
  NAND2_X1 U7016 ( .A1(n5919), .A2(n5966), .ZN(n5920) );
  NAND2_X1 U7017 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5935) );
  XNOR2_X1 U7018 ( .A(n5935), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7757) );
  AOI22_X1 U7019 ( .A1(n5817), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6127), .B2(
        n7757), .ZN(n5921) );
  NAND2_X1 U7020 ( .A1(n5922), .A2(n5921), .ZN(n8010) );
  NAND2_X1 U7021 ( .A1(n6250), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5929) );
  OR2_X1 U7022 ( .A1(n9247), .A2(n7749), .ZN(n5928) );
  NAND2_X1 U7023 ( .A1(n5923), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5924) );
  AND2_X1 U7024 ( .A1(n5940), .A2(n5924), .ZN(n8057) );
  OR2_X1 U7025 ( .A1(n6237), .A2(n8057), .ZN(n5927) );
  INV_X1 U7026 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5925) );
  OR2_X1 U7027 ( .A1(n9251), .A2(n5925), .ZN(n5926) );
  OR2_X1 U7028 ( .A1(n8010), .A2(n8001), .ZN(n9346) );
  NAND2_X1 U7029 ( .A1(n8010), .A2(n8001), .ZN(n9345) );
  NAND2_X1 U7030 ( .A1(n5933), .A2(n5932), .ZN(n7312) );
  OR2_X1 U7031 ( .A1(n7312), .A2(n5851), .ZN(n5938) );
  INV_X1 U7032 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7033 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  NAND2_X1 U7034 ( .A1(n5936), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7035 ( .A(n5949), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7766) );
  AOI22_X1 U7036 ( .A1(n5817), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6127), .B2(
        n7766), .ZN(n5937) );
  NAND2_X1 U7037 ( .A1(n5938), .A2(n5937), .ZN(n8570) );
  NAND2_X1 U7038 ( .A1(n6250), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5945) );
  INV_X1 U7039 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7765) );
  OR2_X1 U7040 ( .A1(n9251), .A2(n7765), .ZN(n5944) );
  INV_X1 U7041 ( .A(n5939), .ZN(n5955) );
  NAND2_X1 U7042 ( .A1(n5940), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5941) );
  AND2_X1 U7043 ( .A1(n5955), .A2(n5941), .ZN(n8571) );
  OR2_X1 U7044 ( .A1(n6237), .A2(n8571), .ZN(n5943) );
  INV_X1 U7045 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7764) );
  OR2_X1 U7046 ( .A1(n6181), .A2(n7764), .ZN(n5942) );
  OR2_X1 U7047 ( .A1(n8570), .A2(n8021), .ZN(n9353) );
  NAND2_X1 U7048 ( .A1(n8570), .A2(n8021), .ZN(n9311) );
  NAND2_X1 U7049 ( .A1(n7995), .A2(n9353), .ZN(n8541) );
  INV_X1 U7050 ( .A(n8541), .ZN(n5961) );
  XNOR2_X1 U7051 ( .A(n5947), .B(n5946), .ZN(n7313) );
  NAND2_X1 U7052 ( .A1(n7313), .A2(n9266), .ZN(n5953) );
  INV_X1 U7053 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U7054 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  NAND2_X1 U7055 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  XNOR2_X1 U7056 ( .A(n5951), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7772) );
  AOI22_X1 U7057 ( .A1(n5817), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6127), .B2(
        n7772), .ZN(n5952) );
  NAND2_X1 U7058 ( .A1(n6250), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5960) );
  INV_X1 U7059 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7770) );
  OR2_X1 U7060 ( .A1(n9247), .A2(n7770), .ZN(n5959) );
  INV_X1 U7061 ( .A(n5954), .ZN(n5974) );
  NAND2_X1 U7062 ( .A1(n5955), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5956) );
  AND2_X1 U7063 ( .A1(n5974), .A2(n5956), .ZN(n11063) );
  OR2_X1 U7064 ( .A1(n6237), .A2(n11063), .ZN(n5958) );
  INV_X1 U7065 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7771) );
  OR2_X1 U7066 ( .A1(n9251), .A2(n7771), .ZN(n5957) );
  NAND4_X1 U7067 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n9646)
         );
  AND2_X1 U7068 ( .A1(n8548), .A2(n9646), .ZN(n9309) );
  INV_X1 U7069 ( .A(n9646), .ZN(n8620) );
  XNOR2_X1 U7070 ( .A(n5963), .B(n5962), .ZN(n7321) );
  NAND2_X1 U7071 ( .A1(n7321), .A2(n9266), .ZN(n5972) );
  INV_X1 U7072 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5967) );
  NAND4_X1 U7073 ( .A1(n5964), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n5968)
         );
  NOR2_X1 U7074 ( .A1(n5969), .A2(n5968), .ZN(n5987) );
  OR2_X1 U7075 ( .A1(n5987), .A2(n5822), .ZN(n5970) );
  XNOR2_X1 U7076 ( .A(n5970), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8927) );
  AOI22_X1 U7077 ( .A1(n5817), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6127), .B2(
        n8927), .ZN(n5971) );
  NAND2_X1 U7078 ( .A1(n6250), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5980) );
  INV_X1 U7079 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5973) );
  OR2_X1 U7080 ( .A1(n9247), .A2(n5973), .ZN(n5979) );
  NAND2_X1 U7081 ( .A1(n5974), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5975) );
  AND2_X1 U7082 ( .A1(n5991), .A2(n5975), .ZN(n8802) );
  OR2_X1 U7083 ( .A1(n6237), .A2(n8802), .ZN(n5978) );
  INV_X1 U7084 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5976) );
  OR2_X1 U7085 ( .A1(n9251), .A2(n5976), .ZN(n5977) );
  NAND4_X1 U7086 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n9645)
         );
  AND2_X1 U7087 ( .A1(n8803), .A2(n9645), .ZN(n9356) );
  INV_X1 U7088 ( .A(n9356), .ZN(n5981) );
  INV_X1 U7089 ( .A(n8803), .ZN(n8622) );
  INV_X1 U7090 ( .A(n9645), .ZN(n8783) );
  AND2_X1 U7091 ( .A1(n8622), .A2(n8783), .ZN(n9313) );
  INV_X1 U7092 ( .A(n9313), .ZN(n9315) );
  NAND2_X1 U7093 ( .A1(n5981), .A2(n9315), .ZN(n8618) );
  NAND2_X1 U7094 ( .A1(n5243), .A2(n5983), .ZN(n5984) );
  NAND2_X1 U7095 ( .A1(n5985), .A2(n5984), .ZN(n7320) );
  OR2_X1 U7096 ( .A1(n7320), .A2(n5851), .ZN(n5990) );
  NAND2_X1 U7097 ( .A1(n5987), .A2(n5986), .ZN(n6000) );
  NAND2_X1 U7098 ( .A1(n6000), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5988) );
  XNOR2_X1 U7099 ( .A(n5988), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U7100 ( .A1(n5817), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6127), .B2(
        n10957), .ZN(n5989) );
  NAND2_X1 U7101 ( .A1(n6250), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5996) );
  INV_X1 U7102 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8936) );
  OR2_X1 U7103 ( .A1(n9247), .A2(n8936), .ZN(n5995) );
  NAND2_X1 U7104 ( .A1(n5991), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5992) );
  AND2_X1 U7105 ( .A1(n6006), .A2(n5992), .ZN(n8846) );
  OR2_X1 U7106 ( .A1(n6237), .A2(n8846), .ZN(n5994) );
  INV_X1 U7107 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8937) );
  OR2_X1 U7108 ( .A1(n9251), .A2(n8937), .ZN(n5993) );
  NOR2_X1 U7109 ( .A1(n8906), .A2(n8836), .ZN(n9355) );
  AND2_X1 U7110 ( .A1(n8906), .A2(n8836), .ZN(n9359) );
  INV_X1 U7111 ( .A(n9359), .ZN(n5997) );
  NAND2_X1 U7112 ( .A1(n7337), .A2(n9266), .ZN(n6004) );
  NAND2_X1 U7113 ( .A1(n6037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7114 ( .A1(n6001), .A2(n6035), .ZN(n6018) );
  OR2_X1 U7115 ( .A1(n6001), .A2(n6035), .ZN(n6002) );
  AOI22_X1 U7116 ( .A1(n5817), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6127), .B2(
        n10975), .ZN(n6003) );
  NAND2_X1 U7117 ( .A1(n6004), .A2(n6003), .ZN(n8915) );
  NAND2_X1 U7118 ( .A1(n6250), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6012) );
  INV_X1 U7119 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6005) );
  OR2_X1 U7120 ( .A1(n9247), .A2(n6005), .ZN(n6011) );
  INV_X1 U7121 ( .A(n6022), .ZN(n6008) );
  NAND2_X1 U7122 ( .A1(n6006), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6007) );
  AND2_X1 U7123 ( .A1(n6008), .A2(n6007), .ZN(n8913) );
  OR2_X1 U7124 ( .A1(n6237), .A2(n8913), .ZN(n6010) );
  INV_X1 U7125 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8797) );
  OR2_X1 U7126 ( .A1(n9251), .A2(n8797), .ZN(n6009) );
  NOR2_X1 U7127 ( .A1(n8915), .A2(n8975), .ZN(n9362) );
  INV_X1 U7128 ( .A(n9362), .ZN(n6013) );
  NAND2_X1 U7129 ( .A1(n8915), .A2(n8975), .ZN(n9361) );
  NAND2_X1 U7130 ( .A1(n8794), .A2(n9361), .ZN(n6028) );
  NAND2_X1 U7131 ( .A1(n6015), .A2(n6014), .ZN(n6017) );
  NAND2_X1 U7132 ( .A1(n6017), .A2(n6016), .ZN(n7468) );
  OR2_X1 U7133 ( .A1(n7468), .A2(n5851), .ZN(n6021) );
  NAND2_X1 U7134 ( .A1(n6018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6019) );
  XNOR2_X1 U7135 ( .A(n6019), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8954) );
  AOI22_X1 U7136 ( .A1(n5817), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6127), .B2(
        n8954), .ZN(n6020) );
  NAND2_X1 U7137 ( .A1(n6250), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7138 ( .A1(n9247), .A2(n9165), .ZN(n6026) );
  OR2_X1 U7139 ( .A1(n6022), .A2(n8943), .ZN(n6023) );
  AND2_X1 U7140 ( .A1(n6042), .A2(n6023), .ZN(n8968) );
  OR2_X1 U7141 ( .A1(n6237), .A2(n8968), .ZN(n6025) );
  INV_X1 U7142 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8984) );
  OR2_X1 U7143 ( .A1(n9251), .A2(n8984), .ZN(n6024) );
  XNOR2_X1 U7144 ( .A(n9367), .B(n8994), .ZN(n9372) );
  NAND2_X1 U7145 ( .A1(n6028), .A2(n9372), .ZN(n8983) );
  AND2_X1 U7146 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  INV_X1 U7147 ( .A(n9368), .ZN(n6029) );
  OR2_X1 U7148 ( .A1(n6031), .A2(n6030), .ZN(n6032) );
  NAND2_X1 U7149 ( .A1(n6033), .A2(n6032), .ZN(n7549) );
  OR2_X1 U7150 ( .A1(n7549), .A2(n5851), .ZN(n6040) );
  INV_X1 U7151 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7152 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  NAND2_X1 U7153 ( .A1(n6051), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6038) );
  XNOR2_X1 U7154 ( .A(n6038), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9668) );
  AOI22_X1 U7155 ( .A1(n5817), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6127), .B2(
        n9668), .ZN(n6039) );
  NAND2_X1 U7156 ( .A1(n6250), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6047) );
  INV_X1 U7157 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6041) );
  OR2_X1 U7158 ( .A1(n9251), .A2(n6041), .ZN(n6046) );
  AOI21_X1 U7159 ( .B1(n6042), .B2(P2_REG3_REG_13__SCAN_IN), .A(n6056), .ZN(
        n9028) );
  OR2_X1 U7160 ( .A1(n6237), .A2(n9028), .ZN(n6045) );
  INV_X1 U7161 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6043) );
  OR2_X1 U7162 ( .A1(n6181), .A2(n6043), .ZN(n6044) );
  NAND2_X1 U7163 ( .A1(n9022), .A2(n9139), .ZN(n9374) );
  INV_X1 U7164 ( .A(n9374), .ZN(n6048) );
  OR2_X1 U7165 ( .A1(n9022), .A2(n9139), .ZN(n9375) );
  XNOR2_X1 U7166 ( .A(n6050), .B(n6049), .ZN(n7574) );
  NAND2_X1 U7167 ( .A1(n7574), .A2(n9266), .ZN(n6053) );
  OAI21_X1 U7168 ( .B1(n6051), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7169 ( .A(n6067), .B(n6066), .ZN(n9689) );
  INV_X1 U7170 ( .A(n9689), .ZN(n9657) );
  AOI22_X1 U7171 ( .A1(n5817), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6127), .B2(
        n9657), .ZN(n6052) );
  NAND2_X1 U7172 ( .A1(n6250), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6061) );
  INV_X1 U7173 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7174 ( .A1(n9251), .A2(n6054), .ZN(n6060) );
  INV_X1 U7175 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6055) );
  OR2_X1 U7176 ( .A1(n9247), .A2(n6055), .ZN(n6059) );
  OAI21_X1 U7177 ( .B1(n9147), .B2(n6056), .A(n6072), .ZN(n9150) );
  INV_X1 U7178 ( .A(n9150), .ZN(n6057) );
  OR2_X1 U7179 ( .A1(n6237), .A2(n6057), .ZN(n6058) );
  XNOR2_X1 U7180 ( .A(n9138), .B(n9197), .ZN(n9377) );
  INV_X1 U7181 ( .A(n9377), .ZN(n9289) );
  NOR2_X1 U7182 ( .A1(n9138), .A2(n9197), .ZN(n9382) );
  NAND2_X1 U7183 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  OR2_X1 U7184 ( .A1(n7652), .A2(n5851), .ZN(n6070) );
  NAND2_X1 U7185 ( .A1(n6067), .A2(n6066), .ZN(n6068) );
  NAND2_X1 U7186 ( .A1(n6068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6081) );
  XNOR2_X1 U7187 ( .A(n6081), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9711) );
  AOI22_X1 U7188 ( .A1(n5817), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6127), .B2(
        n9711), .ZN(n6069) );
  INV_X1 U7189 ( .A(n10028), .ZN(n6295) );
  NAND2_X1 U7190 ( .A1(n6250), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6077) );
  INV_X1 U7191 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6071) );
  OR2_X1 U7192 ( .A1(n6181), .A2(n6071), .ZN(n6076) );
  AOI21_X1 U7193 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(n6072), .A(n6089), .ZN(
        n9120) );
  OR2_X1 U7194 ( .A1(n6237), .A2(n9120), .ZN(n6075) );
  INV_X1 U7195 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7196 ( .A1(n9251), .A2(n6073), .ZN(n6074) );
  NAND4_X1 U7197 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n9640)
         );
  NAND2_X1 U7198 ( .A1(n6295), .A2(n9953), .ZN(n9385) );
  NAND2_X1 U7199 ( .A1(n9119), .A2(n9385), .ZN(n9948) );
  XNOR2_X1 U7200 ( .A(n6079), .B(n6078), .ZN(n7819) );
  NAND2_X1 U7201 ( .A1(n7819), .A2(n9266), .ZN(n6087) );
  INV_X1 U7202 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7203 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  NAND2_X1 U7204 ( .A1(n6082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6084) );
  INV_X1 U7205 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7206 ( .A1(n6084), .A2(n6083), .ZN(n6100) );
  OR2_X1 U7207 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  AOI22_X1 U7208 ( .A1(n6127), .A2(n9714), .B1(n5817), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7209 ( .A1(n6250), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6095) );
  INV_X1 U7210 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6088) );
  OR2_X1 U7211 ( .A1(n9247), .A2(n6088), .ZN(n6094) );
  INV_X1 U7212 ( .A(n6089), .ZN(n6091) );
  INV_X1 U7213 ( .A(n6105), .ZN(n6090) );
  AOI21_X1 U7214 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(n6091), .A(n6090), .ZN(
        n9958) );
  OR2_X1 U7215 ( .A1(n6237), .A2(n9958), .ZN(n6093) );
  INV_X1 U7216 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9959) );
  OR2_X1 U7217 ( .A1(n9251), .A2(n9959), .ZN(n6092) );
  OR2_X1 U7218 ( .A1(n10021), .A2(n9568), .ZN(n9308) );
  NAND2_X1 U7219 ( .A1(n10028), .A2(n9640), .ZN(n9947) );
  NAND2_X1 U7220 ( .A1(n9308), .A2(n9947), .ZN(n9386) );
  INV_X1 U7221 ( .A(n9386), .ZN(n6096) );
  NAND2_X1 U7222 ( .A1(n9948), .A2(n6096), .ZN(n6097) );
  NAND2_X1 U7223 ( .A1(n6097), .A2(n9396), .ZN(n9942) );
  XNOR2_X1 U7224 ( .A(n6099), .B(n6098), .ZN(n8037) );
  NAND2_X1 U7225 ( .A1(n8037), .A2(n9266), .ZN(n6103) );
  NAND2_X1 U7226 ( .A1(n6100), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6101) );
  XNOR2_X1 U7227 ( .A(n6101), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9764) );
  AOI22_X1 U7228 ( .A1(n9764), .A2(n6127), .B1(n5817), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7229 ( .A1(n6250), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6109) );
  INV_X1 U7230 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9940) );
  OR2_X1 U7231 ( .A1(n9251), .A2(n9940), .ZN(n6108) );
  AOI21_X1 U7232 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n6105), .A(n6104), .ZN(
        n9939) );
  OR2_X1 U7233 ( .A1(n6237), .A2(n9939), .ZN(n6107) );
  INV_X1 U7234 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9726) );
  OR2_X1 U7235 ( .A1(n9247), .A2(n9726), .ZN(n6106) );
  OR2_X1 U7236 ( .A1(n10013), .A2(n9955), .ZN(n9401) );
  NAND2_X1 U7237 ( .A1(n10013), .A2(n9955), .ZN(n9392) );
  NAND2_X1 U7238 ( .A1(n9401), .A2(n9392), .ZN(n9390) );
  NAND2_X1 U7239 ( .A1(n5128), .A2(n6110), .ZN(n6111) );
  NAND2_X1 U7240 ( .A1(n6112), .A2(n6111), .ZN(n8054) );
  NAND2_X1 U7241 ( .A1(n6126), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6114) );
  XNOR2_X1 U7242 ( .A(n6114), .B(P2_IR_REG_18__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U7243 ( .A1(n5817), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6127), .B2(
        n11003), .ZN(n6115) );
  NAND2_X1 U7244 ( .A1(n6330), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6123) );
  INV_X1 U7245 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6117) );
  OR2_X1 U7246 ( .A1(n9249), .A2(n6117), .ZN(n6122) );
  AND2_X1 U7247 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(n6118), .ZN(n6119) );
  NOR2_X1 U7248 ( .A1(n6130), .A2(n6119), .ZN(n9921) );
  OR2_X1 U7249 ( .A1(n6237), .A2(n9921), .ZN(n6121) );
  INV_X1 U7250 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9922) );
  OR2_X1 U7251 ( .A1(n9251), .A2(n9922), .ZN(n6120) );
  NAND2_X1 U7252 ( .A1(n10009), .A2(n9906), .ZN(n9399) );
  NAND2_X1 U7253 ( .A1(n9925), .A2(n9394), .ZN(n9909) );
  XNOR2_X1 U7254 ( .A(n6125), .B(n6124), .ZN(n8690) );
  NAND2_X1 U7255 ( .A1(n8690), .A2(n9266), .ZN(n6129) );
  AOI22_X1 U7256 ( .A1(n5817), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9754), .B2(
        n6127), .ZN(n6128) );
  NAND2_X1 U7257 ( .A1(n6250), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6136) );
  INV_X1 U7258 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10006) );
  OR2_X1 U7259 ( .A1(n9247), .A2(n10006), .ZN(n6135) );
  NOR2_X1 U7260 ( .A1(n6130), .A2(n9537), .ZN(n6131) );
  OR2_X1 U7261 ( .A1(n6142), .A2(n6131), .ZN(n9911) );
  INV_X1 U7262 ( .A(n9911), .ZN(n9540) );
  OR2_X1 U7263 ( .A1(n6237), .A2(n9540), .ZN(n6134) );
  INV_X1 U7264 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6132) );
  OR2_X1 U7265 ( .A1(n9251), .A2(n6132), .ZN(n6133) );
  NOR2_X1 U7266 ( .A1(n9910), .A2(n6307), .ZN(n9407) );
  XNOR2_X1 U7267 ( .A(n6137), .B(n6138), .ZN(n8850) );
  NAND2_X1 U7268 ( .A1(n8850), .A2(n9266), .ZN(n6140) );
  INV_X1 U7269 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8851) );
  OR2_X1 U7270 ( .A1(n9267), .A2(n8851), .ZN(n6139) );
  NAND2_X1 U7271 ( .A1(n6330), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6147) );
  INV_X1 U7272 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7273 ( .A1(n9249), .A2(n6141), .ZN(n6146) );
  NOR2_X1 U7274 ( .A1(n6142), .A2(n9591), .ZN(n6143) );
  NOR2_X1 U7275 ( .A1(n6156), .A2(n6143), .ZN(n9895) );
  OR2_X1 U7276 ( .A1(n6237), .A2(n9895), .ZN(n6145) );
  INV_X1 U7277 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9896) );
  OR2_X1 U7278 ( .A1(n9251), .A2(n9896), .ZN(n6144) );
  NAND2_X1 U7279 ( .A1(n10000), .A2(n9907), .ZN(n9412) );
  NAND2_X1 U7280 ( .A1(n9910), .A2(n6307), .ZN(n9898) );
  NAND2_X1 U7281 ( .A1(n9412), .A2(n9898), .ZN(n9405) );
  INV_X1 U7282 ( .A(n9405), .ZN(n6148) );
  NOR2_X1 U7283 ( .A1(n10000), .A2(n9907), .ZN(n9409) );
  INV_X1 U7284 ( .A(n9409), .ZN(n6308) );
  INV_X1 U7285 ( .A(n6149), .ZN(n6151) );
  NAND2_X1 U7286 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  NAND2_X1 U7287 ( .A1(n6153), .A2(n6152), .ZN(n8823) );
  INV_X1 U7288 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8809) );
  OR2_X1 U7289 ( .A1(n9267), .A2(n8809), .ZN(n6154) );
  NAND2_X1 U7290 ( .A1(n5899), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6162) );
  INV_X1 U7291 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9884) );
  OR2_X1 U7292 ( .A1(n9251), .A2(n9884), .ZN(n6161) );
  OR2_X1 U7293 ( .A1(n6156), .A2(n9547), .ZN(n6157) );
  AND2_X1 U7294 ( .A1(n6157), .A2(n6168), .ZN(n9883) );
  OR2_X1 U7295 ( .A1(n6237), .A2(n9883), .ZN(n6160) );
  INV_X1 U7296 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6158) );
  OR2_X1 U7297 ( .A1(n6181), .A2(n6158), .ZN(n6159) );
  NAND2_X1 U7298 ( .A1(n9996), .A2(n9863), .ZN(n9413) );
  NAND2_X1 U7299 ( .A1(n9887), .A2(n9886), .ZN(n9885) );
  NAND2_X1 U7300 ( .A1(n6163), .A2(n8349), .ZN(n6164) );
  NAND2_X1 U7301 ( .A1(n6165), .A2(n6164), .ZN(n9113) );
  OR2_X1 U7302 ( .A1(n9113), .A2(n5851), .ZN(n6167) );
  INV_X1 U7303 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9003) );
  OR2_X1 U7304 ( .A1(n9267), .A2(n9003), .ZN(n6166) );
  NAND2_X1 U7305 ( .A1(n6330), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6173) );
  INV_X1 U7306 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n10055) );
  OR2_X1 U7307 ( .A1(n9249), .A2(n10055), .ZN(n6172) );
  NAND2_X1 U7308 ( .A1(n6168), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6169) );
  AND2_X1 U7309 ( .A1(n6182), .A2(n6169), .ZN(n9866) );
  OR2_X1 U7310 ( .A1(n6237), .A2(n9866), .ZN(n6171) );
  INV_X1 U7311 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9867) );
  OR2_X1 U7312 ( .A1(n9251), .A2(n9867), .ZN(n6170) );
  NOR2_X1 U7313 ( .A1(n9874), .A2(n9548), .ZN(n9419) );
  INV_X1 U7314 ( .A(n9419), .ZN(n6175) );
  AND2_X1 U7315 ( .A1(n9874), .A2(n9548), .ZN(n9418) );
  INV_X1 U7316 ( .A(n9418), .ZN(n6174) );
  NAND2_X1 U7317 ( .A1(n6175), .A2(n6174), .ZN(n9860) );
  INV_X1 U7318 ( .A(n9860), .ZN(n9868) );
  NAND2_X1 U7319 ( .A1(n9134), .A2(n9266), .ZN(n6179) );
  INV_X1 U7320 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9137) );
  OR2_X1 U7321 ( .A1(n9267), .A2(n9137), .ZN(n6178) );
  NAND2_X1 U7322 ( .A1(n6250), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6187) );
  INV_X1 U7323 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6180) );
  OR2_X1 U7324 ( .A1(n6181), .A2(n6180), .ZN(n6186) );
  AND2_X1 U7325 ( .A1(n6182), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6183) );
  NOR2_X1 U7326 ( .A1(n6193), .A2(n6183), .ZN(n9852) );
  OR2_X1 U7327 ( .A1(n6237), .A2(n9852), .ZN(n6185) );
  INV_X1 U7328 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9853) );
  OR2_X1 U7329 ( .A1(n9251), .A2(n9853), .ZN(n6184) );
  XNOR2_X1 U7330 ( .A(n9987), .B(n9639), .ZN(n9855) );
  NOR2_X1 U7331 ( .A1(n9987), .A2(n9862), .ZN(n9423) );
  INV_X1 U7332 ( .A(n9423), .ZN(n6188) );
  XNOR2_X1 U7333 ( .A(n6190), .B(n6189), .ZN(n9232) );
  NAND2_X1 U7334 ( .A1(n9232), .A2(n9266), .ZN(n6192) );
  INV_X1 U7335 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9235) );
  OR2_X1 U7336 ( .A1(n9267), .A2(n9235), .ZN(n6191) );
  NAND2_X1 U7337 ( .A1(n6330), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6199) );
  INV_X1 U7338 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10050) );
  OR2_X1 U7339 ( .A1(n9249), .A2(n10050), .ZN(n6198) );
  NOR2_X1 U7340 ( .A1(n6193), .A2(n9581), .ZN(n6194) );
  OR2_X1 U7341 ( .A1(n6209), .A2(n6194), .ZN(n9584) );
  INV_X1 U7342 ( .A(n9584), .ZN(n9842) );
  OR2_X1 U7343 ( .A1(n6237), .A2(n9842), .ZN(n6197) );
  INV_X1 U7344 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6195) );
  OR2_X1 U7345 ( .A1(n9251), .A2(n6195), .ZN(n6196) );
  AND2_X1 U7346 ( .A1(n9574), .A2(n9830), .ZN(n9427) );
  INV_X1 U7347 ( .A(n9427), .ZN(n6200) );
  NOR2_X1 U7348 ( .A1(n9574), .A2(n9830), .ZN(n9426) );
  INV_X1 U7349 ( .A(n9426), .ZN(n6201) );
  OR2_X1 U7350 ( .A1(n6204), .A2(n6203), .ZN(n6206) );
  NAND2_X1 U7351 ( .A1(n6206), .A2(n6205), .ZN(n9242) );
  INV_X1 U7352 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9239) );
  OR2_X1 U7353 ( .A1(n9267), .A2(n9239), .ZN(n6207) );
  NAND2_X1 U7354 ( .A1(n6330), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6214) );
  INV_X1 U7355 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10046) );
  OR2_X1 U7356 ( .A1(n9249), .A2(n10046), .ZN(n6213) );
  OR2_X1 U7357 ( .A1(n6209), .A2(n9559), .ZN(n6210) );
  AND2_X1 U7358 ( .A1(n6222), .A2(n6210), .ZN(n9832) );
  OR2_X1 U7359 ( .A1(n6237), .A2(n9832), .ZN(n6212) );
  INV_X1 U7360 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9838) );
  OR2_X1 U7361 ( .A1(n9251), .A2(n9838), .ZN(n6211) );
  OR2_X1 U7362 ( .A1(n9554), .A2(n9841), .ZN(n6215) );
  NAND2_X1 U7363 ( .A1(n9554), .A2(n9841), .ZN(n9429) );
  INV_X1 U7364 ( .A(n9834), .ZN(n6216) );
  NOR2_X1 U7365 ( .A1(n9554), .A2(n9841), .ZN(n9430) );
  NAND2_X1 U7366 ( .A1(n10085), .A2(n9266), .ZN(n6221) );
  INV_X1 U7367 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6219) );
  OR2_X1 U7368 ( .A1(n9267), .A2(n6219), .ZN(n6220) );
  NAND2_X1 U7369 ( .A1(n5899), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6227) );
  INV_X1 U7370 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9977) );
  OR2_X1 U7371 ( .A1(n9247), .A2(n9977), .ZN(n6226) );
  NAND2_X1 U7372 ( .A1(n6222), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6223) );
  INV_X1 U7373 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9823) );
  OR2_X1 U7374 ( .A1(n9251), .A2(n9823), .ZN(n6224) );
  NOR2_X1 U7375 ( .A1(n9630), .A2(n9831), .ZN(n6229) );
  NAND2_X1 U7376 ( .A1(n9630), .A2(n9831), .ZN(n6228) );
  NAND2_X1 U7377 ( .A1(n10081), .A2(n9266), .ZN(n6234) );
  INV_X1 U7378 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6232) );
  OR2_X1 U7379 ( .A1(n9267), .A2(n6232), .ZN(n6233) );
  NAND2_X1 U7380 ( .A1(n6330), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6241) );
  INV_X1 U7381 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10037) );
  OR2_X1 U7382 ( .A1(n9249), .A2(n10037), .ZN(n6240) );
  AOI21_X1 U7383 ( .B1(n6236), .B2(P2_REG3_REG_27__SCAN_IN), .A(n6235), .ZN(
        n9809) );
  OR2_X1 U7384 ( .A1(n6237), .A2(n9809), .ZN(n6239) );
  INV_X1 U7385 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9810) );
  OR2_X1 U7386 ( .A1(n9251), .A2(n9810), .ZN(n6238) );
  OR2_X1 U7387 ( .A1(n6268), .A2(n9819), .ZN(n6321) );
  INV_X1 U7388 ( .A(n6321), .ZN(n9435) );
  NAND2_X1 U7389 ( .A1(n6268), .A2(n9819), .ZN(n9434) );
  XNOR2_X1 U7390 ( .A(n9966), .B(n9636), .ZN(n9796) );
  OAI21_X1 U7391 ( .B1(n9441), .B2(n9636), .A(n9795), .ZN(n9264) );
  NAND2_X1 U7392 ( .A1(n6243), .A2(n6242), .ZN(n6247) );
  INV_X1 U7393 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U7394 ( .A1(n6245), .A2(n8138), .ZN(n6246) );
  MUX2_X1 U7395 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7287), .Z(n6974) );
  INV_X1 U7396 ( .A(SI_29_), .ZN(n6248) );
  XNOR2_X1 U7397 ( .A(n6972), .B(n6248), .ZN(n10075) );
  INV_X1 U7398 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U7399 ( .A1(n9267), .A2(n10076), .ZN(n6249) );
  NAND2_X1 U7400 ( .A1(n6250), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6253) );
  INV_X1 U7401 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6388) );
  OR2_X1 U7402 ( .A1(n9247), .A2(n6388), .ZN(n6252) );
  INV_X1 U7403 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9778) );
  OR2_X1 U7404 ( .A1(n9251), .A2(n9778), .ZN(n6251) );
  NAND4_X1 U7405 ( .A1(n9255), .A2(n6253), .A3(n6252), .A4(n6251), .ZN(n9787)
         );
  AND2_X1 U7406 ( .A1(n6390), .A2(n9787), .ZN(n9451) );
  INV_X1 U7407 ( .A(n9451), .ZN(n9265) );
  INV_X1 U7408 ( .A(n6390), .ZN(n9780) );
  INV_X1 U7409 ( .A(n9787), .ZN(n9516) );
  NAND2_X1 U7410 ( .A1(n9780), .A2(n9516), .ZN(n9271) );
  NAND2_X1 U7411 ( .A1(n9265), .A2(n9271), .ZN(n6323) );
  NAND2_X1 U7412 ( .A1(n6255), .A2(n6260), .ZN(n6256) );
  NAND2_X1 U7413 ( .A1(n6265), .A2(n6261), .ZN(n6257) );
  INV_X1 U7414 ( .A(n6258), .ZN(n6262) );
  NAND2_X1 U7415 ( .A1(n6262), .A2(n6338), .ZN(n6263) );
  NAND2_X1 U7416 ( .A1(n6263), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6264) );
  AND2_X1 U7417 ( .A1(n9459), .A2(n9762), .ZN(n6384) );
  INV_X1 U7418 ( .A(n9465), .ZN(n9004) );
  AOI21_X1 U7419 ( .B1(n9004), .B2(n9458), .A(n9754), .ZN(n6266) );
  NAND2_X1 U7420 ( .A1(n10027), .A2(n6266), .ZN(n6267) );
  INV_X1 U7421 ( .A(n7747), .ZN(n7564) );
  NAND2_X1 U7422 ( .A1(n9651), .A2(n7564), .ZN(n6270) );
  INV_X1 U7423 ( .A(n7860), .ZN(n7433) );
  OR2_X1 U7424 ( .A1(n7433), .A2(n6271), .ZN(n6272) );
  NAND2_X1 U7425 ( .A1(n7806), .A2(n9325), .ZN(n6275) );
  OR2_X1 U7426 ( .A1(n5428), .A2(n6273), .ZN(n6274) );
  INV_X1 U7427 ( .A(n7648), .ZN(n7821) );
  NOR2_X1 U7428 ( .A1(n9650), .A2(n7821), .ZN(n6277) );
  NAND2_X1 U7429 ( .A1(n9650), .A2(n7821), .ZN(n6276) );
  INV_X1 U7430 ( .A(n7852), .ZN(n7559) );
  AND2_X1 U7431 ( .A1(n7559), .A2(n7644), .ZN(n6278) );
  AND2_X1 U7432 ( .A1(n8013), .A2(n7826), .ZN(n6280) );
  NAND2_X1 U7433 ( .A1(n7871), .A2(n9649), .ZN(n6279) );
  AND2_X1 U7434 ( .A1(n8010), .A2(n9648), .ZN(n6281) );
  NAND2_X1 U7435 ( .A1(n7999), .A2(n7998), .ZN(n6283) );
  INV_X1 U7436 ( .A(n8021), .ZN(n9647) );
  OR2_X1 U7437 ( .A1(n8570), .A2(n9647), .ZN(n6282) );
  NAND2_X1 U7438 ( .A1(n6283), .A2(n6282), .ZN(n8542) );
  INV_X1 U7439 ( .A(n9309), .ZN(n9354) );
  AND2_X1 U7440 ( .A1(n9354), .A2(n9312), .ZN(n9285) );
  INV_X1 U7441 ( .A(n9285), .ZN(n8543) );
  NAND2_X1 U7442 ( .A1(n8542), .A2(n8543), .ZN(n6285) );
  NAND2_X1 U7443 ( .A1(n8548), .A2(n8620), .ZN(n6284) );
  INV_X1 U7444 ( .A(n8836), .ZN(n9644) );
  INV_X1 U7445 ( .A(n8975), .ZN(n9643) );
  NAND2_X1 U7446 ( .A1(n8792), .A2(n9643), .ZN(n6286) );
  INV_X1 U7447 ( .A(n8915), .ZN(n8921) );
  NAND2_X1 U7448 ( .A1(n6286), .A2(n8921), .ZN(n6289) );
  INV_X1 U7449 ( .A(n8792), .ZN(n6287) );
  NAND2_X1 U7450 ( .A1(n6287), .A2(n8975), .ZN(n6288) );
  NAND2_X1 U7451 ( .A1(n6289), .A2(n6288), .ZN(n8974) );
  INV_X1 U7452 ( .A(n8974), .ZN(n6290) );
  NAND2_X1 U7453 ( .A1(n9367), .A2(n8994), .ZN(n6291) );
  INV_X1 U7454 ( .A(n9139), .ZN(n9642) );
  NAND2_X1 U7455 ( .A1(n9022), .A2(n9642), .ZN(n6292) );
  INV_X1 U7456 ( .A(n9197), .ZN(n9641) );
  NAND2_X1 U7457 ( .A1(n9138), .A2(n9641), .ZN(n6293) );
  NAND2_X1 U7458 ( .A1(n6294), .A2(n6293), .ZN(n9114) );
  NAND2_X1 U7459 ( .A1(n9947), .A2(n9385), .ZN(n9383) );
  NAND2_X1 U7460 ( .A1(n9114), .A2(n9383), .ZN(n6297) );
  NAND2_X1 U7461 ( .A1(n6295), .A2(n9640), .ZN(n6296) );
  NAND2_X1 U7462 ( .A1(n6297), .A2(n6296), .ZN(n9930) );
  NAND2_X1 U7463 ( .A1(n9308), .A2(n9396), .ZN(n9950) );
  INV_X1 U7464 ( .A(n9955), .ZN(n9918) );
  NAND2_X1 U7465 ( .A1(n10013), .A2(n9918), .ZN(n6301) );
  INV_X1 U7466 ( .A(n6301), .ZN(n6298) );
  OR2_X1 U7467 ( .A1(n6298), .A2(n9390), .ZN(n6300) );
  AND2_X1 U7468 ( .A1(n9950), .A2(n6300), .ZN(n6299) );
  NAND2_X1 U7469 ( .A1(n9930), .A2(n6299), .ZN(n6305) );
  INV_X1 U7470 ( .A(n6300), .ZN(n6303) );
  INV_X1 U7471 ( .A(n9568), .ZN(n9935) );
  NAND2_X1 U7472 ( .A1(n10021), .A2(n9935), .ZN(n9931) );
  AND2_X1 U7473 ( .A1(n9931), .A2(n6301), .ZN(n6302) );
  OR2_X1 U7474 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  INV_X1 U7475 ( .A(n9906), .ZN(n9937) );
  NAND2_X1 U7476 ( .A1(n10009), .A2(n9937), .ZN(n6306) );
  NAND2_X1 U7477 ( .A1(n9892), .A2(n9891), .ZN(n9877) );
  INV_X1 U7478 ( .A(n9907), .ZN(n9880) );
  OR2_X1 U7479 ( .A1(n10000), .A2(n9880), .ZN(n9876) );
  INV_X1 U7480 ( .A(n9863), .ZN(n9893) );
  OR2_X1 U7481 ( .A1(n9996), .A2(n9893), .ZN(n6309) );
  AND2_X1 U7482 ( .A1(n9876), .A2(n6309), .ZN(n6311) );
  NOR2_X1 U7483 ( .A1(n9874), .A2(n9881), .ZN(n6312) );
  NAND2_X1 U7484 ( .A1(n9874), .A2(n9881), .ZN(n6313) );
  NAND2_X1 U7485 ( .A1(n6314), .A2(n6313), .ZN(n9849) );
  OR2_X1 U7486 ( .A1(n9987), .A2(n9639), .ZN(n6315) );
  NAND2_X1 U7487 ( .A1(n9828), .A2(n9834), .ZN(n6317) );
  INV_X1 U7488 ( .A(n9841), .ZN(n9638) );
  NAND2_X1 U7489 ( .A1(n9554), .A2(n9638), .ZN(n6316) );
  NAND2_X1 U7490 ( .A1(n6317), .A2(n6316), .ZN(n9817) );
  INV_X1 U7491 ( .A(n9817), .ZN(n6318) );
  NAND2_X1 U7492 ( .A1(n6318), .A2(n5153), .ZN(n6320) );
  OR2_X1 U7493 ( .A1(n9630), .A2(n9637), .ZN(n6319) );
  NAND2_X1 U7494 ( .A1(n6321), .A2(n9434), .ZN(n9812) );
  INV_X1 U7495 ( .A(n9812), .ZN(n9800) );
  NOR2_X1 U7496 ( .A1(n9966), .A2(n9636), .ZN(n6322) );
  XNOR2_X1 U7497 ( .A(n5143), .B(n6323), .ZN(n6326) );
  NAND2_X1 U7498 ( .A1(n9323), .A2(n9458), .ZN(n6324) );
  NAND2_X1 U7499 ( .A1(n9465), .A2(n9754), .ZN(n6365) );
  INV_X1 U7500 ( .A(n9951), .ZN(n6325) );
  NAND2_X1 U7501 ( .A1(n6326), .A2(n6325), .ZN(n6337) );
  OR2_X1 U7502 ( .A1(n9756), .A2(n7359), .ZN(n6328) );
  NAND2_X1 U7503 ( .A1(n5852), .A2(n6328), .ZN(n7429) );
  NOR2_X2 U7504 ( .A1(n7429), .A2(n9449), .ZN(n9934) );
  AND2_X1 U7505 ( .A1(n5852), .A2(P2_B_REG_SCAN_IN), .ZN(n6329) );
  NOR2_X1 U7506 ( .A1(n9956), .A2(n6329), .ZN(n9256) );
  NAND2_X1 U7507 ( .A1(n6330), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6335) );
  INV_X1 U7508 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6331) );
  OR2_X1 U7509 ( .A1(n9249), .A2(n6331), .ZN(n6334) );
  INV_X1 U7510 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6332) );
  OR2_X1 U7511 ( .A1(n9251), .A2(n6332), .ZN(n6333) );
  NAND4_X1 U7512 ( .A1(n9255), .A2(n6335), .A3(n6334), .A4(n6333), .ZN(n9635)
         );
  AOI22_X1 U7513 ( .A1(n9636), .A2(n9934), .B1(n9256), .B2(n9635), .ZN(n6336)
         );
  AND2_X1 U7514 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  OAI21_X1 U7515 ( .B1(n6370), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6342) );
  MUX2_X1 U7516 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6342), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n6343) );
  XNOR2_X1 U7517 ( .A(n6369), .B(n8430), .ZN(n6350) );
  NAND2_X1 U7518 ( .A1(n5146), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6344) );
  MUX2_X1 U7519 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6344), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6346) );
  NAND2_X1 U7520 ( .A1(n6346), .A2(n6345), .ZN(n9240) );
  NAND2_X1 U7521 ( .A1(n6345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6347) );
  MUX2_X1 U7522 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6347), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6349) );
  AOI21_X2 U7523 ( .B1(n6350), .B2(n9240), .A(n10088), .ZN(n7301) );
  INV_X1 U7524 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7306) );
  NAND2_X1 U7525 ( .A1(n7301), .A2(n7306), .ZN(n6351) );
  INV_X1 U7526 ( .A(n6369), .ZN(n9236) );
  NAND2_X1 U7527 ( .A1(n9236), .A2(n10088), .ZN(n7303) );
  NAND2_X1 U7528 ( .A1(n6351), .A2(n7303), .ZN(n6378) );
  INV_X1 U7529 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U7530 ( .A1(n7301), .A2(n7292), .ZN(n6353) );
  NAND2_X1 U7531 ( .A1(n10088), .A2(n9240), .ZN(n6352) );
  INV_X1 U7532 ( .A(n6382), .ZN(n6364) );
  NOR2_X1 U7533 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6357) );
  NOR4_X1 U7534 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6356) );
  NOR4_X1 U7535 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6355) );
  NOR4_X1 U7536 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6354) );
  NAND4_X1 U7537 ( .A1(n6357), .A2(n6356), .A3(n6355), .A4(n6354), .ZN(n6363)
         );
  NOR4_X1 U7538 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6361) );
  NOR4_X1 U7539 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6360) );
  NOR4_X1 U7540 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6359) );
  NOR4_X1 U7541 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6358) );
  NAND4_X1 U7542 ( .A1(n6361), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(n6362)
         );
  OAI21_X1 U7543 ( .B1(n6363), .B2(n6362), .A(n7301), .ZN(n6380) );
  NAND2_X1 U7544 ( .A1(n6364), .A2(n6380), .ZN(n7424) );
  INV_X1 U7545 ( .A(n7418), .ZN(n7407) );
  NOR2_X1 U7546 ( .A1(n7741), .A2(n7407), .ZN(n6367) );
  AND2_X1 U7547 ( .A1(n10027), .A2(n9449), .ZN(n7417) );
  NAND2_X1 U7548 ( .A1(n7417), .A2(n7418), .ZN(n6366) );
  AND2_X1 U7549 ( .A1(n6366), .A2(n9843), .ZN(n7402) );
  NAND3_X1 U7550 ( .A1(n7726), .A2(n7728), .A3(n6380), .ZN(n7431) );
  OAI22_X1 U7551 ( .A1(n7424), .A2(n6367), .B1(n7402), .B2(n7431), .ZN(n6373)
         );
  NOR2_X1 U7552 ( .A1(n10088), .A2(n9240), .ZN(n6368) );
  NAND2_X1 U7553 ( .A1(n6370), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7554 ( .A1(n9780), .A2(n6374), .ZN(n6377) );
  INV_X1 U7555 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6375) );
  OR2_X1 U7556 ( .A1(n11108), .A2(n6375), .ZN(n6376) );
  INV_X1 U7557 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U7558 ( .A1(n6379), .A2(n9302), .ZN(n7413) );
  INV_X1 U7559 ( .A(n7833), .ZN(n8902) );
  AND2_X1 U7560 ( .A1(n6380), .A2(n7425), .ZN(n6381) );
  NAND3_X1 U7561 ( .A1(n9458), .A2(n9465), .A3(n9762), .ZN(n6383) );
  INV_X1 U7562 ( .A(n6385), .ZN(n7727) );
  NAND2_X1 U7563 ( .A1(n7728), .A2(n7727), .ZN(n7730) );
  NOR2_X1 U7564 ( .A1(n9449), .A2(n6384), .ZN(n7725) );
  OAI21_X1 U7565 ( .B1(n7725), .B2(n6385), .A(n7726), .ZN(n6386) );
  OAI211_X4 U7566 ( .C1(n7413), .C2(n8902), .A(n7731), .B(n6387), .ZN(n10023)
         );
  NAND2_X1 U7567 ( .A1(n10023), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6389) );
  OAI21_X1 U7568 ( .B1(n6390), .B2(n10008), .A(n6389), .ZN(n6391) );
  INV_X1 U7569 ( .A(n6391), .ZN(n6392) );
  OAI21_X1 U7570 ( .B1(n6393), .B2(n10023), .A(n6392), .ZN(P2_U3488) );
  NOR2_X1 U7571 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6394) );
  NOR2_X1 U7572 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6398) );
  INV_X1 U7573 ( .A(n6685), .ZN(n6403) );
  INV_X1 U7574 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6419) );
  NOR2_X1 U7575 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6402) );
  NOR2_X1 U7576 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n6401) );
  NAND2_X1 U7577 ( .A1(n6407), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6404) );
  INV_X1 U7578 ( .A(n6449), .ZN(n6405) );
  NAND2_X1 U7579 ( .A1(n6408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6409) );
  OR2_X1 U7580 ( .A1(n7320), .A2(n6872), .ZN(n6417) );
  INV_X2 U7581 ( .A(n6569), .ZN(n6985) );
  INV_X1 U7582 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U7583 ( .A1(n6411), .A2(n6412), .ZN(n6581) );
  NOR2_X1 U7584 ( .A1(n6593), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U7585 ( .A1(n6459), .A2(n8480), .ZN(n6648) );
  NAND2_X1 U7586 ( .A1(n6648), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6610) );
  INV_X1 U7587 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U7588 ( .A1(n6610), .A2(n8488), .ZN(n6413) );
  NAND2_X1 U7589 ( .A1(n6413), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6414) );
  INV_X1 U7590 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8288) );
  NAND2_X1 U7591 ( .A1(n6414), .A2(n8288), .ZN(n6630) );
  OR2_X1 U7592 ( .A1(n6414), .A2(n8288), .ZN(n6415) );
  AOI22_X1 U7593 ( .A1(n6985), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6774), .B2(
        n7531), .ZN(n6416) );
  NOR2_X2 U7594 ( .A1(n6701), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6435) );
  NAND3_X1 U7595 ( .A1(n8511), .A2(n6441), .A3(n6420), .ZN(n6421) );
  OAI21_X1 U7596 ( .B1(n6425), .B2(n6421), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6422) );
  MUX2_X1 U7597 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6422), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6423) );
  NAND2_X1 U7598 ( .A1(n6418), .A2(n6423), .ZN(n9243) );
  NAND2_X1 U7599 ( .A1(n8511), .A2(n6441), .ZN(n6424) );
  XNOR2_X1 U7600 ( .A(n6426), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U7601 ( .A1(n6418), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6427) );
  MUX2_X1 U7602 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6427), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6428) );
  NAND2_X1 U7603 ( .A1(n5163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6432) );
  AND2_X2 U7604 ( .A1(n6483), .A2(n6470), .ZN(n6586) );
  XNOR2_X2 U7605 ( .A(n6438), .B(n6437), .ZN(n8895) );
  INV_X2 U7606 ( .A(n8895), .ZN(n6773) );
  NAND2_X1 U7607 ( .A1(n6470), .A2(n6773), .ZN(n8095) );
  NAND2_X1 U7608 ( .A1(n8095), .A2(n7593), .ZN(n6445) );
  NAND2_X1 U7609 ( .A1(n6439), .A2(n8507), .ZN(n6440) );
  NAND2_X4 U7610 ( .A1(n6446), .A2(n6483), .ZN(n7257) );
  INV_X1 U7611 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6447) );
  OR2_X1 U7612 ( .A1(n6449), .A2(n6447), .ZN(n6448) );
  AND2_X2 U7613 ( .A1(n6452), .A2(n9473), .ZN(n6635) );
  NAND2_X1 U7614 ( .A1(n6635), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6458) );
  INV_X1 U7615 ( .A(n9473), .ZN(n6454) );
  AND2_X2 U7616 ( .A1(n6452), .A2(n6454), .ZN(n6543) );
  NAND2_X1 U7617 ( .A1(n6559), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6574) );
  NOR2_X1 U7618 ( .A1(n6574), .A2(n6573), .ZN(n6597) );
  NAND2_X1 U7619 ( .A1(n6597), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6599) );
  NOR2_X1 U7620 ( .A1(n6616), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U7621 ( .A1(n6995), .A2(n5681), .ZN(n6457) );
  NAND2_X1 U7622 ( .A1(n7090), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6456) );
  AND2_X2 U7623 ( .A1(n6454), .A2(n10791), .ZN(n6519) );
  NAND2_X1 U7624 ( .A1(n6576), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6455) );
  NAND4_X1 U7625 ( .A1(n6458), .A2(n6457), .A3(n6456), .A4(n6455), .ZN(n10248)
         );
  AOI22_X1 U7626 ( .A1(n8646), .A2(n6764), .B1(n6485), .B2(n10248), .ZN(n9090)
         );
  NAND2_X1 U7627 ( .A1(n7313), .A2(n5115), .ZN(n6462) );
  OR2_X1 U7628 ( .A1(n6459), .A2(n6447), .ZN(n6460) );
  XNOR2_X1 U7629 ( .A(n6460), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7487) );
  AOI22_X1 U7630 ( .A1(n6985), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6774), .B2(
        n7487), .ZN(n6461) );
  NAND2_X1 U7631 ( .A1(n6635), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6469) );
  INV_X2 U7632 ( .A(n6463), .ZN(n6995) );
  NAND2_X1 U7633 ( .A1(n6599), .A2(n6464), .ZN(n6465) );
  AND2_X1 U7634 ( .A1(n6614), .A2(n6465), .ZN(n8778) );
  NAND2_X1 U7635 ( .A1(n6995), .A2(n8778), .ZN(n6468) );
  NAND2_X1 U7636 ( .A1(n7090), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7637 ( .A1(n6576), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6466) );
  OAI22_X1 U7638 ( .A1(n8781), .A2(n7262), .B1(n8697), .B2(n7257), .ZN(n6609)
         );
  INV_X1 U7639 ( .A(n6470), .ZN(n6471) );
  NAND2_X1 U7640 ( .A1(n8564), .A2(n5113), .ZN(n6473) );
  OR2_X1 U7641 ( .A1(n8697), .A2(n7262), .ZN(n6472) );
  NAND2_X1 U7642 ( .A1(n6473), .A2(n6472), .ZN(n6474) );
  XNOR2_X1 U7643 ( .A(n6474), .B(n6885), .ZN(n6608) );
  INV_X1 U7644 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8471) );
  NOR2_X1 U7645 ( .A1(n5392), .A2(n6475), .ZN(n6476) );
  XNOR2_X1 U7646 ( .A(n6476), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10801) );
  MUX2_X1 U7647 ( .A(n8471), .B(n10801), .S(n7326), .Z(n8042) );
  INV_X1 U7648 ( .A(n8042), .ZN(n7657) );
  NAND2_X1 U7649 ( .A1(n6497), .A2(n7657), .ZN(n6482) );
  NAND2_X1 U7650 ( .A1(n6543), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U7651 ( .A1(n6635), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U7652 ( .A1(n6600), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U7653 ( .A1(n6519), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U7654 ( .A1(n10258), .A2(n6586), .ZN(n6481) );
  INV_X1 U7655 ( .A(n6483), .ZN(n6486) );
  NAND2_X1 U7656 ( .A1(n6486), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U7657 ( .A1(n10258), .A2(n6485), .ZN(n6488) );
  AOI22_X1 U7658 ( .A1(n6586), .A2(n7657), .B1(n6486), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7659 ( .A1(n6488), .A2(n6487), .ZN(n7654) );
  NAND2_X1 U7660 ( .A1(n7653), .A2(n7654), .ZN(n6491) );
  INV_X1 U7661 ( .A(n6489), .ZN(n6867) );
  NAND2_X1 U7662 ( .A1(n6491), .A2(n6490), .ZN(n6504) );
  NAND2_X1 U7663 ( .A1(n6600), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U7664 ( .A1(n5111), .A2(n6586), .ZN(n6499) );
  NAND2_X1 U7665 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6496) );
  XNOR2_X1 U7666 ( .A(n6496), .B(P1_IR_REG_1__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U7667 ( .A1(n6497), .A2(n7009), .ZN(n6498) );
  NAND2_X1 U7668 ( .A1(n6499), .A2(n6498), .ZN(n6500) );
  NAND2_X1 U7669 ( .A1(n5111), .A2(n6485), .ZN(n6502) );
  NAND2_X1 U7670 ( .A1(n6764), .A2(n7009), .ZN(n6501) );
  NAND2_X1 U7671 ( .A1(n6502), .A2(n6501), .ZN(n7941) );
  NAND2_X1 U7672 ( .A1(n6504), .A2(n6503), .ZN(n7940) );
  NAND2_X1 U7673 ( .A1(n6505), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6508) );
  OR2_X1 U7674 ( .A1(n6506), .A2(n6447), .ZN(n6527) );
  XNOR2_X1 U7675 ( .A(n6527), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U7676 ( .A1(n6635), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U7677 ( .A1(n6543), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U7678 ( .A1(n6600), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U7679 ( .A1(n6519), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6509) );
  OAI22_X1 U7680 ( .A1(n7011), .A2(n7257), .B1(n8103), .B2(n7262), .ZN(n6515)
         );
  XNOR2_X1 U7681 ( .A(n6514), .B(n6515), .ZN(n10196) );
  INV_X1 U7682 ( .A(n6514), .ZN(n6516) );
  OR2_X1 U7683 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  NAND2_X1 U7684 ( .A1(n10194), .A2(n6517), .ZN(n8590) );
  NAND2_X1 U7685 ( .A1(n6635), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6523) );
  INV_X1 U7686 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U7687 ( .A1(n7090), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6521) );
  NAND2_X1 U7688 ( .A1(n6576), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U7689 ( .A1(n10255), .A2(n6764), .ZN(n6534) );
  INV_X1 U7690 ( .A(n7298), .ZN(n6524) );
  NAND2_X1 U7691 ( .A1(n6525), .A2(n6524), .ZN(n6532) );
  NAND2_X1 U7692 ( .A1(n6505), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6531) );
  INV_X1 U7693 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U7694 ( .A1(n6527), .A2(n6526), .ZN(n6528) );
  NAND2_X1 U7695 ( .A1(n6528), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6529) );
  XNOR2_X1 U7696 ( .A(n6529), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U7697 ( .A1(n6774), .A2(n10296), .ZN(n6530) );
  NAND2_X1 U7698 ( .A1(n8748), .A2(n6497), .ZN(n6533) );
  NAND2_X1 U7699 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  XNOR2_X1 U7700 ( .A(n6535), .B(n6489), .ZN(n6540) );
  NAND2_X1 U7701 ( .A1(n10255), .A2(n6485), .ZN(n6537) );
  OR2_X1 U7702 ( .A1(n7919), .A2(n7262), .ZN(n6536) );
  NAND2_X1 U7703 ( .A1(n6537), .A2(n6536), .ZN(n6538) );
  XNOR2_X1 U7704 ( .A(n6540), .B(n6538), .ZN(n8591) );
  INV_X1 U7705 ( .A(n6538), .ZN(n6539) );
  NAND2_X1 U7706 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  NAND2_X1 U7707 ( .A1(n6635), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6547) );
  NOR2_X1 U7708 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6542) );
  NOR2_X1 U7709 ( .A1(n6559), .A2(n6542), .ZN(n8710) );
  NAND2_X1 U7710 ( .A1(n6543), .A2(n8710), .ZN(n6546) );
  NAND2_X1 U7711 ( .A1(n7090), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U7712 ( .A1(n6576), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6544) );
  AND4_X2 U7713 ( .A1(n6547), .A2(n6546), .A3(n6545), .A4(n6544), .ZN(n8634)
         );
  INV_X1 U7714 ( .A(n6548), .ZN(n7294) );
  NAND2_X1 U7715 ( .A1(n6505), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6553) );
  NOR2_X1 U7716 ( .A1(n6549), .A2(n6447), .ZN(n6550) );
  MUX2_X1 U7717 ( .A(n6447), .B(n6550), .S(P1_IR_REG_4__SCAN_IN), .Z(n6551) );
  NOR2_X1 U7718 ( .A1(n6551), .A2(n6411), .ZN(n10309) );
  NAND2_X1 U7719 ( .A1(n6774), .A2(n10309), .ZN(n6552) );
  OAI211_X1 U7720 ( .C1(n6872), .C2(n7294), .A(n6553), .B(n6552), .ZN(n8711)
         );
  OAI22_X1 U7721 ( .A1(n8634), .A2(n7262), .B1(n11036), .B2(n5112), .ZN(n6554)
         );
  XNOR2_X1 U7722 ( .A(n6554), .B(n6885), .ZN(n6557) );
  OAI22_X1 U7723 ( .A1(n8634), .A2(n7257), .B1(n11036), .B2(n7262), .ZN(n6556)
         );
  XNOR2_X1 U7724 ( .A(n6557), .B(n6556), .ZN(n8032) );
  NAND2_X1 U7725 ( .A1(n6557), .A2(n6556), .ZN(n6558) );
  NAND2_X1 U7726 ( .A1(n6839), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6563) );
  OAI21_X1 U7727 ( .B1(n6559), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6574), .ZN(
        n8639) );
  INV_X1 U7728 ( .A(n8639), .ZN(n11045) );
  NAND2_X1 U7729 ( .A1(n6995), .A2(n11045), .ZN(n6562) );
  NAND2_X1 U7730 ( .A1(n7090), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U7731 ( .A1(n6576), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6560) );
  INV_X1 U7732 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7299) );
  NOR2_X1 U7733 ( .A1(n6411), .A2(n6447), .ZN(n6564) );
  MUX2_X1 U7734 ( .A(n6447), .B(n6564), .S(P1_IR_REG_5__SCAN_IN), .Z(n6566) );
  INV_X1 U7735 ( .A(n6581), .ZN(n6565) );
  NOR2_X1 U7736 ( .A1(n6566), .A2(n6565), .ZN(n10323) );
  NAND2_X1 U7737 ( .A1(n6774), .A2(n10323), .ZN(n6567) );
  OAI211_X1 U7738 ( .C1(n6569), .C2(n7299), .A(n6568), .B(n6567), .ZN(n11046)
         );
  OAI22_X1 U7739 ( .A1(n8717), .A2(n7262), .B1(n7946), .B2(n5112), .ZN(n6570)
         );
  XNOR2_X1 U7740 ( .A(n6570), .B(n6489), .ZN(n6571) );
  OAI22_X1 U7741 ( .A1(n8717), .A2(n7257), .B1(n7946), .B2(n7262), .ZN(n8631)
         );
  NAND2_X1 U7742 ( .A1(n6572), .A2(n6571), .ZN(n8629) );
  NAND2_X1 U7743 ( .A1(n6839), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6580) );
  AND2_X1 U7744 ( .A1(n6574), .A2(n6573), .ZN(n6575) );
  NOR2_X1 U7745 ( .A1(n6597), .A2(n6575), .ZN(n8650) );
  NAND2_X1 U7746 ( .A1(n6995), .A2(n8650), .ZN(n6579) );
  NAND2_X1 U7747 ( .A1(n7090), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U7748 ( .A1(n6576), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6577) );
  INV_X1 U7749 ( .A(n8698), .ZN(n10252) );
  OR2_X1 U7750 ( .A1(n7309), .A2(n6872), .ZN(n6584) );
  NAND2_X1 U7751 ( .A1(n6581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6582) );
  XNOR2_X1 U7752 ( .A(n6582), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U7753 ( .A1(n6985), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6774), .B2(
        n10336), .ZN(n6583) );
  NAND2_X1 U7754 ( .A1(n6584), .A2(n6583), .ZN(n8651) );
  AOI22_X1 U7755 ( .A1(n10252), .A2(n6764), .B1(n8651), .B2(n5113), .ZN(n6585)
         );
  XNOR2_X1 U7756 ( .A(n6585), .B(n6867), .ZN(n8606) );
  OR2_X1 U7757 ( .A1(n8698), .A2(n7257), .ZN(n6588) );
  NAND2_X1 U7759 ( .A1(n8651), .A2(n6764), .ZN(n6587) );
  NAND2_X1 U7760 ( .A1(n6588), .A2(n6587), .ZN(n6589) );
  INV_X1 U7761 ( .A(n6589), .ZN(n8605) );
  INV_X1 U7762 ( .A(n8606), .ZN(n6590) );
  NAND2_X1 U7763 ( .A1(n6590), .A2(n6589), .ZN(n6591) );
  OR2_X1 U7764 ( .A1(n7312), .A2(n6872), .ZN(n6596) );
  NAND2_X1 U7765 ( .A1(n6593), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6594) );
  XNOR2_X1 U7766 ( .A(n6594), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U7767 ( .A1(n6985), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6774), .B2(
        n10349), .ZN(n6595) );
  NAND2_X1 U7768 ( .A1(n6839), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6604) );
  OR2_X1 U7769 ( .A1(n6597), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6598) );
  AND2_X1 U7770 ( .A1(n6599), .A2(n6598), .ZN(n8702) );
  NAND2_X1 U7771 ( .A1(n6995), .A2(n8702), .ZN(n6603) );
  NAND2_X1 U7772 ( .A1(n7090), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U7773 ( .A1(n6576), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6601) );
  NAND4_X1 U7774 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n10251)
         );
  AOI22_X1 U7775 ( .A1(n8701), .A2(n5113), .B1(n6764), .B2(n10251), .ZN(n6605)
         );
  XOR2_X1 U7776 ( .A(n6885), .B(n6605), .Z(n6607) );
  INV_X1 U7777 ( .A(n10251), .ZN(n8776) );
  OAI22_X1 U7778 ( .A1(n8110), .A2(n7262), .B1(n8776), .B2(n7257), .ZN(n6606)
         );
  NAND2_X1 U7779 ( .A1(n6607), .A2(n6606), .ZN(n8694) );
  XOR2_X1 U7780 ( .A(n6609), .B(n6608), .Z(n8771) );
  NAND2_X1 U7781 ( .A1(n7321), .A2(n5115), .ZN(n6612) );
  XNOR2_X1 U7782 ( .A(n6610), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7503) );
  AOI22_X1 U7783 ( .A1(n6985), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6774), .B2(
        n7503), .ZN(n6611) );
  NAND2_X1 U7784 ( .A1(n6612), .A2(n6611), .ZN(n8673) );
  INV_X1 U7785 ( .A(n8673), .ZN(n11073) );
  NAND2_X1 U7786 ( .A1(n6635), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6620) );
  AND2_X1 U7787 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  NOR2_X1 U7788 ( .A1(n6616), .A2(n6615), .ZN(n8833) );
  NAND2_X1 U7789 ( .A1(n6995), .A2(n8833), .ZN(n6619) );
  NAND2_X1 U7790 ( .A1(n7090), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U7791 ( .A1(n6576), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6617) );
  OAI22_X1 U7792 ( .A1(n11073), .A2(n7262), .B1(n8121), .B2(n7257), .ZN(n6625)
         );
  NAND2_X1 U7793 ( .A1(n8673), .A2(n5113), .ZN(n6622) );
  OR2_X1 U7794 ( .A1(n8121), .A2(n7262), .ZN(n6621) );
  NAND2_X1 U7795 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  XNOR2_X1 U7796 ( .A(n6623), .B(n6867), .ZN(n6624) );
  XOR2_X1 U7797 ( .A(n6625), .B(n6624), .Z(n8826) );
  INV_X1 U7798 ( .A(n6624), .ZN(n6627) );
  INV_X1 U7799 ( .A(n6625), .ZN(n6626) );
  AOI22_X1 U7800 ( .A1(n8646), .A2(n5113), .B1(n6764), .B2(n10248), .ZN(n6628)
         );
  XOR2_X1 U7801 ( .A(n6867), .B(n6628), .Z(n6629) );
  NAND2_X1 U7802 ( .A1(n6630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6631) );
  XNOR2_X1 U7803 ( .A(n6631), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7517) );
  AOI22_X1 U7804 ( .A1(n6985), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6774), .B2(
        n7517), .ZN(n6632) );
  NAND2_X1 U7805 ( .A1(n6633), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6654) );
  OR2_X1 U7806 ( .A1(n6633), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6634) );
  AND2_X1 U7807 ( .A1(n6654), .A2(n6634), .ZN(n9067) );
  NAND2_X1 U7808 ( .A1(n6995), .A2(n9067), .ZN(n6639) );
  NAND2_X1 U7809 ( .A1(n6635), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U7810 ( .A1(n7090), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U7811 ( .A1(n6576), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6636) );
  NAND4_X1 U7812 ( .A1(n6639), .A2(n6638), .A3(n6637), .A4(n6636), .ZN(n10247)
         );
  OAI22_X1 U7813 ( .A1(n9064), .A2(n5112), .B1(n8727), .B2(n7262), .ZN(n6640)
         );
  XNOR2_X1 U7814 ( .A(n6640), .B(n6489), .ZN(n9058) );
  OR2_X1 U7815 ( .A1(n9064), .A2(n7262), .ZN(n6642) );
  NAND2_X1 U7816 ( .A1(n10247), .A2(n6485), .ZN(n6641) );
  AND2_X1 U7817 ( .A1(n6642), .A2(n6641), .ZN(n6643) );
  NAND2_X1 U7818 ( .A1(n9058), .A2(n6643), .ZN(n6645) );
  INV_X1 U7819 ( .A(n9058), .ZN(n6644) );
  INV_X1 U7820 ( .A(n6643), .ZN(n9057) );
  OR2_X1 U7821 ( .A1(n7468), .A2(n6872), .ZN(n6652) );
  INV_X1 U7822 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8292) );
  NAND3_X1 U7823 ( .A1(n8292), .A2(n8488), .A3(n8288), .ZN(n6647) );
  OAI21_X1 U7824 ( .B1(n6648), .B2(n6647), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6649) );
  MUX2_X1 U7825 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6649), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n6650) );
  AND2_X1 U7826 ( .A1(n6646), .A2(n6650), .ZN(n7669) );
  AOI22_X1 U7827 ( .A1(n6985), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6774), .B2(
        n7669), .ZN(n6651) );
  INV_X2 U7828 ( .A(n6990), .ZN(n6839) );
  NAND2_X1 U7829 ( .A1(n6839), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U7830 ( .A1(n6654), .A2(n6653), .ZN(n6655) );
  AND2_X1 U7831 ( .A1(n6667), .A2(n6655), .ZN(n9193) );
  NAND2_X1 U7832 ( .A1(n6995), .A2(n9193), .ZN(n6658) );
  NAND2_X1 U7833 ( .A1(n7090), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6657) );
  NAND2_X1 U7834 ( .A1(n6576), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6656) );
  AOI22_X1 U7835 ( .A1(n8854), .A2(n5113), .B1(n6764), .B2(n10246), .ZN(n6660)
         );
  XNOR2_X1 U7836 ( .A(n6660), .B(n6867), .ZN(n6679) );
  OAI22_X1 U7837 ( .A1(n11089), .A2(n7262), .B1(n9063), .B2(n7257), .ZN(n6677)
         );
  XNOR2_X1 U7838 ( .A(n6679), .B(n6677), .ZN(n9187) );
  OR2_X1 U7839 ( .A1(n7549), .A2(n6872), .ZN(n6665) );
  NAND2_X1 U7840 ( .A1(n6646), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6662) );
  MUX2_X1 U7841 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6662), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6663) );
  AND2_X1 U7842 ( .A1(n6661), .A2(n6663), .ZN(n10370) );
  AOI22_X1 U7843 ( .A1(n6985), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6774), .B2(
        n10370), .ZN(n6664) );
  NAND2_X1 U7844 ( .A1(n9006), .A2(n5113), .ZN(n6674) );
  NAND2_X1 U7845 ( .A1(n7090), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6672) );
  INV_X1 U7846 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U7847 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  AND2_X1 U7848 ( .A1(n6690), .A2(n6668), .ZN(n10181) );
  NAND2_X1 U7849 ( .A1(n6995), .A2(n10181), .ZN(n6671) );
  NAND2_X1 U7850 ( .A1(n6839), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U7851 ( .A1(n6576), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6669) );
  OR2_X1 U7852 ( .A1(n9191), .A2(n7262), .ZN(n6673) );
  NAND2_X1 U7853 ( .A1(n6674), .A2(n6673), .ZN(n6675) );
  XNOR2_X1 U7854 ( .A(n6675), .B(n6867), .ZN(n6681) );
  NOR2_X1 U7855 ( .A1(n9191), .A2(n7257), .ZN(n6676) );
  AOI21_X1 U7856 ( .B1(n9006), .B2(n6764), .A(n6676), .ZN(n6682) );
  XNOR2_X1 U7857 ( .A(n6681), .B(n6682), .ZN(n10174) );
  INV_X1 U7858 ( .A(n6677), .ZN(n6678) );
  NAND2_X1 U7859 ( .A1(n6679), .A2(n6678), .ZN(n10175) );
  INV_X1 U7860 ( .A(n6681), .ZN(n6683) );
  NOR2_X1 U7861 ( .A1(n6683), .A2(n6682), .ZN(n6700) );
  NAND2_X1 U7862 ( .A1(n7574), .A2(n5115), .ZN(n6688) );
  NAND2_X1 U7863 ( .A1(n6661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6684) );
  MUX2_X1 U7864 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6684), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6686) );
  NAND2_X1 U7865 ( .A1(n6686), .A2(n6685), .ZN(n8073) );
  AOI22_X1 U7866 ( .A1(n6985), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6774), .B2(
        n8065), .ZN(n6687) );
  NAND2_X1 U7867 ( .A1(n10729), .A2(n5113), .ZN(n6697) );
  NAND2_X1 U7868 ( .A1(n6839), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6695) );
  AND2_X1 U7869 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  NOR2_X1 U7870 ( .A1(n6706), .A2(n6691), .ZN(n10097) );
  NAND2_X1 U7871 ( .A1(n6995), .A2(n10097), .ZN(n6694) );
  NAND2_X1 U7872 ( .A1(n7090), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U7873 ( .A1(n6576), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6692) );
  OR2_X1 U7874 ( .A1(n10179), .A2(n7262), .ZN(n6696) );
  NAND2_X1 U7875 ( .A1(n6697), .A2(n6696), .ZN(n6698) );
  XNOR2_X1 U7876 ( .A(n6698), .B(n6885), .ZN(n6699) );
  AOI22_X1 U7877 ( .A1(n10729), .A2(n6764), .B1(n6485), .B2(n10720), .ZN(
        n10092) );
  NAND2_X1 U7878 ( .A1(n6685), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6702) );
  MUX2_X1 U7879 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6702), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6703) );
  AND2_X1 U7880 ( .A1(n6701), .A2(n6703), .ZN(n8080) );
  AOI22_X1 U7881 ( .A1(n6985), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6774), .B2(
        n8080), .ZN(n6704) );
  NAND2_X1 U7882 ( .A1(n6839), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6711) );
  OR2_X1 U7883 ( .A1(n6706), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U7884 ( .A1(n6706), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6723) );
  AND2_X1 U7885 ( .A1(n6707), .A2(n6723), .ZN(n10240) );
  NAND2_X1 U7886 ( .A1(n6995), .A2(n10240), .ZN(n6710) );
  NAND2_X1 U7887 ( .A1(n7090), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U7888 ( .A1(n6576), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6708) );
  NAND4_X1 U7889 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n10730)
         );
  AOI22_X1 U7890 ( .A1(n9053), .A2(n5113), .B1(n6586), .B2(n10730), .ZN(n6712)
         );
  XOR2_X1 U7891 ( .A(n6885), .B(n6712), .Z(n6715) );
  NAND2_X1 U7892 ( .A1(n6714), .A2(n6715), .ZN(n10229) );
  INV_X1 U7893 ( .A(n10730), .ZN(n10138) );
  OAI22_X1 U7894 ( .A1(n10723), .A2(n7262), .B1(n10138), .B2(n7257), .ZN(n6713) );
  INV_X1 U7895 ( .A(n6713), .ZN(n10231) );
  NAND2_X1 U7896 ( .A1(n10229), .A2(n10231), .ZN(n6718) );
  INV_X1 U7897 ( .A(n6715), .ZN(n6716) );
  NAND2_X1 U7898 ( .A1(n6717), .A2(n6716), .ZN(n10230) );
  NAND2_X1 U7899 ( .A1(n7819), .A2(n5115), .ZN(n6721) );
  NAND2_X1 U7900 ( .A1(n6701), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6719) );
  XNOR2_X1 U7901 ( .A(n6719), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8761) );
  AOI22_X1 U7902 ( .A1(n6985), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6774), .B2(
        n8761), .ZN(n6720) );
  NAND2_X1 U7903 ( .A1(n6839), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6728) );
  INV_X1 U7904 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U7905 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  AND2_X1 U7906 ( .A1(n6739), .A2(n6724), .ZN(n10140) );
  NAND2_X1 U7907 ( .A1(n6995), .A2(n10140), .ZN(n6727) );
  NAND2_X1 U7908 ( .A1(n7090), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6726) );
  NAND2_X1 U7909 ( .A1(n6576), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6725) );
  NAND4_X1 U7910 ( .A1(n6728), .A2(n6727), .A3(n6726), .A4(n6725), .ZN(n10719)
         );
  OAI22_X1 U7911 ( .A1(n10714), .A2(n5112), .B1(n10703), .B2(n7262), .ZN(n6729) );
  XNOR2_X1 U7912 ( .A(n6729), .B(n6867), .ZN(n6733) );
  OR2_X1 U7913 ( .A1(n10714), .A2(n7262), .ZN(n6731) );
  NAND2_X1 U7914 ( .A1(n10719), .A2(n6485), .ZN(n6730) );
  NAND2_X1 U7915 ( .A1(n6731), .A2(n6730), .ZN(n6732) );
  NOR2_X1 U7916 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  AOI21_X1 U7917 ( .B1(n6733), .B2(n6732), .A(n6734), .ZN(n10134) );
  INV_X1 U7918 ( .A(n6734), .ZN(n10143) );
  NAND2_X1 U7919 ( .A1(n8037), .A2(n5115), .ZN(n6737) );
  XNOR2_X1 U7920 ( .A(n6735), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8872) );
  AOI22_X1 U7921 ( .A1(n6985), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6774), .B2(
        n8872), .ZN(n6736) );
  NAND2_X1 U7922 ( .A1(n10706), .A2(n5113), .ZN(n6746) );
  INV_X1 U7923 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6738) );
  AND2_X1 U7924 ( .A1(n6739), .A2(n6738), .ZN(n6740) );
  NOR2_X1 U7925 ( .A1(n6758), .A2(n6740), .ZN(n10152) );
  NAND2_X1 U7926 ( .A1(n10152), .A2(n6995), .ZN(n6744) );
  NAND2_X1 U7927 ( .A1(n6839), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6743) );
  NAND2_X1 U7928 ( .A1(n7090), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U7929 ( .A1(n6576), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6741) );
  OR2_X1 U7930 ( .A1(n9219), .A2(n7262), .ZN(n6745) );
  NAND2_X1 U7931 ( .A1(n6746), .A2(n6745), .ZN(n6747) );
  XNOR2_X1 U7932 ( .A(n6747), .B(n6489), .ZN(n6768) );
  NOR2_X1 U7933 ( .A1(n9219), .A2(n7257), .ZN(n6748) );
  AOI21_X1 U7934 ( .B1(n10706), .B2(n6764), .A(n6748), .ZN(n6767) );
  NAND2_X1 U7935 ( .A1(n6768), .A2(n6767), .ZN(n10144) );
  AND2_X1 U7936 ( .A1(n10143), .A2(n10144), .ZN(n6771) );
  OR2_X1 U7937 ( .A1(n8054), .A2(n6872), .ZN(n6757) );
  INV_X1 U7938 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U7939 ( .A1(n6735), .A2(n6749), .ZN(n6750) );
  AND2_X1 U7940 ( .A1(n6750), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U7941 ( .A1(n6751), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6755) );
  AND2_X1 U7942 ( .A1(n6753), .A2(n6752), .ZN(n6754) );
  AND2_X1 U7943 ( .A1(n6755), .A2(n6754), .ZN(n8877) );
  AOI22_X1 U7944 ( .A1(n6985), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6774), .B2(
        n8877), .ZN(n6756) );
  NOR2_X1 U7945 ( .A1(n6758), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6759) );
  OR2_X1 U7946 ( .A1(n6777), .A2(n6759), .ZN(n10213) );
  NAND2_X1 U7947 ( .A1(n7090), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U7948 ( .A1(n6519), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6760) );
  AND2_X1 U7949 ( .A1(n6761), .A2(n6760), .ZN(n6763) );
  NAND2_X1 U7950 ( .A1(n6839), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6762) );
  OAI211_X1 U7951 ( .C1(n10213), .C2(n6463), .A(n6763), .B(n6762), .ZN(n10587)
         );
  AOI22_X1 U7952 ( .A1(n10406), .A2(n5113), .B1(n6764), .B2(n10587), .ZN(n6765) );
  XNOR2_X1 U7953 ( .A(n6765), .B(n6867), .ZN(n6772) );
  INV_X1 U7954 ( .A(n6772), .ZN(n6766) );
  AND2_X1 U7955 ( .A1(n6771), .A2(n6766), .ZN(n6769) );
  OR2_X1 U7956 ( .A1(n6768), .A2(n6767), .ZN(n10145) );
  AOI22_X1 U7957 ( .A1(n10406), .A2(n6764), .B1(n6485), .B2(n10587), .ZN(
        n10206) );
  INV_X1 U7958 ( .A(n10145), .ZN(n6770) );
  NAND2_X1 U7959 ( .A1(n8690), .A2(n5115), .ZN(n6776) );
  AOI22_X1 U7960 ( .A1(n6985), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6773), .B2(
        n6774), .ZN(n6775) );
  NAND2_X1 U7961 ( .A1(n10593), .A2(n5113), .ZN(n6783) );
  OR2_X1 U7962 ( .A1(n6777), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U7963 ( .A1(n6777), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6793) );
  AND2_X1 U7964 ( .A1(n6778), .A2(n6793), .ZN(n10595) );
  NAND2_X1 U7965 ( .A1(n10595), .A2(n6995), .ZN(n6781) );
  AOI22_X1 U7966 ( .A1(n6519), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n7090), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n6780) );
  NAND2_X1 U7967 ( .A1(n6839), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6779) );
  OR2_X1 U7968 ( .A1(n10209), .A2(n7262), .ZN(n6782) );
  NAND2_X1 U7969 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  XNOR2_X1 U7970 ( .A(n6784), .B(n6867), .ZN(n6787) );
  AOI22_X1 U7971 ( .A1(n10593), .A2(n6586), .B1(n6485), .B2(n10694), .ZN(n6785) );
  XNOR2_X1 U7972 ( .A(n6787), .B(n6785), .ZN(n10110) );
  INV_X1 U7973 ( .A(n6785), .ZN(n6786) );
  NAND2_X1 U7974 ( .A1(n6789), .A2(n6788), .ZN(n10165) );
  NAND2_X1 U7975 ( .A1(n8850), .A2(n5115), .ZN(n6791) );
  NAND2_X1 U7976 ( .A1(n6985), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U7977 ( .A1(n10684), .A2(n5113), .ZN(n6801) );
  NAND2_X1 U7978 ( .A1(n6839), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6799) );
  INV_X1 U7979 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6792) );
  NAND2_X1 U7980 ( .A1(n6792), .A2(n6793), .ZN(n6795) );
  INV_X1 U7981 ( .A(n6793), .ZN(n6794) );
  INV_X1 U7982 ( .A(n6809), .ZN(n6811) );
  AND2_X1 U7983 ( .A1(n6795), .A2(n6811), .ZN(n10572) );
  NAND2_X1 U7984 ( .A1(n6995), .A2(n10572), .ZN(n6798) );
  NAND2_X1 U7985 ( .A1(n7090), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U7986 ( .A1(n6519), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6796) );
  NAND4_X1 U7987 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(n10586)
         );
  NAND2_X1 U7988 ( .A1(n10586), .A2(n6586), .ZN(n6800) );
  NAND2_X1 U7989 ( .A1(n6801), .A2(n6800), .ZN(n6802) );
  XNOR2_X1 U7990 ( .A(n6802), .B(n6885), .ZN(n6803) );
  AOI22_X1 U7991 ( .A1(n10684), .A2(n6586), .B1(n6485), .B2(n10586), .ZN(n6804) );
  XNOR2_X1 U7992 ( .A(n6803), .B(n6804), .ZN(n10166) );
  INV_X1 U7993 ( .A(n6803), .ZN(n6805) );
  NAND2_X1 U7994 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  NAND2_X1 U7995 ( .A1(n6985), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6807) );
  NAND2_X1 U7996 ( .A1(n6839), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6816) );
  INV_X1 U7997 ( .A(n6825), .ZN(n6827) );
  INV_X1 U7998 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U7999 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  AND2_X1 U8000 ( .A1(n6827), .A2(n6812), .ZN(n10562) );
  NAND2_X1 U8001 ( .A1(n6995), .A2(n10562), .ZN(n6815) );
  NAND2_X1 U8002 ( .A1(n7090), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U8003 ( .A1(n6519), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6813) );
  OAI22_X1 U8004 ( .A1(n10772), .A2(n7262), .B1(n10669), .B2(n7257), .ZN(n6820) );
  AOI22_X1 U8005 ( .A1(n10561), .A2(n5113), .B1(n6586), .B2(n10577), .ZN(n6817) );
  XNOR2_X1 U8006 ( .A(n6817), .B(n6867), .ZN(n6819) );
  XOR2_X1 U8007 ( .A(n6820), .B(n6819), .Z(n10118) );
  INV_X1 U8008 ( .A(n10118), .ZN(n6818) );
  INV_X1 U8009 ( .A(n6819), .ZN(n6821) );
  NAND2_X1 U8010 ( .A1(n6821), .A2(n6820), .ZN(n6822) );
  NAND2_X1 U8011 ( .A1(n10119), .A2(n6822), .ZN(n6835) );
  OR2_X1 U8012 ( .A1(n9113), .A2(n6872), .ZN(n6824) );
  NAND2_X1 U8013 ( .A1(n6985), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6823) );
  NAND2_X1 U8014 ( .A1(n6839), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6832) );
  INV_X1 U8015 ( .A(n6840), .ZN(n6842) );
  INV_X1 U8016 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U8017 ( .A1(n6827), .A2(n6826), .ZN(n6828) );
  AND2_X1 U8018 ( .A1(n6842), .A2(n6828), .ZN(n10537) );
  NAND2_X1 U8019 ( .A1(n6995), .A2(n10537), .ZN(n6831) );
  NAND2_X1 U8020 ( .A1(n7090), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6830) );
  NAND2_X1 U8021 ( .A1(n6519), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6829) );
  NAND4_X1 U8022 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n10658)
         );
  AOI22_X1 U8023 ( .A1(n10545), .A2(n5113), .B1(n6586), .B2(n10658), .ZN(n6833) );
  XOR2_X1 U8024 ( .A(n6867), .B(n6833), .Z(n6834) );
  OR2_X2 U8025 ( .A1(n6835), .A2(n6834), .ZN(n10186) );
  OAI22_X1 U8026 ( .A1(n10768), .A2(n7262), .B1(n10559), .B2(n7257), .ZN(
        n10188) );
  NAND2_X1 U8027 ( .A1(n6835), .A2(n6834), .ZN(n10185) );
  NAND2_X1 U8028 ( .A1(n9134), .A2(n5115), .ZN(n6838) );
  NAND2_X1 U8029 ( .A1(n6985), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U8030 ( .A1(n6839), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6847) );
  INV_X1 U8031 ( .A(n6858), .ZN(n6860) );
  INV_X1 U8032 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U8033 ( .A1(n6842), .A2(n6841), .ZN(n6843) );
  NAND2_X1 U8034 ( .A1(n6995), .A2(n10522), .ZN(n6846) );
  NAND2_X1 U8035 ( .A1(n7090), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U8036 ( .A1(n6519), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6844) );
  OAI22_X1 U8037 ( .A1(n10764), .A2(n7262), .B1(n10668), .B2(n7257), .ZN(n6852) );
  NAND2_X1 U8038 ( .A1(n10529), .A2(n5113), .ZN(n6849) );
  OR2_X1 U8039 ( .A1(n10668), .A2(n7262), .ZN(n6848) );
  NAND2_X1 U8040 ( .A1(n6849), .A2(n6848), .ZN(n6850) );
  XNOR2_X1 U8041 ( .A(n6850), .B(n6867), .ZN(n6851) );
  XOR2_X1 U8042 ( .A(n6852), .B(n6851), .Z(n10103) );
  INV_X1 U8043 ( .A(n6851), .ZN(n6854) );
  INV_X1 U8044 ( .A(n6852), .ZN(n6853) );
  NAND2_X1 U8045 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  NAND2_X1 U8046 ( .A1(n9232), .A2(n5115), .ZN(n6857) );
  NAND2_X1 U8047 ( .A1(n6985), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8048 ( .A1(n6635), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U8049 ( .A1(n7090), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6864) );
  INV_X1 U8050 ( .A(n6875), .ZN(n6877) );
  INV_X1 U8051 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8052 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  NAND2_X1 U8053 ( .A1(n6995), .A2(n10508), .ZN(n6863) );
  NAND2_X1 U8054 ( .A1(n6519), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6862) );
  AOI22_X1 U8055 ( .A1(n10654), .A2(n5113), .B1(n6586), .B2(n10659), .ZN(n6866) );
  XOR2_X1 U8056 ( .A(n6867), .B(n6866), .Z(n6868) );
  INV_X1 U8057 ( .A(n10654), .ZN(n10510) );
  OAI22_X1 U8058 ( .A1(n10510), .A2(n7262), .B1(n10644), .B2(n7257), .ZN(n6869) );
  NAND2_X1 U8059 ( .A1(n6868), .A2(n6869), .ZN(n10157) );
  INV_X1 U8060 ( .A(n6868), .ZN(n6871) );
  INV_X1 U8061 ( .A(n6869), .ZN(n6870) );
  NAND2_X1 U8062 ( .A1(n6871), .A2(n6870), .ZN(n10156) );
  NAND2_X1 U8063 ( .A1(n6985), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U8064 ( .A1(n6635), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6882) );
  INV_X1 U8065 ( .A(n6889), .ZN(n6891) );
  INV_X1 U8066 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U8067 ( .A1(n6877), .A2(n6876), .ZN(n6878) );
  NAND2_X1 U8068 ( .A1(n6995), .A2(n10497), .ZN(n6881) );
  NAND2_X1 U8069 ( .A1(n7090), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U8070 ( .A1(n6519), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6879) );
  OAI22_X1 U8071 ( .A1(n10496), .A2(n7262), .B1(n10634), .B2(n7257), .ZN(n6901) );
  NAND2_X1 U8072 ( .A1(n10647), .A2(n5113), .ZN(n6884) );
  OR2_X1 U8073 ( .A1(n10634), .A2(n7262), .ZN(n6883) );
  NAND2_X1 U8074 ( .A1(n6884), .A2(n6883), .ZN(n6886) );
  XNOR2_X1 U8075 ( .A(n6886), .B(n6885), .ZN(n6902) );
  XOR2_X1 U8076 ( .A(n6901), .B(n6902), .Z(n10126) );
  NAND2_X1 U8077 ( .A1(n10085), .A2(n5115), .ZN(n6888) );
  NAND2_X1 U8078 ( .A1(n6505), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8079 ( .A1(n10487), .A2(n5113), .ZN(n6898) );
  NAND2_X1 U8080 ( .A1(n7090), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8081 ( .A1(n6635), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6895) );
  INV_X1 U8082 ( .A(n6906), .ZN(n6908) );
  INV_X1 U8083 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U8084 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  NAND2_X1 U8085 ( .A1(n6995), .A2(n10481), .ZN(n6894) );
  NAND2_X1 U8086 ( .A1(n6519), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6893) );
  OR2_X1 U8087 ( .A1(n10643), .A2(n7262), .ZN(n6897) );
  NAND2_X1 U8088 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  XNOR2_X1 U8089 ( .A(n6899), .B(n6489), .ZN(n6923) );
  NOR2_X1 U8090 ( .A1(n10643), .A2(n7257), .ZN(n6900) );
  AOI21_X1 U8091 ( .B1(n10487), .B2(n6586), .A(n6900), .ZN(n6922) );
  XNOR2_X1 U8092 ( .A(n6923), .B(n6922), .ZN(n10219) );
  NOR2_X1 U8093 ( .A1(n6902), .A2(n6901), .ZN(n10220) );
  NOR2_X1 U8094 ( .A1(n10219), .A2(n10220), .ZN(n6903) );
  NAND2_X1 U8095 ( .A1(n10081), .A2(n5115), .ZN(n6905) );
  NAND2_X1 U8096 ( .A1(n6505), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6904) );
  NAND2_X2 U8097 ( .A1(n6905), .A2(n6904), .ZN(n10752) );
  NAND2_X1 U8098 ( .A1(n10752), .A2(n5113), .ZN(n6915) );
  NAND2_X1 U8099 ( .A1(n6635), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U8100 ( .A1(n6906), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6994) );
  INV_X1 U8101 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U8102 ( .A1(n6908), .A2(n6907), .ZN(n6909) );
  NAND2_X1 U8103 ( .A1(n6995), .A2(n10465), .ZN(n6912) );
  NAND2_X1 U8104 ( .A1(n6600), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U8105 ( .A1(n6519), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6910) );
  OR2_X1 U8106 ( .A1(n10633), .A2(n7262), .ZN(n6914) );
  NAND2_X1 U8107 ( .A1(n6915), .A2(n6914), .ZN(n6916) );
  XNOR2_X1 U8108 ( .A(n6916), .B(n6489), .ZN(n6919) );
  INV_X1 U8109 ( .A(n6919), .ZN(n6921) );
  NOR2_X1 U8110 ( .A1(n10633), .A2(n7257), .ZN(n6917) );
  AOI21_X1 U8111 ( .B1(n10752), .B2(n6764), .A(n6917), .ZN(n6918) );
  INV_X1 U8112 ( .A(n6918), .ZN(n6920) );
  AOI21_X1 U8113 ( .B1(n6921), .B2(n6920), .A(n7268), .ZN(n6927) );
  INV_X1 U8114 ( .A(n6927), .ZN(n6925) );
  OR2_X1 U8115 ( .A1(n6923), .A2(n6922), .ZN(n6928) );
  INV_X1 U8116 ( .A(n6928), .ZN(n6924) );
  NOR2_X1 U8117 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  AOI21_X1 U8118 ( .B1(n10222), .B2(n6928), .A(n6927), .ZN(n6950) );
  NAND2_X1 U8119 ( .A1(n9243), .A2(P1_B_REG_SCAN_IN), .ZN(n6930) );
  MUX2_X1 U8120 ( .A(n6930), .B(P1_B_REG_SCAN_IN), .S(n6929), .Z(n6931) );
  OAI22_X1 U8121 ( .A1(n10804), .A2(P1_D_REG_0__SCAN_IN), .B1(n6929), .B2(
        n10797), .ZN(n8039) );
  NOR4_X1 U8122 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6940) );
  NOR4_X1 U8123 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6939) );
  INV_X1 U8124 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10805) );
  INV_X1 U8125 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10807) );
  INV_X1 U8126 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10808) );
  INV_X1 U8127 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10806) );
  NAND4_X1 U8128 ( .A1(n10805), .A2(n10807), .A3(n10808), .A4(n10806), .ZN(
        n6937) );
  NOR4_X1 U8129 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6935) );
  NOR4_X1 U8130 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6934) );
  NOR4_X1 U8131 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6933) );
  NOR4_X1 U8132 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6932) );
  NAND4_X1 U8133 ( .A1(n6935), .A2(n6934), .A3(n6933), .A4(n6932), .ZN(n6936)
         );
  NOR4_X1 U8134 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        n6937), .A4(n6936), .ZN(n6938) );
  AND3_X1 U8135 ( .A1(n6940), .A2(n6939), .A3(n6938), .ZN(n6941) );
  NOR2_X1 U8136 ( .A1(n8039), .A2(n7610), .ZN(n6943) );
  OAI22_X1 U8137 ( .A1(n10804), .A2(P1_D_REG_1__SCAN_IN), .B1(n6942), .B2(
        n10797), .ZN(n7612) );
  INV_X1 U8138 ( .A(n7612), .ZN(n10784) );
  INV_X1 U8139 ( .A(n7599), .ZN(n6958) );
  INV_X1 U8140 ( .A(n7593), .ZN(n6948) );
  AND3_X1 U8141 ( .A1(n10803), .A2(n6958), .A3(n11088), .ZN(n6949) );
  OAI21_X1 U8142 ( .B1(n7277), .B2(n6950), .A(n10223), .ZN(n6971) );
  NOR2_X1 U8143 ( .A1(n8043), .A2(n8920), .ZN(n8099) );
  NAND2_X1 U8144 ( .A1(n10803), .A2(n8099), .ZN(n6952) );
  OR2_X1 U8145 ( .A1(n6963), .A2(n6952), .ZN(n6953) );
  NAND2_X1 U8146 ( .A1(n7090), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6957) );
  NAND2_X1 U8147 ( .A1(n6635), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6956) );
  XNOR2_X1 U8148 ( .A(n6994), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n10456) );
  NAND2_X1 U8149 ( .A1(n6995), .A2(n10456), .ZN(n6955) );
  NAND2_X1 U8150 ( .A1(n6519), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6954) );
  NOR2_X1 U8151 ( .A1(n6958), .A2(n7593), .ZN(n8045) );
  NAND2_X1 U8152 ( .A1(n10803), .A2(n8045), .ZN(n7254) );
  INV_X1 U8153 ( .A(n6961), .ZN(n6960) );
  NOR2_X2 U8154 ( .A1(n6961), .A2(n10271), .ZN(n10233) );
  AOI22_X1 U8155 ( .A1(n10233), .A2(n10464), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n6968) );
  INV_X1 U8156 ( .A(n6962), .ZN(n7611) );
  NAND2_X1 U8157 ( .A1(n6963), .A2(n7611), .ZN(n6964) );
  NAND2_X1 U8158 ( .A1(n7599), .A2(n7593), .ZN(n7608) );
  NAND2_X1 U8159 ( .A1(n6964), .A2(n7608), .ZN(n7655) );
  NAND2_X1 U8160 ( .A1(n7325), .A2(n6483), .ZN(n6965) );
  OR2_X1 U8161 ( .A1(n7655), .A2(n6965), .ZN(n6966) );
  NAND2_X1 U8162 ( .A1(n10241), .A2(n10465), .ZN(n6967) );
  OAI211_X1 U8163 ( .C1(n10626), .C2(n10236), .A(n6968), .B(n6967), .ZN(n6969)
         );
  AOI21_X1 U8164 ( .B1(n10752), .B2(n10215), .A(n6969), .ZN(n6970) );
  NAND2_X1 U8165 ( .A1(n6971), .A2(n6970), .ZN(P1_U3214) );
  NAND2_X1 U8166 ( .A1(n6972), .A2(SI_29_), .ZN(n6977) );
  INV_X1 U8167 ( .A(n6973), .ZN(n6975) );
  NAND2_X1 U8168 ( .A1(n6975), .A2(n6974), .ZN(n6976) );
  INV_X1 U8169 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9470) );
  INV_X1 U8170 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9475) );
  MUX2_X1 U8171 ( .A(n9470), .B(n9475), .S(n7287), .Z(n6978) );
  INV_X1 U8172 ( .A(SI_30_), .ZN(n8139) );
  NAND2_X1 U8173 ( .A1(n6978), .A2(n8139), .ZN(n6981) );
  INV_X1 U8174 ( .A(n6978), .ZN(n6979) );
  NAND2_X1 U8175 ( .A1(n6979), .A2(SI_30_), .ZN(n6980) );
  NAND2_X1 U8176 ( .A1(n6981), .A2(n6980), .ZN(n7087) );
  MUX2_X1 U8177 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7287), .Z(n6982) );
  INV_X1 U8178 ( .A(SI_31_), .ZN(n8335) );
  XNOR2_X1 U8179 ( .A(n6982), .B(n8335), .ZN(n6983) );
  XNOR2_X2 U8180 ( .A(n6984), .B(n6983), .ZN(n10067) );
  NAND2_X1 U8181 ( .A1(n10067), .A2(n5115), .ZN(n6987) );
  NAND2_X1 U8182 ( .A1(n6985), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6986) );
  INV_X1 U8183 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U8184 ( .A1(n6519), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6989) );
  NAND2_X1 U8185 ( .A1(n7090), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6988) );
  OAI211_X1 U8186 ( .C1(n6990), .C2(n10607), .A(n6989), .B(n6988), .ZN(n10383)
         );
  INV_X1 U8187 ( .A(n10383), .ZN(n7102) );
  INV_X1 U8188 ( .A(n7245), .ZN(n7104) );
  NAND2_X1 U8189 ( .A1(n10075), .A2(n5115), .ZN(n6992) );
  NAND2_X1 U8190 ( .A1(n6505), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U8191 ( .A1(n7090), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6999) );
  NAND2_X1 U8192 ( .A1(n6635), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6998) );
  INV_X1 U8193 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6993) );
  NOR2_X1 U8194 ( .A1(n6994), .A2(n6993), .ZN(n10434) );
  NAND2_X1 U8195 ( .A1(n6995), .A2(n10434), .ZN(n6997) );
  NAND2_X1 U8196 ( .A1(n6519), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6996) );
  NAND2_X1 U8197 ( .A1(n10618), .A2(n10450), .ZN(n7178) );
  INV_X1 U8198 ( .A(n7178), .ZN(n7001) );
  INV_X1 U8199 ( .A(n7177), .ZN(n7000) );
  MUX2_X1 U8200 ( .A(n7001), .B(n7000), .S(n7096), .Z(n7101) );
  OR2_X1 U8201 ( .A1(n7070), .A2(n10668), .ZN(n7072) );
  NAND2_X1 U8202 ( .A1(n10768), .A2(n10658), .ZN(n7002) );
  NAND2_X1 U8203 ( .A1(n7072), .A2(n7002), .ZN(n7164) );
  NAND2_X1 U8204 ( .A1(n10545), .A2(n10559), .ZN(n10393) );
  NAND2_X1 U8205 ( .A1(n7002), .A2(n10393), .ZN(n10394) );
  OR2_X1 U8206 ( .A1(n10561), .A2(n10669), .ZN(n7138) );
  NAND2_X1 U8207 ( .A1(n10561), .A2(n10669), .ZN(n7132) );
  NAND2_X1 U8208 ( .A1(n7138), .A2(n7132), .ZN(n10555) );
  NAND2_X1 U8209 ( .A1(n10586), .A2(n7096), .ZN(n7003) );
  NOR2_X1 U8210 ( .A1(n10684), .A2(n7003), .ZN(n7004) );
  NOR2_X1 U8211 ( .A1(n10555), .A2(n7004), .ZN(n7064) );
  INV_X1 U8212 ( .A(n10586), .ZN(n10558) );
  OR2_X1 U8213 ( .A1(n10684), .A2(n10558), .ZN(n7106) );
  OR2_X1 U8214 ( .A1(n10593), .A2(n10209), .ZN(n10551) );
  NAND2_X1 U8215 ( .A1(n7106), .A2(n10551), .ZN(n7136) );
  NAND2_X1 U8216 ( .A1(n10684), .A2(n10558), .ZN(n10554) );
  AND2_X1 U8217 ( .A1(n7136), .A2(n10554), .ZN(n7006) );
  INV_X1 U8218 ( .A(n7138), .ZN(n7005) );
  AOI21_X1 U8219 ( .B1(n7064), .B2(n7006), .A(n7005), .ZN(n7007) );
  NOR2_X1 U8220 ( .A1(n10394), .A2(n7007), .ZN(n7008) );
  OAI21_X1 U8221 ( .B1(n7164), .B2(n7008), .A(n7095), .ZN(n7069) );
  NAND2_X1 U8222 ( .A1(n10729), .A2(n10179), .ZN(n7046) );
  AND2_X1 U8223 ( .A1(n7159), .A2(n7046), .ZN(n7220) );
  NOR2_X1 U8224 ( .A1(n10258), .A2(n8042), .ZN(n7621) );
  INV_X1 U8225 ( .A(n5111), .ZN(n8098) );
  NAND2_X1 U8226 ( .A1(n8098), .A2(n7009), .ZN(n7010) );
  NAND2_X1 U8227 ( .A1(n7619), .A2(n7010), .ZN(n7630) );
  INV_X1 U8228 ( .A(n7011), .ZN(n10256) );
  NAND2_X1 U8229 ( .A1(n8103), .A2(n10256), .ZN(n7013) );
  NAND2_X1 U8230 ( .A1(n7011), .A2(n10198), .ZN(n7194) );
  INV_X1 U8231 ( .A(n7632), .ZN(n7629) );
  INV_X1 U8232 ( .A(n10255), .ZN(n8716) );
  NAND3_X1 U8233 ( .A1(n7139), .A2(n7194), .A3(n7200), .ZN(n7012) );
  NAND2_X1 U8234 ( .A1(n10254), .A2(n11036), .ZN(n7197) );
  NAND2_X1 U8235 ( .A1(n10255), .A2(n7919), .ZN(n7112) );
  NAND3_X1 U8236 ( .A1(n7012), .A2(n7197), .A3(n7112), .ZN(n7018) );
  AND2_X1 U8237 ( .A1(n7112), .A2(n7013), .ZN(n7195) );
  OAI21_X1 U8238 ( .B1(n7630), .B2(n7632), .A(n7195), .ZN(n7016) );
  NAND2_X1 U8239 ( .A1(n8634), .A2(n8711), .ZN(n7926) );
  AND2_X1 U8240 ( .A1(n7926), .A2(n7200), .ZN(n7015) );
  AOI21_X1 U8241 ( .B1(n7016), .B2(n7015), .A(n7014), .ZN(n7017) );
  MUX2_X1 U8242 ( .A(n7018), .B(n7017), .S(n7095), .Z(n7022) );
  NAND2_X1 U8243 ( .A1(n8717), .A2(n11046), .ZN(n7019) );
  NAND2_X1 U8244 ( .A1(n10253), .A2(n7946), .ZN(n7198) );
  NAND2_X1 U8245 ( .A1(n7019), .A2(n7198), .ZN(n7924) );
  NAND2_X1 U8246 ( .A1(n8698), .A2(n8651), .ZN(n7146) );
  INV_X1 U8247 ( .A(n8651), .ZN(n7975) );
  NAND2_X1 U8248 ( .A1(n10252), .A2(n7975), .ZN(n7980) );
  NAND2_X1 U8249 ( .A1(n7926), .A2(n7019), .ZN(n7020) );
  NAND2_X1 U8250 ( .A1(n7020), .A2(n7198), .ZN(n7202) );
  MUX2_X1 U8251 ( .A(n7198), .B(n7202), .S(n7096), .Z(n7021) );
  OAI211_X1 U8252 ( .C1(n7022), .C2(n7924), .A(n7951), .B(n7021), .ZN(n7024)
         );
  XNOR2_X1 U8253 ( .A(n8701), .B(n10251), .ZN(n7978) );
  MUX2_X1 U8254 ( .A(n7980), .B(n7146), .S(n7095), .Z(n7023) );
  NAND3_X1 U8255 ( .A1(n7024), .A2(n7978), .A3(n7023), .ZN(n7026) );
  OR2_X1 U8256 ( .A1(n8564), .A2(n8697), .ZN(n8660) );
  NAND2_X1 U8257 ( .A1(n8564), .A2(n8697), .ZN(n7111) );
  NAND2_X1 U8258 ( .A1(n8701), .A2(n8776), .ZN(n8557) );
  NAND2_X1 U8259 ( .A1(n8110), .A2(n10251), .ZN(n7109) );
  MUX2_X1 U8260 ( .A(n8557), .B(n7109), .S(n7095), .Z(n7025) );
  NAND3_X1 U8261 ( .A1(n7026), .A2(n8560), .A3(n7025), .ZN(n7030) );
  INV_X1 U8262 ( .A(n10248), .ZN(n8830) );
  NAND2_X1 U8263 ( .A1(n8646), .A2(n8830), .ZN(n7151) );
  NAND2_X1 U8264 ( .A1(n7151), .A2(n7111), .ZN(n7027) );
  AND2_X1 U8265 ( .A1(n9092), .A2(n10248), .ZN(n7206) );
  MUX2_X1 U8266 ( .A(n7027), .B(n7206), .S(n7096), .Z(n7028) );
  OR2_X1 U8267 ( .A1(n8673), .A2(n8121), .ZN(n7143) );
  NAND2_X1 U8268 ( .A1(n8673), .A2(n8121), .ZN(n7144) );
  NAND2_X1 U8269 ( .A1(n7143), .A2(n7144), .ZN(n8665) );
  NOR2_X1 U8270 ( .A1(n7028), .A2(n8665), .ZN(n7029) );
  AND2_X1 U8271 ( .A1(n9064), .A2(n10247), .ZN(n7040) );
  AOI21_X1 U8272 ( .B1(n7030), .B2(n7029), .A(n7040), .ZN(n7039) );
  NOR2_X1 U8273 ( .A1(n8660), .A2(n7095), .ZN(n7038) );
  INV_X1 U8274 ( .A(n7143), .ZN(n7031) );
  NAND2_X1 U8275 ( .A1(n7151), .A2(n7031), .ZN(n7032) );
  INV_X1 U8276 ( .A(n7206), .ZN(n7108) );
  AND2_X1 U8277 ( .A1(n7032), .A2(n7108), .ZN(n7036) );
  NAND2_X1 U8278 ( .A1(n8681), .A2(n8727), .ZN(n7153) );
  NAND2_X1 U8279 ( .A1(n7153), .A2(n7151), .ZN(n7209) );
  INV_X1 U8280 ( .A(n7144), .ZN(n7033) );
  AND2_X1 U8281 ( .A1(n7108), .A2(n7033), .ZN(n7034) );
  NOR2_X1 U8282 ( .A1(n7209), .A2(n7034), .ZN(n7035) );
  MUX2_X1 U8283 ( .A(n7036), .B(n7035), .S(n7096), .Z(n7037) );
  OAI21_X1 U8284 ( .B1(n7039), .B2(n7038), .A(n7037), .ZN(n7044) );
  NAND2_X1 U8285 ( .A1(n8854), .A2(n9063), .ZN(n8863) );
  NAND2_X1 U8286 ( .A1(n8863), .A2(n7153), .ZN(n7041) );
  INV_X1 U8287 ( .A(n7040), .ZN(n8721) );
  NAND2_X1 U8288 ( .A1(n7107), .A2(n8721), .ZN(n7212) );
  MUX2_X1 U8289 ( .A(n7041), .B(n7212), .S(n7096), .Z(n7042) );
  INV_X1 U8290 ( .A(n7042), .ZN(n7043) );
  NAND2_X1 U8291 ( .A1(n7044), .A2(n7043), .ZN(n7050) );
  AND2_X1 U8292 ( .A1(n10184), .A2(n10733), .ZN(n7049) );
  INV_X1 U8293 ( .A(n7049), .ZN(n7214) );
  NAND3_X1 U8294 ( .A1(n7050), .A2(n7214), .A3(n7107), .ZN(n7045) );
  NAND2_X1 U8295 ( .A1(n9006), .A2(n9191), .ZN(n7158) );
  NAND2_X1 U8296 ( .A1(n7045), .A2(n7158), .ZN(n7047) );
  NAND2_X1 U8297 ( .A1(n9045), .A2(n7046), .ZN(n9017) );
  INV_X1 U8298 ( .A(n9017), .ZN(n9070) );
  NAND2_X1 U8299 ( .A1(n7047), .A2(n9070), .ZN(n7048) );
  NAND2_X1 U8300 ( .A1(n7220), .A2(n7048), .ZN(n7053) );
  AND2_X1 U8301 ( .A1(n7158), .A2(n8863), .ZN(n7213) );
  AOI21_X1 U8302 ( .B1(n7050), .B2(n7213), .A(n7049), .ZN(n7051) );
  NAND2_X1 U8303 ( .A1(n10723), .A2(n10730), .ZN(n7217) );
  OAI211_X1 U8304 ( .C1(n7051), .C2(n9017), .A(n9045), .B(n7217), .ZN(n7052)
         );
  INV_X1 U8305 ( .A(n10714), .ZN(n9086) );
  NAND2_X1 U8306 ( .A1(n9086), .A2(n10703), .ZN(n7190) );
  AND2_X1 U8307 ( .A1(n10714), .A2(n10719), .ZN(n7054) );
  XNOR2_X1 U8308 ( .A(n10706), .B(n9219), .ZN(n9159) );
  NOR2_X1 U8309 ( .A1(n7055), .A2(n9159), .ZN(n7058) );
  INV_X1 U8310 ( .A(n10587), .ZN(n10150) );
  OR2_X1 U8311 ( .A1(n10406), .A2(n10150), .ZN(n7224) );
  OR2_X1 U8312 ( .A1(n10706), .A2(n9219), .ZN(n7161) );
  AND2_X1 U8313 ( .A1(n7224), .A2(n7161), .ZN(n7222) );
  NAND2_X1 U8314 ( .A1(n10406), .A2(n10150), .ZN(n7162) );
  NAND2_X1 U8315 ( .A1(n10593), .A2(n10209), .ZN(n7227) );
  INV_X1 U8316 ( .A(n7227), .ZN(n7163) );
  AND2_X1 U8317 ( .A1(n10554), .A2(n7227), .ZN(n7056) );
  MUX2_X1 U8318 ( .A(n7163), .B(n7056), .S(n7096), .Z(n7060) );
  NAND2_X1 U8319 ( .A1(n10706), .A2(n9219), .ZN(n7057) );
  NAND2_X1 U8320 ( .A1(n7162), .A2(n7057), .ZN(n7225) );
  XNOR2_X1 U8321 ( .A(n10593), .B(n10694), .ZN(n10583) );
  OAI211_X1 U8322 ( .C1(n7058), .C2(n7225), .A(n7224), .B(n10583), .ZN(n7059)
         );
  NAND2_X1 U8323 ( .A1(n7060), .A2(n7059), .ZN(n7062) );
  OR2_X1 U8324 ( .A1(n10554), .A2(n7096), .ZN(n7061) );
  NAND4_X1 U8325 ( .A1(n7064), .A2(n7063), .A3(n7062), .A4(n7061), .ZN(n7066)
         );
  NAND3_X1 U8326 ( .A1(n10561), .A2(n10669), .A3(n7096), .ZN(n7065) );
  NAND2_X1 U8327 ( .A1(n7066), .A2(n7065), .ZN(n7067) );
  NAND2_X1 U8328 ( .A1(n10535), .A2(n7067), .ZN(n7068) );
  NAND2_X1 U8329 ( .A1(n7070), .A2(n10668), .ZN(n10395) );
  NAND2_X1 U8330 ( .A1(n10395), .A2(n7095), .ZN(n7071) );
  NAND2_X1 U8331 ( .A1(n10395), .A2(n10393), .ZN(n7134) );
  NAND3_X1 U8332 ( .A1(n7134), .A2(n7096), .A3(n7072), .ZN(n7073) );
  OR2_X1 U8333 ( .A1(n10654), .A2(n10644), .ZN(n10397) );
  NAND2_X1 U8334 ( .A1(n10654), .A2(n10644), .ZN(n7165) );
  NAND2_X1 U8335 ( .A1(n10397), .A2(n7165), .ZN(n10511) );
  NAND2_X1 U8336 ( .A1(n10647), .A2(n10634), .ZN(n10399) );
  NAND2_X1 U8337 ( .A1(n10487), .A2(n10643), .ZN(n10400) );
  OR2_X1 U8338 ( .A1(n10487), .A2(n10643), .ZN(n7170) );
  OAI21_X1 U8339 ( .B1(n7074), .B2(n10476), .A(n7170), .ZN(n7080) );
  NAND2_X1 U8340 ( .A1(n10399), .A2(n7165), .ZN(n7075) );
  OAI21_X1 U8341 ( .B1(n7076), .B2(n7075), .A(n7105), .ZN(n7078) );
  INV_X1 U8342 ( .A(n7170), .ZN(n7077) );
  AOI21_X1 U8343 ( .B1(n7078), .B2(n10400), .A(n7077), .ZN(n7079) );
  MUX2_X1 U8344 ( .A(n7080), .B(n7079), .S(n7096), .Z(n7084) );
  OR2_X1 U8345 ( .A1(n10752), .A2(n10633), .ZN(n7171) );
  NAND2_X1 U8346 ( .A1(n10752), .A2(n10633), .ZN(n10402) );
  NAND2_X1 U8347 ( .A1(n9471), .A2(n5115), .ZN(n7082) );
  NAND2_X1 U8348 ( .A1(n6505), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8349 ( .A1(n10620), .A2(n10626), .ZN(n10403) );
  MUX2_X1 U8350 ( .A(n10402), .B(n7171), .S(n7096), .Z(n7083) );
  OAI211_X1 U8351 ( .C1(n7084), .C2(n5563), .A(n10447), .B(n7083), .ZN(n7086)
         );
  MUX2_X1 U8352 ( .A(n7172), .B(n10403), .S(n7096), .Z(n7085) );
  NAND2_X1 U8353 ( .A1(n7086), .A2(n7085), .ZN(n7094) );
  NAND2_X1 U8354 ( .A1(n6505), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U8355 ( .A1(n6635), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7093) );
  NAND2_X1 U8356 ( .A1(n6519), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7092) );
  NAND2_X1 U8357 ( .A1(n7090), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7091) );
  AND3_X1 U8358 ( .A1(n7093), .A2(n7092), .A3(n7091), .ZN(n10245) );
  OAI21_X1 U8359 ( .B1(n10245), .B2(n7102), .A(n7124), .ZN(n7182) );
  OAI211_X1 U8360 ( .C1(n10429), .C2(n7094), .A(n7180), .B(n7182), .ZN(n7100)
         );
  NAND2_X1 U8361 ( .A1(n10379), .A2(n7102), .ZN(n7243) );
  NAND2_X1 U8362 ( .A1(n7129), .A2(n6947), .ZN(n7103) );
  AOI211_X1 U8363 ( .C1(n6773), .C2(n7104), .A(n6444), .B(n7103), .ZN(n7252)
         );
  NAND2_X1 U8364 ( .A1(n7105), .A2(n10399), .ZN(n10398) );
  INV_X1 U8365 ( .A(n7222), .ZN(n7120) );
  NAND2_X1 U8366 ( .A1(n7214), .A2(n7158), .ZN(n8862) );
  NAND2_X1 U8367 ( .A1(n7107), .A2(n8863), .ZN(n8728) );
  NAND2_X1 U8368 ( .A1(n8721), .A2(n7153), .ZN(n8687) );
  AND3_X1 U8369 ( .A1(n8660), .A2(n7980), .A3(n7109), .ZN(n7110) );
  NAND2_X1 U8370 ( .A1(n7111), .A2(n8557), .ZN(n7142) );
  NAND2_X1 U8371 ( .A1(n7200), .A2(n7112), .ZN(n7591) );
  INV_X1 U8372 ( .A(n7621), .ZN(n7113) );
  NAND2_X1 U8373 ( .A1(n10258), .A2(n8042), .ZN(n7192) );
  AND2_X1 U8374 ( .A1(n7113), .A2(n7192), .ZN(n11019) );
  NAND4_X1 U8375 ( .A1(n7629), .A2(n7601), .A3(n11019), .A4(n8824), .ZN(n7115)
         );
  AND2_X1 U8376 ( .A1(n7926), .A2(n7197), .ZN(n7922) );
  INV_X1 U8377 ( .A(n7924), .ZN(n7928) );
  NAND3_X1 U8378 ( .A1(n7922), .A2(n7928), .A3(n7620), .ZN(n7114) );
  INV_X1 U8379 ( .A(n7146), .ZN(n7981) );
  NOR4_X1 U8380 ( .A1(n7142), .A2(n7115), .A3(n7114), .A4(n7981), .ZN(n7116)
         );
  NAND4_X1 U8381 ( .A1(n8123), .A2(n7203), .A3(n7116), .A4(n7144), .ZN(n7117)
         );
  NOR4_X1 U8382 ( .A1(n8862), .A2(n8728), .A3(n8687), .A4(n7117), .ZN(n7118)
         );
  NAND4_X1 U8383 ( .A1(n9078), .A2(n9070), .A3(n9073), .A4(n7118), .ZN(n7119)
         );
  NOR4_X1 U8384 ( .A1(n10555), .A2(n7120), .A3(n7225), .A4(n7119), .ZN(n7121)
         );
  NAND4_X1 U8385 ( .A1(n10535), .A2(n10576), .A3(n7121), .A4(n10583), .ZN(
        n7122) );
  NOR4_X1 U8386 ( .A1(n10398), .A2(n10511), .A3(n10521), .A4(n7122), .ZN(n7123) );
  NAND4_X1 U8387 ( .A1(n10447), .A2(n10471), .A3(n10479), .A4(n7123), .ZN(
        n7125) );
  AND2_X1 U8388 ( .A1(n7124), .A2(n10245), .ZN(n7238) );
  NOR3_X1 U8389 ( .A1(n7125), .A2(n7241), .A3(n7238), .ZN(n7126) );
  INV_X1 U8390 ( .A(n7126), .ZN(n7127) );
  NOR2_X1 U8391 ( .A1(n10429), .A2(n7127), .ZN(n7128) );
  NAND3_X1 U8392 ( .A1(n7128), .A2(n7245), .A3(n7243), .ZN(n7186) );
  OAI211_X1 U8393 ( .C1(n6444), .C2(n8824), .A(n7186), .B(n6773), .ZN(n7130)
         );
  INV_X1 U8394 ( .A(n10554), .ZN(n7131) );
  NAND2_X1 U8395 ( .A1(n7138), .A2(n7131), .ZN(n7133) );
  NAND2_X1 U8396 ( .A1(n7133), .A2(n7132), .ZN(n10390) );
  NOR2_X1 U8397 ( .A1(n7134), .A2(n10390), .ZN(n7135) );
  AND2_X1 U8398 ( .A1(n7135), .A2(n7165), .ZN(n7189) );
  INV_X1 U8399 ( .A(n7136), .ZN(n7137) );
  NAND2_X1 U8400 ( .A1(n7138), .A2(n7137), .ZN(n7230) );
  NAND2_X1 U8401 ( .A1(n7139), .A2(n7194), .ZN(n7602) );
  NAND2_X1 U8402 ( .A1(n7602), .A2(n7601), .ZN(n7140) );
  INV_X1 U8403 ( .A(n7198), .ZN(n7141) );
  NAND2_X1 U8404 ( .A1(n7982), .A2(n7203), .ZN(n7150) );
  NAND3_X1 U8405 ( .A1(n7143), .A2(n8660), .A3(n7142), .ZN(n7145) );
  AND2_X1 U8406 ( .A1(n7145), .A2(n7144), .ZN(n7149) );
  INV_X1 U8407 ( .A(n7203), .ZN(n7147) );
  NAND2_X1 U8408 ( .A1(n7150), .A2(n7208), .ZN(n8126) );
  NAND2_X1 U8409 ( .A1(n8126), .A2(n8123), .ZN(n7152) );
  INV_X1 U8410 ( .A(n7153), .ZN(n7154) );
  INV_X1 U8411 ( .A(n7212), .ZN(n7155) );
  INV_X1 U8412 ( .A(n8862), .ZN(n7156) );
  NAND2_X1 U8413 ( .A1(n7157), .A2(n7156), .ZN(n8866) );
  NAND2_X1 U8414 ( .A1(n8866), .A2(n7158), .ZN(n9018) );
  INV_X1 U8415 ( .A(n9159), .ZN(n7160) );
  NAND2_X1 U8416 ( .A1(n7224), .A2(n7162), .ZN(n9222) );
  NAND3_X1 U8417 ( .A1(n7165), .A2(n10395), .A3(n7164), .ZN(n7166) );
  NAND2_X1 U8418 ( .A1(n5151), .A2(n7166), .ZN(n7234) );
  AOI21_X1 U8419 ( .B1(n7189), .B2(n10391), .A(n7234), .ZN(n7181) );
  INV_X1 U8420 ( .A(n7175), .ZN(n7168) );
  NAND2_X1 U8421 ( .A1(n10400), .A2(n10399), .ZN(n7167) );
  NOR2_X1 U8422 ( .A1(n7168), .A2(n7167), .ZN(n7169) );
  NAND2_X1 U8423 ( .A1(n7178), .A2(n7169), .ZN(n7237) );
  NAND2_X1 U8424 ( .A1(n7171), .A2(n7170), .ZN(n7174) );
  INV_X1 U8425 ( .A(n7172), .ZN(n7173) );
  AOI21_X1 U8426 ( .B1(n7175), .B2(n7174), .A(n7173), .ZN(n7176) );
  NAND2_X1 U8427 ( .A1(n7177), .A2(n7176), .ZN(n7179) );
  NAND2_X1 U8428 ( .A1(n7179), .A2(n7178), .ZN(n7235) );
  OAI211_X1 U8429 ( .C1(n7181), .C2(n7237), .A(n7180), .B(n7235), .ZN(n7183)
         );
  NAND3_X1 U8430 ( .A1(n7183), .A2(n7182), .A3(n7245), .ZN(n7184) );
  NAND3_X1 U8431 ( .A1(n7184), .A2(n7599), .A3(n7243), .ZN(n7185) );
  AOI21_X1 U8432 ( .B1(n7186), .B2(n7185), .A(n6773), .ZN(n7187) );
  INV_X1 U8433 ( .A(n7189), .ZN(n7232) );
  NAND2_X1 U8434 ( .A1(n5111), .A2(n7815), .ZN(n7191) );
  NAND3_X1 U8435 ( .A1(n7192), .A2(n6947), .A3(n7191), .ZN(n7193) );
  NAND2_X1 U8436 ( .A1(n7194), .A2(n7193), .ZN(n7196) );
  OAI21_X1 U8437 ( .B1(n7630), .B2(n7196), .A(n7195), .ZN(n7201) );
  NAND2_X1 U8438 ( .A1(n7198), .A2(n7197), .ZN(n7199) );
  AOI21_X1 U8439 ( .B1(n7201), .B2(n7200), .A(n7199), .ZN(n7205) );
  INV_X1 U8440 ( .A(n7202), .ZN(n7204) );
  OAI21_X1 U8441 ( .B1(n7205), .B2(n7204), .A(n7203), .ZN(n7207) );
  AOI21_X1 U8442 ( .B1(n7208), .B2(n7207), .A(n7206), .ZN(n7210) );
  NOR2_X1 U8443 ( .A1(n7210), .A2(n7209), .ZN(n7211) );
  NOR2_X1 U8444 ( .A1(n7212), .A2(n7211), .ZN(n7216) );
  INV_X1 U8445 ( .A(n7213), .ZN(n7215) );
  OAI211_X1 U8446 ( .C1(n7216), .C2(n7215), .A(n9045), .B(n7214), .ZN(n7219)
         );
  INV_X1 U8447 ( .A(n7217), .ZN(n7218) );
  AOI21_X1 U8448 ( .B1(n7220), .B2(n7219), .A(n7218), .ZN(n7223) );
  OAI211_X1 U8449 ( .C1(n5320), .C2(n7223), .A(n7222), .B(n7221), .ZN(n7228)
         );
  NAND2_X1 U8450 ( .A1(n7225), .A2(n7224), .ZN(n7226) );
  AND3_X1 U8451 ( .A1(n7228), .A2(n7227), .A3(n7226), .ZN(n7229) );
  NOR2_X1 U8452 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  NOR2_X1 U8453 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  NOR2_X1 U8454 ( .A1(n7234), .A2(n7233), .ZN(n7236) );
  OAI21_X1 U8455 ( .B1(n7237), .B2(n7236), .A(n7235), .ZN(n7240) );
  INV_X1 U8456 ( .A(n7238), .ZN(n7239) );
  NAND2_X1 U8457 ( .A1(n7240), .A2(n7239), .ZN(n7244) );
  INV_X1 U8458 ( .A(n7241), .ZN(n7242) );
  NAND3_X1 U8459 ( .A1(n7244), .A2(n7243), .A3(n7242), .ZN(n7246) );
  NAND2_X1 U8460 ( .A1(n7246), .A2(n7245), .ZN(n7248) );
  NAND3_X1 U8461 ( .A1(n7248), .A2(n6773), .A3(n8920), .ZN(n7247) );
  AND2_X1 U8462 ( .A1(n7328), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9130) );
  OAI211_X1 U8463 ( .C1(n7248), .C2(n7593), .A(n7247), .B(n9130), .ZN(n7249)
         );
  OAI21_X1 U8464 ( .B1(n7252), .B2(n7251), .A(n7250), .ZN(n7256) );
  INV_X1 U8465 ( .A(n10271), .ZN(n7598) );
  INV_X1 U8466 ( .A(n10795), .ZN(n10272) );
  NAND2_X1 U8467 ( .A1(n7598), .A2(n10272), .ZN(n10274) );
  NAND2_X1 U8468 ( .A1(n9130), .A2(n6946), .ZN(n7253) );
  OAI211_X1 U8469 ( .C1(n7254), .C2(n10274), .A(P1_B_REG_SCAN_IN), .B(n7253), 
        .ZN(n7255) );
  NAND2_X1 U8470 ( .A1(n7256), .A2(n7255), .ZN(P1_U3242) );
  NAND2_X1 U8471 ( .A1(n10620), .A2(n6764), .ZN(n7259) );
  OR2_X1 U8472 ( .A1(n10626), .A2(n7257), .ZN(n7258) );
  NAND2_X1 U8473 ( .A1(n7259), .A2(n7258), .ZN(n7260) );
  XNOR2_X1 U8474 ( .A(n7260), .B(n6489), .ZN(n7264) );
  NAND2_X1 U8475 ( .A1(n10620), .A2(n5113), .ZN(n7261) );
  OAI21_X1 U8476 ( .B1(n10626), .B2(n7262), .A(n7261), .ZN(n7263) );
  XNOR2_X1 U8477 ( .A(n7264), .B(n7263), .ZN(n7269) );
  INV_X1 U8478 ( .A(n7269), .ZN(n7266) );
  INV_X1 U8479 ( .A(n7268), .ZN(n7265) );
  NAND4_X1 U8480 ( .A1(n7267), .A2(n7266), .A3(n10223), .A4(n7265), .ZN(n7279)
         );
  NAND3_X1 U8481 ( .A1(n7269), .A2(n10223), .A3(n7268), .ZN(n7274) );
  INV_X1 U8482 ( .A(n10633), .ZN(n10425) );
  AOI22_X1 U8483 ( .A1(n10233), .A2(n10425), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n7271) );
  NAND2_X1 U8484 ( .A1(n10241), .A2(n10456), .ZN(n7270) );
  OAI211_X1 U8485 ( .C1(n10450), .C2(n10236), .A(n7271), .B(n7270), .ZN(n7272)
         );
  AOI21_X1 U8486 ( .B1(n10620), .B2(n10215), .A(n7272), .ZN(n7273) );
  NAND2_X1 U8487 ( .A1(n7274), .A2(n7273), .ZN(n7275) );
  AOI21_X1 U8488 ( .B1(n7277), .B2(n7276), .A(n7275), .ZN(n7278) );
  NOR2_X1 U8489 ( .A1(n6483), .A2(P1_U3086), .ZN(n7280) );
  INV_X1 U8490 ( .A(n7305), .ZN(n7281) );
  NAND2_X1 U8491 ( .A1(n7405), .A2(n9449), .ZN(n7282) );
  NAND2_X1 U8492 ( .A1(n7282), .A2(n7404), .ZN(n7340) );
  NAND2_X1 U8493 ( .A1(n7340), .A2(n5852), .ZN(n7283) );
  NAND2_X1 U8494 ( .A1(n7283), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X2 U8495 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U8496 ( .A(n10266), .ZN(n7383) );
  NAND2_X1 U8497 ( .A1(n7287), .A2(P1_U3086), .ZN(n9234) );
  INV_X1 U8498 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7285) );
  NAND2_X1 U8499 ( .A1(n5392), .A2(P1_U3086), .ZN(n10792) );
  OAI222_X1 U8500 ( .A1(P1_U3086), .A2(n7383), .B1(n9234), .B2(n7288), .C1(
        n7285), .C2(n10792), .ZN(P1_U3354) );
  INV_X1 U8501 ( .A(n10283), .ZN(n7385) );
  INV_X1 U8502 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7286) );
  OAI222_X1 U8503 ( .A1(P1_U3086), .A2(n7385), .B1(n9234), .B2(n7295), .C1(
        n7286), .C2(n10792), .ZN(P1_U3353) );
  INV_X1 U8504 ( .A(n10296), .ZN(n7388) );
  OAI222_X1 U8505 ( .A1(P1_U3086), .A2(n7388), .B1(n9234), .B2(n7298), .C1(
        n5707), .C2(n10792), .ZN(P1_U3352) );
  NAND2_X1 U8506 ( .A1(n7287), .A2(P2_U3151), .ZN(n10086) );
  NAND2_X1 U8507 ( .A1(n5392), .A2(P2_U3151), .ZN(n10087) );
  OAI222_X1 U8508 ( .A1(n10086), .A2(n7289), .B1(n7441), .B2(P2_U3151), .C1(
        n10087), .C2(n7288), .ZN(P2_U3294) );
  INV_X1 U8509 ( .A(n7728), .ZN(n7290) );
  NAND2_X1 U8510 ( .A1(n7290), .A2(n7425), .ZN(n7291) );
  OAI21_X1 U8511 ( .B1(n7425), .B2(n7292), .A(n7291), .ZN(P2_U3377) );
  INV_X1 U8512 ( .A(n10086), .ZN(n10083) );
  AOI22_X1 U8513 ( .A1(n10934), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n10083), .ZN(n7293) );
  OAI21_X1 U8514 ( .B1(n7294), .B2(n10087), .A(n7293), .ZN(P2_U3291) );
  INV_X1 U8515 ( .A(n10309), .ZN(n7389) );
  INV_X1 U8516 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7317) );
  OAI222_X1 U8517 ( .A1(n7389), .A2(P1_U3086), .B1(n9234), .B2(n7294), .C1(
        n10792), .C2(n7317), .ZN(P1_U3351) );
  INV_X1 U8518 ( .A(n10083), .ZN(n10070) );
  INV_X1 U8519 ( .A(n7453), .ZN(n10912) );
  OAI222_X1 U8520 ( .A1(n10070), .A2(n7296), .B1(n10912), .B2(P2_U3151), .C1(
        n10087), .C2(n7295), .ZN(P2_U3293) );
  INV_X1 U8521 ( .A(n10944), .ZN(n7705) );
  INV_X1 U8522 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7297) );
  OAI222_X1 U8523 ( .A1(n10087), .A2(n7300), .B1(n7705), .B2(P2_U3151), .C1(
        n7297), .C2(n10086), .ZN(P2_U3290) );
  INV_X1 U8524 ( .A(n10087), .ZN(n9133) );
  INV_X1 U8525 ( .A(n7708), .ZN(n7696) );
  OAI222_X1 U8526 ( .A1(n10077), .A2(n7298), .B1(n7696), .B2(P2_U3151), .C1(
        n5709), .C2(n10086), .ZN(P2_U3292) );
  INV_X1 U8527 ( .A(n10323), .ZN(n7391) );
  OAI222_X1 U8528 ( .A1(P1_U3086), .A2(n7391), .B1(n9234), .B2(n7300), .C1(
        n7299), .C2(n10792), .ZN(P1_U3350) );
  INV_X1 U8529 ( .A(n7425), .ZN(n7302) );
  INV_X1 U8530 ( .A(n7303), .ZN(n7304) );
  AOI22_X1 U8531 ( .A1(n9238), .A2(n7306), .B1(n7305), .B2(n7304), .ZN(
        P2_U3376) );
  INV_X1 U8532 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7307) );
  OAI222_X1 U8533 ( .A1(n10087), .A2(n7309), .B1(n7748), .B2(P2_U3151), .C1(
        n7307), .C2(n10086), .ZN(P2_U3289) );
  INV_X1 U8534 ( .A(n10336), .ZN(n7393) );
  INV_X1 U8535 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7308) );
  OAI222_X1 U8536 ( .A1(P1_U3086), .A2(n7393), .B1(n9234), .B2(n7309), .C1(
        n7308), .C2(n10792), .ZN(P1_U3349) );
  INV_X1 U8537 ( .A(n7766), .ZN(n7846) );
  INV_X1 U8538 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7310) );
  OAI222_X1 U8539 ( .A1(n10077), .A2(n7312), .B1(n7846), .B2(P2_U3151), .C1(
        n7310), .C2(n10086), .ZN(P2_U3288) );
  INV_X1 U8540 ( .A(n10349), .ZN(n7394) );
  INV_X1 U8541 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7311) );
  OAI222_X1 U8542 ( .A1(P1_U3086), .A2(n7394), .B1(n9234), .B2(n7312), .C1(
        n7311), .C2(n10792), .ZN(P1_U3348) );
  INV_X1 U8543 ( .A(n7313), .ZN(n7315) );
  AOI22_X1 U8544 ( .A1(n7487), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10796), .ZN(n7314) );
  OAI21_X1 U8545 ( .B1(n7315), .B2(n9234), .A(n7314), .ZN(P1_U3347) );
  OAI222_X1 U8546 ( .A1(n10070), .A2(n5247), .B1(n10087), .B2(n7315), .C1(
        P2_U3151), .C2(n7877), .ZN(P2_U3287) );
  NAND2_X1 U8547 ( .A1(n7644), .A2(P2_U3893), .ZN(n7316) );
  OAI21_X1 U8548 ( .B1(P2_U3893), .B2(n7317), .A(n7316), .ZN(P2_U3495) );
  AOI22_X1 U8549 ( .A1(n7531), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10796), .ZN(n7318) );
  OAI21_X1 U8550 ( .B1(n7320), .B2(n10799), .A(n7318), .ZN(P1_U3345) );
  INV_X1 U8551 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7319) );
  OAI222_X1 U8552 ( .A1(n10077), .A2(n7320), .B1(n8945), .B2(P2_U3151), .C1(
        n7319), .C2(n10086), .ZN(P2_U3285) );
  INV_X1 U8553 ( .A(n7321), .ZN(n7324) );
  INV_X1 U8554 ( .A(n8927), .ZN(n8947) );
  INV_X1 U8555 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7322) );
  OAI222_X1 U8556 ( .A1(n10077), .A2(n7324), .B1(n8947), .B2(P2_U3151), .C1(
        n7322), .C2(n10086), .ZN(P2_U3286) );
  INV_X1 U8557 ( .A(n7503), .ZN(n7478) );
  INV_X1 U8558 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7323) );
  OAI222_X1 U8559 ( .A1(P1_U3086), .A2(n7478), .B1(n9234), .B2(n7324), .C1(
        n7323), .C2(n10792), .ZN(P1_U3346) );
  NAND2_X1 U8560 ( .A1(n7325), .A2(n7599), .ZN(n7327) );
  NAND2_X1 U8561 ( .A1(n7327), .A2(n7326), .ZN(n7330) );
  INV_X1 U8562 ( .A(n7330), .ZN(n7329) );
  OAI21_X1 U8563 ( .B1(n6483), .B2(n7328), .A(P1_STATE_REG_SCAN_IN), .ZN(n7331) );
  NOR2_X1 U8564 ( .A1(n10265), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8565 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7336) );
  INV_X1 U8566 ( .A(n7396), .ZN(n7334) );
  INV_X1 U8567 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8052) );
  AOI21_X1 U8568 ( .B1(n10272), .B2(n8052), .A(n10271), .ZN(n10276) );
  OAI21_X1 U8569 ( .B1(n10272), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10276), .ZN(
        n7332) );
  XNOR2_X1 U8570 ( .A(n7332), .B(P1_IR_REG_0__SCAN_IN), .ZN(n7333) );
  AOI22_X1 U8571 ( .A1(n7334), .A2(n7333), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n7335) );
  OAI21_X1 U8572 ( .B1(n10367), .B2(n7336), .A(n7335), .ZN(P1_U3243) );
  INV_X1 U8573 ( .A(n7337), .ZN(n7363) );
  AOI22_X1 U8574 ( .A1(n7517), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10796), .ZN(n7338) );
  OAI21_X1 U8575 ( .B1(n7363), .B2(n10799), .A(n7338), .ZN(P1_U3344) );
  NOR2_X1 U8576 ( .A1(n9756), .A2(P2_U3151), .ZN(n10082) );
  NAND2_X1 U8577 ( .A1(n7340), .A2(n10082), .ZN(n7339) );
  INV_X1 U8578 ( .A(n7359), .ZN(n9462) );
  MUX2_X1 U8579 ( .A(n7339), .B(n11001), .S(n9462), .Z(n11000) );
  NOR2_X1 U8580 ( .A1(n7359), .A2(P2_U3151), .ZN(n10078) );
  AND2_X1 U8581 ( .A1(n7340), .A2(n10078), .ZN(n10895) );
  INV_X1 U8582 ( .A(n9756), .ZN(n7341) );
  NAND2_X1 U8583 ( .A1(n10895), .A2(n7341), .ZN(n11008) );
  AND2_X1 U8584 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n7347), .ZN(n7343) );
  OAI22_X1 U8585 ( .A1(n7441), .A2(n7343), .B1(n7342), .B2(n7358), .ZN(n7345)
         );
  NAND2_X1 U8586 ( .A1(n7345), .A2(n7344), .ZN(n7346) );
  NAND2_X1 U8587 ( .A1(n7451), .A2(n7346), .ZN(n7355) );
  AND2_X1 U8588 ( .A1(n7347), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7348) );
  NAND2_X1 U8589 ( .A1(n7449), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7454) );
  OAI21_X1 U8590 ( .B1(n7441), .B2(n7348), .A(n7454), .ZN(n7349) );
  INV_X1 U8591 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7573) );
  OR2_X1 U8592 ( .A1(n7349), .A2(n7573), .ZN(n7455) );
  NAND2_X1 U8593 ( .A1(n7349), .A2(n7573), .ZN(n7350) );
  AND2_X1 U8594 ( .A1(n7455), .A2(n7350), .ZN(n7351) );
  OAI22_X1 U8595 ( .A1(n11011), .A2(n7351), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7859), .ZN(n7354) );
  INV_X1 U8596 ( .A(n7404), .ZN(n9135) );
  NOR2_X1 U8597 ( .A1(n7405), .A2(n9135), .ZN(n7352) );
  INV_X1 U8598 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10840) );
  NOR2_X1 U8599 ( .A1(n10940), .A2(n10840), .ZN(n7353) );
  AOI211_X1 U8600 ( .C1(n10983), .C2(n7355), .A(n7354), .B(n7353), .ZN(n7362)
         );
  MUX2_X1 U8601 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n9756), .Z(n7442) );
  XNOR2_X1 U8602 ( .A(n7442), .B(n7356), .ZN(n7443) );
  MUX2_X1 U8603 ( .A(n7358), .B(n7357), .S(n9756), .Z(n10893) );
  NAND2_X1 U8604 ( .A1(n10893), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10892) );
  XOR2_X1 U8605 ( .A(n7443), .B(n10892), .Z(n7360) );
  NAND2_X1 U8606 ( .A1(n7360), .A2(n10996), .ZN(n7361) );
  OAI211_X1 U8607 ( .C1(n11000), .C2(n7441), .A(n7362), .B(n7361), .ZN(
        P2_U3183) );
  INV_X1 U8608 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7364) );
  INV_X1 U8609 ( .A(n10975), .ZN(n8951) );
  OAI222_X1 U8610 ( .A1(n10070), .A2(n7364), .B1(n10087), .B2(n7363), .C1(
        P2_U3151), .C2(n8951), .ZN(P2_U3284) );
  INV_X1 U8611 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8581) );
  MUX2_X1 U8612 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n8581), .S(n7487), .Z(n7378)
         );
  INV_X1 U8613 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7365) );
  XNOR2_X1 U8614 ( .A(n10283), .B(n7365), .ZN(n10286) );
  INV_X1 U8615 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7366) );
  XNOR2_X1 U8616 ( .A(n10266), .B(n7366), .ZN(n10263) );
  NAND2_X1 U8617 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10275) );
  INV_X1 U8618 ( .A(n10275), .ZN(n10264) );
  NAND2_X1 U8619 ( .A1(n10263), .A2(n10264), .ZN(n10262) );
  NAND2_X1 U8620 ( .A1(n10266), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7367) );
  NAND2_X1 U8621 ( .A1(n10262), .A2(n7367), .ZN(n10285) );
  NAND2_X1 U8622 ( .A1(n10286), .A2(n10285), .ZN(n10284) );
  NAND2_X1 U8623 ( .A1(n10283), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7368) );
  NAND2_X1 U8624 ( .A1(n10284), .A2(n7368), .ZN(n10298) );
  INV_X1 U8625 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n8746) );
  XNOR2_X1 U8626 ( .A(n10296), .B(n8746), .ZN(n10299) );
  NAND2_X1 U8627 ( .A1(n10298), .A2(n10299), .ZN(n10297) );
  NAND2_X1 U8628 ( .A1(n10296), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7369) );
  NAND2_X1 U8629 ( .A1(n10297), .A2(n7369), .ZN(n10314) );
  INV_X1 U8630 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7370) );
  MUX2_X1 U8631 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7370), .S(n10309), .Z(n10315) );
  NAND2_X1 U8632 ( .A1(n10314), .A2(n10315), .ZN(n10313) );
  NAND2_X1 U8633 ( .A1(n10309), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7371) );
  NAND2_X1 U8634 ( .A1(n10313), .A2(n7371), .ZN(n10325) );
  INV_X1 U8635 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7372) );
  XNOR2_X1 U8636 ( .A(n10323), .B(n7372), .ZN(n10326) );
  NAND2_X1 U8637 ( .A1(n10325), .A2(n10326), .ZN(n10324) );
  NAND2_X1 U8638 ( .A1(n10323), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7373) );
  NAND2_X1 U8639 ( .A1(n10324), .A2(n7373), .ZN(n10338) );
  INV_X1 U8640 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7374) );
  XNOR2_X1 U8641 ( .A(n10336), .B(n7374), .ZN(n10339) );
  NAND2_X1 U8642 ( .A1(n10338), .A2(n10339), .ZN(n10337) );
  NAND2_X1 U8643 ( .A1(n10336), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7375) );
  NAND2_X1 U8644 ( .A1(n10337), .A2(n7375), .ZN(n10351) );
  INV_X1 U8645 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7376) );
  MUX2_X1 U8646 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7376), .S(n10349), .Z(n10352) );
  NAND2_X1 U8647 ( .A1(n10351), .A2(n10352), .ZN(n10350) );
  NAND2_X1 U8648 ( .A1(n10349), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7377) );
  NAND2_X1 U8649 ( .A1(n10350), .A2(n7377), .ZN(n7379) );
  NOR2_X2 U8650 ( .A1(n7396), .A2(n10274), .ZN(n10372) );
  OAI21_X1 U8651 ( .B1(n7378), .B2(n7379), .A(n10372), .ZN(n7401) );
  AND2_X1 U8652 ( .A1(n7379), .A2(n7378), .ZN(n7477) );
  NOR2_X2 U8653 ( .A1(n7396), .A2(n7598), .ZN(n10369) );
  INV_X1 U8654 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7380) );
  NAND2_X1 U8655 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8773) );
  OAI21_X1 U8656 ( .B1(n10367), .B2(n7380), .A(n8773), .ZN(n7381) );
  AOI21_X1 U8657 ( .B1(n7487), .B2(n10369), .A(n7381), .ZN(n7400) );
  INV_X1 U8658 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7382) );
  MUX2_X1 U8659 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7382), .S(n7487), .Z(n7398)
         );
  INV_X1 U8660 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7395) );
  INV_X1 U8661 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7392) );
  INV_X1 U8662 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7390) );
  INV_X1 U8663 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7387) );
  INV_X1 U8664 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7386) );
  XOR2_X1 U8665 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10283), .Z(n10289) );
  INV_X1 U8666 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7384) );
  XOR2_X1 U8667 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10266), .Z(n10261) );
  INV_X1 U8668 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n11026) );
  NAND3_X1 U8669 ( .A1(n10261), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10259) );
  OAI21_X1 U8670 ( .B1(n7384), .B2(n7383), .A(n10259), .ZN(n10288) );
  NAND2_X1 U8671 ( .A1(n10289), .A2(n10288), .ZN(n10287) );
  OAI21_X1 U8672 ( .B1(n7386), .B2(n7385), .A(n10287), .ZN(n10301) );
  XOR2_X1 U8673 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10296), .Z(n10302) );
  NAND2_X1 U8674 ( .A1(n10301), .A2(n10302), .ZN(n10300) );
  OAI21_X1 U8675 ( .B1(n7388), .B2(n7387), .A(n10300), .ZN(n10311) );
  MUX2_X1 U8676 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7390), .S(n10309), .Z(n10312) );
  NAND2_X1 U8677 ( .A1(n10311), .A2(n10312), .ZN(n10310) );
  OAI21_X1 U8678 ( .B1(n7390), .B2(n7389), .A(n10310), .ZN(n10328) );
  XOR2_X1 U8679 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10323), .Z(n10329) );
  NAND2_X1 U8680 ( .A1(n10328), .A2(n10329), .ZN(n10327) );
  OAI21_X1 U8681 ( .B1(n7392), .B2(n7391), .A(n10327), .ZN(n10341) );
  XOR2_X1 U8682 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10336), .Z(n10342) );
  NAND2_X1 U8683 ( .A1(n10341), .A2(n10342), .ZN(n10340) );
  OAI21_X1 U8684 ( .B1(n7958), .B2(n7393), .A(n10340), .ZN(n10355) );
  MUX2_X1 U8685 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7395), .S(n10349), .Z(n10356) );
  NAND2_X1 U8686 ( .A1(n10355), .A2(n10356), .ZN(n10353) );
  OAI21_X1 U8687 ( .B1(n7395), .B2(n7394), .A(n10353), .ZN(n7397) );
  NOR2_X2 U8688 ( .A1(n7396), .A2(n10272), .ZN(n10354) );
  NAND2_X1 U8689 ( .A1(n7397), .A2(n7398), .ZN(n7485) );
  OAI211_X1 U8690 ( .C1(n7398), .C2(n7397), .A(n10354), .B(n7485), .ZN(n7399)
         );
  OAI211_X1 U8691 ( .C1(n7401), .C2(n7477), .A(n7400), .B(n7399), .ZN(P1_U3251) );
  INV_X1 U8692 ( .A(n7402), .ZN(n7403) );
  NAND2_X1 U8693 ( .A1(n7424), .A2(n7403), .ZN(n7409) );
  NAND2_X1 U8694 ( .A1(n7405), .A2(n7404), .ZN(n7406) );
  NOR2_X1 U8695 ( .A1(n7725), .A2(n7406), .ZN(n7408) );
  NAND2_X1 U8696 ( .A1(n7431), .A2(n7407), .ZN(n7420) );
  NAND3_X1 U8697 ( .A1(n7409), .A2(n7408), .A3(n7420), .ZN(n7410) );
  NAND2_X1 U8698 ( .A1(n7410), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7412) );
  NAND2_X1 U8699 ( .A1(n7431), .A2(n9463), .ZN(n7411) );
  NOR2_X1 U8700 ( .A1(n9606), .A2(P2_U3151), .ZN(n7476) );
  NAND2_X1 U8701 ( .A1(n7413), .A2(n9458), .ZN(n7415) );
  NAND2_X1 U8702 ( .A1(n9302), .A2(n7734), .ZN(n7414) );
  NAND2_X4 U8703 ( .A1(n7415), .A2(n7414), .ZN(n9513) );
  OAI21_X1 U8704 ( .B1(n9510), .B2(n7564), .A(n7436), .ZN(n7416) );
  OAI21_X1 U8705 ( .B1(n5145), .B2(n7416), .A(n7469), .ZN(n7423) );
  INV_X1 U8706 ( .A(n7417), .ZN(n7419) );
  OAI21_X1 U8707 ( .B1(n7424), .B2(n7419), .A(n7418), .ZN(n7422) );
  AND2_X1 U8708 ( .A1(n7420), .A2(n7425), .ZN(n7421) );
  NAND2_X1 U8709 ( .A1(n7423), .A2(n9600), .ZN(n7435) );
  NAND2_X1 U8710 ( .A1(n7424), .A2(n9026), .ZN(n7426) );
  INV_X1 U8711 ( .A(n9651), .ZN(n7568) );
  INV_X1 U8712 ( .A(n7429), .ZN(n7427) );
  NAND2_X1 U8713 ( .A1(n9463), .A2(n7427), .ZN(n7428) );
  NAND2_X1 U8714 ( .A1(n9463), .A2(n7429), .ZN(n7430) );
  OAI22_X1 U8715 ( .A1(n7568), .A2(n9613), .B1(n9626), .B2(n5427), .ZN(n7432)
         );
  AOI21_X1 U8716 ( .B1(n9629), .B2(n7433), .A(n7432), .ZN(n7434) );
  OAI211_X1 U8717 ( .C1(n7476), .C2(n7859), .A(n7435), .B(n7434), .ZN(P2_U3162) );
  NAND2_X1 U8718 ( .A1(n9651), .A2(n7747), .ZN(n9322) );
  AND2_X1 U8719 ( .A1(n7436), .A2(n9322), .ZN(n9278) );
  INV_X1 U8720 ( .A(n9278), .ZN(n7438) );
  INV_X1 U8721 ( .A(n9629), .ZN(n9609) );
  OAI22_X1 U8722 ( .A1(n9609), .A2(n7747), .B1(n5573), .B2(n9626), .ZN(n7437)
         );
  AOI21_X1 U8723 ( .B1(n9600), .B2(n7438), .A(n7437), .ZN(n7439) );
  OAI21_X1 U8724 ( .B1(n7476), .B2(n10898), .A(n7439), .ZN(P2_U3172) );
  AOI22_X1 U8725 ( .A1(n7669), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10796), .ZN(n7440) );
  OAI21_X1 U8726 ( .B1(n7468), .B2(n10799), .A(n7440), .ZN(P1_U3343) );
  AOI22_X1 U8727 ( .A1(n7443), .A2(n10892), .B1(n7442), .B2(n7441), .ZN(n10914) );
  MUX2_X1 U8728 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9756), .Z(n7444) );
  XNOR2_X1 U8729 ( .A(n7444), .B(n10912), .ZN(n10915) );
  INV_X1 U8730 ( .A(n7444), .ZN(n7445) );
  OAI22_X1 U8731 ( .A1(n10914), .A2(n10915), .B1(n7453), .B2(n7445), .ZN(n7448) );
  MUX2_X1 U8732 ( .A(n7736), .B(n7446), .S(n9756), .Z(n7709) );
  XNOR2_X1 U8733 ( .A(n7709), .B(n7708), .ZN(n7447) );
  NOR2_X1 U8734 ( .A1(n7447), .A2(n7448), .ZN(n7707) );
  AOI21_X1 U8735 ( .B1(n7448), .B2(n7447), .A(n7707), .ZN(n7466) );
  INV_X1 U8736 ( .A(n10996), .ZN(n7890) );
  INV_X1 U8737 ( .A(n11000), .ZN(n10976) );
  INV_X1 U8738 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U8739 ( .A1(n7449), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U8740 ( .A1(n7451), .A2(n7450), .ZN(n10900) );
  XNOR2_X1 U8741 ( .A(n7695), .B(n7708), .ZN(n7452) );
  NAND2_X1 U8742 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(n7452), .ZN(n7697) );
  OAI21_X1 U8743 ( .B1(n7452), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7697), .ZN(
        n7461) );
  INV_X1 U8744 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7737) );
  NOR2_X1 U8745 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7737), .ZN(n7542) );
  NAND2_X1 U8746 ( .A1(n7455), .A2(n7454), .ZN(n10905) );
  NAND2_X1 U8747 ( .A1(n7456), .A2(n7708), .ZN(n7457) );
  AOI21_X1 U8748 ( .B1(n7458), .B2(n7446), .A(n7688), .ZN(n7459) );
  NOR2_X1 U8749 ( .A1(n7459), .A2(n11011), .ZN(n7460) );
  AOI211_X1 U8750 ( .C1(n10983), .C2(n7461), .A(n7542), .B(n7460), .ZN(n7462)
         );
  OAI21_X1 U8751 ( .B1(n7463), .B2(n10940), .A(n7462), .ZN(n7464) );
  AOI21_X1 U8752 ( .B1(n7708), .B2(n10976), .A(n7464), .ZN(n7465) );
  OAI21_X1 U8753 ( .B1(n7466), .B2(n7890), .A(n7465), .ZN(P2_U3185) );
  INV_X1 U8754 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7467) );
  OAI222_X1 U8755 ( .A1(n10077), .A2(n7468), .B1(n9175), .B2(P2_U3151), .C1(
        n7467), .C2(n10070), .ZN(P2_U3283) );
  XNOR2_X1 U8756 ( .A(n9513), .B(n7805), .ZN(n7537) );
  XNOR2_X1 U8757 ( .A(n7537), .B(n6273), .ZN(n7471) );
  NAND2_X1 U8758 ( .A1(n7469), .A2(n5127), .ZN(n7470) );
  NAND2_X1 U8759 ( .A1(n7470), .A2(n7471), .ZN(n7539) );
  OAI21_X1 U8760 ( .B1(n7471), .B2(n7470), .A(n7539), .ZN(n7472) );
  NAND2_X1 U8761 ( .A1(n7472), .A2(n9600), .ZN(n7475) );
  INV_X1 U8762 ( .A(n9650), .ZN(n7789) );
  OAI22_X1 U8763 ( .A1(n5573), .A2(n9613), .B1(n9626), .B2(n7789), .ZN(n7473)
         );
  AOI21_X1 U8764 ( .B1(n9629), .B2(n5428), .A(n7473), .ZN(n7474) );
  OAI211_X1 U8765 ( .C1(n7476), .C2(n10902), .A(n7475), .B(n7474), .ZN(
        P2_U3177) );
  AOI21_X1 U8766 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7487), .A(n7477), .ZN(
        n7480) );
  INV_X1 U8767 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8671) );
  AOI22_X1 U8768 ( .A1(n7503), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8671), .B2(
        n7478), .ZN(n7479) );
  NAND2_X1 U8769 ( .A1(n7479), .A2(n7480), .ZN(n7502) );
  OAI21_X1 U8770 ( .B1(n7480), .B2(n7479), .A(n7502), .ZN(n7484) );
  INV_X1 U8771 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7482) );
  NAND2_X1 U8772 ( .A1(n10369), .A2(n7503), .ZN(n7481) );
  NAND2_X1 U8773 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n8828) );
  OAI211_X1 U8774 ( .C1(n7482), .C2(n10367), .A(n7481), .B(n8828), .ZN(n7483)
         );
  AOI21_X1 U8775 ( .B1(n10372), .B2(n7484), .A(n7483), .ZN(n7493) );
  INV_X1 U8776 ( .A(n7485), .ZN(n7486) );
  AOI21_X1 U8777 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7487), .A(n7486), .ZN(
        n7490) );
  INV_X1 U8778 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7488) );
  MUX2_X1 U8779 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7488), .S(n7503), .Z(n7489)
         );
  NAND2_X1 U8780 ( .A1(n7489), .A2(n7490), .ZN(n7495) );
  OAI21_X1 U8781 ( .B1(n7490), .B2(n7489), .A(n7495), .ZN(n7491) );
  NAND2_X1 U8782 ( .A1(n7491), .A2(n10354), .ZN(n7492) );
  NAND2_X1 U8783 ( .A1(n7493), .A2(n7492), .ZN(P1_U3252) );
  INV_X1 U8784 ( .A(n7669), .ZN(n7509) );
  INV_X1 U8785 ( .A(n10369), .ZN(n8896) );
  INV_X1 U8786 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7494) );
  MUX2_X1 U8787 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7494), .S(n7531), .Z(n7526)
         );
  OR2_X1 U8788 ( .A1(n7503), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7496) );
  AND2_X1 U8789 ( .A1(n7496), .A2(n7495), .ZN(n7527) );
  AND2_X1 U8790 ( .A1(n7526), .A2(n7527), .ZN(n7528) );
  AND2_X1 U8791 ( .A1(n7531), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7497) );
  INV_X1 U8792 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8815) );
  MUX2_X1 U8793 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n8815), .S(n7517), .Z(n7513)
         );
  AOI21_X1 U8794 ( .B1(n7517), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7516), .ZN(
        n7500) );
  INV_X1 U8795 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7498) );
  MUX2_X1 U8796 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7498), .S(n7669), .Z(n7499)
         );
  NAND2_X1 U8797 ( .A1(n7499), .A2(n7500), .ZN(n7668) );
  OAI21_X1 U8798 ( .B1(n7500), .B2(n7499), .A(n7668), .ZN(n7506) );
  INV_X1 U8799 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7501) );
  XNOR2_X1 U8800 ( .A(n7669), .B(n7501), .ZN(n7662) );
  XNOR2_X1 U8801 ( .A(n7531), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7524) );
  OAI21_X1 U8802 ( .B1(n7503), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7502), .ZN(
        n7525) );
  NOR2_X1 U8803 ( .A1(n7524), .A2(n7525), .ZN(n7523) );
  AOI21_X1 U8804 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7531), .A(n7523), .ZN(
        n7512) );
  NAND2_X1 U8805 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7517), .ZN(n7504) );
  OAI21_X1 U8806 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7517), .A(n7504), .ZN(
        n7511) );
  NOR2_X1 U8807 ( .A1(n7512), .A2(n7511), .ZN(n7510) );
  AOI21_X1 U8808 ( .B1(n7517), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7510), .ZN(
        n7661) );
  XNOR2_X1 U8809 ( .A(n7662), .B(n7661), .ZN(n7505) );
  AOI22_X1 U8810 ( .A1(n10354), .A2(n7506), .B1(n10372), .B2(n7505), .ZN(n7508) );
  AND2_X1 U8811 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9189) );
  AOI21_X1 U8812 ( .B1(n10265), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9189), .ZN(
        n7507) );
  OAI211_X1 U8813 ( .C1(n7509), .C2(n8896), .A(n7508), .B(n7507), .ZN(P1_U3255) );
  INV_X1 U8814 ( .A(n10372), .ZN(n8901) );
  AOI211_X1 U8815 ( .C1(n7512), .C2(n7511), .A(n7510), .B(n8901), .ZN(n7522)
         );
  INV_X1 U8816 ( .A(n10354), .ZN(n10360) );
  NOR2_X1 U8817 ( .A1(n7514), .A2(n7513), .ZN(n7515) );
  NOR3_X1 U8818 ( .A1(n10360), .A2(n7516), .A3(n7515), .ZN(n7521) );
  INV_X1 U8819 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U8820 ( .A1(n10369), .A2(n7517), .ZN(n7518) );
  NAND2_X1 U8821 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9061) );
  OAI211_X1 U8822 ( .C1(n7519), .C2(n10367), .A(n7518), .B(n9061), .ZN(n7520)
         );
  OR3_X1 U8823 ( .A1(n7522), .A2(n7521), .A3(n7520), .ZN(P1_U3254) );
  AOI211_X1 U8824 ( .C1(n7525), .C2(n7524), .A(n7523), .B(n8901), .ZN(n7536)
         );
  INV_X1 U8825 ( .A(n7526), .ZN(n7530) );
  INV_X1 U8826 ( .A(n7527), .ZN(n7529) );
  AOI211_X1 U8827 ( .C1(n7530), .C2(n7529), .A(n7528), .B(n10360), .ZN(n7535)
         );
  INV_X1 U8828 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U8829 ( .A1(n10369), .A2(n7531), .ZN(n7532) );
  NAND2_X1 U8830 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9093) );
  OAI211_X1 U8831 ( .C1(n7533), .C2(n10367), .A(n7532), .B(n9093), .ZN(n7534)
         );
  OR3_X1 U8832 ( .A1(n7536), .A2(n7535), .A3(n7534), .ZN(P1_U3253) );
  NAND2_X1 U8833 ( .A1(n7537), .A2(n5427), .ZN(n7538) );
  AND2_X1 U8834 ( .A1(n7539), .A2(n7538), .ZN(n7541) );
  XNOR2_X1 U8835 ( .A(n9513), .B(n7648), .ZN(n7551) );
  XNOR2_X1 U8836 ( .A(n7551), .B(n9650), .ZN(n7540) );
  OAI211_X1 U8837 ( .C1(n7541), .C2(n7540), .A(n9600), .B(n7550), .ZN(n7546)
         );
  AOI21_X1 U8838 ( .B1(n9624), .B2(n6273), .A(n7542), .ZN(n7543) );
  OAI21_X1 U8839 ( .B1(n7828), .B2(n9626), .A(n7543), .ZN(n7544) );
  AOI21_X1 U8840 ( .B1(n9629), .B2(n7821), .A(n7544), .ZN(n7545) );
  OAI211_X1 U8841 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9623), .A(n7546), .B(
        n7545), .ZN(P2_U3158) );
  AOI22_X1 U8842 ( .A1(n10370), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10796), .ZN(n7547) );
  OAI21_X1 U8843 ( .B1(n7549), .B2(n10799), .A(n7547), .ZN(P1_U3342) );
  INV_X1 U8844 ( .A(n9668), .ZN(n9658) );
  INV_X1 U8845 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7548) );
  OAI222_X1 U8846 ( .A1(n10077), .A2(n7549), .B1(n9658), .B2(P2_U3151), .C1(
        n7548), .C2(n10070), .ZN(P2_U3282) );
  XNOR2_X1 U8847 ( .A(n9513), .B(n7852), .ZN(n7552) );
  NAND2_X1 U8848 ( .A1(n7552), .A2(n7828), .ZN(n7579) );
  OAI21_X1 U8849 ( .B1(n7552), .B2(n7828), .A(n7579), .ZN(n7553) );
  AOI21_X1 U8850 ( .B1(n7554), .B2(n7553), .A(n5194), .ZN(n7561) );
  INV_X1 U8851 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7555) );
  NOR2_X1 U8852 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7555), .ZN(n10929) );
  AOI21_X1 U8853 ( .B1(n9615), .B2(n9649), .A(n10929), .ZN(n7556) );
  OAI21_X1 U8854 ( .B1(n7789), .B2(n9613), .A(n7556), .ZN(n7558) );
  NOR2_X1 U8855 ( .A1(n9623), .A2(n7851), .ZN(n7557) );
  AOI211_X1 U8856 ( .C1(n9629), .C2(n7559), .A(n7558), .B(n7557), .ZN(n7560)
         );
  OAI21_X1 U8857 ( .B1(n7561), .B2(n9632), .A(n7560), .ZN(P2_U3170) );
  NAND2_X1 U8858 ( .A1(n6271), .A2(n9936), .ZN(n7744) );
  INV_X1 U8859 ( .A(n7744), .ZN(n7563) );
  AOI21_X1 U8860 ( .B1(n9951), .B2(n10017), .A(n9278), .ZN(n7562) );
  AOI211_X1 U8861 ( .C1(n10022), .C2(n7564), .A(n7563), .B(n7562), .ZN(n11030)
         );
  OR2_X1 U8862 ( .A1(n11030), .A2(n10023), .ZN(n7565) );
  OAI21_X1 U8863 ( .B1(n10033), .B2(n7357), .A(n7565), .ZN(P2_U3459) );
  OAI21_X1 U8864 ( .B1(n9280), .B2(n9324), .A(n7566), .ZN(n7858) );
  NOR2_X1 U8865 ( .A1(n7860), .A2(n10027), .ZN(n7571) );
  NOR3_X1 U8866 ( .A1(n6269), .A2(n9951), .A3(n7747), .ZN(n7567) );
  NOR2_X1 U8867 ( .A1(n7567), .A2(n9934), .ZN(n7569) );
  OAI222_X1 U8868 ( .A1(n9956), .A2(n5427), .B1(n7570), .B2(n9951), .C1(n7569), 
        .C2(n7568), .ZN(n7863) );
  AOI211_X1 U8869 ( .C1(n10025), .C2(n7858), .A(n7571), .B(n7863), .ZN(n11032)
         );
  OR2_X1 U8870 ( .A1(n11032), .A2(n10023), .ZN(n7572) );
  OAI21_X1 U8871 ( .B1(n10033), .B2(n7573), .A(n7572), .ZN(P2_U3460) );
  INV_X1 U8872 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7575) );
  INV_X1 U8873 ( .A(n7574), .ZN(n7577) );
  OAI222_X1 U8874 ( .A1(n10070), .A2(n7575), .B1(n10087), .B2(n7577), .C1(
        P2_U3151), .C2(n9689), .ZN(P2_U3281) );
  INV_X1 U8875 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7576) );
  OAI222_X1 U8876 ( .A1(n8073), .A2(P1_U3086), .B1(n9234), .B2(n7577), .C1(
        n7576), .C2(n10792), .ZN(P1_U3341) );
  INV_X1 U8877 ( .A(P1_U3973), .ZN(n10278) );
  NAND2_X1 U8878 ( .A1(n10278), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7578) );
  OAI21_X1 U8879 ( .B1(n10450), .B2(n10278), .A(n7578), .ZN(P1_U3583) );
  INV_X1 U8880 ( .A(n7579), .ZN(n7580) );
  XNOR2_X1 U8881 ( .A(n9513), .B(n7826), .ZN(n7677) );
  XNOR2_X1 U8882 ( .A(n7677), .B(n8013), .ZN(n7581) );
  AOI21_X1 U8883 ( .B1(n7582), .B2(n7581), .A(n7681), .ZN(n7588) );
  INV_X1 U8884 ( .A(n7583), .ZN(n7870) );
  NOR2_X1 U8885 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8211), .ZN(n10950) );
  NOR2_X1 U8886 ( .A1(n9626), .A2(n8001), .ZN(n7584) );
  AOI211_X1 U8887 ( .C1(n9624), .C2(n7644), .A(n10950), .B(n7584), .ZN(n7585)
         );
  OAI21_X1 U8888 ( .B1(n7826), .B2(n9609), .A(n7585), .ZN(n7586) );
  AOI21_X1 U8889 ( .B1(n7870), .B2(n9606), .A(n7586), .ZN(n7587) );
  OAI21_X1 U8890 ( .B1(n7588), .B2(n9632), .A(n7587), .ZN(P2_U3167) );
  NAND2_X1 U8891 ( .A1(n10258), .A2(n7657), .ZN(n7617) );
  NAND2_X1 U8892 ( .A1(n7617), .A2(n7618), .ZN(n7616) );
  NAND2_X1 U8893 ( .A1(n8098), .A2(n7815), .ZN(n7589) );
  NAND2_X1 U8894 ( .A1(n7616), .A2(n7589), .ZN(n7633) );
  NAND2_X1 U8895 ( .A1(n7633), .A2(n7632), .ZN(n7631) );
  NAND2_X1 U8896 ( .A1(n7011), .A2(n8103), .ZN(n7590) );
  OAI21_X1 U8897 ( .B1(n7592), .B2(n7591), .A(n7921), .ZN(n8752) );
  NAND2_X1 U8898 ( .A1(n7594), .A2(n7593), .ZN(n7595) );
  NAND2_X1 U8899 ( .A1(n7595), .A2(n8043), .ZN(n7596) );
  OR2_X1 U8900 ( .A1(n7596), .A2(n8045), .ZN(n8094) );
  OAI22_X1 U8901 ( .A1(n8634), .A2(n10667), .B1(n7011), .B2(n10702), .ZN(n7600) );
  AOI211_X1 U8902 ( .C1(n8748), .C2(n7635), .A(n10591), .B(n8709), .ZN(n8745)
         );
  AOI211_X1 U8903 ( .C1(n8752), .C2(n11091), .A(n7600), .B(n8745), .ZN(n7607)
         );
  XNOR2_X1 U8904 ( .A(n7602), .B(n7601), .ZN(n7606) );
  OR2_X1 U8905 ( .A1(n6946), .A2(n8895), .ZN(n7605) );
  NAND2_X1 U8906 ( .A1(n6947), .A2(n7603), .ZN(n7604) );
  NAND2_X1 U8907 ( .A1(n7606), .A2(n10725), .ZN(n8754) );
  NAND2_X1 U8908 ( .A1(n7607), .A2(n8754), .ZN(n7800) );
  NAND2_X1 U8909 ( .A1(n10803), .A2(n7608), .ZN(n7609) );
  AND2_X1 U8910 ( .A1(n7612), .A2(n7611), .ZN(n7613) );
  INV_X1 U8911 ( .A(n8039), .ZN(n10785) );
  OAI22_X1 U8912 ( .A1(n10693), .A2(n7919), .B1(n11094), .B2(n7387), .ZN(n7614) );
  AOI21_X1 U8913 ( .B1(n7800), .B2(n11094), .A(n7614), .ZN(n7615) );
  INV_X1 U8914 ( .A(n7615), .ZN(P1_U3525) );
  OAI21_X1 U8915 ( .B1(n7618), .B2(n7617), .A(n7616), .ZN(n8737) );
  NAND2_X1 U8916 ( .A1(n8737), .A2(n11091), .ZN(n7625) );
  AOI22_X1 U8917 ( .A1(n10256), .A2(n10731), .B1(n10732), .B2(n10258), .ZN(
        n7624) );
  OAI21_X1 U8918 ( .B1(n7621), .B2(n7620), .A(n7619), .ZN(n7622) );
  NAND2_X1 U8919 ( .A1(n7622), .A2(n10725), .ZN(n8736) );
  AOI21_X1 U8920 ( .B1(n7657), .B2(n7009), .A(n10591), .ZN(n7623) );
  NAND2_X1 U8921 ( .A1(n7623), .A2(n7634), .ZN(n8740) );
  NAND4_X1 U8922 ( .A1(n7625), .A2(n7624), .A3(n8736), .A4(n8740), .ZN(n7817)
         );
  OAI22_X1 U8923 ( .A1(n10693), .A2(n7815), .B1(n11094), .B2(n7384), .ZN(n7626) );
  AOI21_X1 U8924 ( .B1(n11094), .B2(n7817), .A(n7626), .ZN(n7627) );
  INV_X1 U8925 ( .A(n7627), .ZN(P1_U3523) );
  AOI22_X1 U8926 ( .A1(n8080), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10796), .ZN(n7628) );
  OAI21_X1 U8927 ( .B1(n7652), .B2(n10799), .A(n7628), .ZN(P1_U3340) );
  XNOR2_X1 U8928 ( .A(n7630), .B(n7629), .ZN(n8093) );
  OAI21_X1 U8929 ( .B1(n7633), .B2(n7632), .A(n7631), .ZN(n8106) );
  INV_X1 U8930 ( .A(n8106), .ZN(n7638) );
  AOI22_X1 U8931 ( .A1(n10731), .A2(n10255), .B1(n5111), .B2(n10732), .ZN(
        n7637) );
  AOI21_X1 U8932 ( .B1(n7634), .B2(n10198), .A(n10591), .ZN(n7636) );
  NAND2_X1 U8933 ( .A1(n7636), .A2(n7635), .ZN(n8097) );
  OAI211_X1 U8934 ( .C1(n7638), .C2(n11021), .A(n7637), .B(n8097), .ZN(n7639)
         );
  AOI21_X1 U8935 ( .B1(n8093), .B2(n10725), .A(n7639), .ZN(n7797) );
  INV_X1 U8936 ( .A(n10693), .ZN(n10631) );
  AOI22_X1 U8937 ( .A1(n10631), .A2(n10198), .B1(P1_REG1_REG_2__SCAN_IN), .B2(
        n11093), .ZN(n7640) );
  OAI21_X1 U8938 ( .B1(n7797), .B2(n11093), .A(n7640), .ZN(P1_U3524) );
  OAI21_X1 U8939 ( .B1(n7642), .B2(n9279), .A(n7641), .ZN(n7724) );
  XOR2_X1 U8940 ( .A(n7643), .B(n9279), .Z(n7645) );
  AOI222_X1 U8941 ( .A1(n6325), .A2(n7645), .B1(n6273), .B2(n9934), .C1(n7644), 
        .C2(n9936), .ZN(n7735) );
  INV_X1 U8942 ( .A(n7735), .ZN(n7646) );
  AOI21_X1 U8943 ( .B1(n10025), .B2(n7724), .A(n7646), .ZN(n7823) );
  INV_X1 U8944 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7647) );
  OAI22_X1 U8945 ( .A1(n10063), .A2(n7648), .B1(n11108), .B2(n7647), .ZN(n7649) );
  INV_X1 U8946 ( .A(n7649), .ZN(n7650) );
  OAI21_X1 U8947 ( .B1(n7823), .B2(n11105), .A(n7650), .ZN(P2_U3399) );
  INV_X1 U8948 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7651) );
  OAI222_X1 U8949 ( .A1(n10077), .A2(n7652), .B1(n5213), .B2(P2_U3151), .C1(
        n7651), .C2(n10070), .ZN(P2_U3280) );
  XOR2_X1 U8950 ( .A(n7653), .B(n7654), .Z(n10273) );
  INV_X1 U8951 ( .A(n7655), .ZN(n7656) );
  NAND2_X1 U8952 ( .A1(n7656), .A2(n10803), .ZN(n10199) );
  AOI22_X1 U8953 ( .A1(n10223), .A2(n10273), .B1(n10199), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7659) );
  AOI22_X1 U8954 ( .A1(n10200), .A2(n5111), .B1(n7657), .B2(n10215), .ZN(n7658) );
  NAND2_X1 U8955 ( .A1(n7659), .A2(n7658), .ZN(P1_U3232) );
  NOR2_X1 U8956 ( .A1(n7669), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7660) );
  AOI21_X1 U8957 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n10373) );
  INV_X1 U8958 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7663) );
  XNOR2_X1 U8959 ( .A(n10370), .B(n7663), .ZN(n10374) );
  NAND2_X1 U8960 ( .A1(n10373), .A2(n10374), .ZN(n10371) );
  INV_X1 U8961 ( .A(n10371), .ZN(n7664) );
  AOI21_X1 U8962 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n10370), .A(n7664), .ZN(
        n7667) );
  NAND2_X1 U8963 ( .A1(n8065), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7665) );
  OAI21_X1 U8964 ( .B1(n8065), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7665), .ZN(
        n7666) );
  NOR2_X1 U8965 ( .A1(n7667), .A2(n7666), .ZN(n8070) );
  AOI211_X1 U8966 ( .C1(n7667), .C2(n7666), .A(n8070), .B(n8901), .ZN(n7676)
         );
  OAI21_X1 U8967 ( .B1(n7669), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7668), .ZN(
        n10362) );
  XNOR2_X1 U8968 ( .A(n10370), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n10363) );
  NOR2_X1 U8969 ( .A1(n10362), .A2(n10363), .ZN(n10361) );
  AOI21_X1 U8970 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n10370), .A(n10361), .ZN(
        n7671) );
  XNOR2_X1 U8971 ( .A(n8065), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7670) );
  NOR2_X1 U8972 ( .A1(n7671), .A2(n7670), .ZN(n8064) );
  AOI211_X1 U8973 ( .C1(n7671), .C2(n7670), .A(n8064), .B(n10360), .ZN(n7675)
         );
  INV_X1 U8974 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U8975 ( .A1(n10369), .A2(n8065), .ZN(n7672) );
  NAND2_X1 U8976 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10094) );
  OAI211_X1 U8977 ( .C1(n7673), .C2(n10367), .A(n7672), .B(n10094), .ZN(n7674)
         );
  OR3_X1 U8978 ( .A1(n7676), .A2(n7675), .A3(n7674), .ZN(P1_U3257) );
  INV_X1 U8979 ( .A(n7677), .ZN(n7678) );
  NOR2_X1 U8980 ( .A1(n7678), .A2(n9649), .ZN(n7680) );
  XNOR2_X1 U8981 ( .A(n8010), .B(n9513), .ZN(n7966) );
  XNOR2_X1 U8982 ( .A(n7966), .B(n9648), .ZN(n7679) );
  INV_X1 U8983 ( .A(n7965), .ZN(n7683) );
  OAI21_X1 U8984 ( .B1(n7681), .B2(n7680), .A(n7679), .ZN(n7682) );
  NAND3_X1 U8985 ( .A1(n7683), .A2(n9600), .A3(n7682), .ZN(n7687) );
  INV_X1 U8986 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8236) );
  NOR2_X1 U8987 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8236), .ZN(n7717) );
  AOI21_X1 U8988 ( .B1(n9624), .B2(n9649), .A(n7717), .ZN(n7684) );
  OAI21_X1 U8989 ( .B1(n8021), .B2(n9626), .A(n7684), .ZN(n7685) );
  AOI21_X1 U8990 ( .B1(n9629), .B2(n8010), .A(n7685), .ZN(n7686) );
  OAI211_X1 U8991 ( .C1(n8057), .C2(n9623), .A(n7687), .B(n7686), .ZN(P2_U3179) );
  INV_X1 U8992 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7792) );
  MUX2_X1 U8993 ( .A(n7792), .B(P2_REG1_REG_4__SCAN_IN), .S(n10934), .Z(n10920) );
  INV_X1 U8994 ( .A(n10934), .ZN(n7689) );
  NAND2_X1 U8995 ( .A1(n7689), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7690) );
  NOR2_X1 U8996 ( .A1(n10944), .A2(n7691), .ZN(n7692) );
  NOR2_X1 U8997 ( .A1(n10947), .A2(n5900), .ZN(n10946) );
  NOR2_X1 U8998 ( .A1(n7692), .A2(n10946), .ZN(n7694) );
  AOI22_X1 U8999 ( .A1(n7757), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n7749), .B2(
        n7748), .ZN(n7693) );
  NOR2_X1 U9000 ( .A1(n7694), .A2(n7693), .ZN(n7751) );
  AOI21_X1 U9001 ( .B1(n7694), .B2(n7693), .A(n7751), .ZN(n7722) );
  AOI22_X1 U9002 ( .A1(n7757), .A2(n5925), .B1(P2_REG2_REG_6__SCAN_IN), .B2(
        n7748), .ZN(n7702) );
  MUX2_X1 U9003 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n5890), .S(n10934), .Z(n10927) );
  NAND2_X1 U9004 ( .A1(n7696), .A2(n7695), .ZN(n7698) );
  NAND2_X1 U9005 ( .A1(n7705), .A2(n7699), .ZN(n7700) );
  NAND2_X1 U9006 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(n10943), .ZN(n10942) );
  OAI21_X1 U9007 ( .B1(n7702), .B2(n7701), .A(n7756), .ZN(n7720) );
  MUX2_X1 U9008 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9756), .Z(n7703) );
  NOR2_X1 U9009 ( .A1(n7703), .A2(n7748), .ZN(n7763) );
  AOI21_X1 U9010 ( .B1(n7703), .B2(n7748), .A(n7763), .ZN(n7704) );
  INV_X1 U9011 ( .A(n7704), .ZN(n7714) );
  MUX2_X1 U9012 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9756), .Z(n7711) );
  NAND2_X1 U9013 ( .A1(n7711), .A2(n7705), .ZN(n7712) );
  MUX2_X1 U9014 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9756), .Z(n7706) );
  INV_X1 U9015 ( .A(n7706), .ZN(n7710) );
  XNOR2_X1 U9016 ( .A(n7706), .B(n10934), .ZN(n10937) );
  AOI21_X1 U9017 ( .B1(n7709), .B2(n7708), .A(n7707), .ZN(n10936) );
  NAND2_X1 U9018 ( .A1(n10937), .A2(n10936), .ZN(n10935) );
  OAI21_X1 U9019 ( .B1(n10934), .B2(n7710), .A(n10935), .ZN(n10953) );
  XNOR2_X1 U9020 ( .A(n7711), .B(n10944), .ZN(n10952) );
  NAND2_X1 U9021 ( .A1(n10953), .A2(n10952), .ZN(n10951) );
  NAND2_X1 U9022 ( .A1(n7712), .A2(n10951), .ZN(n7713) );
  NOR2_X1 U9023 ( .A1(n7714), .A2(n7713), .ZN(n7762) );
  AOI21_X1 U9024 ( .B1(n7714), .B2(n7713), .A(n7762), .ZN(n7715) );
  NOR2_X1 U9025 ( .A1(n7715), .A2(n7890), .ZN(n7716) );
  AOI211_X1 U9026 ( .C1(n10999), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7717), .B(
        n7716), .ZN(n7718) );
  OAI21_X1 U9027 ( .B1(n7748), .B2(n11000), .A(n7718), .ZN(n7719) );
  AOI21_X1 U9028 ( .B1(n10983), .B2(n7720), .A(n7719), .ZN(n7721) );
  OAI21_X1 U9029 ( .B1(n7722), .B2(n11011), .A(n7721), .ZN(P2_U3188) );
  NAND2_X1 U9030 ( .A1(n10464), .A2(P1_U3973), .ZN(n7723) );
  OAI21_X1 U9031 ( .B1(n6219), .B2(P1_U3973), .A(n7723), .ZN(P1_U3580) );
  INV_X1 U9032 ( .A(n7724), .ZN(n7740) );
  OR2_X1 U9033 ( .A1(n7726), .A2(n7725), .ZN(n7729) );
  OAI22_X1 U9034 ( .A1(n7730), .A2(n7729), .B1(n7728), .B2(n7727), .ZN(n7732)
         );
  AND2_X1 U9035 ( .A1(n7734), .A2(n9323), .ZN(n7804) );
  OR2_X1 U9036 ( .A1(n8840), .A2(n7804), .ZN(n11059) );
  MUX2_X1 U9037 ( .A(n7736), .B(n7735), .S(n11069), .Z(n7739) );
  NOR2_X2 U9038 ( .A1(n7742), .A2(n9843), .ZN(n11064) );
  AOI22_X1 U9039 ( .A1(n11064), .A2(n7821), .B1(n11066), .B2(n7737), .ZN(n7738) );
  OAI211_X1 U9040 ( .C1(n7740), .C2(n9963), .A(n7739), .B(n7738), .ZN(P2_U3230) );
  NOR4_X1 U9041 ( .A1(n9278), .A2(n7742), .A3(n7741), .A4(n10022), .ZN(n7743)
         );
  AOI21_X1 U9042 ( .B1(n11066), .B2(P2_REG3_REG_0__SCAN_IN), .A(n7743), .ZN(
        n7746) );
  MUX2_X1 U9043 ( .A(n7358), .B(n7744), .S(n11069), .Z(n7745) );
  OAI211_X1 U9044 ( .C1(n7747), .C2(n9913), .A(n7746), .B(n7745), .ZN(P2_U3233) );
  NOR2_X1 U9045 ( .A1(n7766), .A2(n7752), .ZN(n7753) );
  NAND2_X1 U9046 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7877), .ZN(n7754) );
  OAI21_X1 U9047 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7877), .A(n7754), .ZN(
        n7755) );
  AOI21_X1 U9048 ( .B1(n5190), .B2(n7755), .A(n7875), .ZN(n7784) );
  AOI22_X1 U9049 ( .A1(n7772), .A2(n7771), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n7877), .ZN(n7761) );
  NAND2_X1 U9050 ( .A1(n7846), .A2(n7758), .ZN(n7759) );
  NAND2_X1 U9051 ( .A1(P2_REG2_REG_7__SCAN_IN), .A2(n7838), .ZN(n7837) );
  OAI21_X1 U9052 ( .B1(n7761), .B2(n7760), .A(n7878), .ZN(n7782) );
  NOR2_X1 U9053 ( .A1(n7763), .A2(n7762), .ZN(n7841) );
  MUX2_X1 U9054 ( .A(n7765), .B(n7764), .S(n9756), .Z(n7767) );
  NAND2_X1 U9055 ( .A1(n7767), .A2(n7766), .ZN(n7777) );
  INV_X1 U9056 ( .A(n7767), .ZN(n7768) );
  NAND2_X1 U9057 ( .A1(n7768), .A2(n7846), .ZN(n7769) );
  NAND2_X1 U9058 ( .A1(n7777), .A2(n7769), .ZN(n7840) );
  OR2_X1 U9059 ( .A1(n7841), .A2(n7840), .ZN(n7843) );
  MUX2_X1 U9060 ( .A(n7771), .B(n7770), .S(n9756), .Z(n7773) );
  NAND2_X1 U9061 ( .A1(n7773), .A2(n7772), .ZN(n7881) );
  INV_X1 U9062 ( .A(n7773), .ZN(n7774) );
  NAND2_X1 U9063 ( .A1(n7774), .A2(n7877), .ZN(n7775) );
  NAND2_X1 U9064 ( .A1(n7881), .A2(n7775), .ZN(n7776) );
  AOI21_X1 U9065 ( .B1(n7843), .B2(n7777), .A(n7776), .ZN(n7883) );
  AND3_X1 U9066 ( .A1(n7843), .A2(n7777), .A3(n7776), .ZN(n7778) );
  OAI21_X1 U9067 ( .B1(n7883), .B2(n7778), .A(n10996), .ZN(n7780) );
  NOR2_X1 U9068 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8401), .ZN(n8023) );
  AOI21_X1 U9069 ( .B1(n10999), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8023), .ZN(
        n7779) );
  OAI211_X1 U9070 ( .C1(n11000), .C2(n7877), .A(n7780), .B(n7779), .ZN(n7781)
         );
  AOI21_X1 U9071 ( .B1(n7782), .B2(n10983), .A(n7781), .ZN(n7783) );
  OAI21_X1 U9072 ( .B1(n7784), .B2(n11011), .A(n7783), .ZN(P2_U3190) );
  OAI21_X1 U9073 ( .B1(n7786), .B2(n9331), .A(n7785), .ZN(n7856) );
  NOR2_X1 U9074 ( .A1(n7852), .A2(n10027), .ZN(n7790) );
  INV_X1 U9075 ( .A(n9331), .ZN(n9282) );
  XNOR2_X1 U9076 ( .A(n7787), .B(n9282), .ZN(n7788) );
  OAI222_X1 U9077 ( .A1(n9954), .A2(n7789), .B1(n9956), .B2(n8013), .C1(n7788), 
        .C2(n9951), .ZN(n7853) );
  AOI211_X1 U9078 ( .C1(n10025), .C2(n7856), .A(n7790), .B(n7853), .ZN(n11034)
         );
  OR2_X1 U9079 ( .A1(n11034), .A2(n10023), .ZN(n7791) );
  OAI21_X1 U9080 ( .B1(n10033), .B2(n7792), .A(n7791), .ZN(P2_U3463) );
  INV_X1 U9081 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7794) );
  OAI22_X1 U9082 ( .A1(n10777), .A2(n8103), .B1(n11079), .B2(n7794), .ZN(n7795) );
  INV_X1 U9083 ( .A(n7795), .ZN(n7796) );
  OAI21_X1 U9084 ( .B1(n7797), .B2(n11095), .A(n7796), .ZN(P1_U3459) );
  INV_X1 U9085 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7798) );
  OAI22_X1 U9086 ( .A1(n10777), .A2(n7919), .B1(n11079), .B2(n7798), .ZN(n7799) );
  AOI21_X1 U9087 ( .B1(n7800), .B2(n11079), .A(n7799), .ZN(n7801) );
  INV_X1 U9088 ( .A(n7801), .ZN(P1_U3462) );
  OAI21_X1 U9089 ( .B1(n7803), .B2(n5426), .A(n7802), .ZN(n8536) );
  INV_X1 U9090 ( .A(n8536), .ZN(n7813) );
  NAND2_X1 U9091 ( .A1(n11069), .A2(n7804), .ZN(n9783) );
  OAI22_X1 U9092 ( .A1(n7805), .A2(n9843), .B1(n9957), .B2(n10902), .ZN(n7809)
         );
  XNOR2_X1 U9093 ( .A(n7806), .B(n9325), .ZN(n7807) );
  AOI222_X1 U9094 ( .A1(n6325), .A2(n7807), .B1(n9650), .B2(n9936), .C1(n6271), 
        .C2(n9934), .ZN(n8538) );
  INV_X1 U9095 ( .A(n8538), .ZN(n7808) );
  AOI211_X1 U9096 ( .C1(n8840), .C2(n8536), .A(n7809), .B(n7808), .ZN(n7810)
         );
  MUX2_X1 U9097 ( .A(n7811), .B(n7810), .S(n11069), .Z(n7812) );
  OAI21_X1 U9098 ( .B1(n7813), .B2(n9783), .A(n7812), .ZN(P2_U3231) );
  INV_X1 U9099 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7814) );
  OAI22_X1 U9100 ( .A1(n10777), .A2(n7815), .B1(n11079), .B2(n7814), .ZN(n7816) );
  AOI21_X1 U9101 ( .B1(n11079), .B2(n7817), .A(n7816), .ZN(n7818) );
  INV_X1 U9102 ( .A(n7818), .ZN(P1_U3456) );
  INV_X1 U9103 ( .A(n7819), .ZN(n7896) );
  AOI22_X1 U9104 ( .A1(n8761), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10796), .ZN(n7820) );
  OAI21_X1 U9105 ( .B1(n7896), .B2(n10799), .A(n7820), .ZN(P1_U3339) );
  INV_X1 U9106 ( .A(n10008), .ZN(n8621) );
  AOI22_X1 U9107 ( .A1(n8621), .A2(n7821), .B1(n10023), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7822) );
  OAI21_X1 U9108 ( .B1(n7823), .B2(n10023), .A(n7822), .ZN(P2_U3462) );
  OR2_X1 U9109 ( .A1(n7824), .A2(n9281), .ZN(n7825) );
  NAND2_X1 U9110 ( .A1(n8007), .A2(n7825), .ZN(n7866) );
  NOR2_X1 U9111 ( .A1(n7826), .A2(n10027), .ZN(n7832) );
  XNOR2_X1 U9112 ( .A(n7827), .B(n9281), .ZN(n7831) );
  OAI22_X1 U9113 ( .A1(n7828), .A2(n9954), .B1(n8001), .B2(n9956), .ZN(n7829)
         );
  AOI21_X1 U9114 ( .B1(n7866), .B2(n8840), .A(n7829), .ZN(n7830) );
  OAI21_X1 U9115 ( .B1(n7831), .B2(n9951), .A(n7830), .ZN(n7867) );
  AOI211_X1 U9116 ( .C1(n7833), .C2(n7866), .A(n7832), .B(n7867), .ZN(n11043)
         );
  NAND2_X1 U9117 ( .A1(n10023), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7834) );
  OAI21_X1 U9118 ( .B1(n11043), .B2(n10023), .A(n7834), .ZN(P2_U3464) );
  AOI21_X1 U9119 ( .B1(n7764), .B2(n7836), .A(n7835), .ZN(n7850) );
  OAI21_X1 U9120 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7838), .A(n7837), .ZN(
        n7848) );
  INV_X1 U9121 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7839) );
  NOR2_X1 U9122 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7839), .ZN(n7970) );
  NAND2_X1 U9123 ( .A1(n7841), .A2(n7840), .ZN(n7842) );
  AOI21_X1 U9124 ( .B1(n7843), .B2(n7842), .A(n7890), .ZN(n7844) );
  AOI211_X1 U9125 ( .C1(n10999), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7970), .B(
        n7844), .ZN(n7845) );
  OAI21_X1 U9126 ( .B1(n7846), .B2(n11000), .A(n7845), .ZN(n7847) );
  AOI21_X1 U9127 ( .B1(n7848), .B2(n10983), .A(n7847), .ZN(n7849) );
  OAI21_X1 U9128 ( .B1(n7850), .B2(n11011), .A(n7849), .ZN(P2_U3189) );
  OAI22_X1 U9129 ( .A1(n9913), .A2(n7852), .B1(n7851), .B2(n9957), .ZN(n7855)
         );
  MUX2_X1 U9130 ( .A(n7853), .B(P2_REG2_REG_4__SCAN_IN), .S(n9946), .Z(n7854)
         );
  AOI211_X1 U9131 ( .C1(n9943), .C2(n7856), .A(n7855), .B(n7854), .ZN(n7857)
         );
  INV_X1 U9132 ( .A(n7857), .ZN(P2_U3229) );
  INV_X1 U9133 ( .A(n7858), .ZN(n7865) );
  NOR2_X1 U9134 ( .A1(n11069), .A2(n7344), .ZN(n7862) );
  OAI22_X1 U9135 ( .A1(n9913), .A2(n7860), .B1(n9957), .B2(n7859), .ZN(n7861)
         );
  AOI211_X1 U9136 ( .C1(n7863), .C2(n11069), .A(n7862), .B(n7861), .ZN(n7864)
         );
  OAI21_X1 U9137 ( .B1(n7865), .B2(n9963), .A(n7864), .ZN(P2_U3232) );
  INV_X1 U9138 ( .A(n7866), .ZN(n7874) );
  INV_X1 U9139 ( .A(n7867), .ZN(n7868) );
  MUX2_X1 U9140 ( .A(n7869), .B(n7868), .S(n11069), .Z(n7873) );
  AOI22_X1 U9141 ( .A1(n11064), .A2(n7871), .B1(n11066), .B2(n7870), .ZN(n7872) );
  OAI211_X1 U9142 ( .C1(n7874), .C2(n9783), .A(n7873), .B(n7872), .ZN(P2_U3228) );
  AOI21_X1 U9143 ( .B1(n5973), .B2(n7876), .A(n8928), .ZN(n7895) );
  NAND2_X1 U9144 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7877), .ZN(n7879) );
  NAND2_X1 U9145 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n7880), .ZN(n8948) );
  OAI21_X1 U9146 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7880), .A(n8948), .ZN(
        n7893) );
  INV_X1 U9147 ( .A(n7881), .ZN(n7882) );
  NOR2_X1 U9148 ( .A1(n7883), .A2(n7882), .ZN(n7887) );
  MUX2_X1 U9149 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9756), .Z(n7884) );
  NOR2_X1 U9150 ( .A1(n7884), .A2(n8947), .ZN(n8935) );
  AOI21_X1 U9151 ( .B1(n7884), .B2(n8947), .A(n8935), .ZN(n7885) );
  INV_X1 U9152 ( .A(n7885), .ZN(n7886) );
  NOR2_X1 U9153 ( .A1(n7887), .A2(n7886), .ZN(n8934) );
  AOI21_X1 U9154 ( .B1(n7887), .B2(n7886), .A(n8934), .ZN(n7891) );
  AND2_X1 U9155 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8087) );
  NOR2_X1 U9156 ( .A1(n11000), .A2(n8947), .ZN(n7888) );
  AOI211_X1 U9157 ( .C1(n10999), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n8087), .B(
        n7888), .ZN(n7889) );
  OAI21_X1 U9158 ( .B1(n7891), .B2(n7890), .A(n7889), .ZN(n7892) );
  AOI21_X1 U9159 ( .B1(n7893), .B2(n10983), .A(n7892), .ZN(n7894) );
  OAI21_X1 U9160 ( .B1(n7895), .B2(n11011), .A(n7894), .ZN(P2_U3191) );
  INV_X1 U9161 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7897) );
  OAI222_X1 U9162 ( .A1(n10070), .A2(n7897), .B1(n10087), .B2(n7896), .C1(
        P2_U3151), .C2(n9736), .ZN(P2_U3279) );
  NOR2_X1 U9163 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7898) );
  AOI21_X1 U9164 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7898), .ZN(n10891) );
  INV_X1 U9165 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n8766) );
  INV_X1 U9166 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7899) );
  AOI22_X1 U9167 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n8766), .B2(n7899), .ZN(n10888) );
  NOR2_X1 U9168 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7900) );
  AOI21_X1 U9169 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7900), .ZN(n10885) );
  NOR2_X1 U9170 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7901) );
  AOI21_X1 U9171 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7901), .ZN(n10882) );
  NOR2_X1 U9172 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7902) );
  AOI21_X1 U9173 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7902), .ZN(n10879) );
  NOR2_X1 U9174 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7903) );
  AOI21_X1 U9175 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7903), .ZN(n10876) );
  NOR2_X1 U9176 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7904) );
  AOI21_X1 U9177 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7904), .ZN(n10873) );
  NOR2_X1 U9178 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7905) );
  AOI21_X1 U9179 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7905), .ZN(n10870) );
  NOR2_X1 U9180 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7906) );
  AOI21_X1 U9181 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7906), .ZN(n10867) );
  NOR2_X1 U9182 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7907) );
  AOI21_X1 U9183 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7907), .ZN(n10864) );
  NOR2_X1 U9184 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7908) );
  AOI21_X1 U9185 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7908), .ZN(n10861) );
  NOR2_X1 U9186 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7909) );
  AOI21_X1 U9187 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7909), .ZN(n10858) );
  NOR2_X1 U9188 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7910) );
  AOI21_X1 U9189 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7910), .ZN(n10855) );
  NOR2_X1 U9190 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7911) );
  AOI21_X1 U9191 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7911), .ZN(n10852) );
  AND2_X1 U9192 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7912) );
  NOR2_X1 U9193 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7912), .ZN(n10837) );
  INV_X1 U9194 ( .A(n10837), .ZN(n10838) );
  NAND3_X1 U9195 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10839) );
  NAND2_X1 U9196 ( .A1(n10840), .A2(n10839), .ZN(n10836) );
  NAND2_X1 U9197 ( .A1(n10838), .A2(n10836), .ZN(n10843) );
  NAND2_X1 U9198 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7913) );
  OAI21_X1 U9199 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7913), .ZN(n10842) );
  NOR2_X1 U9200 ( .A1(n10843), .A2(n10842), .ZN(n10841) );
  AOI21_X1 U9201 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10841), .ZN(n10846) );
  NAND2_X1 U9202 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7914) );
  OAI21_X1 U9203 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7914), .ZN(n10845) );
  NOR2_X1 U9204 ( .A1(n10846), .A2(n10845), .ZN(n10844) );
  AOI21_X1 U9205 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10844), .ZN(n10849) );
  NOR2_X1 U9206 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7915) );
  AOI21_X1 U9207 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7915), .ZN(n10848) );
  NAND2_X1 U9208 ( .A1(n10849), .A2(n10848), .ZN(n10847) );
  OAI21_X1 U9209 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10847), .ZN(n10851) );
  NAND2_X1 U9210 ( .A1(n10852), .A2(n10851), .ZN(n10850) );
  OAI21_X1 U9211 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10850), .ZN(n10854) );
  NAND2_X1 U9212 ( .A1(n10855), .A2(n10854), .ZN(n10853) );
  OAI21_X1 U9213 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10853), .ZN(n10857) );
  NAND2_X1 U9214 ( .A1(n10858), .A2(n10857), .ZN(n10856) );
  OAI21_X1 U9215 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10856), .ZN(n10860) );
  NAND2_X1 U9216 ( .A1(n10861), .A2(n10860), .ZN(n10859) );
  OAI21_X1 U9217 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10859), .ZN(n10863) );
  NAND2_X1 U9218 ( .A1(n10864), .A2(n10863), .ZN(n10862) );
  OAI21_X1 U9219 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10862), .ZN(n10866) );
  NAND2_X1 U9220 ( .A1(n10867), .A2(n10866), .ZN(n10865) );
  OAI21_X1 U9221 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10865), .ZN(n10869) );
  NAND2_X1 U9222 ( .A1(n10870), .A2(n10869), .ZN(n10868) );
  OAI21_X1 U9223 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10868), .ZN(n10872) );
  NAND2_X1 U9224 ( .A1(n10873), .A2(n10872), .ZN(n10871) );
  OAI21_X1 U9225 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10871), .ZN(n10875) );
  NAND2_X1 U9226 ( .A1(n10876), .A2(n10875), .ZN(n10874) );
  OAI21_X1 U9227 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10874), .ZN(n10878) );
  NAND2_X1 U9228 ( .A1(n10879), .A2(n10878), .ZN(n10877) );
  OAI21_X1 U9229 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10877), .ZN(n10881) );
  NAND2_X1 U9230 ( .A1(n10882), .A2(n10881), .ZN(n10880) );
  OAI21_X1 U9231 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10880), .ZN(n10884) );
  NAND2_X1 U9232 ( .A1(n10885), .A2(n10884), .ZN(n10883) );
  OAI21_X1 U9233 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10883), .ZN(n10887) );
  NAND2_X1 U9234 ( .A1(n10888), .A2(n10887), .ZN(n10886) );
  OAI21_X1 U9235 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10886), .ZN(n10890) );
  NAND2_X1 U9236 ( .A1(n10891), .A2(n10890), .ZN(n10889) );
  OAI21_X1 U9237 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10889), .ZN(n7918) );
  XNOR2_X1 U9238 ( .A(n7916), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7917) );
  XNOR2_X1 U9239 ( .A(n7918), .B(n7917), .ZN(ADD_1068_U4) );
  NAND2_X1 U9240 ( .A1(n8716), .A2(n7919), .ZN(n7920) );
  NAND2_X1 U9241 ( .A1(n8634), .A2(n11036), .ZN(n7923) );
  OAI21_X1 U9242 ( .B1(n7925), .B2(n7924), .A(n7948), .ZN(n11054) );
  INV_X1 U9243 ( .A(n11054), .ZN(n7932) );
  NAND2_X1 U9244 ( .A1(n7927), .A2(n7926), .ZN(n7929) );
  XNOR2_X1 U9245 ( .A(n7929), .B(n7928), .ZN(n7930) );
  AOI222_X1 U9246 ( .A1(n10725), .A2(n7930), .B1(n10254), .B2(n10732), .C1(
        n10252), .C2(n10731), .ZN(n11056) );
  NAND2_X1 U9247 ( .A1(n8709), .A2(n11036), .ZN(n8708) );
  INV_X1 U9248 ( .A(n8708), .ZN(n7931) );
  OAI211_X1 U9249 ( .C1(n7931), .C2(n7946), .A(n10542), .B(n7953), .ZN(n11051)
         );
  OAI211_X1 U9250 ( .C1(n11021), .C2(n7932), .A(n11056), .B(n11051), .ZN(n7937) );
  INV_X1 U9251 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7933) );
  OAI22_X1 U9252 ( .A1(n10777), .A2(n7946), .B1(n11079), .B2(n7933), .ZN(n7934) );
  AOI21_X1 U9253 ( .B1(n7937), .B2(n11079), .A(n7934), .ZN(n7935) );
  INV_X1 U9254 ( .A(n7935), .ZN(P1_U3468) );
  OAI22_X1 U9255 ( .A1(n10693), .A2(n7946), .B1(n11094), .B2(n7392), .ZN(n7936) );
  AOI21_X1 U9256 ( .B1(n7937), .B2(n11094), .A(n7936), .ZN(n7938) );
  INV_X1 U9257 ( .A(n7938), .ZN(P1_U3527) );
  NAND2_X1 U9258 ( .A1(n7939), .A2(n7940), .ZN(n7942) );
  XOR2_X1 U9259 ( .A(n7942), .B(n7941), .Z(n7945) );
  AOI22_X1 U9260 ( .A1(n10233), .A2(n10258), .B1(n7009), .B2(n10215), .ZN(
        n7944) );
  AOI22_X1 U9261 ( .A1(n10200), .A2(n10256), .B1(n10199), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7943) );
  OAI211_X1 U9262 ( .C1(n7945), .C2(n10243), .A(n7944), .B(n7943), .ZN(
        P1_U3222) );
  NAND2_X1 U9263 ( .A1(n8717), .A2(n7946), .ZN(n7947) );
  NAND2_X1 U9264 ( .A1(n7948), .A2(n7947), .ZN(n7950) );
  INV_X1 U9265 ( .A(n7951), .ZN(n7949) );
  NAND2_X1 U9266 ( .A1(n7950), .A2(n7949), .ZN(n7977) );
  OAI21_X1 U9267 ( .B1(n7950), .B2(n7949), .A(n7977), .ZN(n8657) );
  NAND2_X1 U9268 ( .A1(n8657), .A2(n11091), .ZN(n7957) );
  AOI22_X1 U9269 ( .A1(n10253), .A2(n10732), .B1(n10731), .B2(n10251), .ZN(
        n7956) );
  XNOR2_X1 U9270 ( .A(n7982), .B(n7951), .ZN(n7952) );
  NAND2_X1 U9271 ( .A1(n7952), .A2(n10725), .ZN(n8659) );
  NAND2_X1 U9272 ( .A1(n7953), .A2(n8651), .ZN(n7954) );
  NAND2_X1 U9273 ( .A1(n7954), .A2(n10542), .ZN(n7955) );
  OR2_X1 U9274 ( .A1(n7985), .A2(n7955), .ZN(n8654) );
  NAND4_X1 U9275 ( .A1(n7957), .A2(n7956), .A3(n8659), .A4(n8654), .ZN(n7963)
         );
  INV_X1 U9276 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7958) );
  OAI22_X1 U9277 ( .A1(n10693), .A2(n7975), .B1(n11094), .B2(n7958), .ZN(n7959) );
  AOI21_X1 U9278 ( .B1(n7963), .B2(n11094), .A(n7959), .ZN(n7960) );
  INV_X1 U9279 ( .A(n7960), .ZN(P1_U3528) );
  INV_X1 U9280 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7961) );
  OAI22_X1 U9281 ( .A1(n10777), .A2(n7975), .B1(n11079), .B2(n7961), .ZN(n7962) );
  AOI21_X1 U9282 ( .B1(n7963), .B2(n11079), .A(n7962), .ZN(n7964) );
  INV_X1 U9283 ( .A(n7964), .ZN(P1_U3471) );
  XNOR2_X1 U9284 ( .A(n8570), .B(n9513), .ZN(n8016) );
  XNOR2_X1 U9285 ( .A(n8016), .B(n8021), .ZN(n7968) );
  OAI21_X1 U9286 ( .B1(n7968), .B2(n7967), .A(n8018), .ZN(n7969) );
  NAND2_X1 U9287 ( .A1(n7969), .A2(n9600), .ZN(n7974) );
  AOI21_X1 U9288 ( .B1(n9624), .B2(n9648), .A(n7970), .ZN(n7971) );
  OAI21_X1 U9289 ( .B1(n8620), .B2(n9626), .A(n7971), .ZN(n7972) );
  AOI21_X1 U9290 ( .B1(n9629), .B2(n8570), .A(n7972), .ZN(n7973) );
  OAI211_X1 U9291 ( .C1(n8571), .C2(n9623), .A(n7974), .B(n7973), .ZN(P2_U3153) );
  NAND2_X1 U9292 ( .A1(n8698), .A2(n7975), .ZN(n7976) );
  NAND2_X1 U9293 ( .A1(n7977), .A2(n7976), .ZN(n7979) );
  NAND2_X1 U9294 ( .A1(n7979), .A2(n7984), .ZN(n8119) );
  OAI21_X1 U9295 ( .B1(n7979), .B2(n7984), .A(n8119), .ZN(n8114) );
  OAI21_X1 U9296 ( .B1(n7982), .B2(n7981), .A(n7980), .ZN(n7983) );
  NOR2_X1 U9297 ( .A1(n7983), .A2(n7984), .ZN(n8559) );
  AOI21_X1 U9298 ( .B1(n7984), .B2(n7983), .A(n8559), .ZN(n8117) );
  INV_X1 U9299 ( .A(n7985), .ZN(n7986) );
  AOI211_X1 U9300 ( .C1(n8701), .C2(n7986), .A(n10591), .B(n8555), .ZN(n8113)
         );
  OAI22_X1 U9301 ( .A1(n8698), .A2(n10702), .B1(n8697), .B2(n10667), .ZN(n7987) );
  NOR2_X1 U9302 ( .A1(n8113), .A2(n7987), .ZN(n7988) );
  OAI21_X1 U9303 ( .B1(n8117), .B2(n11020), .A(n7988), .ZN(n7989) );
  AOI21_X1 U9304 ( .B1(n11091), .B2(n8114), .A(n7989), .ZN(n7994) );
  AOI22_X1 U9305 ( .A1(n10631), .A2(n8701), .B1(n11093), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7990) );
  OAI21_X1 U9306 ( .B1(n7994), .B2(n11093), .A(n7990), .ZN(P1_U3529) );
  INV_X1 U9307 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7991) );
  OAI22_X1 U9308 ( .A1(n10777), .A2(n8110), .B1(n11079), .B2(n7991), .ZN(n7992) );
  INV_X1 U9309 ( .A(n7992), .ZN(n7993) );
  OAI21_X1 U9310 ( .B1(n7994), .B2(n11095), .A(n7993), .ZN(P1_U3474) );
  INV_X1 U9311 ( .A(n7995), .ZN(n7996) );
  AOI21_X1 U9312 ( .B1(n7998), .B2(n7997), .A(n7996), .ZN(n8576) );
  XNOR2_X1 U9313 ( .A(n7999), .B(n9348), .ZN(n8000) );
  OAI222_X1 U9314 ( .A1(n9956), .A2(n8620), .B1(n9954), .B2(n8001), .C1(n9951), 
        .C2(n8000), .ZN(n8573) );
  AOI21_X1 U9315 ( .B1(n8576), .B2(n10025), .A(n8573), .ZN(n8006) );
  INV_X1 U9316 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8002) );
  NOR2_X1 U9317 ( .A1(n11108), .A2(n8002), .ZN(n8003) );
  AOI21_X1 U9318 ( .B1(n6374), .B2(n8570), .A(n8003), .ZN(n8004) );
  OAI21_X1 U9319 ( .B1(n8006), .B2(n11105), .A(n8004), .ZN(P2_U3411) );
  AOI22_X1 U9320 ( .A1(n8621), .A2(n8570), .B1(n10023), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n8005) );
  OAI21_X1 U9321 ( .B1(n8006), .B2(n10023), .A(n8005), .ZN(P2_U3466) );
  NAND3_X1 U9322 ( .A1(n8007), .A2(n9338), .A3(n5167), .ZN(n8008) );
  NAND2_X1 U9323 ( .A1(n8009), .A2(n8008), .ZN(n8062) );
  INV_X1 U9324 ( .A(n8010), .ZN(n8058) );
  NOR2_X1 U9325 ( .A1(n8058), .A2(n10027), .ZN(n8014) );
  XNOR2_X1 U9326 ( .A(n8011), .B(n5167), .ZN(n8012) );
  OAI222_X1 U9327 ( .A1(n9956), .A2(n8021), .B1(n9954), .B2(n8013), .C1(n8012), 
        .C2(n9951), .ZN(n8059) );
  AOI211_X1 U9328 ( .C1(n10025), .C2(n8062), .A(n8014), .B(n8059), .ZN(n11058)
         );
  OR2_X1 U9329 ( .A1(n11058), .A2(n10023), .ZN(n8015) );
  OAI21_X1 U9330 ( .B1(n10033), .B2(n7749), .A(n8015), .ZN(P2_U3465) );
  XNOR2_X1 U9331 ( .A(n8548), .B(n9510), .ZN(n8019) );
  NAND2_X1 U9332 ( .A1(n8019), .A2(n9646), .ZN(n8083) );
  NAND2_X1 U9333 ( .A1(n5193), .A2(n8083), .ZN(n8020) );
  XNOR2_X1 U9334 ( .A(n8084), .B(n8020), .ZN(n8027) );
  NOR2_X1 U9335 ( .A1(n9613), .A2(n8021), .ZN(n8022) );
  AOI211_X1 U9336 ( .C1(n9615), .C2(n9645), .A(n8023), .B(n8022), .ZN(n8024)
         );
  OAI21_X1 U9337 ( .B1(n11063), .B2(n9623), .A(n8024), .ZN(n8025) );
  AOI21_X1 U9338 ( .B1(n9629), .B2(n11065), .A(n8025), .ZN(n8026) );
  OAI21_X1 U9339 ( .B1(n8027), .B2(n9632), .A(n8026), .ZN(P2_U3161) );
  AOI22_X1 U9340 ( .A1(n10200), .A2(n10253), .B1(n10233), .B2(n10255), .ZN(
        n8028) );
  NAND2_X1 U9341 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10306) );
  OAI211_X1 U9342 ( .C1(n11036), .C2(n10237), .A(n8028), .B(n10306), .ZN(n8034) );
  INV_X1 U9343 ( .A(n8030), .ZN(n8031) );
  AOI211_X1 U9344 ( .C1(n8032), .C2(n8029), .A(n10243), .B(n8031), .ZN(n8033)
         );
  AOI211_X1 U9345 ( .C1(n10241), .C2(n8710), .A(n8034), .B(n8033), .ZN(n8035)
         );
  INV_X1 U9346 ( .A(n8035), .ZN(P1_U3230) );
  AOI22_X1 U9347 ( .A1(n8877), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10796), .ZN(n8036) );
  OAI21_X1 U9348 ( .B1(n8054), .B2(n10799), .A(n8036), .ZN(P1_U3337) );
  INV_X1 U9349 ( .A(n8037), .ZN(n8056) );
  AOI22_X1 U9350 ( .A1(n8872), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10796), .ZN(n8038) );
  OAI21_X1 U9351 ( .B1(n8056), .B2(n10799), .A(n8038), .ZN(P1_U3338) );
  NAND3_X1 U9352 ( .A1(n8040), .A2(n10784), .A3(n8039), .ZN(n8041) );
  NOR2_X1 U9353 ( .A1(n8042), .A2(n8043), .ZN(n11024) );
  NAND2_X1 U9354 ( .A1(n10594), .A2(n11024), .ZN(n8051) );
  INV_X1 U9355 ( .A(n8043), .ZN(n8044) );
  NOR3_X1 U9356 ( .A1(n11019), .A2(n8045), .A3(n8044), .ZN(n8049) );
  INV_X1 U9357 ( .A(n11024), .ZN(n8047) );
  INV_X2 U9358 ( .A(n10435), .ZN(n11044) );
  NAND2_X1 U9359 ( .A1(n11044), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U9360 ( .A1(n5111), .A2(n10731), .ZN(n11022) );
  OAI211_X1 U9361 ( .C1(n8047), .C2(n8920), .A(n8046), .B(n11022), .ZN(n8048)
         );
  OAI21_X1 U9362 ( .B1(n8049), .B2(n8048), .A(n10601), .ZN(n8050) );
  OAI211_X1 U9363 ( .C1(n8052), .C2(n10601), .A(n8051), .B(n8050), .ZN(
        P1_U3293) );
  INV_X1 U9364 ( .A(n11003), .ZN(n10995) );
  INV_X1 U9365 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8053) );
  OAI222_X1 U9366 ( .A1(n10077), .A2(n8054), .B1(n10995), .B2(P2_U3151), .C1(
        n8053), .C2(n10070), .ZN(P2_U3277) );
  INV_X1 U9367 ( .A(n9764), .ZN(n9734) );
  INV_X1 U9368 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8055) );
  OAI222_X1 U9369 ( .A1(n10077), .A2(n8056), .B1(n9734), .B2(P2_U3151), .C1(
        n8055), .C2(n10070), .ZN(P2_U3278) );
  OAI22_X1 U9370 ( .A1(n9913), .A2(n8058), .B1(n8057), .B2(n9957), .ZN(n8061)
         );
  MUX2_X1 U9371 ( .A(n8059), .B(P2_REG2_REG_6__SCAN_IN), .S(n9946), .Z(n8060)
         );
  AOI211_X1 U9372 ( .C1(n9943), .C2(n8062), .A(n8061), .B(n8060), .ZN(n8063)
         );
  INV_X1 U9373 ( .A(n8063), .ZN(P2_U3227) );
  AOI21_X1 U9374 ( .B1(n8065), .B2(P1_REG1_REG_14__SCAN_IN), .A(n8064), .ZN(
        n8067) );
  INV_X1 U9375 ( .A(n8080), .ZN(n8066) );
  NOR2_X1 U9376 ( .A1(n8067), .A2(n8066), .ZN(n8596) );
  AOI21_X1 U9377 ( .B1(n8067), .B2(n8066), .A(n8596), .ZN(n8068) );
  OAI21_X1 U9378 ( .B1(n8068), .B2(P1_REG1_REG_15__SCAN_IN), .A(n10354), .ZN(
        n8082) );
  AND2_X1 U9379 ( .A1(n8068), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8595) );
  INV_X1 U9380 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U9381 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n10234) );
  OAI21_X1 U9382 ( .B1(n10367), .B2(n8069), .A(n10234), .ZN(n8079) );
  INV_X1 U9383 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8077) );
  INV_X1 U9384 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8072) );
  INV_X1 U9385 ( .A(n8070), .ZN(n8071) );
  OAI21_X1 U9386 ( .B1(n8073), .B2(n8072), .A(n8071), .ZN(n8075) );
  AND2_X1 U9387 ( .A1(n8075), .A2(n8080), .ZN(n8598) );
  INV_X1 U9388 ( .A(n8598), .ZN(n8074) );
  OAI21_X1 U9389 ( .B1(n8080), .B2(n8075), .A(n8074), .ZN(n8076) );
  NOR2_X1 U9390 ( .A1(n8077), .A2(n8076), .ZN(n8597) );
  AOI211_X1 U9391 ( .C1(n8077), .C2(n8076), .A(n8597), .B(n8901), .ZN(n8078)
         );
  AOI211_X1 U9392 ( .C1(n10369), .C2(n8080), .A(n8079), .B(n8078), .ZN(n8081)
         );
  OAI21_X1 U9393 ( .B1(n8082), .B2(n8595), .A(n8081), .ZN(P1_U3258) );
  XNOR2_X1 U9394 ( .A(n8803), .B(n9513), .ZN(n8782) );
  XNOR2_X1 U9395 ( .A(n8782), .B(n9645), .ZN(n8085) );
  NAND2_X1 U9396 ( .A1(n8086), .A2(n8085), .ZN(n8786) );
  OAI211_X1 U9397 ( .C1(n8086), .C2(n8085), .A(n8786), .B(n9600), .ZN(n8092)
         );
  INV_X1 U9398 ( .A(n8802), .ZN(n8090) );
  AOI21_X1 U9399 ( .B1(n9624), .B2(n9646), .A(n8087), .ZN(n8088) );
  OAI21_X1 U9400 ( .B1(n8836), .B2(n9626), .A(n8088), .ZN(n8089) );
  AOI21_X1 U9401 ( .B1(n9606), .B2(n8090), .A(n8089), .ZN(n8091) );
  OAI211_X1 U9402 ( .C1(n8803), .C2(n9609), .A(n8092), .B(n8091), .ZN(P2_U3171) );
  INV_X1 U9403 ( .A(n8093), .ZN(n8108) );
  AND2_X1 U9404 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  OR2_X1 U9405 ( .A1(n10596), .A2(n10702), .ZN(n10440) );
  OAI22_X1 U9406 ( .A1(n8098), .A2(n10440), .B1(n11050), .B2(n8097), .ZN(n8105) );
  INV_X1 U9407 ( .A(n8099), .ZN(n8100) );
  INV_X1 U9408 ( .A(n10540), .ZN(n8744) );
  NAND2_X1 U9409 ( .A1(n8744), .A2(n10255), .ZN(n8102) );
  AOI22_X1 U9410 ( .A1(n10596), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n11044), .ZN(n8101) );
  OAI211_X1 U9411 ( .C1(n8103), .C2(n10599), .A(n8102), .B(n8101), .ZN(n8104)
         );
  AOI211_X1 U9412 ( .C1(n11053), .C2(n8106), .A(n8105), .B(n8104), .ZN(n8107)
         );
  OAI21_X1 U9413 ( .B1(n10548), .B2(n8108), .A(n8107), .ZN(P1_U3291) );
  AOI22_X1 U9414 ( .A1(n10596), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n8702), .B2(
        n11044), .ZN(n8109) );
  OAI21_X1 U9415 ( .B1(n10599), .B2(n8110), .A(n8109), .ZN(n8112) );
  OAI22_X1 U9416 ( .A1(n8698), .A2(n10440), .B1(n10540), .B2(n8697), .ZN(n8111) );
  AOI211_X1 U9417 ( .C1(n8113), .C2(n10594), .A(n8112), .B(n8111), .ZN(n8116)
         );
  NAND2_X1 U9418 ( .A1(n8114), .A2(n11053), .ZN(n8115) );
  OAI211_X1 U9419 ( .C1(n8117), .C2(n10548), .A(n8116), .B(n8115), .ZN(
        P1_U3286) );
  OR2_X1 U9420 ( .A1(n10251), .A2(n8701), .ZN(n8118) );
  NAND2_X1 U9421 ( .A1(n8119), .A2(n8118), .ZN(n8554) );
  INV_X1 U9422 ( .A(n8560), .ZN(n8553) );
  NAND2_X1 U9423 ( .A1(n8554), .A2(n8553), .ZN(n8552) );
  INV_X1 U9424 ( .A(n8697), .ZN(n10250) );
  OR2_X1 U9425 ( .A1(n8564), .A2(n10250), .ZN(n8120) );
  NAND2_X1 U9426 ( .A1(n8552), .A2(n8120), .ZN(n8666) );
  NAND2_X1 U9427 ( .A1(n8666), .A2(n8665), .ZN(n8664) );
  OR2_X1 U9428 ( .A1(n8673), .A2(n10249), .ZN(n8122) );
  OAI21_X1 U9429 ( .B1(n8124), .B2(n8125), .A(n8679), .ZN(n8640) );
  XNOR2_X1 U9430 ( .A(n8126), .B(n8125), .ZN(n8649) );
  AOI22_X1 U9431 ( .A1(n10249), .A2(n10732), .B1(n10731), .B2(n10247), .ZN(
        n8128) );
  OAI21_X1 U9432 ( .B1(n8667), .B2(n8673), .A(n8646), .ZN(n8127) );
  NAND3_X1 U9433 ( .A1(n8127), .A2(n10542), .A3(n8680), .ZN(n8643) );
  OAI211_X1 U9434 ( .C1(n8649), .C2(n11020), .A(n8128), .B(n8643), .ZN(n8129)
         );
  AOI21_X1 U9435 ( .B1(n8640), .B2(n11091), .A(n8129), .ZN(n8134) );
  AOI22_X1 U9436 ( .A1(n8646), .A2(n10631), .B1(n11093), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n8130) );
  OAI21_X1 U9437 ( .B1(n8134), .B2(n11093), .A(n8130), .ZN(P1_U3532) );
  INV_X1 U9438 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8131) );
  OAI22_X1 U9439 ( .A1(n9092), .A2(n10777), .B1(n11079), .B2(n8131), .ZN(n8132) );
  INV_X1 U9440 ( .A(n8132), .ZN(n8133) );
  OAI21_X1 U9441 ( .B1(n8134), .B2(n11095), .A(n8133), .ZN(P1_U3483) );
  XOR2_X1 U9442 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .Z(n8137) );
  XNOR2_X1 U9443 ( .A(n8335), .B(keyinput_129), .ZN(n8136) );
  XNOR2_X1 U9444 ( .A(SI_29_), .B(keyinput_131), .ZN(n8135) );
  AOI21_X1 U9445 ( .B1(n8137), .B2(n8136), .A(n8135), .ZN(n8142) );
  XNOR2_X1 U9446 ( .A(n8138), .B(keyinput_132), .ZN(n8141) );
  XNOR2_X1 U9447 ( .A(n8139), .B(keyinput_130), .ZN(n8140) );
  NAND3_X1 U9448 ( .A1(n8142), .A2(n8141), .A3(n8140), .ZN(n8146) );
  XNOR2_X1 U9449 ( .A(SI_27_), .B(keyinput_133), .ZN(n8145) );
  XNOR2_X1 U9450 ( .A(n8143), .B(keyinput_134), .ZN(n8144) );
  AOI21_X1 U9451 ( .B1(n8146), .B2(n8145), .A(n8144), .ZN(n8154) );
  XNOR2_X1 U9452 ( .A(n8147), .B(keyinput_135), .ZN(n8153) );
  XNOR2_X1 U9453 ( .A(n8349), .B(keyinput_138), .ZN(n8151) );
  XNOR2_X1 U9454 ( .A(n8347), .B(keyinput_139), .ZN(n8150) );
  XNOR2_X1 U9455 ( .A(SI_23_), .B(keyinput_137), .ZN(n8149) );
  XNOR2_X1 U9456 ( .A(SI_24_), .B(keyinput_136), .ZN(n8148) );
  NOR4_X1 U9457 ( .A1(n8151), .A2(n8150), .A3(n8149), .A4(n8148), .ZN(n8152)
         );
  OAI21_X1 U9458 ( .B1(n8154), .B2(n8153), .A(n8152), .ZN(n8158) );
  XNOR2_X1 U9459 ( .A(n8354), .B(keyinput_140), .ZN(n8157) );
  XNOR2_X1 U9460 ( .A(n8155), .B(keyinput_141), .ZN(n8156) );
  NAND3_X1 U9461 ( .A1(n8158), .A2(n8157), .A3(n8156), .ZN(n8171) );
  XNOR2_X1 U9462 ( .A(n8159), .B(keyinput_142), .ZN(n8170) );
  XNOR2_X1 U9463 ( .A(n8160), .B(keyinput_146), .ZN(n8163) );
  XNOR2_X1 U9464 ( .A(SI_15_), .B(keyinput_145), .ZN(n8162) );
  XNOR2_X1 U9465 ( .A(SI_16_), .B(keyinput_144), .ZN(n8161) );
  NOR3_X1 U9466 ( .A1(n8163), .A2(n8162), .A3(n8161), .ZN(n8168) );
  XNOR2_X1 U9467 ( .A(n8164), .B(keyinput_147), .ZN(n8167) );
  XNOR2_X1 U9468 ( .A(n8165), .B(keyinput_143), .ZN(n8166) );
  NAND3_X1 U9469 ( .A1(n8168), .A2(n8167), .A3(n8166), .ZN(n8169) );
  AOI21_X1 U9470 ( .B1(n8171), .B2(n8170), .A(n8169), .ZN(n8175) );
  XOR2_X1 U9471 ( .A(SI_12_), .B(keyinput_148), .Z(n8174) );
  XNOR2_X1 U9472 ( .A(n8172), .B(keyinput_149), .ZN(n8173) );
  OAI21_X1 U9473 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(n8179) );
  XNOR2_X1 U9474 ( .A(SI_10_), .B(keyinput_150), .ZN(n8178) );
  XNOR2_X1 U9475 ( .A(n8176), .B(keyinput_151), .ZN(n8177) );
  AOI21_X1 U9476 ( .B1(n8179), .B2(n8178), .A(n8177), .ZN(n8182) );
  XNOR2_X1 U9477 ( .A(SI_8_), .B(keyinput_152), .ZN(n8181) );
  XNOR2_X1 U9478 ( .A(SI_7_), .B(keyinput_153), .ZN(n8180) );
  OAI21_X1 U9479 ( .B1(n8182), .B2(n8181), .A(n8180), .ZN(n8190) );
  XOR2_X1 U9480 ( .A(SI_4_), .B(keyinput_156), .Z(n8186) );
  XNOR2_X1 U9481 ( .A(n8379), .B(keyinput_157), .ZN(n8185) );
  XNOR2_X1 U9482 ( .A(n8378), .B(keyinput_155), .ZN(n8184) );
  XNOR2_X1 U9483 ( .A(SI_6_), .B(keyinput_154), .ZN(n8183) );
  NOR4_X1 U9484 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(n8189)
         );
  XOR2_X1 U9485 ( .A(SI_2_), .B(keyinput_158), .Z(n8188) );
  XNOR2_X1 U9486 ( .A(SI_1_), .B(keyinput_159), .ZN(n8187) );
  AOI211_X1 U9487 ( .C1(n8190), .C2(n8189), .A(n8188), .B(n8187), .ZN(n8197)
         );
  XNOR2_X1 U9488 ( .A(SI_0_), .B(keyinput_160), .ZN(n8196) );
  XOR2_X1 U9489 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .Z(n8194) );
  XNOR2_X1 U9490 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n8193) );
  XNOR2_X1 U9491 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n8192)
         );
  XNOR2_X1 U9492 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_162), .ZN(n8191) );
  NOR4_X1 U9493 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n8195)
         );
  OAI21_X1 U9494 ( .B1(n8197), .B2(n8196), .A(n8195), .ZN(n8200) );
  XOR2_X1 U9495 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n8199) );
  XNOR2_X1 U9496 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n8198)
         );
  NAND3_X1 U9497 ( .A1(n8200), .A2(n8199), .A3(n8198), .ZN(n8203) );
  XNOR2_X1 U9498 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n8202)
         );
  XNOR2_X1 U9499 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n8201) );
  AOI21_X1 U9500 ( .B1(n8203), .B2(n8202), .A(n8201), .ZN(n8210) );
  XNOR2_X1 U9501 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n8209)
         );
  XNOR2_X1 U9502 ( .A(n8204), .B(keyinput_170), .ZN(n8207) );
  XNOR2_X1 U9503 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n8206) );
  XNOR2_X1 U9504 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n8205) );
  NOR3_X1 U9505 ( .A1(n8207), .A2(n8206), .A3(n8205), .ZN(n8208) );
  OAI21_X1 U9506 ( .B1(n8210), .B2(n8209), .A(n8208), .ZN(n8218) );
  XNOR2_X1 U9507 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_173), .ZN(n8217)
         );
  XNOR2_X1 U9508 ( .A(n9559), .B(keyinput_175), .ZN(n8215) );
  XNOR2_X1 U9509 ( .A(n8211), .B(keyinput_177), .ZN(n8214) );
  XNOR2_X1 U9510 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n8213)
         );
  XNOR2_X1 U9511 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n8212)
         );
  NAND4_X1 U9512 ( .A1(n8215), .A2(n8214), .A3(n8213), .A4(n8212), .ZN(n8216)
         );
  AOI21_X1 U9513 ( .B1(n8218), .B2(n8217), .A(n8216), .ZN(n8222) );
  XNOR2_X1 U9514 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n8221)
         );
  XNOR2_X1 U9515 ( .A(n9581), .B(keyinput_179), .ZN(n8220) );
  XNOR2_X1 U9516 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n8219) );
  OAI211_X1 U9517 ( .C1(n8222), .C2(n8221), .A(n8220), .B(n8219), .ZN(n8226)
         );
  XOR2_X1 U9518 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .Z(n8225) );
  XNOR2_X1 U9519 ( .A(n8419), .B(keyinput_181), .ZN(n8224) );
  XNOR2_X1 U9520 ( .A(n9591), .B(keyinput_183), .ZN(n8223) );
  NAND4_X1 U9521 ( .A1(n8226), .A2(n8225), .A3(n8224), .A4(n8223), .ZN(n8229)
         );
  XOR2_X1 U9522 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_185), .Z(n8228) );
  XNOR2_X1 U9523 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n8227)
         );
  NAND3_X1 U9524 ( .A1(n8229), .A2(n8228), .A3(n8227), .ZN(n8232) );
  XOR2_X1 U9525 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .Z(n8231) );
  XOR2_X1 U9526 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n8230) );
  NAND3_X1 U9527 ( .A1(n8232), .A2(n8231), .A3(n8230), .ZN(n8240) );
  INV_X1 U9528 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8234) );
  OAI22_X1 U9529 ( .A1(n8234), .A2(keyinput_190), .B1(keyinput_191), .B2(
        P2_REG3_REG_15__SCAN_IN), .ZN(n8233) );
  AOI221_X1 U9530 ( .B1(n8234), .B2(keyinput_190), .C1(P2_REG3_REG_15__SCAN_IN), .C2(keyinput_191), .A(n8233), .ZN(n8239) );
  XNOR2_X1 U9531 ( .A(n8430), .B(keyinput_192), .ZN(n8238) );
  OAI22_X1 U9532 ( .A1(n8236), .A2(keyinput_189), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(keyinput_188), .ZN(n8235) );
  AOI221_X1 U9533 ( .B1(n8236), .B2(keyinput_189), .C1(keyinput_188), .C2(
        P2_REG3_REG_18__SCAN_IN), .A(n8235), .ZN(n8237) );
  NAND4_X1 U9534 ( .A1(n8240), .A2(n8239), .A3(n8238), .A4(n8237), .ZN(n8244)
         );
  XOR2_X1 U9535 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .Z(n8243) );
  XNOR2_X1 U9536 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n8242)
         );
  XNOR2_X1 U9537 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .ZN(n8241)
         );
  NAND4_X1 U9538 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n8248)
         );
  XOR2_X1 U9539 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .Z(n8247) );
  XOR2_X1 U9540 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .Z(n8246) );
  XOR2_X1 U9541 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .Z(n8245) );
  NAND4_X1 U9542 ( .A1(n8248), .A2(n8247), .A3(n8246), .A4(n8245), .ZN(n8251)
         );
  XNOR2_X1 U9543 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n8250)
         );
  XNOR2_X1 U9544 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n8249)
         );
  AOI21_X1 U9545 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8258) );
  XOR2_X1 U9546 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_201), .Z(n8257) );
  XOR2_X1 U9547 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n8255) );
  XOR2_X1 U9548 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .Z(n8254) );
  XNOR2_X1 U9549 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_204), .ZN(n8253)
         );
  XNOR2_X1 U9550 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .ZN(n8252)
         );
  NOR4_X1 U9551 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n8256)
         );
  OAI21_X1 U9552 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8262) );
  XOR2_X1 U9553 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .Z(n8261) );
  XOR2_X1 U9554 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_208), .Z(n8260) );
  XNOR2_X1 U9555 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n8259)
         );
  AOI211_X1 U9556 ( .C1(n8262), .C2(n8261), .A(n8260), .B(n8259), .ZN(n8269)
         );
  XOR2_X1 U9557 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .Z(n8266) );
  XNOR2_X1 U9558 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .ZN(n8265)
         );
  XNOR2_X1 U9559 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n8264)
         );
  XNOR2_X1 U9560 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n8263)
         );
  NAND4_X1 U9561 ( .A1(n8266), .A2(n8265), .A3(n8264), .A4(n8263), .ZN(n8268)
         );
  XOR2_X1 U9562 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .Z(n8267) );
  OAI21_X1 U9563 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8273) );
  XNOR2_X1 U9564 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n8272)
         );
  XOR2_X1 U9565 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .Z(n8271) );
  XNOR2_X1 U9566 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n8270)
         );
  AOI211_X1 U9567 ( .C1(n8273), .C2(n8272), .A(n8271), .B(n8270), .ZN(n8276)
         );
  XNOR2_X1 U9568 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n8275)
         );
  XNOR2_X1 U9569 ( .A(n8471), .B(keyinput_218), .ZN(n8274) );
  OAI21_X1 U9570 ( .B1(n8276), .B2(n8275), .A(n8274), .ZN(n8280) );
  XOR2_X1 U9571 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_219), .Z(n8279) );
  XNOR2_X1 U9572 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_220), .ZN(n8278) );
  XNOR2_X1 U9573 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_221), .ZN(n8277) );
  AOI211_X1 U9574 ( .C1(n8280), .C2(n8279), .A(n8278), .B(n8277), .ZN(n8287)
         );
  XNOR2_X1 U9575 ( .A(n8479), .B(keyinput_222), .ZN(n8286) );
  XNOR2_X1 U9576 ( .A(n8480), .B(keyinput_226), .ZN(n8284) );
  XNOR2_X1 U9577 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_225), .ZN(n8283) );
  XNOR2_X1 U9578 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_223), .ZN(n8282) );
  XNOR2_X1 U9579 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_224), .ZN(n8281) );
  NOR4_X1 U9580 ( .A1(n8284), .A2(n8283), .A3(n8282), .A4(n8281), .ZN(n8285)
         );
  OAI21_X1 U9581 ( .B1(n8287), .B2(n8286), .A(n8285), .ZN(n8291) );
  XNOR2_X1 U9582 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_227), .ZN(n8290) );
  XNOR2_X1 U9583 ( .A(n8288), .B(keyinput_228), .ZN(n8289) );
  AOI21_X1 U9584 ( .B1(n8291), .B2(n8290), .A(n8289), .ZN(n8295) );
  XNOR2_X1 U9585 ( .A(n8292), .B(keyinput_229), .ZN(n8294) );
  XNOR2_X1 U9586 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_230), .ZN(n8293) );
  OAI21_X1 U9587 ( .B1(n8295), .B2(n8294), .A(n8293), .ZN(n8299) );
  XOR2_X1 U9588 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .Z(n8298) );
  XNOR2_X1 U9589 ( .A(n8495), .B(keyinput_232), .ZN(n8297) );
  XNOR2_X1 U9590 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_233), .ZN(n8296) );
  AOI211_X1 U9591 ( .C1(n8299), .C2(n8298), .A(n8297), .B(n8296), .ZN(n8302)
         );
  XOR2_X1 U9592 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_234), .Z(n8301) );
  XNOR2_X1 U9593 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_235), .ZN(n8300) );
  NOR3_X1 U9594 ( .A1(n8302), .A2(n8301), .A3(n8300), .ZN(n8307) );
  XNOR2_X1 U9595 ( .A(n8303), .B(keyinput_236), .ZN(n8306) );
  XNOR2_X1 U9596 ( .A(n6437), .B(keyinput_237), .ZN(n8305) );
  XNOR2_X1 U9597 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_238), .ZN(n8304) );
  OAI211_X1 U9598 ( .C1(n8307), .C2(n8306), .A(n8305), .B(n8304), .ZN(n8310)
         );
  XNOR2_X1 U9599 ( .A(n8507), .B(keyinput_239), .ZN(n8309) );
  XNOR2_X1 U9600 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_240), .ZN(n8308) );
  NAND3_X1 U9601 ( .A1(n8310), .A2(n8309), .A3(n8308), .ZN(n8315) );
  XNOR2_X1 U9602 ( .A(n8511), .B(keyinput_241), .ZN(n8314) );
  XNOR2_X1 U9603 ( .A(n8311), .B(keyinput_243), .ZN(n8313) );
  XNOR2_X1 U9604 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_242), .ZN(n8312) );
  NAND4_X1 U9605 ( .A1(n8315), .A2(n8314), .A3(n8313), .A4(n8312), .ZN(n8319)
         );
  XNOR2_X1 U9606 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_244), .ZN(n8318) );
  XNOR2_X1 U9607 ( .A(n8316), .B(keyinput_245), .ZN(n8317) );
  AOI21_X1 U9608 ( .B1(n8319), .B2(n8318), .A(n8317), .ZN(n8322) );
  XNOR2_X1 U9609 ( .A(n8518), .B(keyinput_247), .ZN(n8321) );
  XNOR2_X1 U9610 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_246), .ZN(n8320) );
  NOR3_X1 U9611 ( .A1(n8322), .A2(n8321), .A3(n8320), .ZN(n8326) );
  XNOR2_X1 U9612 ( .A(n8323), .B(keyinput_248), .ZN(n8325) );
  XOR2_X1 U9613 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .Z(n8324) );
  NOR3_X1 U9614 ( .A1(n8326), .A2(n8325), .A3(n8324), .ZN(n8334) );
  XNOR2_X1 U9615 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_250), .ZN(n8333) );
  XNOR2_X1 U9616 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_254), .ZN(n8332) );
  XNOR2_X1 U9617 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_252), .ZN(n8330) );
  XNOR2_X1 U9618 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_251), .ZN(n8329) );
  XNOR2_X1 U9619 ( .A(P1_D_REG_5__SCAN_IN), .B(keyinput_255), .ZN(n8328) );
  XNOR2_X1 U9620 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_253), .ZN(n8327) );
  NAND4_X1 U9621 ( .A1(n8330), .A2(n8329), .A3(n8328), .A4(n8327), .ZN(n8331)
         );
  NOR4_X1 U9622 ( .A1(n8334), .A2(n8333), .A3(n8332), .A4(n8331), .ZN(n8535)
         );
  XOR2_X1 U9623 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n8338) );
  XNOR2_X1 U9624 ( .A(n8335), .B(keyinput_1), .ZN(n8337) );
  XNOR2_X1 U9625 ( .A(SI_28_), .B(keyinput_4), .ZN(n8336) );
  AOI21_X1 U9626 ( .B1(n8338), .B2(n8337), .A(n8336), .ZN(n8341) );
  XNOR2_X1 U9627 ( .A(SI_29_), .B(keyinput_3), .ZN(n8340) );
  XNOR2_X1 U9628 ( .A(SI_30_), .B(keyinput_2), .ZN(n8339) );
  NAND3_X1 U9629 ( .A1(n8341), .A2(n8340), .A3(n8339), .ZN(n8344) );
  XNOR2_X1 U9630 ( .A(SI_27_), .B(keyinput_5), .ZN(n8343) );
  XNOR2_X1 U9631 ( .A(SI_26_), .B(keyinput_6), .ZN(n8342) );
  AOI21_X1 U9632 ( .B1(n8344), .B2(n8343), .A(n8342), .ZN(n8346) );
  XNOR2_X1 U9633 ( .A(SI_25_), .B(keyinput_7), .ZN(n8345) );
  NOR2_X1 U9634 ( .A1(n8346), .A2(n8345), .ZN(n8358) );
  XNOR2_X1 U9635 ( .A(n8347), .B(keyinput_11), .ZN(n8353) );
  XNOR2_X1 U9636 ( .A(n8348), .B(keyinput_9), .ZN(n8352) );
  XNOR2_X1 U9637 ( .A(n8349), .B(keyinput_10), .ZN(n8351) );
  XNOR2_X1 U9638 ( .A(SI_24_), .B(keyinput_8), .ZN(n8350) );
  NAND4_X1 U9639 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n8357)
         );
  XNOR2_X1 U9640 ( .A(n8354), .B(keyinput_12), .ZN(n8356) );
  XNOR2_X1 U9641 ( .A(SI_19_), .B(keyinput_13), .ZN(n8355) );
  OAI211_X1 U9642 ( .C1(n8358), .C2(n8357), .A(n8356), .B(n8355), .ZN(n8367)
         );
  XNOR2_X1 U9643 ( .A(SI_18_), .B(keyinput_14), .ZN(n8366) );
  OAI22_X1 U9644 ( .A1(SI_17_), .A2(keyinput_15), .B1(SI_14_), .B2(keyinput_18), .ZN(n8359) );
  AOI221_X1 U9645 ( .B1(SI_17_), .B2(keyinput_15), .C1(keyinput_18), .C2(
        SI_14_), .A(n8359), .ZN(n8364) );
  OAI22_X1 U9646 ( .A1(n8361), .A2(keyinput_16), .B1(SI_13_), .B2(keyinput_19), 
        .ZN(n8360) );
  AOI221_X1 U9647 ( .B1(n8361), .B2(keyinput_16), .C1(keyinput_19), .C2(SI_13_), .A(n8360), .ZN(n8363) );
  XOR2_X1 U9648 ( .A(SI_15_), .B(keyinput_17), .Z(n8362) );
  NAND3_X1 U9649 ( .A1(n8364), .A2(n8363), .A3(n8362), .ZN(n8365) );
  AOI21_X1 U9650 ( .B1(n8367), .B2(n8366), .A(n8365), .ZN(n8370) );
  XOR2_X1 U9651 ( .A(SI_12_), .B(keyinput_20), .Z(n8369) );
  XNOR2_X1 U9652 ( .A(SI_11_), .B(keyinput_21), .ZN(n8368) );
  OAI21_X1 U9653 ( .B1(n8370), .B2(n8369), .A(n8368), .ZN(n8373) );
  XNOR2_X1 U9654 ( .A(SI_10_), .B(keyinput_22), .ZN(n8372) );
  XNOR2_X1 U9655 ( .A(SI_9_), .B(keyinput_23), .ZN(n8371) );
  AOI21_X1 U9656 ( .B1(n8373), .B2(n8372), .A(n8371), .ZN(n8377) );
  XNOR2_X1 U9657 ( .A(SI_8_), .B(keyinput_24), .ZN(n8376) );
  XNOR2_X1 U9658 ( .A(n8374), .B(keyinput_25), .ZN(n8375) );
  OAI21_X1 U9659 ( .B1(n8377), .B2(n8376), .A(n8375), .ZN(n8387) );
  XNOR2_X1 U9660 ( .A(n8378), .B(keyinput_27), .ZN(n8383) );
  XNOR2_X1 U9661 ( .A(n8379), .B(keyinput_29), .ZN(n8382) );
  XNOR2_X1 U9662 ( .A(SI_4_), .B(keyinput_28), .ZN(n8381) );
  XNOR2_X1 U9663 ( .A(SI_6_), .B(keyinput_26), .ZN(n8380) );
  NOR4_X1 U9664 ( .A1(n8383), .A2(n8382), .A3(n8381), .A4(n8380), .ZN(n8386)
         );
  XNOR2_X1 U9665 ( .A(SI_2_), .B(keyinput_30), .ZN(n8385) );
  XNOR2_X1 U9666 ( .A(SI_1_), .B(keyinput_31), .ZN(n8384) );
  AOI211_X1 U9667 ( .C1(n8387), .C2(n8386), .A(n8385), .B(n8384), .ZN(n8394)
         );
  XOR2_X1 U9668 ( .A(SI_0_), .B(keyinput_32), .Z(n8393) );
  XOR2_X1 U9669 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .Z(n8391) );
  XNOR2_X1 U9670 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n8390) );
  XNOR2_X1 U9671 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n8389) );
  XNOR2_X1 U9672 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n8388) );
  NOR4_X1 U9673 ( .A1(n8391), .A2(n8390), .A3(n8389), .A4(n8388), .ZN(n8392)
         );
  OAI21_X1 U9674 ( .B1(n8394), .B2(n8393), .A(n8392), .ZN(n8397) );
  XOR2_X1 U9675 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .Z(n8396) );
  XNOR2_X1 U9676 ( .A(keyinput_37), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n8395) );
  NAND3_X1 U9677 ( .A1(n8397), .A2(n8396), .A3(n8395), .ZN(n8400) );
  XNOR2_X1 U9678 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n8399) );
  XNOR2_X1 U9679 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n8398) );
  AOI21_X1 U9680 ( .B1(n8400), .B2(n8399), .A(n8398), .ZN(n8407) );
  XNOR2_X1 U9681 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n8406) );
  XOR2_X1 U9682 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n8404) );
  XNOR2_X1 U9683 ( .A(n8401), .B(keyinput_43), .ZN(n8403) );
  XNOR2_X1 U9684 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n8402) );
  NOR3_X1 U9685 ( .A1(n8404), .A2(n8403), .A3(n8402), .ZN(n8405) );
  OAI21_X1 U9686 ( .B1(n8407), .B2(n8406), .A(n8405), .ZN(n8414) );
  XNOR2_X1 U9687 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n8413) );
  XOR2_X1 U9688 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .Z(n8411) );
  XNOR2_X1 U9689 ( .A(n9559), .B(keyinput_47), .ZN(n8410) );
  XNOR2_X1 U9690 ( .A(n8943), .B(keyinput_46), .ZN(n8409) );
  XNOR2_X1 U9691 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n8408) );
  NAND4_X1 U9692 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(n8412)
         );
  AOI21_X1 U9693 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(n8418) );
  XNOR2_X1 U9694 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n8417) );
  XOR2_X1 U9695 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .Z(n8416) );
  XNOR2_X1 U9696 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n8415) );
  OAI211_X1 U9697 ( .C1(n8418), .C2(n8417), .A(n8416), .B(n8415), .ZN(n8423)
         );
  XOR2_X1 U9698 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n8422) );
  XNOR2_X1 U9699 ( .A(n8419), .B(keyinput_53), .ZN(n8421) );
  XNOR2_X1 U9700 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n8420) );
  NAND4_X1 U9701 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n8426)
         );
  XOR2_X1 U9702 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .Z(n8425) );
  XOR2_X1 U9703 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .Z(n8424) );
  NAND3_X1 U9704 ( .A1(n8426), .A2(n8425), .A3(n8424), .ZN(n8429) );
  XOR2_X1 U9705 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .Z(n8428) );
  XNOR2_X1 U9706 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n8427) );
  NAND3_X1 U9707 ( .A1(n8429), .A2(n8428), .A3(n8427), .ZN(n8437) );
  XOR2_X1 U9708 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .Z(n8433) );
  XOR2_X1 U9709 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_63), .Z(n8432) );
  XNOR2_X1 U9710 ( .A(n8430), .B(keyinput_64), .ZN(n8431) );
  NOR3_X1 U9711 ( .A1(n8433), .A2(n8432), .A3(n8431), .ZN(n8436) );
  XNOR2_X1 U9712 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n8435) );
  XNOR2_X1 U9713 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n8434) );
  NAND4_X1 U9714 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .ZN(n8441)
         );
  XNOR2_X1 U9715 ( .A(n9475), .B(keyinput_66), .ZN(n8440) );
  XOR2_X1 U9716 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n8439) );
  XNOR2_X1 U9717 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n8438)
         );
  NAND4_X1 U9718 ( .A1(n8441), .A2(n8440), .A3(n8439), .A4(n8438), .ZN(n8445)
         );
  XOR2_X1 U9719 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .Z(n8444) );
  XOR2_X1 U9720 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n8443) );
  XOR2_X1 U9721 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .Z(n8442) );
  NAND4_X1 U9722 ( .A1(n8445), .A2(n8444), .A3(n8443), .A4(n8442), .ZN(n8448)
         );
  XOR2_X1 U9723 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .Z(n8447) );
  XNOR2_X1 U9724 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .ZN(n8446)
         );
  AOI21_X1 U9725 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(n8455) );
  XNOR2_X1 U9726 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n8454)
         );
  XOR2_X1 U9727 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .Z(n8452) );
  XOR2_X1 U9728 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .Z(n8451) );
  XOR2_X1 U9729 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n8450) );
  XNOR2_X1 U9730 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n8449)
         );
  NOR4_X1 U9731 ( .A1(n8452), .A2(n8451), .A3(n8450), .A4(n8449), .ZN(n8453)
         );
  OAI21_X1 U9732 ( .B1(n8455), .B2(n8454), .A(n8453), .ZN(n8459) );
  XOR2_X1 U9733 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n8458) );
  XOR2_X1 U9734 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n8457) );
  XOR2_X1 U9735 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .Z(n8456) );
  AOI211_X1 U9736 ( .C1(n8459), .C2(n8458), .A(n8457), .B(n8456), .ZN(n8466)
         );
  XNOR2_X1 U9737 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n8463)
         );
  XNOR2_X1 U9738 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n8462)
         );
  XNOR2_X1 U9739 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n8461)
         );
  XNOR2_X1 U9740 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n8460)
         );
  NAND4_X1 U9741 ( .A1(n8463), .A2(n8462), .A3(n8461), .A4(n8460), .ZN(n8465)
         );
  XNOR2_X1 U9742 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n8464)
         );
  OAI21_X1 U9743 ( .B1(n8466), .B2(n8465), .A(n8464), .ZN(n8470) );
  XNOR2_X1 U9744 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n8469)
         );
  XOR2_X1 U9745 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .Z(n8468) );
  XNOR2_X1 U9746 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n8467) );
  AOI211_X1 U9747 ( .C1(n8470), .C2(n8469), .A(n8468), .B(n8467), .ZN(n8474)
         );
  XOR2_X1 U9748 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n8473) );
  XNOR2_X1 U9749 ( .A(n8471), .B(keyinput_90), .ZN(n8472) );
  OAI21_X1 U9750 ( .B1(n8474), .B2(n8473), .A(n8472), .ZN(n8478) );
  XOR2_X1 U9751 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_91), .Z(n8477) );
  XNOR2_X1 U9752 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_92), .ZN(n8476) );
  XNOR2_X1 U9753 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n8475) );
  AOI211_X1 U9754 ( .C1(n8478), .C2(n8477), .A(n8476), .B(n8475), .ZN(n8487)
         );
  XNOR2_X1 U9755 ( .A(n8479), .B(keyinput_94), .ZN(n8486) );
  XNOR2_X1 U9756 ( .A(n8480), .B(keyinput_98), .ZN(n8484) );
  XNOR2_X1 U9757 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_96), .ZN(n8483) );
  XNOR2_X1 U9758 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_95), .ZN(n8482) );
  XNOR2_X1 U9759 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_97), .ZN(n8481) );
  NOR4_X1 U9760 ( .A1(n8484), .A2(n8483), .A3(n8482), .A4(n8481), .ZN(n8485)
         );
  OAI21_X1 U9761 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8491) );
  XNOR2_X1 U9762 ( .A(n8488), .B(keyinput_99), .ZN(n8490) );
  XNOR2_X1 U9763 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_100), .ZN(n8489) );
  AOI21_X1 U9764 ( .B1(n8491), .B2(n8490), .A(n8489), .ZN(n8494) );
  XNOR2_X1 U9765 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_101), .ZN(n8493) );
  XNOR2_X1 U9766 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .ZN(n8492) );
  OAI21_X1 U9767 ( .B1(n8494), .B2(n8493), .A(n8492), .ZN(n8499) );
  XNOR2_X1 U9768 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .ZN(n8498) );
  XOR2_X1 U9769 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_105), .Z(n8497) );
  XNOR2_X1 U9770 ( .A(n8495), .B(keyinput_104), .ZN(n8496) );
  AOI211_X1 U9771 ( .C1(n8499), .C2(n8498), .A(n8497), .B(n8496), .ZN(n8502)
         );
  XNOR2_X1 U9772 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_106), .ZN(n8501) );
  XNOR2_X1 U9773 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_107), .ZN(n8500) );
  NOR3_X1 U9774 ( .A1(n8502), .A2(n8501), .A3(n8500), .ZN(n8506) );
  XNOR2_X1 U9775 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_108), .ZN(n8505) );
  XNOR2_X1 U9776 ( .A(n6437), .B(keyinput_109), .ZN(n8504) );
  XNOR2_X1 U9777 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_110), .ZN(n8503) );
  OAI211_X1 U9778 ( .C1(n8506), .C2(n8505), .A(n8504), .B(n8503), .ZN(n8510)
         );
  XNOR2_X1 U9779 ( .A(n8507), .B(keyinput_111), .ZN(n8509) );
  XNOR2_X1 U9780 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_112), .ZN(n8508) );
  NAND3_X1 U9781 ( .A1(n8510), .A2(n8509), .A3(n8508), .ZN(n8517) );
  XNOR2_X1 U9782 ( .A(n8511), .B(keyinput_113), .ZN(n8514) );
  XNOR2_X1 U9783 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_115), .ZN(n8513) );
  XNOR2_X1 U9784 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_114), .ZN(n8512) );
  NOR3_X1 U9785 ( .A1(n8514), .A2(n8513), .A3(n8512), .ZN(n8516) );
  XNOR2_X1 U9786 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .ZN(n8515) );
  AOI21_X1 U9787 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8522) );
  XNOR2_X1 U9788 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_117), .ZN(n8521) );
  XNOR2_X1 U9789 ( .A(n8518), .B(keyinput_119), .ZN(n8520) );
  XNOR2_X1 U9790 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_118), .ZN(n8519) );
  OAI211_X1 U9791 ( .C1(n8522), .C2(n8521), .A(n8520), .B(n8519), .ZN(n8525)
         );
  XNOR2_X1 U9792 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_120), .ZN(n8524) );
  XNOR2_X1 U9793 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_121), .ZN(n8523) );
  NAND3_X1 U9794 ( .A1(n8525), .A2(n8524), .A3(n8523), .ZN(n8533) );
  XOR2_X1 U9795 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_125), .Z(n8532) );
  XOR2_X1 U9796 ( .A(P1_D_REG_5__SCAN_IN), .B(keyinput_127), .Z(n8531) );
  XOR2_X1 U9797 ( .A(keyinput_126), .B(P1_D_REG_4__SCAN_IN), .Z(n8529) );
  XOR2_X1 U9798 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_124), .Z(n8528) );
  XOR2_X1 U9799 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_123), .Z(n8527) );
  XNOR2_X1 U9800 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_122), .ZN(n8526) );
  NOR4_X1 U9801 ( .A1(n8529), .A2(n8528), .A3(n8527), .A4(n8526), .ZN(n8530)
         );
  NAND4_X1 U9802 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n8534)
         );
  NAND2_X1 U9803 ( .A1(n8535), .A2(n8534), .ZN(n8540) );
  AOI22_X1 U9804 ( .A1(n8536), .A2(n10025), .B1(n10022), .B2(n5428), .ZN(n8537) );
  NAND2_X1 U9805 ( .A1(n8538), .A2(n8537), .ZN(n11033) );
  MUX2_X1 U9806 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n11033), .S(n10033), .Z(n8539) );
  XNOR2_X1 U9807 ( .A(n8540), .B(n8539), .ZN(P2_U3461) );
  XNOR2_X1 U9808 ( .A(n8541), .B(n9285), .ZN(n11061) );
  XNOR2_X1 U9809 ( .A(n8542), .B(n8543), .ZN(n8544) );
  AOI222_X1 U9810 ( .A1(n6325), .A2(n8544), .B1(n9645), .B2(n9936), .C1(n9647), 
        .C2(n9934), .ZN(n11060) );
  OAI21_X1 U9811 ( .B1(n10017), .B2(n11061), .A(n11060), .ZN(n8550) );
  INV_X1 U9812 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8545) );
  OAI22_X1 U9813 ( .A1(n8548), .A2(n10063), .B1(n11108), .B2(n8545), .ZN(n8546) );
  AOI21_X1 U9814 ( .B1(n8550), .B2(n11108), .A(n8546), .ZN(n8547) );
  INV_X1 U9815 ( .A(n8547), .ZN(P2_U3414) );
  OAI22_X1 U9816 ( .A1(n8548), .A2(n10008), .B1(n10033), .B2(n7770), .ZN(n8549) );
  AOI21_X1 U9817 ( .B1(n8550), .B2(n10033), .A(n8549), .ZN(n8551) );
  INV_X1 U9818 ( .A(n8551), .ZN(P2_U3467) );
  OAI21_X1 U9819 ( .B1(n8554), .B2(n8553), .A(n8552), .ZN(n8578) );
  OR2_X1 U9820 ( .A1(n8555), .A2(n8781), .ZN(n8556) );
  AND3_X1 U9821 ( .A1(n8667), .A2(n10542), .A3(n8556), .ZN(n8584) );
  INV_X1 U9822 ( .A(n8557), .ZN(n8558) );
  NOR2_X1 U9823 ( .A1(n8559), .A2(n8558), .ZN(n8561) );
  NAND2_X1 U9824 ( .A1(n8561), .A2(n8560), .ZN(n8661) );
  OAI211_X1 U9825 ( .C1(n8561), .C2(n8560), .A(n8661), .B(n10725), .ZN(n8563)
         );
  AOI22_X1 U9826 ( .A1(n10249), .A2(n10731), .B1(n10732), .B2(n10251), .ZN(
        n8562) );
  NAND2_X1 U9827 ( .A1(n8563), .A2(n8562), .ZN(n8579) );
  AOI211_X1 U9828 ( .C1(n11091), .C2(n8578), .A(n8584), .B(n8579), .ZN(n8569)
         );
  AOI22_X1 U9829 ( .A1(n10631), .A2(n8564), .B1(n11093), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n8565) );
  OAI21_X1 U9830 ( .B1(n8569), .B2(n11093), .A(n8565), .ZN(P1_U3530) );
  INV_X1 U9831 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8566) );
  OAI22_X1 U9832 ( .A1(n10777), .A2(n8781), .B1(n11079), .B2(n8566), .ZN(n8567) );
  INV_X1 U9833 ( .A(n8567), .ZN(n8568) );
  OAI21_X1 U9834 ( .B1(n8569), .B2(n11095), .A(n8568), .ZN(P1_U3477) );
  INV_X1 U9835 ( .A(n8570), .ZN(n8572) );
  OAI22_X1 U9836 ( .A1(n9913), .A2(n8572), .B1(n8571), .B2(n9957), .ZN(n8575)
         );
  MUX2_X1 U9837 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n8573), .S(n11069), .Z(n8574)
         );
  AOI211_X1 U9838 ( .C1(n9943), .C2(n8576), .A(n8575), .B(n8574), .ZN(n8577)
         );
  INV_X1 U9839 ( .A(n8577), .ZN(P2_U3226) );
  INV_X1 U9840 ( .A(n8578), .ZN(n8587) );
  NAND2_X1 U9841 ( .A1(n8579), .A2(n10601), .ZN(n8586) );
  NOR2_X1 U9842 ( .A1(n10599), .A2(n8781), .ZN(n8583) );
  INV_X1 U9843 ( .A(n8778), .ZN(n8580) );
  OAI22_X1 U9844 ( .A1(n10601), .A2(n8581), .B1(n8580), .B2(n10435), .ZN(n8582) );
  AOI211_X1 U9845 ( .C1(n8584), .C2(n10594), .A(n8583), .B(n8582), .ZN(n8585)
         );
  OAI211_X1 U9846 ( .C1(n8587), .C2(n10603), .A(n8586), .B(n8585), .ZN(
        P1_U3285) );
  INV_X1 U9847 ( .A(n10241), .ZN(n10212) );
  NAND2_X1 U9848 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10293) );
  INV_X1 U9849 ( .A(n10293), .ZN(n8589) );
  OAI22_X1 U9850 ( .A1(n10169), .A2(n7011), .B1(n8634), .B2(n10236), .ZN(n8588) );
  AOI211_X1 U9851 ( .C1(n8748), .C2(n10215), .A(n8589), .B(n8588), .ZN(n8594)
         );
  XNOR2_X1 U9852 ( .A(n8590), .B(n8591), .ZN(n8592) );
  NAND2_X1 U9853 ( .A1(n8592), .A2(n10223), .ZN(n8593) );
  OAI211_X1 U9854 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10212), .A(n8594), .B(
        n8593), .ZN(P1_U3218) );
  INV_X1 U9855 ( .A(n8761), .ZN(n8756) );
  NOR2_X1 U9856 ( .A1(n8596), .A2(n8595), .ZN(n8758) );
  XNOR2_X1 U9857 ( .A(n8761), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n8755) );
  XOR2_X1 U9858 ( .A(n8758), .B(n8755), .Z(n8602) );
  NOR2_X1 U9859 ( .A1(n8598), .A2(n8597), .ZN(n8600) );
  XNOR2_X1 U9860 ( .A(n8761), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n8599) );
  NOR2_X1 U9861 ( .A1(n8599), .A2(n8600), .ZN(n8760) );
  AOI211_X1 U9862 ( .C1(n8600), .C2(n8599), .A(n8760), .B(n8901), .ZN(n8601)
         );
  AOI21_X1 U9863 ( .B1(n10354), .B2(n8602), .A(n8601), .ZN(n8604) );
  AND2_X1 U9864 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10136) );
  AOI21_X1 U9865 ( .B1(n10265), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10136), .ZN(
        n8603) );
  OAI211_X1 U9866 ( .C1(n8756), .C2(n8896), .A(n8604), .B(n8603), .ZN(P1_U3259) );
  XNOR2_X1 U9867 ( .A(n8606), .B(n8605), .ZN(n8607) );
  XNOR2_X1 U9868 ( .A(n8608), .B(n8607), .ZN(n8613) );
  NAND2_X1 U9869 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10333) );
  INV_X1 U9870 ( .A(n10333), .ZN(n8610) );
  OAI22_X1 U9871 ( .A1(n10169), .A2(n8717), .B1(n8776), .B2(n10236), .ZN(n8609) );
  AOI211_X1 U9872 ( .C1(n8651), .C2(n10215), .A(n8610), .B(n8609), .ZN(n8612)
         );
  NAND2_X1 U9873 ( .A1(n10241), .A2(n8650), .ZN(n8611) );
  OAI211_X1 U9874 ( .C1(n8613), .C2(n10243), .A(n8612), .B(n8611), .ZN(
        P1_U3239) );
  INV_X1 U9875 ( .A(n8615), .ZN(n8616) );
  AOI21_X1 U9876 ( .B1(n8618), .B2(n8614), .A(n8616), .ZN(n8807) );
  XNOR2_X1 U9877 ( .A(n8617), .B(n5458), .ZN(n8619) );
  OAI222_X1 U9878 ( .A1(n9956), .A2(n8836), .B1(n9954), .B2(n8620), .C1(n9951), 
        .C2(n8619), .ZN(n8804) );
  AOI21_X1 U9879 ( .B1(n8807), .B2(n10025), .A(n8804), .ZN(n8627) );
  AOI22_X1 U9880 ( .A1(n8622), .A2(n8621), .B1(n10023), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n8623) );
  OAI21_X1 U9881 ( .B1(n8627), .B2(n10023), .A(n8623), .ZN(P2_U3468) );
  INV_X1 U9882 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8624) );
  OAI22_X1 U9883 ( .A1(n8803), .A2(n10063), .B1(n11108), .B2(n8624), .ZN(n8625) );
  INV_X1 U9884 ( .A(n8625), .ZN(n8626) );
  OAI21_X1 U9885 ( .B1(n8627), .B2(n11105), .A(n8626), .ZN(P2_U3417) );
  INV_X1 U9886 ( .A(n8628), .ZN(n8630) );
  NAND2_X1 U9887 ( .A1(n8630), .A2(n8629), .ZN(n8632) );
  XNOR2_X1 U9888 ( .A(n8632), .B(n8631), .ZN(n8633) );
  NAND2_X1 U9889 ( .A1(n8633), .A2(n10223), .ZN(n8638) );
  NAND2_X1 U9890 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10320) );
  INV_X1 U9891 ( .A(n10320), .ZN(n8636) );
  OAI22_X1 U9892 ( .A1(n10169), .A2(n8634), .B1(n8698), .B2(n10236), .ZN(n8635) );
  AOI211_X1 U9893 ( .C1(n11046), .C2(n10215), .A(n8636), .B(n8635), .ZN(n8637)
         );
  OAI211_X1 U9894 ( .C1(n10212), .C2(n8639), .A(n8638), .B(n8637), .ZN(
        P1_U3227) );
  NAND2_X1 U9895 ( .A1(n8640), .A2(n11053), .ZN(n8648) );
  NAND2_X1 U9896 ( .A1(n10536), .A2(n10249), .ZN(n8642) );
  AOI22_X1 U9897 ( .A1(n10596), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n5681), .B2(
        n11044), .ZN(n8641) );
  OAI211_X1 U9898 ( .C1(n8727), .C2(n10540), .A(n8642), .B(n8641), .ZN(n8645)
         );
  NOR2_X1 U9899 ( .A1(n8643), .A2(n11050), .ZN(n8644) );
  AOI211_X1 U9900 ( .C1(n11047), .C2(n8646), .A(n8645), .B(n8644), .ZN(n8647)
         );
  OAI211_X1 U9901 ( .C1(n8649), .C2(n10548), .A(n8648), .B(n8647), .ZN(
        P1_U3283) );
  OAI22_X1 U9902 ( .A1(n8776), .A2(n10540), .B1(n10440), .B2(n8717), .ZN(n8656) );
  AOI22_X1 U9903 ( .A1(n10596), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n8650), .B2(
        n11044), .ZN(n8653) );
  NAND2_X1 U9904 ( .A1(n11047), .A2(n8651), .ZN(n8652) );
  OAI211_X1 U9905 ( .C1(n8654), .C2(n11050), .A(n8653), .B(n8652), .ZN(n8655)
         );
  AOI211_X1 U9906 ( .C1(n8657), .C2(n11053), .A(n8656), .B(n8655), .ZN(n8658)
         );
  OAI21_X1 U9907 ( .B1(n10596), .B2(n8659), .A(n8658), .ZN(P1_U3287) );
  NAND2_X1 U9908 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  XOR2_X1 U9909 ( .A(n8665), .B(n8662), .Z(n8663) );
  OAI22_X1 U9910 ( .A1(n8663), .A2(n11020), .B1(n8697), .B2(n10702), .ZN(
        n11074) );
  INV_X1 U9911 ( .A(n11074), .ZN(n8677) );
  OAI21_X1 U9912 ( .B1(n8666), .B2(n8665), .A(n8664), .ZN(n11076) );
  XNOR2_X1 U9913 ( .A(n8667), .B(n11073), .ZN(n8669) );
  AND2_X1 U9914 ( .A1(n10248), .A2(n10731), .ZN(n8668) );
  AOI21_X1 U9915 ( .B1(n8669), .B2(n10542), .A(n8668), .ZN(n11072) );
  INV_X1 U9916 ( .A(n8833), .ZN(n8670) );
  OAI22_X1 U9917 ( .A1(n10601), .A2(n8671), .B1(n8670), .B2(n10435), .ZN(n8672) );
  AOI21_X1 U9918 ( .B1(n11047), .B2(n8673), .A(n8672), .ZN(n8674) );
  OAI21_X1 U9919 ( .B1(n11072), .B2(n11050), .A(n8674), .ZN(n8675) );
  AOI21_X1 U9920 ( .B1(n11076), .B2(n11053), .A(n8675), .ZN(n8676) );
  OAI21_X1 U9921 ( .B1(n8677), .B2(n10596), .A(n8676), .ZN(P1_U3284) );
  NAND2_X1 U9922 ( .A1(n9092), .A2(n8830), .ZN(n8678) );
  XOR2_X1 U9923 ( .A(n8726), .B(n8687), .Z(n8814) );
  NOR2_X4 U9924 ( .A1(n8680), .A2(n8681), .ZN(n8729) );
  AOI211_X1 U9925 ( .C1(n8681), .C2(n8680), .A(n10591), .B(n8729), .ZN(n8810)
         );
  NOR2_X1 U9926 ( .A1(n9064), .A2(n10599), .ZN(n8685) );
  NAND2_X1 U9927 ( .A1(n10536), .A2(n10248), .ZN(n8683) );
  AOI22_X1 U9928 ( .A1(n10596), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9067), .B2(
        n11044), .ZN(n8682) );
  OAI211_X1 U9929 ( .C1(n9063), .C2(n10540), .A(n8683), .B(n8682), .ZN(n8684)
         );
  AOI211_X1 U9930 ( .C1(n8810), .C2(n10594), .A(n8685), .B(n8684), .ZN(n8689)
         );
  XOR2_X1 U9931 ( .A(n8687), .B(n8686), .Z(n8812) );
  NAND2_X1 U9932 ( .A1(n8812), .A2(n10473), .ZN(n8688) );
  OAI211_X1 U9933 ( .C1(n8814), .C2(n10603), .A(n8689), .B(n8688), .ZN(
        P1_U3282) );
  INV_X1 U9934 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8691) );
  INV_X1 U9935 ( .A(n8690), .ZN(n8693) );
  OAI222_X1 U9936 ( .A1(n10070), .A2(n8691), .B1(n10087), .B2(n8693), .C1(
        n9762), .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U9937 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U9938 ( .A1(n5189), .A2(n8694), .ZN(n8695) );
  XNOR2_X1 U9939 ( .A(n8696), .B(n8695), .ZN(n8705) );
  NAND2_X1 U9940 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10346) );
  INV_X1 U9941 ( .A(n10346), .ZN(n8700) );
  OAI22_X1 U9942 ( .A1(n10169), .A2(n8698), .B1(n8697), .B2(n10236), .ZN(n8699) );
  AOI211_X1 U9943 ( .C1(n8701), .C2(n10215), .A(n8700), .B(n8699), .ZN(n8704)
         );
  NAND2_X1 U9944 ( .A1(n10241), .A2(n8702), .ZN(n8703) );
  OAI211_X1 U9945 ( .C1(n8705), .C2(n10243), .A(n8704), .B(n8703), .ZN(
        P1_U3213) );
  OAI21_X1 U9946 ( .B1(n8707), .B2(n8713), .A(n8706), .ZN(n11039) );
  OAI211_X1 U9947 ( .C1(n8709), .C2(n11036), .A(n8708), .B(n10542), .ZN(n11035) );
  AOI22_X1 U9948 ( .A1(n11047), .A2(n8711), .B1(n11044), .B2(n8710), .ZN(n8712) );
  OAI21_X1 U9949 ( .B1(n11050), .B2(n11035), .A(n8712), .ZN(n8719) );
  XNOR2_X1 U9950 ( .A(n8714), .B(n8713), .ZN(n8715) );
  OAI222_X1 U9951 ( .A1(n10667), .A2(n8717), .B1(n10702), .B2(n8716), .C1(
        n8715), .C2(n11020), .ZN(n11037) );
  MUX2_X1 U9952 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11037), .S(n10601), .Z(n8718) );
  AOI211_X1 U9953 ( .C1(n11053), .C2(n11039), .A(n8719), .B(n8718), .ZN(n8720)
         );
  INV_X1 U9954 ( .A(n8720), .ZN(P1_U3289) );
  NAND2_X1 U9955 ( .A1(n8722), .A2(n8721), .ZN(n8723) );
  XNOR2_X1 U9956 ( .A(n8723), .B(n8728), .ZN(n8724) );
  AOI222_X1 U9957 ( .A1(n10725), .A2(n8724), .B1(n10733), .B2(n10731), .C1(
        n10247), .C2(n10732), .ZN(n11087) );
  OR2_X1 U9958 ( .A1(n9064), .A2(n8727), .ZN(n8725) );
  XNOR2_X1 U9959 ( .A(n8852), .B(n8728), .ZN(n11092) );
  NAND2_X1 U9960 ( .A1(n11092), .A2(n11053), .ZN(n8734) );
  OAI211_X1 U9961 ( .C1(n8729), .C2(n11089), .A(n8857), .B(n10542), .ZN(n11086) );
  INV_X1 U9962 ( .A(n11086), .ZN(n8732) );
  AOI22_X1 U9963 ( .A1(n10596), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9193), .B2(
        n11044), .ZN(n8730) );
  OAI21_X1 U9964 ( .B1(n11089), .B2(n10599), .A(n8730), .ZN(n8731) );
  AOI21_X1 U9965 ( .B1(n8732), .B2(n10594), .A(n8731), .ZN(n8733) );
  OAI211_X1 U9966 ( .C1(n10596), .C2(n11087), .A(n8734), .B(n8733), .ZN(
        P1_U3281) );
  AOI22_X1 U9967 ( .A1(n10596), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n11044), .ZN(n8735) );
  OAI21_X1 U9968 ( .B1(n10596), .B2(n8736), .A(n8735), .ZN(n8742) );
  AOI22_X1 U9969 ( .A1(n11053), .A2(n8737), .B1(n11047), .B2(n7009), .ZN(n8739) );
  NAND2_X1 U9970 ( .A1(n8744), .A2(n10256), .ZN(n8738) );
  OAI211_X1 U9971 ( .C1(n8740), .C2(n11050), .A(n8739), .B(n8738), .ZN(n8741)
         );
  AOI211_X1 U9972 ( .C1(n10536), .C2(n10258), .A(n8742), .B(n8741), .ZN(n8743)
         );
  INV_X1 U9973 ( .A(n8743), .ZN(P1_U3292) );
  AOI22_X1 U9974 ( .A1(n8745), .A2(n10594), .B1(n8744), .B2(n10254), .ZN(n8750) );
  OAI22_X1 U9975 ( .A1(n10601), .A2(n8746), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10435), .ZN(n8747) );
  AOI21_X1 U9976 ( .B1(n11047), .B2(n8748), .A(n8747), .ZN(n8749) );
  OAI211_X1 U9977 ( .C1(n7011), .C2(n10440), .A(n8750), .B(n8749), .ZN(n8751)
         );
  AOI21_X1 U9978 ( .B1(n11053), .B2(n8752), .A(n8751), .ZN(n8753) );
  OAI21_X1 U9979 ( .B1(n10596), .B2(n8754), .A(n8753), .ZN(P1_U3290) );
  INV_X1 U9980 ( .A(n8755), .ZN(n8759) );
  INV_X1 U9981 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8757) );
  AOI22_X1 U9982 ( .A1(n8759), .A2(n8758), .B1(n8757), .B2(n8756), .ZN(n8874)
         );
  XNOR2_X1 U9983 ( .A(n8872), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8873) );
  XNOR2_X1 U9984 ( .A(n8874), .B(n8873), .ZN(n8765) );
  XOR2_X1 U9985 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n8872), .Z(n8763) );
  AOI21_X1 U9986 ( .B1(n8761), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8760), .ZN(
        n8762) );
  NAND2_X1 U9987 ( .A1(n8762), .A2(n8763), .ZN(n8869) );
  OAI21_X1 U9988 ( .B1(n8763), .B2(n8762), .A(n8869), .ZN(n8764) );
  AOI22_X1 U9989 ( .A1(n10354), .A2(n8765), .B1(n10372), .B2(n8764), .ZN(n8769) );
  NAND2_X1 U9990 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10148) );
  OAI21_X1 U9991 ( .B1(n10367), .B2(n8766), .A(n10148), .ZN(n8767) );
  AOI21_X1 U9992 ( .B1(n8872), .B2(n10369), .A(n8767), .ZN(n8768) );
  NAND2_X1 U9993 ( .A1(n8769), .A2(n8768), .ZN(P1_U3260) );
  OAI211_X1 U9994 ( .C1(n8772), .C2(n8771), .A(n8770), .B(n10223), .ZN(n8780)
         );
  INV_X1 U9995 ( .A(n8773), .ZN(n8774) );
  AOI21_X1 U9996 ( .B1(n10200), .B2(n10249), .A(n8774), .ZN(n8775) );
  OAI21_X1 U9997 ( .B1(n8776), .B2(n10169), .A(n8775), .ZN(n8777) );
  AOI21_X1 U9998 ( .B1(n8778), .B2(n10241), .A(n8777), .ZN(n8779) );
  OAI211_X1 U9999 ( .C1(n8781), .C2(n10237), .A(n8780), .B(n8779), .ZN(
        P1_U3221) );
  INV_X1 U10000 ( .A(n8782), .ZN(n8784) );
  NAND2_X1 U10001 ( .A1(n8784), .A2(n9645), .ZN(n8785) );
  XNOR2_X1 U10002 ( .A(n8906), .B(n9513), .ZN(n8908) );
  XNOR2_X1 U10003 ( .A(n8910), .B(n8836), .ZN(n8791) );
  AOI22_X1 U10004 ( .A1(n9615), .A2(n9643), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3151), .ZN(n8788) );
  NAND2_X1 U10005 ( .A1(n9624), .A2(n9645), .ZN(n8787) );
  OAI211_X1 U10006 ( .C1(n9623), .C2(n8846), .A(n8788), .B(n8787), .ZN(n8789)
         );
  AOI21_X1 U10007 ( .B1(n8906), .B2(n9629), .A(n8789), .ZN(n8790) );
  OAI21_X1 U10008 ( .B1(n8791), .B2(n9632), .A(n8790), .ZN(P2_U3157) );
  INV_X1 U10009 ( .A(n8795), .ZN(n9287) );
  XNOR2_X1 U10010 ( .A(n8792), .B(n9287), .ZN(n8793) );
  OAI222_X1 U10011 ( .A1(n9954), .A2(n8836), .B1(n9956), .B2(n9366), .C1(n8793), .C2(n9951), .ZN(n8922) );
  INV_X1 U10012 ( .A(n8922), .ZN(n8801) );
  OAI21_X1 U10013 ( .B1(n8796), .B2(n8795), .A(n8794), .ZN(n8924) );
  NOR2_X1 U10014 ( .A1(n8921), .A2(n9913), .ZN(n8799) );
  OAI22_X1 U10015 ( .A1(n11071), .A2(n8797), .B1(n8913), .B2(n9957), .ZN(n8798) );
  AOI211_X1 U10016 ( .C1(n8924), .C2(n9943), .A(n8799), .B(n8798), .ZN(n8800)
         );
  OAI21_X1 U10017 ( .B1(n8801), .B2(n9946), .A(n8800), .ZN(P2_U3222) );
  OAI22_X1 U10018 ( .A1(n8803), .A2(n9913), .B1(n8802), .B2(n9957), .ZN(n8806)
         );
  MUX2_X1 U10019 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8804), .S(n11069), .Z(n8805) );
  AOI211_X1 U10020 ( .C1(n9943), .C2(n8807), .A(n8806), .B(n8805), .ZN(n8808)
         );
  INV_X1 U10021 ( .A(n8808), .ZN(P2_U3224) );
  OAI222_X1 U10022 ( .A1(n10077), .A2(n8823), .B1(P2_U3151), .B2(n9302), .C1(
        n8809), .C2(n10070), .ZN(P2_U3274) );
  OAI22_X1 U10023 ( .A1(n8830), .A2(n10702), .B1(n9063), .B2(n10667), .ZN(
        n8811) );
  AOI211_X1 U10024 ( .C1(n8812), .C2(n10725), .A(n8811), .B(n8810), .ZN(n8813)
         );
  OAI21_X1 U10025 ( .B1(n8814), .B2(n11021), .A(n8813), .ZN(n8820) );
  OAI22_X1 U10026 ( .A1(n9064), .A2(n10693), .B1(n11094), .B2(n8815), .ZN(
        n8816) );
  AOI21_X1 U10027 ( .B1(n8820), .B2(n11094), .A(n8816), .ZN(n8817) );
  INV_X1 U10028 ( .A(n8817), .ZN(P1_U3533) );
  INV_X1 U10029 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8818) );
  OAI22_X1 U10030 ( .A1(n9064), .A2(n10777), .B1(n11079), .B2(n8818), .ZN(
        n8819) );
  AOI21_X1 U10031 ( .B1(n8820), .B2(n11079), .A(n8819), .ZN(n8821) );
  INV_X1 U10032 ( .A(n8821), .ZN(P1_U3486) );
  INV_X1 U10033 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8822) );
  OAI222_X1 U10034 ( .A1(P1_U3086), .A2(n8824), .B1(n10799), .B2(n8823), .C1(
        n8822), .C2(n10792), .ZN(P1_U3334) );
  OAI211_X1 U10035 ( .C1(n8827), .C2(n8826), .A(n8825), .B(n10223), .ZN(n8835)
         );
  NOR2_X1 U10036 ( .A1(n10237), .A2(n11073), .ZN(n8832) );
  NAND2_X1 U10037 ( .A1(n10233), .A2(n10250), .ZN(n8829) );
  OAI211_X1 U10038 ( .C1(n8830), .C2(n10236), .A(n8829), .B(n8828), .ZN(n8831)
         );
  AOI211_X1 U10039 ( .C1(n10241), .C2(n8833), .A(n8832), .B(n8831), .ZN(n8834)
         );
  NAND2_X1 U10040 ( .A1(n8835), .A2(n8834), .ZN(P1_U3231) );
  XNOR2_X1 U10041 ( .A(n8906), .B(n8836), .ZN(n9288) );
  XNOR2_X1 U10042 ( .A(n8837), .B(n9288), .ZN(n8841) );
  INV_X1 U10043 ( .A(n8841), .ZN(n8903) );
  INV_X1 U10044 ( .A(n9288), .ZN(n8838) );
  XNOR2_X1 U10045 ( .A(n8839), .B(n8838), .ZN(n8844) );
  NAND2_X1 U10046 ( .A1(n8841), .A2(n8840), .ZN(n8843) );
  AOI22_X1 U10047 ( .A1(n9643), .A2(n9936), .B1(n9934), .B2(n9645), .ZN(n8842)
         );
  OAI211_X1 U10048 ( .C1(n8844), .C2(n9951), .A(n8843), .B(n8842), .ZN(n8904)
         );
  MUX2_X1 U10049 ( .A(n8904), .B(P2_REG2_REG_10__SCAN_IN), .S(n9946), .Z(n8845) );
  INV_X1 U10050 ( .A(n8845), .ZN(n8849) );
  INV_X1 U10051 ( .A(n8846), .ZN(n8847) );
  AOI22_X1 U10052 ( .A1(n8906), .A2(n11064), .B1(n11066), .B2(n8847), .ZN(
        n8848) );
  OAI211_X1 U10053 ( .C1(n8903), .C2(n9783), .A(n8849), .B(n8848), .ZN(
        P2_U3223) );
  INV_X1 U10054 ( .A(n8850), .ZN(n8919) );
  OAI222_X1 U10055 ( .A1(n10087), .A2(n8919), .B1(P2_U3151), .B2(n9459), .C1(
        n8851), .C2(n10070), .ZN(P2_U3275) );
  INV_X1 U10056 ( .A(n8852), .ZN(n8853) );
  NAND2_X1 U10057 ( .A1(n8854), .A2(n10246), .ZN(n8855) );
  XNOR2_X1 U10058 ( .A(n9005), .B(n8862), .ZN(n9036) );
  INV_X1 U10059 ( .A(n9012), .ZN(n8856) );
  AOI211_X1 U10060 ( .C1(n9006), .C2(n8857), .A(n10591), .B(n8856), .ZN(n9032)
         );
  NOR2_X1 U10061 ( .A1(n10184), .A2(n10599), .ZN(n8861) );
  NAND2_X1 U10062 ( .A1(n10536), .A2(n10246), .ZN(n8859) );
  AOI22_X1 U10063 ( .A1(n10596), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n10181), 
        .B2(n11044), .ZN(n8858) );
  OAI211_X1 U10064 ( .C1(n10179), .C2(n10540), .A(n8859), .B(n8858), .ZN(n8860) );
  AOI211_X1 U10065 ( .C1(n9032), .C2(n10594), .A(n8861), .B(n8860), .ZN(n8868)
         );
  NAND3_X1 U10066 ( .A1(n8864), .A2(n8863), .A3(n8862), .ZN(n8865) );
  NAND2_X1 U10067 ( .A1(n8866), .A2(n8865), .ZN(n9034) );
  NAND2_X1 U10068 ( .A1(n9034), .A2(n10473), .ZN(n8867) );
  OAI211_X1 U10069 ( .C1(n9036), .C2(n10603), .A(n8868), .B(n8867), .ZN(
        P1_U3280) );
  NAND2_X1 U10070 ( .A1(n8877), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8883) );
  OAI21_X1 U10071 ( .B1(n8877), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8883), .ZN(
        n8871) );
  OAI21_X1 U10072 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n8872), .A(n8869), .ZN(
        n8870) );
  NOR2_X1 U10073 ( .A1(n8870), .A2(n8871), .ZN(n8885) );
  AOI211_X1 U10074 ( .C1(n8871), .C2(n8870), .A(n8885), .B(n8901), .ZN(n8882)
         );
  NAND2_X1 U10075 ( .A1(n8877), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8889) );
  OAI21_X1 U10076 ( .B1(n8877), .B2(P1_REG1_REG_18__SCAN_IN), .A(n8889), .ZN(
        n8876) );
  OAI22_X1 U10077 ( .A1(n8874), .A2(n8873), .B1(P1_REG1_REG_17__SCAN_IN), .B2(
        n8872), .ZN(n8875) );
  NOR2_X1 U10078 ( .A1(n8875), .A2(n8876), .ZN(n8891) );
  AOI211_X1 U10079 ( .C1(n8876), .C2(n8875), .A(n8891), .B(n10360), .ZN(n8881)
         );
  INV_X1 U10080 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U10081 ( .A1(n10369), .A2(n8877), .ZN(n8878) );
  NAND2_X1 U10082 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10208)
         );
  OAI211_X1 U10083 ( .C1(n8879), .C2(n10367), .A(n8878), .B(n10208), .ZN(n8880) );
  OR3_X1 U10084 ( .A1(n8882), .A2(n8881), .A3(n8880), .ZN(P1_U3261) );
  INV_X1 U10085 ( .A(n8883), .ZN(n8884) );
  NOR2_X1 U10086 ( .A1(n8885), .A2(n8884), .ZN(n8888) );
  INV_X1 U10087 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8886) );
  MUX2_X1 U10088 ( .A(n8886), .B(P1_REG2_REG_19__SCAN_IN), .S(n6773), .Z(n8887) );
  XNOR2_X1 U10089 ( .A(n8888), .B(n8887), .ZN(n8900) );
  INV_X1 U10090 ( .A(n8889), .ZN(n8890) );
  NOR2_X1 U10091 ( .A1(n8891), .A2(n8890), .ZN(n8893) );
  INV_X1 U10092 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10691) );
  XNOR2_X1 U10093 ( .A(n6773), .B(n10691), .ZN(n8892) );
  XNOR2_X1 U10094 ( .A(n8893), .B(n8892), .ZN(n8898) );
  NAND2_X1 U10095 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10111)
         );
  NAND2_X1 U10096 ( .A1(n10265), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n8894) );
  OAI211_X1 U10097 ( .C1(n8896), .C2(n8895), .A(n10111), .B(n8894), .ZN(n8897)
         );
  AOI21_X1 U10098 ( .B1(n10354), .B2(n8898), .A(n8897), .ZN(n8899) );
  OAI21_X1 U10099 ( .B1(n8901), .B2(n8900), .A(n8899), .ZN(P1_U3262) );
  NOR2_X1 U10100 ( .A1(n8903), .A2(n8902), .ZN(n8905) );
  AOI211_X1 U10101 ( .C1(n10022), .C2(n8906), .A(n8905), .B(n8904), .ZN(n11081) );
  OR2_X1 U10102 ( .A1(n11081), .A2(n10023), .ZN(n8907) );
  OAI21_X1 U10103 ( .B1(n10033), .B2(n8936), .A(n8907), .ZN(P2_U3469) );
  XNOR2_X1 U10104 ( .A(n8915), .B(n9513), .ZN(n8962) );
  XNOR2_X1 U10105 ( .A(n8962), .B(n8975), .ZN(n8964) );
  XOR2_X1 U10106 ( .A(n8965), .B(n8964), .Z(n8917) );
  AOI22_X1 U10107 ( .A1(n9615), .A2(n8994), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3151), .ZN(n8912) );
  NAND2_X1 U10108 ( .A1(n9624), .A2(n9644), .ZN(n8911) );
  OAI211_X1 U10109 ( .C1(n9623), .C2(n8913), .A(n8912), .B(n8911), .ZN(n8914)
         );
  AOI21_X1 U10110 ( .B1(n8915), .B2(n9629), .A(n8914), .ZN(n8916) );
  OAI21_X1 U10111 ( .B1(n8917), .B2(n9632), .A(n8916), .ZN(P2_U3176) );
  INV_X1 U10112 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8918) );
  OAI222_X1 U10113 ( .A1(P1_U3086), .A2(n8920), .B1(n9234), .B2(n8919), .C1(
        n8918), .C2(n10792), .ZN(P1_U3335) );
  NOR2_X1 U10114 ( .A1(n8921), .A2(n10027), .ZN(n8923) );
  AOI211_X1 U10115 ( .C1(n10025), .C2(n8924), .A(n8923), .B(n8922), .ZN(n11083) );
  OR2_X1 U10116 ( .A1(n11083), .A2(n10023), .ZN(n8925) );
  OAI21_X1 U10117 ( .B1(n10033), .B2(n6005), .A(n8925), .ZN(P2_U3470) );
  NOR2_X1 U10118 ( .A1(n8927), .A2(n8926), .ZN(n8929) );
  NAND2_X1 U10119 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n8945), .ZN(n8930) );
  OAI21_X1 U10120 ( .B1(n8945), .B2(P2_REG1_REG_10__SCAN_IN), .A(n8930), .ZN(
        n10969) );
  NOR2_X1 U10121 ( .A1(n10975), .A2(n8931), .ZN(n8932) );
  XNOR2_X1 U10122 ( .A(n10975), .B(n8931), .ZN(n10986) );
  AOI22_X1 U10123 ( .A1(n8954), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n9165), .B2(
        n9175), .ZN(n8933) );
  AOI21_X1 U10124 ( .B1(n5185), .B2(n8933), .A(n9166), .ZN(n8961) );
  MUX2_X1 U10125 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9756), .Z(n9168) );
  XNOR2_X1 U10126 ( .A(n9168), .B(n8954), .ZN(n8942) );
  MUX2_X1 U10127 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9756), .Z(n8939) );
  OR2_X1 U10128 ( .A1(n8939), .A2(n8951), .ZN(n8940) );
  NOR2_X1 U10129 ( .A1(n8935), .A2(n8934), .ZN(n10962) );
  MUX2_X1 U10130 ( .A(n8937), .B(n8936), .S(n9756), .Z(n8938) );
  NAND2_X1 U10131 ( .A1(n8938), .A2(n10957), .ZN(n10959) );
  NOR2_X1 U10132 ( .A1(n8938), .A2(n10957), .ZN(n10958) );
  AOI21_X1 U10133 ( .B1(n10962), .B2(n10959), .A(n10958), .ZN(n10979) );
  XNOR2_X1 U10134 ( .A(n8939), .B(n10975), .ZN(n10978) );
  NAND2_X1 U10135 ( .A1(n10979), .A2(n10978), .ZN(n10977) );
  NAND2_X1 U10136 ( .A1(n8940), .A2(n10977), .ZN(n8941) );
  NAND2_X1 U10137 ( .A1(n8942), .A2(n8941), .ZN(n9169) );
  OAI21_X1 U10138 ( .B1(n8942), .B2(n8941), .A(n9169), .ZN(n8959) );
  NOR2_X1 U10139 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8943), .ZN(n8969) );
  AOI21_X1 U10140 ( .B1(n10999), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8969), .ZN(
        n8944) );
  OAI21_X1 U10141 ( .B1(n9175), .B2(n11000), .A(n8944), .ZN(n8958) );
  NAND2_X1 U10142 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8945), .ZN(n8950) );
  AOI22_X1 U10143 ( .A1(n10957), .A2(n8937), .B1(P2_REG2_REG_10__SCAN_IN), 
        .B2(n8945), .ZN(n10965) );
  NAND2_X1 U10144 ( .A1(n8947), .A2(n8946), .ZN(n8949) );
  NAND2_X1 U10145 ( .A1(n8949), .A2(n8948), .ZN(n10964) );
  NAND2_X1 U10146 ( .A1(n10965), .A2(n10964), .ZN(n10963) );
  NAND2_X1 U10147 ( .A1(n8950), .A2(n10963), .ZN(n8952) );
  NAND2_X1 U10148 ( .A1(n8951), .A2(n8952), .ZN(n8953) );
  XNOR2_X1 U10149 ( .A(n10975), .B(n8952), .ZN(n10981) );
  NAND2_X1 U10150 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n10981), .ZN(n10980) );
  NAND2_X1 U10151 ( .A1(n8954), .A2(n8984), .ZN(n9174) );
  OAI21_X1 U10152 ( .B1(n8954), .B2(n8984), .A(n9174), .ZN(n8955) );
  XNOR2_X1 U10153 ( .A(n9173), .B(n8955), .ZN(n8956) );
  NOR2_X1 U10154 ( .A1(n8956), .A2(n11008), .ZN(n8957) );
  AOI211_X1 U10155 ( .C1(n10996), .C2(n8959), .A(n8958), .B(n8957), .ZN(n8960)
         );
  OAI21_X1 U10156 ( .B1(n8961), .B2(n11011), .A(n8960), .ZN(P2_U3194) );
  INV_X1 U10157 ( .A(n9367), .ZN(n8989) );
  INV_X1 U10158 ( .A(n8962), .ZN(n8963) );
  XNOR2_X1 U10159 ( .A(n9367), .B(n9513), .ZN(n8993) );
  XNOR2_X1 U10160 ( .A(n8993), .B(n9366), .ZN(n8966) );
  OAI211_X1 U10161 ( .C1(n8967), .C2(n8966), .A(n8995), .B(n9600), .ZN(n8973)
         );
  INV_X1 U10162 ( .A(n8968), .ZN(n8980) );
  AOI21_X1 U10163 ( .B1(n9624), .B2(n9643), .A(n8969), .ZN(n8970) );
  OAI21_X1 U10164 ( .B1(n9139), .B2(n9626), .A(n8970), .ZN(n8971) );
  AOI21_X1 U10165 ( .B1(n9606), .B2(n8980), .A(n8971), .ZN(n8972) );
  OAI211_X1 U10166 ( .C1(n8989), .C2(n9609), .A(n8973), .B(n8972), .ZN(
        P2_U3164) );
  AOI21_X1 U10167 ( .B1(n8974), .B2(n9372), .A(n9951), .ZN(n8978) );
  OAI22_X1 U10168 ( .A1(n9139), .A2(n9956), .B1(n8975), .B2(n9954), .ZN(n8976)
         );
  AOI21_X1 U10169 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n8988) );
  INV_X1 U10170 ( .A(n8988), .ZN(n8979) );
  AOI21_X1 U10171 ( .B1(n11066), .B2(n8980), .A(n8979), .ZN(n8987) );
  INV_X1 U10172 ( .A(n9372), .ZN(n8981) );
  NAND3_X1 U10173 ( .A1(n8794), .A2(n8981), .A3(n9361), .ZN(n8982) );
  NAND2_X1 U10174 ( .A1(n8983), .A2(n8982), .ZN(n8991) );
  OAI22_X1 U10175 ( .A1(n8989), .A2(n9913), .B1(n8984), .B2(n11069), .ZN(n8985) );
  AOI21_X1 U10176 ( .B1(n8991), .B2(n9943), .A(n8985), .ZN(n8986) );
  OAI21_X1 U10177 ( .B1(n8987), .B2(n9946), .A(n8986), .ZN(P2_U3221) );
  OAI21_X1 U10178 ( .B1(n8989), .B2(n10027), .A(n8988), .ZN(n8990) );
  AOI21_X1 U10179 ( .B1(n10025), .B2(n8991), .A(n8990), .ZN(n11085) );
  OR2_X1 U10180 ( .A1(n10033), .A2(n9165), .ZN(n8992) );
  OAI21_X1 U10181 ( .B1(n11085), .B2(n10023), .A(n8992), .ZN(P2_U3471) );
  XNOR2_X1 U10182 ( .A(n9022), .B(n9510), .ZN(n9140) );
  XNOR2_X1 U10183 ( .A(n9140), .B(n9642), .ZN(n8996) );
  XNOR2_X1 U10184 ( .A(n9143), .B(n8996), .ZN(n9002) );
  INV_X1 U10185 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8997) );
  NOR2_X1 U10186 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8997), .ZN(n9179) );
  NOR2_X1 U10187 ( .A1(n9626), .A2(n9197), .ZN(n8998) );
  AOI211_X1 U10188 ( .C1(n9624), .C2(n8994), .A(n9179), .B(n8998), .ZN(n8999)
         );
  OAI21_X1 U10189 ( .B1(n9028), .B2(n9623), .A(n8999), .ZN(n9000) );
  AOI21_X1 U10190 ( .B1(n9022), .B2(n9629), .A(n9000), .ZN(n9001) );
  OAI21_X1 U10191 ( .B1(n9002), .B2(n9632), .A(n9001), .ZN(P2_U3174) );
  OAI222_X1 U10192 ( .A1(n10077), .A2(n9113), .B1(P2_U3151), .B2(n9004), .C1(
        n9003), .C2(n10070), .ZN(P2_U3273) );
  OR2_X1 U10193 ( .A1(n9006), .A2(n10733), .ZN(n9007) );
  NAND2_X1 U10194 ( .A1(n9008), .A2(n9007), .ZN(n9077) );
  INV_X1 U10195 ( .A(n9077), .ZN(n9009) );
  NAND2_X1 U10196 ( .A1(n9009), .A2(n9017), .ZN(n9043) );
  OAI21_X1 U10197 ( .B1(n9009), .B2(n9017), .A(n9043), .ZN(n10739) );
  NAND2_X1 U10198 ( .A1(n10536), .A2(n10733), .ZN(n9011) );
  AOI22_X1 U10199 ( .A1(n10596), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n10097), 
        .B2(n11044), .ZN(n9010) );
  OAI211_X1 U10200 ( .C1(n10138), .C2(n10540), .A(n9011), .B(n9010), .ZN(n9016) );
  NAND2_X1 U10201 ( .A1(n9012), .A2(n10729), .ZN(n9013) );
  NAND2_X1 U10202 ( .A1(n9013), .A2(n10542), .ZN(n9014) );
  OR2_X1 U10203 ( .A1(n5187), .A2(n9014), .ZN(n10735) );
  NOR2_X1 U10204 ( .A1(n10735), .A2(n11050), .ZN(n9015) );
  AOI211_X1 U10205 ( .C1(n11047), .C2(n10729), .A(n9016), .B(n9015), .ZN(n9021) );
  AOI21_X1 U10206 ( .B1(n9018), .B2(n9017), .A(n11020), .ZN(n9019) );
  NAND2_X1 U10207 ( .A1(n9019), .A2(n9046), .ZN(n10737) );
  OR2_X1 U10208 ( .A1(n10737), .A2(n10596), .ZN(n9020) );
  OAI211_X1 U10209 ( .C1(n10739), .C2(n10603), .A(n9021), .B(n9020), .ZN(
        P1_U3279) );
  INV_X1 U10210 ( .A(n9022), .ZN(n9023) );
  NOR2_X1 U10211 ( .A1(n9023), .A2(n10027), .ZN(n9103) );
  NAND2_X1 U10212 ( .A1(n9375), .A2(n9374), .ZN(n9370) );
  XNOR2_X1 U10213 ( .A(n9024), .B(n9370), .ZN(n9025) );
  OAI222_X1 U10214 ( .A1(n9954), .A2(n9366), .B1(n9956), .B2(n9197), .C1(n9025), .C2(n9951), .ZN(n9102) );
  AOI21_X1 U10215 ( .B1(n9103), .B2(n9026), .A(n9102), .ZN(n9031) );
  XOR2_X1 U10216 ( .A(n9027), .B(n9370), .Z(n9104) );
  OAI22_X1 U10217 ( .A1(n11071), .A2(n6041), .B1(n9028), .B2(n9957), .ZN(n9029) );
  AOI21_X1 U10218 ( .B1(n9104), .B2(n9943), .A(n9029), .ZN(n9030) );
  OAI21_X1 U10219 ( .B1(n9031), .B2(n9946), .A(n9030), .ZN(P2_U3220) );
  INV_X1 U10220 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9038) );
  OAI22_X1 U10221 ( .A1(n9063), .A2(n10702), .B1(n10179), .B2(n10667), .ZN(
        n9033) );
  AOI211_X1 U10222 ( .C1(n10725), .C2(n9034), .A(n9033), .B(n9032), .ZN(n9035)
         );
  OAI21_X1 U10223 ( .B1(n9036), .B2(n11021), .A(n9035), .ZN(n9037) );
  INV_X1 U10224 ( .A(n9037), .ZN(n9040) );
  MUX2_X1 U10225 ( .A(n9038), .B(n9040), .S(n11094), .Z(n9039) );
  OAI21_X1 U10226 ( .B1(n10184), .B2(n10693), .A(n9039), .ZN(P1_U3535) );
  INV_X1 U10227 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9041) );
  MUX2_X1 U10228 ( .A(n9041), .B(n9040), .S(n11079), .Z(n9042) );
  OAI21_X1 U10229 ( .B1(n10184), .B2(n10777), .A(n9042), .ZN(P1_U3492) );
  NAND2_X1 U10230 ( .A1(n10729), .A2(n10720), .ZN(n9072) );
  NAND2_X1 U10231 ( .A1(n9043), .A2(n9072), .ZN(n9044) );
  XOR2_X1 U10232 ( .A(n9073), .B(n9044), .Z(n10728) );
  AND2_X1 U10233 ( .A1(n9046), .A2(n9045), .ZN(n9048) );
  OAI21_X1 U10234 ( .B1(n9048), .B2(n9073), .A(n9047), .ZN(n10726) );
  INV_X1 U10235 ( .A(n9082), .ZN(n9049) );
  OAI211_X1 U10236 ( .C1(n10723), .C2(n5187), .A(n9049), .B(n10542), .ZN(
        n10722) );
  NAND2_X1 U10237 ( .A1(n10536), .A2(n10720), .ZN(n9051) );
  AOI22_X1 U10238 ( .A1(n10596), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10240), 
        .B2(n11044), .ZN(n9050) );
  OAI211_X1 U10239 ( .C1(n10703), .C2(n10540), .A(n9051), .B(n9050), .ZN(n9052) );
  AOI21_X1 U10240 ( .B1(n9053), .B2(n11047), .A(n9052), .ZN(n9054) );
  OAI21_X1 U10241 ( .B1(n10722), .B2(n11050), .A(n9054), .ZN(n9055) );
  AOI21_X1 U10242 ( .B1(n10726), .B2(n10473), .A(n9055), .ZN(n9056) );
  OAI21_X1 U10243 ( .B1(n10728), .B2(n10603), .A(n9056), .ZN(P1_U3278) );
  XNOR2_X1 U10244 ( .A(n9058), .B(n9057), .ZN(n9059) );
  XNOR2_X1 U10245 ( .A(n9060), .B(n9059), .ZN(n9069) );
  NAND2_X1 U10246 ( .A1(n10233), .A2(n10248), .ZN(n9062) );
  OAI211_X1 U10247 ( .C1(n9063), .C2(n10236), .A(n9062), .B(n9061), .ZN(n9066)
         );
  NOR2_X1 U10248 ( .A1(n9064), .A2(n10237), .ZN(n9065) );
  AOI211_X1 U10249 ( .C1(n10241), .C2(n9067), .A(n9066), .B(n9065), .ZN(n9068)
         );
  OAI21_X1 U10250 ( .B1(n9069), .B2(n10243), .A(n9068), .ZN(P1_U3236) );
  INV_X1 U10251 ( .A(n9073), .ZN(n9071) );
  NAND2_X1 U10252 ( .A1(n9071), .A2(n9017), .ZN(n9076) );
  OAI22_X1 U10253 ( .A1(n9073), .A2(n9072), .B1(n10723), .B2(n10138), .ZN(
        n9074) );
  INV_X1 U10254 ( .A(n9074), .ZN(n9075) );
  OAI21_X2 U10255 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9079) );
  NAND2_X1 U10256 ( .A1(n9079), .A2(n9080), .ZN(n9154) );
  OAI21_X1 U10257 ( .B1(n9079), .B2(n9080), .A(n9154), .ZN(n10718) );
  XNOR2_X1 U10258 ( .A(n9081), .B(n9080), .ZN(n10716) );
  NAND2_X1 U10259 ( .A1(n10714), .A2(n9082), .ZN(n9156) );
  OAI211_X1 U10260 ( .C1(n10714), .C2(n9082), .A(n10542), .B(n9156), .ZN(
        n10713) );
  NAND2_X1 U10261 ( .A1(n10536), .A2(n10730), .ZN(n9084) );
  AOI22_X1 U10262 ( .A1(n10596), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10140), 
        .B2(n11044), .ZN(n9083) );
  OAI211_X1 U10263 ( .C1(n9219), .C2(n10540), .A(n9084), .B(n9083), .ZN(n9085)
         );
  AOI21_X1 U10264 ( .B1(n9086), .B2(n11047), .A(n9085), .ZN(n9087) );
  OAI21_X1 U10265 ( .B1(n10713), .B2(n11050), .A(n9087), .ZN(n9088) );
  AOI21_X1 U10266 ( .B1(n10716), .B2(n10473), .A(n9088), .ZN(n9089) );
  OAI21_X1 U10267 ( .B1(n10718), .B2(n10603), .A(n9089), .ZN(P1_U3277) );
  NOR2_X1 U10268 ( .A1(n5184), .A2(n5131), .ZN(n9091) );
  XNOR2_X1 U10269 ( .A(n9091), .B(n9090), .ZN(n9100) );
  NOR2_X1 U10270 ( .A1(n9092), .A2(n10237), .ZN(n9099) );
  INV_X1 U10271 ( .A(n9093), .ZN(n9094) );
  AOI21_X1 U10272 ( .B1(n10200), .B2(n10247), .A(n9094), .ZN(n9097) );
  NAND2_X1 U10273 ( .A1(n10241), .A2(n5681), .ZN(n9096) );
  NAND2_X1 U10274 ( .A1(n10233), .A2(n10249), .ZN(n9095) );
  NAND3_X1 U10275 ( .A1(n9097), .A2(n9096), .A3(n9095), .ZN(n9098) );
  AOI211_X1 U10276 ( .C1(n9100), .C2(n10223), .A(n9099), .B(n9098), .ZN(n9101)
         );
  INV_X1 U10277 ( .A(n9101), .ZN(P1_U3217) );
  AOI211_X1 U10278 ( .C1(n9104), .C2(n10025), .A(n9103), .B(n9102), .ZN(n11099) );
  NAND2_X1 U10279 ( .A1(n10023), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9105) );
  OAI21_X1 U10280 ( .B1(n11099), .B2(n10023), .A(n9105), .ZN(P2_U3472) );
  XNOR2_X1 U10281 ( .A(n9106), .B(n9377), .ZN(n9107) );
  OAI222_X1 U10282 ( .A1(n9956), .A2(n9953), .B1(n9954), .B2(n9139), .C1(n9951), .C2(n9107), .ZN(n9126) );
  OAI21_X1 U10283 ( .B1(n9109), .B2(n9289), .A(n9108), .ZN(n9129) );
  INV_X1 U10284 ( .A(n9138), .ZN(n9380) );
  OAI22_X1 U10285 ( .A1(n9129), .A2(n10017), .B1(n9380), .B2(n10027), .ZN(
        n9110) );
  NOR2_X1 U10286 ( .A1(n9126), .A2(n9110), .ZN(n11101) );
  OR2_X1 U10287 ( .A1(n10033), .A2(n6055), .ZN(n9111) );
  OAI21_X1 U10288 ( .B1(n11101), .B2(n10023), .A(n9111), .ZN(P2_U3473) );
  INV_X1 U10289 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9112) );
  OAI222_X1 U10290 ( .A1(P1_U3086), .A2(n6946), .B1(n10799), .B2(n9113), .C1(
        n9112), .C2(n10792), .ZN(P1_U3333) );
  INV_X1 U10291 ( .A(n9383), .ZN(n9291) );
  XNOR2_X1 U10292 ( .A(n9114), .B(n9291), .ZN(n9115) );
  NAND2_X1 U10293 ( .A1(n9115), .A2(n6325), .ZN(n9118) );
  OAI22_X1 U10294 ( .A1(n9197), .A2(n9954), .B1(n9568), .B2(n9956), .ZN(n9116)
         );
  INV_X1 U10295 ( .A(n9116), .ZN(n9117) );
  NAND2_X1 U10296 ( .A1(n9118), .A2(n9117), .ZN(n10031) );
  INV_X1 U10297 ( .A(n10031), .ZN(n9124) );
  XNOR2_X1 U10298 ( .A(n9119), .B(n9383), .ZN(n10026) );
  INV_X1 U10299 ( .A(n9120), .ZN(n9207) );
  AOI22_X1 U10300 ( .A1(n9946), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11066), 
        .B2(n9207), .ZN(n9121) );
  OAI21_X1 U10301 ( .B1(n10028), .B2(n9913), .A(n9121), .ZN(n9122) );
  AOI21_X1 U10302 ( .B1(n10026), .B2(n9943), .A(n9122), .ZN(n9123) );
  OAI21_X1 U10303 ( .B1(n9124), .B2(n9946), .A(n9123), .ZN(P2_U3218) );
  NOR2_X1 U10304 ( .A1(n9380), .A2(n9843), .ZN(n9125) );
  OAI21_X1 U10305 ( .B1(n9126), .B2(n9125), .A(n11069), .ZN(n9128) );
  AOI22_X1 U10306 ( .A1(n9946), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9150), .B2(
        n11066), .ZN(n9127) );
  OAI211_X1 U10307 ( .C1(n9129), .C2(n9963), .A(n9128), .B(n9127), .ZN(
        P2_U3219) );
  INV_X1 U10308 ( .A(n9134), .ZN(n9132) );
  AOI21_X1 U10309 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10796), .A(n9130), 
        .ZN(n9131) );
  OAI21_X1 U10310 ( .B1(n9132), .B2(n9234), .A(n9131), .ZN(P1_U3332) );
  NAND2_X1 U10311 ( .A1(n9134), .A2(n9133), .ZN(n9136) );
  NAND2_X1 U10312 ( .A1(n9135), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9467) );
  OAI211_X1 U10313 ( .C1(n9137), .C2(n10070), .A(n9136), .B(n9467), .ZN(
        P2_U3272) );
  XNOR2_X1 U10314 ( .A(n9138), .B(n9513), .ZN(n9196) );
  XNOR2_X1 U10315 ( .A(n9196), .B(n9197), .ZN(n9145) );
  NAND2_X1 U10316 ( .A1(n9140), .A2(n9139), .ZN(n9142) );
  INV_X1 U10317 ( .A(n9140), .ZN(n9141) );
  NAND2_X1 U10318 ( .A1(n9144), .A2(n9145), .ZN(n9201) );
  OAI21_X1 U10319 ( .B1(n9145), .B2(n9144), .A(n9201), .ZN(n9146) );
  NAND2_X1 U10320 ( .A1(n9146), .A2(n9600), .ZN(n9152) );
  NOR2_X1 U10321 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9147), .ZN(n9664) );
  AOI21_X1 U10322 ( .B1(n9624), .B2(n9642), .A(n9664), .ZN(n9148) );
  OAI21_X1 U10323 ( .B1(n9953), .B2(n9626), .A(n9148), .ZN(n9149) );
  AOI21_X1 U10324 ( .B1(n9606), .B2(n9150), .A(n9149), .ZN(n9151) );
  OAI211_X1 U10325 ( .C1(n9380), .C2(n9609), .A(n9152), .B(n9151), .ZN(
        P2_U3155) );
  OR2_X1 U10326 ( .A1(n10714), .A2(n10703), .ZN(n9153) );
  OAI21_X1 U10327 ( .B1(n9155), .B2(n9159), .A(n9220), .ZN(n10710) );
  NOR2_X2 U10328 ( .A1(n10706), .A2(n9156), .ZN(n9224) );
  AOI211_X1 U10329 ( .C1(n10706), .C2(n9156), .A(n10591), .B(n9224), .ZN(
        n10704) );
  NAND2_X1 U10330 ( .A1(n10706), .A2(n11047), .ZN(n9158) );
  AOI22_X1 U10331 ( .A1(n10596), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10152), 
        .B2(n11044), .ZN(n9157) );
  OAI211_X1 U10332 ( .C1(n10703), .C2(n10440), .A(n9158), .B(n9157), .ZN(n9163) );
  XNOR2_X1 U10333 ( .A(n9160), .B(n9159), .ZN(n9161) );
  AOI22_X1 U10334 ( .A1(n9161), .A2(n10725), .B1(n10731), .B2(n10587), .ZN(
        n10709) );
  NOR2_X1 U10335 ( .A1(n10709), .A2(n10596), .ZN(n9162) );
  AOI211_X1 U10336 ( .C1(n10704), .C2(n10594), .A(n9163), .B(n9162), .ZN(n9164) );
  OAI21_X1 U10337 ( .B1(n10710), .B2(n10603), .A(n9164), .ZN(P1_U3276) );
  XNOR2_X1 U10338 ( .A(n9652), .B(n9668), .ZN(n9167) );
  AOI21_X1 U10339 ( .B1(n6043), .B2(n9167), .A(n9653), .ZN(n9184) );
  MUX2_X1 U10340 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9756), .Z(n9659) );
  XNOR2_X1 U10341 ( .A(n9659), .B(n9668), .ZN(n9172) );
  OR2_X1 U10342 ( .A1(n9168), .A2(n9175), .ZN(n9170) );
  NAND2_X1 U10343 ( .A1(n9170), .A2(n9169), .ZN(n9171) );
  NAND2_X1 U10344 ( .A1(n9172), .A2(n9171), .ZN(n9660) );
  OAI21_X1 U10345 ( .B1(n9172), .B2(n9171), .A(n9660), .ZN(n9182) );
  XNOR2_X1 U10346 ( .A(n9668), .B(n9667), .ZN(n9176) );
  NOR2_X1 U10347 ( .A1(n6041), .A2(n9176), .ZN(n9669) );
  AOI21_X1 U10348 ( .B1(n9176), .B2(n6041), .A(n9669), .ZN(n9177) );
  NOR2_X1 U10349 ( .A1(n11008), .A2(n9177), .ZN(n9178) );
  AOI211_X1 U10350 ( .C1(n10999), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n9179), .B(
        n9178), .ZN(n9180) );
  OAI21_X1 U10351 ( .B1(n9658), .B2(n11000), .A(n9180), .ZN(n9181) );
  AOI21_X1 U10352 ( .B1(n10996), .B2(n9182), .A(n9181), .ZN(n9183) );
  OAI21_X1 U10353 ( .B1(n9184), .B2(n11011), .A(n9183), .ZN(P2_U3195) );
  OAI21_X1 U10354 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(n9188) );
  NAND2_X1 U10355 ( .A1(n9188), .A2(n10223), .ZN(n9195) );
  AOI21_X1 U10356 ( .B1(n10233), .B2(n10247), .A(n9189), .ZN(n9190) );
  OAI21_X1 U10357 ( .B1(n9191), .B2(n10236), .A(n9190), .ZN(n9192) );
  AOI21_X1 U10358 ( .B1(n9193), .B2(n10241), .A(n9192), .ZN(n9194) );
  OAI211_X1 U10359 ( .C1(n11089), .C2(n10237), .A(n9195), .B(n9194), .ZN(
        P1_U3224) );
  INV_X1 U10360 ( .A(n9196), .ZN(n9198) );
  NAND2_X1 U10361 ( .A1(n9198), .A2(n9197), .ZN(n9199) );
  AND2_X1 U10362 ( .A1(n9201), .A2(n9199), .ZN(n9203) );
  XNOR2_X1 U10363 ( .A(n10028), .B(n9513), .ZN(n9210) );
  XNOR2_X1 U10364 ( .A(n9210), .B(n9640), .ZN(n9202) );
  AND2_X1 U10365 ( .A1(n9202), .A2(n9199), .ZN(n9200) );
  OAI211_X1 U10366 ( .C1(n9203), .C2(n9202), .A(n9600), .B(n9212), .ZN(n9209)
         );
  INV_X1 U10367 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9204) );
  NOR2_X1 U10368 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9204), .ZN(n9691) );
  AOI21_X1 U10369 ( .B1(n9624), .B2(n9641), .A(n9691), .ZN(n9205) );
  OAI21_X1 U10370 ( .B1(n9568), .B2(n9626), .A(n9205), .ZN(n9206) );
  AOI21_X1 U10371 ( .B1(n9606), .B2(n9207), .A(n9206), .ZN(n9208) );
  OAI211_X1 U10372 ( .C1(n10028), .C2(n9609), .A(n9209), .B(n9208), .ZN(
        P2_U3181) );
  XNOR2_X1 U10373 ( .A(n10021), .B(n9513), .ZN(n9478) );
  XNOR2_X1 U10374 ( .A(n9478), .B(n9568), .ZN(n9476) );
  XNOR2_X1 U10375 ( .A(n9477), .B(n9476), .ZN(n9218) );
  OR2_X1 U10376 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9213), .ZN(n9708) );
  OAI21_X1 U10377 ( .B1(n9613), .B2(n9953), .A(n9708), .ZN(n9214) );
  AOI21_X1 U10378 ( .B1(n9615), .B2(n9918), .A(n9214), .ZN(n9215) );
  OAI21_X1 U10379 ( .B1(n9623), .B2(n9958), .A(n9215), .ZN(n9216) );
  AOI21_X1 U10380 ( .B1(n10021), .B2(n9629), .A(n9216), .ZN(n9217) );
  OAI21_X1 U10381 ( .B1(n9218), .B2(n9632), .A(n9217), .ZN(P2_U3166) );
  INV_X1 U10382 ( .A(n9219), .ZN(n10711) );
  OAI21_X1 U10383 ( .B1(n9221), .B2(n9222), .A(n10408), .ZN(n10701) );
  XNOR2_X1 U10384 ( .A(n9223), .B(n9222), .ZN(n10699) );
  INV_X1 U10385 ( .A(n10406), .ZN(n10697) );
  NAND2_X1 U10386 ( .A1(n10697), .A2(n9224), .ZN(n10592) );
  OAI211_X1 U10387 ( .C1(n10697), .C2(n9224), .A(n10542), .B(n10592), .ZN(
        n10696) );
  INV_X1 U10388 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9225) );
  OAI22_X1 U10389 ( .A1(n10601), .A2(n9225), .B1(n10213), .B2(n10435), .ZN(
        n9226) );
  AOI21_X1 U10390 ( .B1(n10536), .B2(n10711), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10391 ( .B1(n10209), .B2(n10540), .A(n9227), .ZN(n9228) );
  AOI21_X1 U10392 ( .B1(n10406), .B2(n11047), .A(n9228), .ZN(n9229) );
  OAI21_X1 U10393 ( .B1(n10696), .B2(n11050), .A(n9229), .ZN(n9230) );
  AOI21_X1 U10394 ( .B1(n10699), .B2(n10473), .A(n9230), .ZN(n9231) );
  OAI21_X1 U10395 ( .B1(n10701), .B2(n10603), .A(n9231), .ZN(P1_U3275) );
  INV_X1 U10396 ( .A(n9232), .ZN(n9237) );
  AOI22_X1 U10397 ( .A1(n6929), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10796), .ZN(n9233) );
  OAI21_X1 U10398 ( .B1(n9237), .B2(n9234), .A(n9233), .ZN(P1_U3331) );
  OAI222_X1 U10399 ( .A1(n10077), .A2(n9237), .B1(P2_U3151), .B2(n9236), .C1(
        n9235), .C2(n10086), .ZN(P2_U3271) );
  AND2_X1 U10400 ( .A1(n9238), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U10401 ( .A1(n9238), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U10402 ( .A1(n9238), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U10403 ( .A1(n9238), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U10404 ( .A1(n9238), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U10405 ( .A1(n9238), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U10406 ( .A1(n9238), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U10407 ( .A1(n9238), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U10408 ( .A1(n9238), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U10409 ( .A1(n9238), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U10410 ( .A1(n9238), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U10411 ( .A1(n9238), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U10412 ( .A1(n9238), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U10413 ( .A1(n9238), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U10414 ( .A1(n9238), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U10415 ( .A1(n9238), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U10416 ( .A1(n9238), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U10417 ( .A1(n9238), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U10418 ( .A1(n9238), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U10419 ( .A1(n9238), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U10420 ( .A1(n9238), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U10421 ( .A1(n9238), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U10422 ( .A1(n9238), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U10423 ( .A1(n9238), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U10424 ( .A1(n9238), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U10425 ( .A1(n9238), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U10426 ( .A1(n9238), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U10427 ( .A1(n9238), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U10428 ( .A1(n9238), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U10429 ( .A1(n9238), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  OAI222_X1 U10430 ( .A1(n10077), .A2(n9242), .B1(P2_U3151), .B2(n9240), .C1(
        n9239), .C2(n10086), .ZN(P2_U3270) );
  INV_X1 U10431 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9241) );
  OAI222_X1 U10432 ( .A1(P1_U3086), .A2(n9243), .B1(n10799), .B2(n9242), .C1(
        n9241), .C2(n10792), .ZN(P1_U3330) );
  NOR2_X1 U10433 ( .A1(n9267), .A2(n9470), .ZN(n9245) );
  AOI21_X2 U10434 ( .B1(n9244), .B2(n9266), .A(n9245), .ZN(n9277) );
  INV_X1 U10435 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9246) );
  OR2_X1 U10436 ( .A1(n9247), .A2(n9246), .ZN(n9254) );
  INV_X1 U10437 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9248) );
  OR2_X1 U10438 ( .A1(n9249), .A2(n9248), .ZN(n9253) );
  INV_X1 U10439 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9250) );
  OR2_X1 U10440 ( .A1(n9251), .A2(n9250), .ZN(n9252) );
  INV_X1 U10441 ( .A(n9256), .ZN(n9257) );
  NOR2_X1 U10442 ( .A1(n11105), .A2(n9262), .ZN(n10034) );
  AOI21_X1 U10443 ( .B1(n11105), .B2(P2_REG0_REG_30__SCAN_IN), .A(n10034), 
        .ZN(n9258) );
  OAI21_X1 U10444 ( .B1(n9277), .B2(n10063), .A(n9258), .ZN(P2_U3457) );
  NOR2_X1 U10445 ( .A1(n10023), .A2(n9262), .ZN(n9964) );
  AOI21_X1 U10446 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10023), .A(n9964), .ZN(
        n9259) );
  OAI21_X1 U10447 ( .B1(n9277), .B2(n10008), .A(n9259), .ZN(P2_U3489) );
  INV_X1 U10448 ( .A(n9260), .ZN(n9261) );
  NAND2_X1 U10449 ( .A1(n11066), .A2(n9261), .ZN(n9777) );
  NAND3_X1 U10450 ( .A1(n11071), .A2(n9777), .A3(n9262), .ZN(n9773) );
  OAI21_X1 U10451 ( .B1(n11069), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9773), .ZN(
        n9263) );
  OAI21_X1 U10452 ( .B1(n9277), .B2(n9913), .A(n9263), .ZN(P2_U3203) );
  INV_X1 U10453 ( .A(n9264), .ZN(n9276) );
  NAND2_X1 U10454 ( .A1(n10067), .A2(n9266), .ZN(n9269) );
  INV_X1 U10455 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10071) );
  OR2_X1 U10456 ( .A1(n9267), .A2(n10071), .ZN(n9268) );
  INV_X1 U10457 ( .A(n9277), .ZN(n9270) );
  NAND2_X1 U10458 ( .A1(n5683), .A2(n9270), .ZN(n9274) );
  OR2_X1 U10459 ( .A1(n9277), .A2(n9635), .ZN(n9450) );
  NAND2_X1 U10460 ( .A1(n9450), .A2(n9271), .ZN(n9455) );
  INV_X1 U10461 ( .A(n9304), .ZN(n9634) );
  NAND2_X1 U10462 ( .A1(n5683), .A2(n9634), .ZN(n9457) );
  INV_X1 U10463 ( .A(n9457), .ZN(n9272) );
  AND2_X1 U10464 ( .A1(n9277), .A2(n9635), .ZN(n9452) );
  INV_X1 U10465 ( .A(n9452), .ZN(n9299) );
  INV_X1 U10466 ( .A(n9455), .ZN(n9301) );
  INV_X1 U10467 ( .A(n9855), .ZN(n9295) );
  NAND4_X1 U10468 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n5426), .ZN(n9283)
         );
  NOR4_X1 U10469 ( .A1(n9283), .A2(n5167), .A3(n9282), .A4(n5289), .ZN(n9284)
         );
  NAND4_X1 U10470 ( .A1(n5458), .A2(n9348), .A3(n9285), .A4(n9284), .ZN(n9286)
         );
  NOR4_X1 U10471 ( .A1(n9370), .A2(n9288), .A3(n9287), .A4(n9286), .ZN(n9290)
         );
  NAND4_X1 U10472 ( .A1(n9291), .A2(n9290), .A3(n9372), .A4(n9289), .ZN(n9292)
         );
  NOR4_X1 U10473 ( .A1(n9927), .A2(n9390), .A3(n9950), .A4(n9292), .ZN(n9293)
         );
  XNOR2_X1 U10474 ( .A(n9910), .B(n9919), .ZN(n9908) );
  NAND4_X1 U10475 ( .A1(n9886), .A2(n9900), .A3(n9293), .A4(n9908), .ZN(n9294)
         );
  NOR4_X1 U10476 ( .A1(n9834), .A2(n9295), .A3(n9860), .A4(n9294), .ZN(n9297)
         );
  XNOR2_X1 U10477 ( .A(n9630), .B(n9831), .ZN(n9820) );
  INV_X1 U10478 ( .A(n9820), .ZN(n9296) );
  XNOR2_X1 U10479 ( .A(n9574), .B(n9850), .ZN(n9845) );
  NAND4_X1 U10480 ( .A1(n9800), .A2(n9297), .A3(n9296), .A4(n9845), .ZN(n9298)
         );
  NOR3_X1 U10481 ( .A1(n9451), .A2(n5276), .A3(n9298), .ZN(n9300) );
  NAND4_X1 U10482 ( .A1(n9457), .A2(n9301), .A3(n9300), .A4(n9299), .ZN(n9303)
         );
  NAND2_X1 U10483 ( .A1(n9305), .A2(n9304), .ZN(n9454) );
  INV_X1 U10484 ( .A(n9308), .ZN(n9391) );
  NOR2_X1 U10485 ( .A1(n9356), .A2(n9309), .ZN(n9310) );
  MUX2_X1 U10486 ( .A(n9310), .B(n9312), .S(n9449), .Z(n9316) );
  NAND2_X1 U10487 ( .A1(n9312), .A2(n9311), .ZN(n9314) );
  AOI211_X1 U10488 ( .C1(n9316), .C2(n9314), .A(n9359), .B(n9313), .ZN(n9349)
         );
  NAND2_X1 U10489 ( .A1(n9316), .A2(n9315), .ZN(n9352) );
  INV_X1 U10490 ( .A(n9322), .ZN(n9318) );
  INV_X1 U10491 ( .A(n9321), .ZN(n9317) );
  AOI21_X1 U10492 ( .B1(n9318), .B2(n9326), .A(n9317), .ZN(n9320) );
  OAI211_X1 U10493 ( .C1(n9320), .C2(n9325), .A(n9336), .B(n9319), .ZN(n9330)
         );
  OAI211_X1 U10494 ( .C1(n9324), .C2(n9323), .A(n9322), .B(n9321), .ZN(n9327)
         );
  NAND2_X1 U10495 ( .A1(n9332), .A2(n9331), .ZN(n9340) );
  OAI211_X1 U10496 ( .C1(n9340), .C2(n9334), .A(n9341), .B(n9333), .ZN(n9335)
         );
  NAND3_X1 U10497 ( .A1(n9335), .A2(n9338), .A3(n9345), .ZN(n9344) );
  INV_X1 U10498 ( .A(n9336), .ZN(n9339) );
  OAI211_X1 U10499 ( .C1(n9340), .C2(n9339), .A(n9338), .B(n9337), .ZN(n9342)
         );
  NAND3_X1 U10500 ( .A1(n9342), .A2(n9346), .A3(n9341), .ZN(n9343) );
  MUX2_X1 U10501 ( .A(n9346), .B(n9345), .S(n9449), .Z(n9347) );
  NOR2_X1 U10502 ( .A1(n9362), .A2(n9355), .ZN(n9351) );
  INV_X1 U10503 ( .A(n9361), .ZN(n9350) );
  AOI21_X1 U10504 ( .B1(n9358), .B2(n9351), .A(n9350), .ZN(n9365) );
  AOI21_X1 U10505 ( .B1(n9354), .B2(n9353), .A(n9352), .ZN(n9357) );
  NOR2_X1 U10506 ( .A1(n9360), .A2(n9359), .ZN(n9363) );
  OAI21_X1 U10507 ( .B1(n9363), .B2(n9362), .A(n9361), .ZN(n9364) );
  NOR2_X1 U10508 ( .A1(n9367), .A2(n9366), .ZN(n9369) );
  MUX2_X1 U10509 ( .A(n9369), .B(n9368), .S(n9449), .Z(n9371) );
  INV_X1 U10510 ( .A(n9375), .ZN(n9376) );
  MUX2_X1 U10511 ( .A(n6048), .B(n9376), .S(n9449), .Z(n9378) );
  NOR2_X1 U10512 ( .A1(n9380), .A2(n9641), .ZN(n9381) );
  MUX2_X1 U10513 ( .A(n9382), .B(n9381), .S(n9449), .Z(n9384) );
  INV_X1 U10514 ( .A(n9385), .ZN(n9387) );
  MUX2_X1 U10515 ( .A(n9387), .B(n9386), .S(n9449), .Z(n9388) );
  INV_X1 U10516 ( .A(n9392), .ZN(n9393) );
  INV_X1 U10517 ( .A(n9394), .ZN(n9397) );
  NOR2_X1 U10518 ( .A1(n9395), .A2(n9397), .ZN(n9404) );
  OAI22_X1 U10519 ( .A1(n9398), .A2(n9927), .B1(n9397), .B2(n9396), .ZN(n9402)
         );
  INV_X1 U10520 ( .A(n9399), .ZN(n9400) );
  AOI21_X1 U10521 ( .B1(n9402), .B2(n9401), .A(n9400), .ZN(n9403) );
  MUX2_X1 U10522 ( .A(n9404), .B(n9403), .S(n9449), .Z(n9406) );
  AOI22_X1 U10523 ( .A1(n9406), .A2(n9908), .B1(n5422), .B2(n9405), .ZN(n9410)
         );
  OAI21_X1 U10524 ( .B1(n9409), .B2(n9407), .A(n9449), .ZN(n9408) );
  OAI21_X1 U10525 ( .B1(n9410), .B2(n9409), .A(n9408), .ZN(n9411) );
  INV_X1 U10526 ( .A(n9413), .ZN(n9416) );
  INV_X1 U10527 ( .A(n9414), .ZN(n9415) );
  MUX2_X1 U10528 ( .A(n9416), .B(n9415), .S(n9449), .Z(n9417) );
  NOR2_X1 U10529 ( .A1(n9860), .A2(n9417), .ZN(n9421) );
  MUX2_X1 U10530 ( .A(n9419), .B(n9418), .S(n9449), .Z(n9420) );
  INV_X1 U10531 ( .A(n9987), .ZN(n9422) );
  NOR2_X1 U10532 ( .A1(n9422), .A2(n9639), .ZN(n9424) );
  MUX2_X1 U10533 ( .A(n9424), .B(n9423), .S(n9449), .Z(n9425) );
  MUX2_X1 U10534 ( .A(n9427), .B(n9426), .S(n5422), .Z(n9428) );
  INV_X1 U10535 ( .A(n9429), .ZN(n9431) );
  MUX2_X1 U10536 ( .A(n9431), .B(n9430), .S(n9449), .Z(n9432) );
  NOR3_X1 U10537 ( .A1(n9433), .A2(n9820), .A3(n9432), .ZN(n9440) );
  NAND3_X1 U10538 ( .A1(n5124), .A2(n5677), .A3(n9800), .ZN(n9439) );
  INV_X1 U10539 ( .A(n9434), .ZN(n9436) );
  MUX2_X1 U10540 ( .A(n9436), .B(n9435), .S(n9449), .Z(n9437) );
  INV_X1 U10541 ( .A(n9444), .ZN(n9447) );
  MUX2_X1 U10542 ( .A(n9805), .B(n9441), .S(n9449), .Z(n9443) );
  INV_X1 U10543 ( .A(n9443), .ZN(n9446) );
  MUX2_X1 U10544 ( .A(n9966), .B(n9636), .S(n9449), .Z(n9442) );
  AOI21_X1 U10545 ( .B1(n9444), .B2(n9443), .A(n9442), .ZN(n9445) );
  AOI21_X1 U10546 ( .B1(n9447), .B2(n9446), .A(n9445), .ZN(n9448) );
  XOR2_X1 U10547 ( .A(n9449), .B(n9448), .Z(n9456) );
  OAI21_X1 U10548 ( .B1(n9452), .B2(n9451), .A(n9450), .ZN(n9453) );
  XNOR2_X1 U10549 ( .A(n9461), .B(n9754), .ZN(n9468) );
  NAND3_X1 U10550 ( .A1(n9463), .A2(n9462), .A3(n9756), .ZN(n9464) );
  OAI211_X1 U10551 ( .C1(n9465), .C2(n9467), .A(n9464), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9466) );
  OAI21_X1 U10552 ( .B1(n9468), .B2(n9467), .A(n9466), .ZN(P2_U3296) );
  INV_X1 U10553 ( .A(n9244), .ZN(n9474) );
  OAI222_X1 U10554 ( .A1(n10070), .A2(n9470), .B1(n10087), .B2(n9474), .C1(
        P2_U3151), .C2(n5828), .ZN(P2_U3265) );
  INV_X1 U10555 ( .A(n9471), .ZN(n10080) );
  INV_X1 U10556 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9472) );
  OAI222_X1 U10557 ( .A1(P1_U3086), .A2(n10271), .B1(n10799), .B2(n10080), 
        .C1(n9472), .C2(n10792), .ZN(P1_U3327) );
  OAI222_X1 U10558 ( .A1(n10792), .A2(n9475), .B1(n10799), .B2(n9474), .C1(
        n9473), .C2(P1_U3086), .ZN(P1_U3325) );
  INV_X1 U10559 ( .A(n9478), .ZN(n9479) );
  XNOR2_X1 U10560 ( .A(n10013), .B(n9513), .ZN(n9564) );
  NAND2_X1 U10561 ( .A1(n9566), .A2(n9480), .ZN(n9482) );
  INV_X1 U10562 ( .A(n9564), .ZN(n9481) );
  NAND2_X1 U10563 ( .A1(n9482), .A2(n5682), .ZN(n9610) );
  XNOR2_X1 U10564 ( .A(n10009), .B(n9513), .ZN(n9483) );
  XNOR2_X1 U10565 ( .A(n9483), .B(n9906), .ZN(n9611) );
  NAND2_X1 U10566 ( .A1(n9610), .A2(n9611), .ZN(n9485) );
  NAND2_X1 U10567 ( .A1(n9483), .A2(n9937), .ZN(n9484) );
  NAND2_X1 U10568 ( .A1(n9485), .A2(n9484), .ZN(n9535) );
  XOR2_X1 U10569 ( .A(n9513), .B(n9908), .Z(n9536) );
  NAND2_X1 U10570 ( .A1(n9535), .A2(n9536), .ZN(n9487) );
  NAND2_X1 U10571 ( .A1(n9487), .A2(n9486), .ZN(n9589) );
  XNOR2_X1 U10572 ( .A(n10000), .B(n9510), .ZN(n9488) );
  NAND2_X1 U10573 ( .A1(n9488), .A2(n9907), .ZN(n9490) );
  OAI21_X1 U10574 ( .B1(n9488), .B2(n9907), .A(n9490), .ZN(n9590) );
  XNOR2_X1 U10575 ( .A(n9996), .B(n9513), .ZN(n9491) );
  XNOR2_X1 U10576 ( .A(n9491), .B(n9863), .ZN(n9545) );
  XNOR2_X1 U10577 ( .A(n9874), .B(n9513), .ZN(n9494) );
  XNOR2_X1 U10578 ( .A(n9494), .B(n9548), .ZN(n9601) );
  INV_X1 U10579 ( .A(n9491), .ZN(n9492) );
  NAND2_X1 U10580 ( .A1(n9492), .A2(n9863), .ZN(n9597) );
  NAND2_X1 U10581 ( .A1(n9598), .A2(n9493), .ZN(n9599) );
  NAND2_X1 U10582 ( .A1(n9494), .A2(n9881), .ZN(n9495) );
  NAND2_X1 U10583 ( .A1(n9599), .A2(n9495), .ZN(n9497) );
  XNOR2_X1 U10584 ( .A(n9987), .B(n9513), .ZN(n9496) );
  NAND2_X1 U10585 ( .A1(n9497), .A2(n9496), .ZN(n9498) );
  XNOR2_X1 U10586 ( .A(n9574), .B(n9510), .ZN(n9499) );
  NAND2_X1 U10587 ( .A1(n9499), .A2(n9830), .ZN(n9503) );
  INV_X1 U10588 ( .A(n9499), .ZN(n9500) );
  NAND2_X1 U10589 ( .A1(n9500), .A2(n9850), .ZN(n9501) );
  NAND2_X1 U10590 ( .A1(n9502), .A2(n9576), .ZN(n9578) );
  XNOR2_X1 U10591 ( .A(n9554), .B(n9513), .ZN(n9504) );
  XNOR2_X1 U10592 ( .A(n9504), .B(n9841), .ZN(n9557) );
  INV_X1 U10593 ( .A(n9504), .ZN(n9505) );
  NAND2_X1 U10594 ( .A1(n9505), .A2(n9841), .ZN(n9506) );
  XNOR2_X1 U10595 ( .A(n9630), .B(n9513), .ZN(n9508) );
  NAND2_X1 U10596 ( .A1(n9507), .A2(n5135), .ZN(n9509) );
  NAND2_X1 U10597 ( .A1(n9508), .A2(n9637), .ZN(n9620) );
  XNOR2_X1 U10598 ( .A(n6268), .B(n9510), .ZN(n9511) );
  NOR2_X1 U10599 ( .A1(n9511), .A2(n9819), .ZN(n9512) );
  AOI21_X1 U10600 ( .B1(n9511), .B2(n9819), .A(n9512), .ZN(n9522) );
  XNOR2_X1 U10601 ( .A(n5276), .B(n9513), .ZN(n9514) );
  NOR2_X1 U10602 ( .A1(n9623), .A2(n9792), .ZN(n9518) );
  AOI22_X1 U10603 ( .A1(n9624), .A2(n9786), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n9515) );
  OAI21_X1 U10604 ( .B1(n9516), .B2(n9626), .A(n9515), .ZN(n9517) );
  AOI211_X1 U10605 ( .C1(n9966), .C2(n9629), .A(n9518), .B(n9517), .ZN(n9519)
         );
  OAI21_X1 U10606 ( .B1(n9520), .B2(n9632), .A(n9519), .ZN(P2_U3160) );
  OAI211_X1 U10607 ( .C1(n9523), .C2(n9522), .A(n9521), .B(n9600), .ZN(n9528)
         );
  INV_X1 U10608 ( .A(n9809), .ZN(n9526) );
  AOI22_X1 U10609 ( .A1(n9624), .A2(n9637), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n9524) );
  OAI21_X1 U10610 ( .B1(n9805), .B2(n9626), .A(n9524), .ZN(n9525) );
  AOI21_X1 U10611 ( .B1(n9606), .B2(n9526), .A(n9525), .ZN(n9527) );
  OAI211_X1 U10612 ( .C1(n10040), .C2(n9609), .A(n9528), .B(n9527), .ZN(
        P2_U3154) );
  AOI21_X1 U10613 ( .B1(n9639), .B2(n9529), .A(n5134), .ZN(n9534) );
  AOI22_X1 U10614 ( .A1(n9615), .A2(n9850), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n9531) );
  NAND2_X1 U10615 ( .A1(n9624), .A2(n9881), .ZN(n9530) );
  OAI211_X1 U10616 ( .C1(n9623), .C2(n9852), .A(n9531), .B(n9530), .ZN(n9532)
         );
  AOI21_X1 U10617 ( .B1(n9987), .B2(n9629), .A(n9532), .ZN(n9533) );
  OAI21_X1 U10618 ( .B1(n9534), .B2(n9632), .A(n9533), .ZN(P2_U3156) );
  XNOR2_X1 U10619 ( .A(n9535), .B(n9536), .ZN(n9543) );
  NOR2_X1 U10620 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9537), .ZN(n9760) );
  NOR2_X1 U10621 ( .A1(n9613), .A2(n9906), .ZN(n9538) );
  AOI211_X1 U10622 ( .C1(n9615), .C2(n9880), .A(n9760), .B(n9538), .ZN(n9539)
         );
  OAI21_X1 U10623 ( .B1(n9540), .B2(n9623), .A(n9539), .ZN(n9541) );
  AOI21_X1 U10624 ( .B1(n9910), .B2(n9629), .A(n9541), .ZN(n9542) );
  OAI21_X1 U10625 ( .B1(n9543), .B2(n9632), .A(n9542), .ZN(P2_U3159) );
  INV_X1 U10626 ( .A(n9996), .ZN(n9553) );
  OAI21_X1 U10627 ( .B1(n9545), .B2(n9544), .A(n9598), .ZN(n9546) );
  NAND2_X1 U10628 ( .A1(n9546), .A2(n9600), .ZN(n9552) );
  OAI22_X1 U10629 ( .A1(n9626), .A2(n9548), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9547), .ZN(n9550) );
  NOR2_X1 U10630 ( .A1(n9623), .A2(n9883), .ZN(n9549) );
  AOI211_X1 U10631 ( .C1(n9624), .C2(n9880), .A(n9550), .B(n9549), .ZN(n9551)
         );
  OAI211_X1 U10632 ( .C1(n9553), .C2(n9609), .A(n9552), .B(n9551), .ZN(
        P2_U3163) );
  OAI21_X1 U10633 ( .B1(n9557), .B2(n9556), .A(n9555), .ZN(n9558) );
  NAND2_X1 U10634 ( .A1(n9558), .A2(n9600), .ZN(n9563) );
  OAI22_X1 U10635 ( .A1(n9626), .A2(n9831), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9559), .ZN(n9561) );
  NOR2_X1 U10636 ( .A1(n9623), .A2(n9832), .ZN(n9560) );
  AOI211_X1 U10637 ( .C1(n9624), .C2(n9850), .A(n9561), .B(n9560), .ZN(n9562)
         );
  OAI211_X1 U10638 ( .C1(n10048), .C2(n9609), .A(n9563), .B(n9562), .ZN(
        P2_U3165) );
  XNOR2_X1 U10639 ( .A(n9564), .B(n9955), .ZN(n9565) );
  XNOR2_X1 U10640 ( .A(n9566), .B(n9565), .ZN(n9573) );
  INV_X1 U10641 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9567) );
  NOR2_X1 U10642 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9567), .ZN(n9732) );
  NOR2_X1 U10643 ( .A1(n9613), .A2(n9568), .ZN(n9569) );
  AOI211_X1 U10644 ( .C1(n9615), .C2(n9937), .A(n9732), .B(n9569), .ZN(n9570)
         );
  OAI21_X1 U10645 ( .B1(n9939), .B2(n9623), .A(n9570), .ZN(n9571) );
  AOI21_X1 U10646 ( .B1(n10013), .B2(n9629), .A(n9571), .ZN(n9572) );
  OAI21_X1 U10647 ( .B1(n9573), .B2(n9632), .A(n9572), .ZN(P2_U3168) );
  INV_X1 U10648 ( .A(n9575), .ZN(n9577) );
  NOR3_X1 U10649 ( .A1(n5134), .A2(n9577), .A3(n9576), .ZN(n9580) );
  INV_X1 U10650 ( .A(n9578), .ZN(n9579) );
  OAI21_X1 U10651 ( .B1(n9580), .B2(n9579), .A(n9600), .ZN(n9586) );
  NOR2_X1 U10652 ( .A1(n9613), .A2(n9862), .ZN(n9583) );
  OAI22_X1 U10653 ( .A1(n9626), .A2(n9841), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9581), .ZN(n9582) );
  AOI211_X1 U10654 ( .C1(n9606), .C2(n9584), .A(n9583), .B(n9582), .ZN(n9585)
         );
  OAI211_X1 U10655 ( .C1(n10052), .C2(n9609), .A(n9586), .B(n9585), .ZN(
        P2_U3169) );
  INV_X1 U10656 ( .A(n9587), .ZN(n9588) );
  AOI21_X1 U10657 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9596) );
  OAI22_X1 U10658 ( .A1(n9626), .A2(n9863), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9591), .ZN(n9592) );
  AOI21_X1 U10659 ( .B1(n9624), .B2(n9919), .A(n9592), .ZN(n9593) );
  OAI21_X1 U10660 ( .B1(n9623), .B2(n9895), .A(n9593), .ZN(n9594) );
  AOI21_X1 U10661 ( .B1(n10000), .B2(n9629), .A(n9594), .ZN(n9595) );
  OAI21_X1 U10662 ( .B1(n9596), .B2(n9632), .A(n9595), .ZN(P2_U3173) );
  AND2_X1 U10663 ( .A1(n9598), .A2(n9597), .ZN(n9602) );
  OAI211_X1 U10664 ( .C1(n9602), .C2(n9601), .A(n9600), .B(n9599), .ZN(n9608)
         );
  INV_X1 U10665 ( .A(n9866), .ZN(n9605) );
  AOI22_X1 U10666 ( .A1(n9624), .A2(n9893), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9603) );
  OAI21_X1 U10667 ( .B1(n9862), .B2(n9626), .A(n9603), .ZN(n9604) );
  AOI21_X1 U10668 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9607) );
  OAI211_X1 U10669 ( .C1(n10057), .C2(n9609), .A(n9608), .B(n9607), .ZN(
        P2_U3175) );
  XNOR2_X1 U10670 ( .A(n9610), .B(n9611), .ZN(n9619) );
  INV_X1 U10671 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9612) );
  NOR2_X1 U10672 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9612), .ZN(n10998) );
  NOR2_X1 U10673 ( .A1(n9613), .A2(n9955), .ZN(n9614) );
  AOI211_X1 U10674 ( .C1(n9615), .C2(n9919), .A(n10998), .B(n9614), .ZN(n9616)
         );
  OAI21_X1 U10675 ( .B1(n9921), .B2(n9623), .A(n9616), .ZN(n9617) );
  AOI21_X1 U10676 ( .B1(n10009), .B2(n9629), .A(n9617), .ZN(n9618) );
  OAI21_X1 U10677 ( .B1(n9619), .B2(n9632), .A(n9618), .ZN(P2_U3178) );
  NAND2_X1 U10678 ( .A1(n5135), .A2(n9620), .ZN(n9621) );
  XNOR2_X1 U10679 ( .A(n9622), .B(n9621), .ZN(n9633) );
  NOR2_X1 U10680 ( .A1(n9623), .A2(n9822), .ZN(n9628) );
  AOI22_X1 U10681 ( .A1(n9624), .A2(n9638), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9625) );
  OAI21_X1 U10682 ( .B1(n9819), .B2(n9626), .A(n9625), .ZN(n9627) );
  AOI211_X1 U10683 ( .C1(n9630), .C2(n9629), .A(n9628), .B(n9627), .ZN(n9631)
         );
  OAI21_X1 U10684 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(P2_U3180) );
  MUX2_X1 U10685 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9634), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10686 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9635), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10687 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9787), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10688 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9636), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10689 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9786), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10690 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9637), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10691 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9638), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10692 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9850), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10693 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9639), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10694 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9881), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10695 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9893), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10696 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9880), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10697 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9919), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10698 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9937), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10699 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9918), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10700 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9935), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10701 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9640), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10702 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9641), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10703 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9642), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10704 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8994), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10705 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9643), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10706 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9644), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10707 ( .A(n9645), .B(P2_DATAO_REG_9__SCAN_IN), .S(n11001), .Z(
        P2_U3500) );
  MUX2_X1 U10708 ( .A(n9646), .B(P2_DATAO_REG_8__SCAN_IN), .S(n11001), .Z(
        P2_U3499) );
  MUX2_X1 U10709 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n9647), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10710 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9648), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10711 ( .A(n9649), .B(P2_DATAO_REG_5__SCAN_IN), .S(n11001), .Z(
        P2_U3496) );
  MUX2_X1 U10712 ( .A(n9650), .B(P2_DATAO_REG_3__SCAN_IN), .S(n11001), .Z(
        P2_U3494) );
  MUX2_X1 U10713 ( .A(n6273), .B(P2_DATAO_REG_2__SCAN_IN), .S(n11001), .Z(
        P2_U3493) );
  MUX2_X1 U10714 ( .A(n6271), .B(P2_DATAO_REG_1__SCAN_IN), .S(n11001), .Z(
        P2_U3492) );
  MUX2_X1 U10715 ( .A(n9651), .B(P2_DATAO_REG_0__SCAN_IN), .S(n11001), .Z(
        P2_U3491) );
  NOR2_X1 U10716 ( .A1(n9668), .A2(n9652), .ZN(n9654) );
  NAND2_X1 U10717 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9689), .ZN(n9655) );
  OAI21_X1 U10718 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9689), .A(n9655), .ZN(
        n9656) );
  AOI21_X1 U10719 ( .B1(n5182), .B2(n9656), .A(n9681), .ZN(n9679) );
  MUX2_X1 U10720 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9756), .Z(n9683) );
  XNOR2_X1 U10721 ( .A(n9683), .B(n9657), .ZN(n9663) );
  OR2_X1 U10722 ( .A1(n9659), .A2(n9658), .ZN(n9661) );
  NAND2_X1 U10723 ( .A1(n9661), .A2(n9660), .ZN(n9662) );
  NAND2_X1 U10724 ( .A1(n9663), .A2(n9662), .ZN(n9684) );
  OAI21_X1 U10725 ( .B1(n9663), .B2(n9662), .A(n9684), .ZN(n9677) );
  NAND2_X1 U10726 ( .A1(n10999), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n9666) );
  INV_X1 U10727 ( .A(n9664), .ZN(n9665) );
  OAI211_X1 U10728 ( .C1(n11000), .C2(n9689), .A(n9666), .B(n9665), .ZN(n9676)
         );
  NOR2_X1 U10729 ( .A1(n9668), .A2(n9667), .ZN(n9670) );
  NAND2_X1 U10730 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9689), .ZN(n9671) );
  OAI21_X1 U10731 ( .B1(n9689), .B2(P2_REG2_REG_14__SCAN_IN), .A(n9671), .ZN(
        n9672) );
  AOI21_X1 U10732 ( .B1(n9673), .B2(n9672), .A(n9688), .ZN(n9674) );
  NOR2_X1 U10733 ( .A1(n9674), .A2(n11008), .ZN(n9675) );
  AOI211_X1 U10734 ( .C1(n10996), .C2(n9677), .A(n9676), .B(n9675), .ZN(n9678)
         );
  OAI21_X1 U10735 ( .B1(n9679), .B2(n11011), .A(n9678), .ZN(P2_U3196) );
  AND2_X1 U10736 ( .A1(n9689), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9680) );
  AOI21_X1 U10737 ( .B1(n6071), .B2(n9682), .A(n9700), .ZN(n9698) );
  MUX2_X1 U10738 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9756), .Z(n9703) );
  XNOR2_X1 U10739 ( .A(n9703), .B(n9711), .ZN(n9687) );
  OR2_X1 U10740 ( .A1(n9683), .A2(n9689), .ZN(n9685) );
  NAND2_X1 U10741 ( .A1(n9685), .A2(n9684), .ZN(n9686) );
  NAND2_X1 U10742 ( .A1(n9687), .A2(n9686), .ZN(n9704) );
  OAI21_X1 U10743 ( .B1(n9687), .B2(n9686), .A(n9704), .ZN(n9696) );
  NOR2_X1 U10744 ( .A1(n6073), .A2(n9690), .ZN(n9712) );
  AOI21_X1 U10745 ( .B1(n9690), .B2(n6073), .A(n9712), .ZN(n9694) );
  NAND2_X1 U10746 ( .A1(n10976), .A2(n9711), .ZN(n9693) );
  AOI21_X1 U10747 ( .B1(n10999), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n9691), .ZN(
        n9692) );
  OAI211_X1 U10748 ( .C1(n9694), .C2(n11008), .A(n9693), .B(n9692), .ZN(n9695)
         );
  AOI21_X1 U10749 ( .B1(n10996), .B2(n9696), .A(n9695), .ZN(n9697) );
  OAI21_X1 U10750 ( .B1(n9698), .B2(n11011), .A(n9697), .ZN(P2_U3197) );
  NOR2_X1 U10751 ( .A1(n9711), .A2(n9699), .ZN(n9701) );
  AOI22_X1 U10752 ( .A1(n9714), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n6088), .B2(
        n9736), .ZN(n9702) );
  AOI21_X1 U10753 ( .B1(n5177), .B2(n9702), .A(n9724), .ZN(n9723) );
  MUX2_X1 U10754 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9756), .Z(n9727) );
  XNOR2_X1 U10755 ( .A(n9714), .B(n9727), .ZN(n9707) );
  OR2_X1 U10756 ( .A1(n9703), .A2(n5213), .ZN(n9705) );
  NAND2_X1 U10757 ( .A1(n9705), .A2(n9704), .ZN(n9706) );
  NAND2_X1 U10758 ( .A1(n9707), .A2(n9706), .ZN(n9728) );
  OAI21_X1 U10759 ( .B1(n9707), .B2(n9706), .A(n9728), .ZN(n9721) );
  NAND2_X1 U10760 ( .A1(n10999), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9709) );
  OAI211_X1 U10761 ( .C1(n11000), .C2(n9736), .A(n9709), .B(n9708), .ZN(n9720)
         );
  NOR2_X1 U10762 ( .A1(n9711), .A2(n9710), .ZN(n9713) );
  MUX2_X1 U10763 ( .A(n9959), .B(P2_REG2_REG_16__SCAN_IN), .S(n9714), .Z(n9715) );
  INV_X1 U10764 ( .A(n9715), .ZN(n9716) );
  AOI21_X1 U10765 ( .B1(n9717), .B2(n9716), .A(n9735), .ZN(n9718) );
  NOR2_X1 U10766 ( .A1(n9718), .A2(n11008), .ZN(n9719) );
  AOI211_X1 U10767 ( .C1(n10996), .C2(n9721), .A(n9720), .B(n9719), .ZN(n9722)
         );
  OAI21_X1 U10768 ( .B1(n9723), .B2(n11011), .A(n9722), .ZN(P2_U3198) );
  AOI21_X1 U10769 ( .B1(n9726), .B2(n9725), .A(n9745), .ZN(n9743) );
  MUX2_X1 U10770 ( .A(n9940), .B(n9726), .S(n9756), .Z(n9751) );
  XNOR2_X1 U10771 ( .A(n9734), .B(n9751), .ZN(n9731) );
  OR2_X1 U10772 ( .A1(n9727), .A2(n9736), .ZN(n9729) );
  NAND2_X1 U10773 ( .A1(n9729), .A2(n9728), .ZN(n9730) );
  NAND2_X1 U10774 ( .A1(n9731), .A2(n9730), .ZN(n9749) );
  OAI21_X1 U10775 ( .B1(n9731), .B2(n9730), .A(n9749), .ZN(n9741) );
  AOI21_X1 U10776 ( .B1(n10999), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n9732), .ZN(
        n9733) );
  OAI21_X1 U10777 ( .B1(n9734), .B2(n11000), .A(n9733), .ZN(n9740) );
  AOI21_X1 U10778 ( .B1(n9737), .B2(n9940), .A(n9765), .ZN(n9738) );
  NOR2_X1 U10779 ( .A1(n9738), .A2(n11008), .ZN(n9739) );
  AOI211_X1 U10780 ( .C1(n10996), .C2(n9741), .A(n9740), .B(n9739), .ZN(n9742)
         );
  OAI21_X1 U10781 ( .B1(n9743), .B2(n11011), .A(n9742), .ZN(P2_U3199) );
  NOR2_X1 U10782 ( .A1(n9764), .A2(n9744), .ZN(n9746) );
  NAND2_X1 U10783 ( .A1(n10995), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9747) );
  OAI21_X1 U10784 ( .B1(n10995), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9747), .ZN(
        n11010) );
  XNOR2_X1 U10785 ( .A(n9754), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9755) );
  XNOR2_X1 U10786 ( .A(n9748), .B(n9755), .ZN(n9772) );
  INV_X1 U10787 ( .A(n9749), .ZN(n9750) );
  AOI21_X1 U10788 ( .B1(n9764), .B2(n9751), .A(n9750), .ZN(n9753) );
  MUX2_X1 U10789 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n9756), .Z(n9752) );
  NOR2_X1 U10790 ( .A1(n9753), .A2(n9752), .ZN(n10992) );
  NAND2_X1 U10791 ( .A1(n9753), .A2(n9752), .ZN(n10993) );
  OAI21_X1 U10792 ( .B1(n10992), .B2(n11003), .A(n10993), .ZN(n9759) );
  MUX2_X1 U10793 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n6132), .S(n9754), .Z(n9769) );
  INV_X1 U10794 ( .A(n9755), .ZN(n9757) );
  MUX2_X1 U10795 ( .A(n9769), .B(n9757), .S(n9756), .Z(n9758) );
  XNOR2_X1 U10796 ( .A(n9759), .B(n9758), .ZN(n9771) );
  AOI21_X1 U10797 ( .B1(n10999), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9760), .ZN(
        n9761) );
  OAI21_X1 U10798 ( .B1(n9762), .B2(n11000), .A(n9761), .ZN(n9770) );
  NOR2_X1 U10799 ( .A1(n9764), .A2(n9763), .ZN(n9766) );
  NOR2_X1 U10800 ( .A1(n9766), .A2(n9765), .ZN(n11007) );
  NAND2_X1 U10801 ( .A1(n10995), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9767) );
  OAI21_X1 U10802 ( .B1(n10995), .B2(P2_REG2_REG_18__SCAN_IN), .A(n9767), .ZN(
        n11006) );
  INV_X1 U10803 ( .A(n9767), .ZN(n9768) );
  OAI21_X1 U10804 ( .B1(n11069), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9773), .ZN(
        n9774) );
  OAI21_X1 U10805 ( .B1(n5683), .B2(n9913), .A(n9774), .ZN(P2_U3202) );
  INV_X1 U10806 ( .A(n9775), .ZN(n9784) );
  NAND2_X1 U10807 ( .A1(n9776), .A2(n11069), .ZN(n9782) );
  OAI21_X1 U10808 ( .B1(n11069), .B2(n9778), .A(n9777), .ZN(n9779) );
  AOI21_X1 U10809 ( .B1(n9780), .B2(n11064), .A(n9779), .ZN(n9781) );
  OAI211_X1 U10810 ( .C1(n9784), .C2(n9783), .A(n9782), .B(n9781), .ZN(
        P2_U3204) );
  XNOR2_X1 U10811 ( .A(n9785), .B(n5276), .ZN(n9791) );
  NAND2_X1 U10812 ( .A1(n9786), .A2(n9934), .ZN(n9789) );
  OAI22_X1 U10813 ( .A1(n11069), .A2(n9793), .B1(n9792), .B2(n9957), .ZN(n9794) );
  AOI21_X1 U10814 ( .B1(n9966), .B2(n11064), .A(n9794), .ZN(n9799) );
  OAI21_X1 U10815 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(n9967) );
  NAND2_X1 U10816 ( .A1(n9967), .A2(n9943), .ZN(n9798) );
  OAI211_X1 U10817 ( .C1(n9968), .C2(n9946), .A(n9799), .B(n9798), .ZN(
        P2_U3205) );
  NAND2_X1 U10818 ( .A1(n9801), .A2(n9800), .ZN(n9802) );
  NAND2_X1 U10819 ( .A1(n9802), .A2(n6325), .ZN(n9804) );
  OR2_X1 U10820 ( .A1(n9804), .A2(n9803), .ZN(n9808) );
  OAI22_X1 U10821 ( .A1(n9831), .A2(n9954), .B1(n9805), .B2(n9956), .ZN(n9806)
         );
  INV_X1 U10822 ( .A(n9806), .ZN(n9807) );
  NAND2_X1 U10823 ( .A1(n9808), .A2(n9807), .ZN(n9972) );
  INV_X1 U10824 ( .A(n9972), .ZN(n9816) );
  OAI22_X1 U10825 ( .A1(n11069), .A2(n9810), .B1(n9809), .B2(n9957), .ZN(n9811) );
  AOI21_X1 U10826 ( .B1(n6268), .B2(n11064), .A(n9811), .ZN(n9815) );
  XNOR2_X1 U10827 ( .A(n9813), .B(n9812), .ZN(n9970) );
  NAND2_X1 U10828 ( .A1(n9970), .A2(n9943), .ZN(n9814) );
  OAI211_X1 U10829 ( .C1(n9816), .C2(n9946), .A(n9815), .B(n9814), .ZN(
        P2_U3206) );
  XNOR2_X1 U10830 ( .A(n9817), .B(n9820), .ZN(n9818) );
  OAI222_X1 U10831 ( .A1(n9954), .A2(n9841), .B1(n9956), .B2(n9819), .C1(n9951), .C2(n9818), .ZN(n9975) );
  INV_X1 U10832 ( .A(n9975), .ZN(n9827) );
  XNOR2_X1 U10833 ( .A(n9821), .B(n9820), .ZN(n9976) );
  NOR2_X1 U10834 ( .A1(n10044), .A2(n9913), .ZN(n9825) );
  OAI22_X1 U10835 ( .A1(n11071), .A2(n9823), .B1(n9822), .B2(n9957), .ZN(n9824) );
  AOI211_X1 U10836 ( .C1(n9976), .C2(n9943), .A(n9825), .B(n9824), .ZN(n9826)
         );
  OAI21_X1 U10837 ( .B1(n9827), .B2(n9946), .A(n9826), .ZN(P2_U3207) );
  XNOR2_X1 U10838 ( .A(n9828), .B(n9834), .ZN(n9829) );
  OAI222_X1 U10839 ( .A1(n9956), .A2(n9831), .B1(n9954), .B2(n9830), .C1(n9829), .C2(n9951), .ZN(n9979) );
  OAI22_X1 U10840 ( .A1(n10048), .A2(n9843), .B1(n9832), .B2(n9957), .ZN(n9833) );
  OAI21_X1 U10841 ( .B1(n9979), .B2(n9833), .A(n11071), .ZN(n9837) );
  XNOR2_X1 U10842 ( .A(n9835), .B(n9834), .ZN(n9980) );
  NAND2_X1 U10843 ( .A1(n9980), .A2(n9943), .ZN(n9836) );
  OAI211_X1 U10844 ( .C1(n11069), .C2(n9838), .A(n9837), .B(n9836), .ZN(
        P2_U3208) );
  XNOR2_X1 U10845 ( .A(n9839), .B(n9845), .ZN(n9840) );
  OAI222_X1 U10846 ( .A1(n9954), .A2(n9862), .B1(n9956), .B2(n9841), .C1(n9840), .C2(n9951), .ZN(n9983) );
  OAI22_X1 U10847 ( .A1(n10052), .A2(n9843), .B1(n9842), .B2(n9957), .ZN(n9844) );
  OAI21_X1 U10848 ( .B1(n9983), .B2(n9844), .A(n11069), .ZN(n9848) );
  XOR2_X1 U10849 ( .A(n9846), .B(n9845), .Z(n9984) );
  AOI22_X1 U10850 ( .A1(n9984), .A2(n9943), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9946), .ZN(n9847) );
  NAND2_X1 U10851 ( .A1(n9848), .A2(n9847), .ZN(P2_U3209) );
  XNOR2_X1 U10852 ( .A(n9849), .B(n9855), .ZN(n9851) );
  AOI222_X1 U10853 ( .A1(n6325), .A2(n9851), .B1(n9850), .B2(n9936), .C1(n9881), .C2(n9934), .ZN(n9989) );
  OAI22_X1 U10854 ( .A1(n11071), .A2(n9853), .B1(n9852), .B2(n9957), .ZN(n9858) );
  OAI21_X1 U10855 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(n9990) );
  NOR2_X1 U10856 ( .A1(n9990), .A2(n9963), .ZN(n9857) );
  AOI211_X1 U10857 ( .C1(n11064), .C2(n9987), .A(n9858), .B(n9857), .ZN(n9859)
         );
  OAI21_X1 U10858 ( .B1(n9989), .B2(n9946), .A(n9859), .ZN(P2_U3210) );
  XNOR2_X1 U10859 ( .A(n9861), .B(n9860), .ZN(n9865) );
  OAI22_X1 U10860 ( .A1(n9863), .A2(n9954), .B1(n9862), .B2(n9956), .ZN(n9864)
         );
  AOI21_X1 U10861 ( .B1(n9865), .B2(n6325), .A(n9864), .ZN(n9993) );
  OAI22_X1 U10862 ( .A1(n11071), .A2(n9867), .B1(n9866), .B2(n9957), .ZN(n9873) );
  OR2_X1 U10863 ( .A1(n9869), .A2(n9868), .ZN(n9870) );
  NAND2_X1 U10864 ( .A1(n9871), .A2(n9870), .ZN(n9991) );
  NOR2_X1 U10865 ( .A1(n9991), .A2(n9963), .ZN(n9872) );
  AOI211_X1 U10866 ( .C1(n11064), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9875)
         );
  OAI21_X1 U10867 ( .B1(n9946), .B2(n9993), .A(n9875), .ZN(P2_U3211) );
  NAND2_X1 U10868 ( .A1(n9877), .A2(n9876), .ZN(n9879) );
  INV_X1 U10869 ( .A(n9886), .ZN(n9878) );
  XNOR2_X1 U10870 ( .A(n9879), .B(n9878), .ZN(n9882) );
  AOI222_X1 U10871 ( .A1(n6325), .A2(n9882), .B1(n9881), .B2(n9936), .C1(n9880), .C2(n9934), .ZN(n9998) );
  OAI22_X1 U10872 ( .A1(n11071), .A2(n9884), .B1(n9883), .B2(n9957), .ZN(n9889) );
  OAI21_X1 U10873 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(n9999) );
  NOR2_X1 U10874 ( .A1(n9999), .A2(n9963), .ZN(n9888) );
  AOI211_X1 U10875 ( .C1(n11064), .C2(n9996), .A(n9889), .B(n9888), .ZN(n9890)
         );
  OAI21_X1 U10876 ( .B1(n9998), .B2(n9946), .A(n9890), .ZN(P2_U3212) );
  XNOR2_X1 U10877 ( .A(n9892), .B(n9891), .ZN(n9894) );
  AOI222_X1 U10878 ( .A1(n6325), .A2(n9894), .B1(n9919), .B2(n9934), .C1(n9893), .C2(n9936), .ZN(n10003) );
  OAI22_X1 U10879 ( .A1(n11071), .A2(n9896), .B1(n9895), .B2(n9957), .ZN(n9897) );
  AOI21_X1 U10880 ( .B1(n10000), .B2(n11064), .A(n9897), .ZN(n9903) );
  NAND2_X1 U10881 ( .A1(n9899), .A2(n9898), .ZN(n9901) );
  XNOR2_X1 U10882 ( .A(n9901), .B(n9900), .ZN(n10001) );
  NAND2_X1 U10883 ( .A1(n10001), .A2(n9943), .ZN(n9902) );
  OAI211_X1 U10884 ( .C1(n10003), .C2(n9946), .A(n9903), .B(n9902), .ZN(
        P2_U3213) );
  XOR2_X1 U10885 ( .A(n9908), .B(n9904), .Z(n9905) );
  OAI222_X1 U10886 ( .A1(n9956), .A2(n9907), .B1(n9954), .B2(n9906), .C1(n9951), .C2(n9905), .ZN(n10004) );
  INV_X1 U10887 ( .A(n10004), .ZN(n9916) );
  XOR2_X1 U10888 ( .A(n9909), .B(n9908), .Z(n10005) );
  INV_X1 U10889 ( .A(n9910), .ZN(n10064) );
  AOI22_X1 U10890 ( .A1(n9946), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n11066), 
        .B2(n9911), .ZN(n9912) );
  OAI21_X1 U10891 ( .B1(n10064), .B2(n9913), .A(n9912), .ZN(n9914) );
  AOI21_X1 U10892 ( .B1(n10005), .B2(n9943), .A(n9914), .ZN(n9915) );
  OAI21_X1 U10893 ( .B1(n9916), .B2(n9946), .A(n9915), .ZN(P2_U3214) );
  XOR2_X1 U10894 ( .A(n9917), .B(n9927), .Z(n9920) );
  AOI222_X1 U10895 ( .A1(n6325), .A2(n9920), .B1(n9919), .B2(n9936), .C1(n9918), .C2(n9934), .ZN(n10012) );
  OAI22_X1 U10896 ( .A1(n11071), .A2(n9922), .B1(n9921), .B2(n9957), .ZN(n9923) );
  AOI21_X1 U10897 ( .B1(n10009), .B2(n11064), .A(n9923), .ZN(n9929) );
  INV_X1 U10898 ( .A(n9925), .ZN(n9926) );
  AOI21_X1 U10899 ( .B1(n9927), .B2(n9924), .A(n9926), .ZN(n10010) );
  NAND2_X1 U10900 ( .A1(n10010), .A2(n9943), .ZN(n9928) );
  OAI211_X1 U10901 ( .C1(n10012), .C2(n9946), .A(n9929), .B(n9928), .ZN(
        P2_U3215) );
  NAND2_X1 U10902 ( .A1(n9930), .A2(n9950), .ZN(n9932) );
  NAND2_X1 U10903 ( .A1(n9932), .A2(n9931), .ZN(n9933) );
  XNOR2_X1 U10904 ( .A(n9933), .B(n5432), .ZN(n9938) );
  AOI222_X1 U10905 ( .A1(n6325), .A2(n9938), .B1(n9937), .B2(n9936), .C1(n9935), .C2(n9934), .ZN(n10016) );
  OAI22_X1 U10906 ( .A1(n11071), .A2(n9940), .B1(n9939), .B2(n9957), .ZN(n9941) );
  AOI21_X1 U10907 ( .B1(n10013), .B2(n11064), .A(n9941), .ZN(n9945) );
  XNOR2_X1 U10908 ( .A(n9942), .B(n5432), .ZN(n10014) );
  NAND2_X1 U10909 ( .A1(n10014), .A2(n9943), .ZN(n9944) );
  OAI211_X1 U10910 ( .C1(n10016), .C2(n9946), .A(n9945), .B(n9944), .ZN(
        P2_U3216) );
  NAND2_X1 U10911 ( .A1(n9948), .A2(n9947), .ZN(n9949) );
  XOR2_X1 U10912 ( .A(n9950), .B(n9949), .Z(n10018) );
  XNOR2_X1 U10913 ( .A(n9930), .B(n9950), .ZN(n9952) );
  OAI222_X1 U10914 ( .A1(n9956), .A2(n9955), .B1(n9954), .B2(n9953), .C1(n9952), .C2(n9951), .ZN(n10019) );
  NAND2_X1 U10915 ( .A1(n10019), .A2(n11069), .ZN(n9962) );
  OAI22_X1 U10916 ( .A1(n11071), .A2(n9959), .B1(n9958), .B2(n9957), .ZN(n9960) );
  AOI21_X1 U10917 ( .B1(n10021), .B2(n11064), .A(n9960), .ZN(n9961) );
  OAI211_X1 U10918 ( .C1(n10018), .C2(n9963), .A(n9962), .B(n9961), .ZN(
        P2_U3217) );
  AOI21_X1 U10919 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10023), .A(n9964), .ZN(
        n9965) );
  OAI21_X1 U10920 ( .B1(n5683), .B2(n10008), .A(n9965), .ZN(P2_U3490) );
  AOI22_X1 U10921 ( .A1(n9967), .A2(n10025), .B1(n10022), .B2(n9966), .ZN(
        n9969) );
  MUX2_X1 U10922 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n10036), .S(n10033), .Z(
        P2_U3487) );
  INV_X1 U10923 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9973) );
  AND2_X1 U10924 ( .A1(n9970), .A2(n10025), .ZN(n9971) );
  NOR2_X1 U10925 ( .A1(n9972), .A2(n9971), .ZN(n10038) );
  MUX2_X1 U10926 ( .A(n9973), .B(n10038), .S(n10033), .Z(n9974) );
  OAI21_X1 U10927 ( .B1(n10040), .B2(n10008), .A(n9974), .ZN(P2_U3486) );
  AOI21_X1 U10928 ( .B1(n9976), .B2(n10025), .A(n9975), .ZN(n10041) );
  MUX2_X1 U10929 ( .A(n9977), .B(n10041), .S(n10033), .Z(n9978) );
  OAI21_X1 U10930 ( .B1(n10044), .B2(n10008), .A(n9978), .ZN(P2_U3485) );
  INV_X1 U10931 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9981) );
  AOI21_X1 U10932 ( .B1(n10025), .B2(n9980), .A(n9979), .ZN(n10045) );
  MUX2_X1 U10933 ( .A(n9981), .B(n10045), .S(n10033), .Z(n9982) );
  OAI21_X1 U10934 ( .B1(n10048), .B2(n10008), .A(n9982), .ZN(P2_U3484) );
  INV_X1 U10935 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9985) );
  AOI21_X1 U10936 ( .B1(n9984), .B2(n10025), .A(n9983), .ZN(n10049) );
  MUX2_X1 U10937 ( .A(n9985), .B(n10049), .S(n10033), .Z(n9986) );
  OAI21_X1 U10938 ( .B1(n10052), .B2(n10008), .A(n9986), .ZN(P2_U3483) );
  NAND2_X1 U10939 ( .A1(n9987), .A2(n10022), .ZN(n9988) );
  OAI211_X1 U10940 ( .C1(n10017), .C2(n9990), .A(n9989), .B(n9988), .ZN(n10053) );
  MUX2_X1 U10941 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n10053), .S(n10033), .Z(
        P2_U3482) );
  INV_X1 U10942 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9994) );
  OR2_X1 U10943 ( .A1(n9991), .A2(n10017), .ZN(n9992) );
  AND2_X1 U10944 ( .A1(n9993), .A2(n9992), .ZN(n10054) );
  MUX2_X1 U10945 ( .A(n9994), .B(n10054), .S(n10033), .Z(n9995) );
  OAI21_X1 U10946 ( .B1(n10057), .B2(n10008), .A(n9995), .ZN(P2_U3481) );
  NAND2_X1 U10947 ( .A1(n9996), .A2(n10022), .ZN(n9997) );
  OAI211_X1 U10948 ( .C1(n10017), .C2(n9999), .A(n9998), .B(n9997), .ZN(n10058) );
  MUX2_X1 U10949 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n10058), .S(n10033), .Z(
        P2_U3480) );
  AOI22_X1 U10950 ( .A1(n10001), .A2(n10025), .B1(n10022), .B2(n10000), .ZN(
        n10002) );
  NAND2_X1 U10951 ( .A1(n10003), .A2(n10002), .ZN(n10059) );
  MUX2_X1 U10952 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n10059), .S(n10033), .Z(
        P2_U3479) );
  AOI21_X1 U10953 ( .B1(n10005), .B2(n10025), .A(n10004), .ZN(n10060) );
  MUX2_X1 U10954 ( .A(n10006), .B(n10060), .S(n10033), .Z(n10007) );
  OAI21_X1 U10955 ( .B1(n10064), .B2(n10008), .A(n10007), .ZN(P2_U3478) );
  AOI22_X1 U10956 ( .A1(n10010), .A2(n10025), .B1(n10022), .B2(n10009), .ZN(
        n10011) );
  NAND2_X1 U10957 ( .A1(n10012), .A2(n10011), .ZN(n10065) );
  MUX2_X1 U10958 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n10065), .S(n10033), .Z(
        P2_U3477) );
  AOI22_X1 U10959 ( .A1(n10014), .A2(n10025), .B1(n10022), .B2(n10013), .ZN(
        n10015) );
  NAND2_X1 U10960 ( .A1(n10016), .A2(n10015), .ZN(n10066) );
  MUX2_X1 U10961 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n10066), .S(n10033), .Z(
        P2_U3476) );
  NOR2_X1 U10962 ( .A1(n10018), .A2(n10017), .ZN(n10020) );
  AOI211_X1 U10963 ( .C1(n10022), .C2(n10021), .A(n10020), .B(n10019), .ZN(
        n11107) );
  OR2_X1 U10964 ( .A1(n11107), .A2(n10023), .ZN(n10024) );
  OAI21_X1 U10965 ( .B1(n10033), .B2(n6088), .A(n10024), .ZN(P2_U3475) );
  AND2_X1 U10966 ( .A1(n10026), .A2(n10025), .ZN(n10030) );
  NOR2_X1 U10967 ( .A1(n10028), .A2(n10027), .ZN(n10029) );
  NAND2_X1 U10968 ( .A1(n11102), .A2(n10033), .ZN(n10032) );
  OAI21_X1 U10969 ( .B1(n10033), .B2(n6071), .A(n10032), .ZN(P2_U3474) );
  AOI21_X1 U10970 ( .B1(n11105), .B2(P2_REG0_REG_31__SCAN_IN), .A(n10034), 
        .ZN(n10035) );
  OAI21_X1 U10971 ( .B1(n5683), .B2(n10063), .A(n10035), .ZN(P2_U3458) );
  MUX2_X1 U10972 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n10036), .S(n11108), .Z(
        P2_U3455) );
  MUX2_X1 U10973 ( .A(n10038), .B(n10037), .S(n11105), .Z(n10039) );
  OAI21_X1 U10974 ( .B1(n10040), .B2(n10063), .A(n10039), .ZN(P2_U3454) );
  INV_X1 U10975 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10042) );
  MUX2_X1 U10976 ( .A(n10042), .B(n10041), .S(n11108), .Z(n10043) );
  OAI21_X1 U10977 ( .B1(n10044), .B2(n10063), .A(n10043), .ZN(P2_U3453) );
  MUX2_X1 U10978 ( .A(n10046), .B(n10045), .S(n11108), .Z(n10047) );
  OAI21_X1 U10979 ( .B1(n10048), .B2(n10063), .A(n10047), .ZN(P2_U3452) );
  MUX2_X1 U10980 ( .A(n10050), .B(n10049), .S(n11108), .Z(n10051) );
  OAI21_X1 U10981 ( .B1(n10052), .B2(n10063), .A(n10051), .ZN(P2_U3451) );
  MUX2_X1 U10982 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n10053), .S(n11108), .Z(
        P2_U3450) );
  MUX2_X1 U10983 ( .A(n10055), .B(n10054), .S(n11108), .Z(n10056) );
  OAI21_X1 U10984 ( .B1(n10057), .B2(n10063), .A(n10056), .ZN(P2_U3449) );
  MUX2_X1 U10985 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n10058), .S(n11108), .Z(
        P2_U3448) );
  MUX2_X1 U10986 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n10059), .S(n11108), .Z(
        P2_U3447) );
  INV_X1 U10987 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U10988 ( .A(n10061), .B(n10060), .S(n11108), .Z(n10062) );
  OAI21_X1 U10989 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(P2_U3446) );
  MUX2_X1 U10990 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n10065), .S(n11108), .Z(
        P2_U3444) );
  MUX2_X1 U10991 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n10066), .S(n11108), .Z(
        P2_U3441) );
  INV_X1 U10992 ( .A(n10067), .ZN(n10788) );
  NAND3_X1 U10993 ( .A1(n10069), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n10072) );
  OAI22_X1 U10994 ( .A1(n10068), .A2(n10072), .B1(n10071), .B2(n10070), .ZN(
        n10073) );
  INV_X1 U10995 ( .A(n10073), .ZN(n10074) );
  OAI21_X1 U10996 ( .B1(n10788), .B2(n10087), .A(n10074), .ZN(P2_U3264) );
  INV_X1 U10997 ( .A(n10075), .ZN(n10790) );
  OAI222_X1 U10998 ( .A1(n10077), .A2(n10790), .B1(n5826), .B2(P2_U3151), .C1(
        n10076), .C2(n10086), .ZN(P2_U3266) );
  AOI21_X1 U10999 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n10083), .A(n10078), 
        .ZN(n10079) );
  OAI21_X1 U11000 ( .B1(n10080), .B2(n10087), .A(n10079), .ZN(P2_U3267) );
  INV_X1 U11001 ( .A(n10081), .ZN(n10794) );
  AOI21_X1 U11002 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n10083), .A(n10082), 
        .ZN(n10084) );
  OAI21_X1 U11003 ( .B1(n10794), .B2(n10087), .A(n10084), .ZN(P2_U3268) );
  INV_X1 U11004 ( .A(n10085), .ZN(n10800) );
  OAI222_X1 U11005 ( .A1(P2_U3151), .A2(n10088), .B1(n10087), .B2(n10800), 
        .C1(n10086), .C2(n6219), .ZN(P2_U3269) );
  INV_X1 U11006 ( .A(n10089), .ZN(n10090) );
  MUX2_X1 U11007 ( .A(n10090), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U11008 ( .A1(n5181), .A2(n10091), .ZN(n10093) );
  XNOR2_X1 U11009 ( .A(n10093), .B(n10092), .ZN(n10100) );
  NAND2_X1 U11010 ( .A1(n10233), .A2(n10733), .ZN(n10095) );
  OAI211_X1 U11011 ( .C1(n10138), .C2(n10236), .A(n10095), .B(n10094), .ZN(
        n10096) );
  AOI21_X1 U11012 ( .B1(n10097), .B2(n10241), .A(n10096), .ZN(n10099) );
  NAND2_X1 U11013 ( .A1(n10729), .A2(n10215), .ZN(n10098) );
  OAI211_X1 U11014 ( .C1(n10100), .C2(n10243), .A(n10099), .B(n10098), .ZN(
        P1_U3215) );
  OAI21_X1 U11015 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(n10104) );
  NAND2_X1 U11016 ( .A1(n10104), .A2(n10223), .ZN(n10108) );
  AOI22_X1 U11017 ( .A1(n10200), .A2(n10659), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10105) );
  OAI21_X1 U11018 ( .B1(n10559), .B2(n10169), .A(n10105), .ZN(n10106) );
  AOI21_X1 U11019 ( .B1(n10522), .B2(n10241), .A(n10106), .ZN(n10107) );
  OAI211_X1 U11020 ( .C1(n10764), .C2(n10237), .A(n10108), .B(n10107), .ZN(
        P1_U3216) );
  XOR2_X1 U11021 ( .A(n10109), .B(n10110), .Z(n10116) );
  NAND2_X1 U11022 ( .A1(n10233), .A2(n10587), .ZN(n10112) );
  OAI211_X1 U11023 ( .C1(n10558), .C2(n10236), .A(n10112), .B(n10111), .ZN(
        n10113) );
  AOI21_X1 U11024 ( .B1(n10595), .B2(n10241), .A(n10113), .ZN(n10115) );
  NAND2_X1 U11025 ( .A1(n10593), .A2(n10215), .ZN(n10114) );
  OAI211_X1 U11026 ( .C1(n10116), .C2(n10243), .A(n10115), .B(n10114), .ZN(
        P1_U3219) );
  AOI21_X1 U11027 ( .B1(n10117), .B2(n10118), .A(n10243), .ZN(n10120) );
  NAND2_X1 U11028 ( .A1(n10120), .A2(n10119), .ZN(n10124) );
  AOI22_X1 U11029 ( .A1(n10233), .A2(n10586), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10121) );
  OAI21_X1 U11030 ( .B1(n10559), .B2(n10236), .A(n10121), .ZN(n10122) );
  AOI21_X1 U11031 ( .B1(n10562), .B2(n10241), .A(n10122), .ZN(n10123) );
  OAI211_X1 U11032 ( .C1(n10772), .C2(n10237), .A(n10124), .B(n10123), .ZN(
        P1_U3223) );
  OAI21_X1 U11033 ( .B1(n10126), .B2(n10125), .A(n10218), .ZN(n10127) );
  NAND2_X1 U11034 ( .A1(n10127), .A2(n10223), .ZN(n10131) );
  AOI22_X1 U11035 ( .A1(n10200), .A2(n10464), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10128) );
  OAI21_X1 U11036 ( .B1(n10644), .B2(n10169), .A(n10128), .ZN(n10129) );
  AOI21_X1 U11037 ( .B1(n10497), .B2(n10241), .A(n10129), .ZN(n10130) );
  OAI211_X1 U11038 ( .C1(n10496), .C2(n10237), .A(n10131), .B(n10130), .ZN(
        P1_U3225) );
  OAI21_X1 U11039 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10135) );
  NAND2_X1 U11040 ( .A1(n10135), .A2(n10223), .ZN(n10142) );
  AOI21_X1 U11041 ( .B1(n10200), .B2(n10711), .A(n10136), .ZN(n10137) );
  OAI21_X1 U11042 ( .B1(n10138), .B2(n10169), .A(n10137), .ZN(n10139) );
  AOI21_X1 U11043 ( .B1(n10140), .B2(n10241), .A(n10139), .ZN(n10141) );
  OAI211_X1 U11044 ( .C1(n10714), .C2(n10237), .A(n10142), .B(n10141), .ZN(
        P1_U3226) );
  NAND2_X1 U11045 ( .A1(n10132), .A2(n10143), .ZN(n10147) );
  NAND2_X1 U11046 ( .A1(n10145), .A2(n10144), .ZN(n10146) );
  XNOR2_X1 U11047 ( .A(n10147), .B(n10146), .ZN(n10155) );
  NAND2_X1 U11048 ( .A1(n10233), .A2(n10719), .ZN(n10149) );
  OAI211_X1 U11049 ( .C1(n10150), .C2(n10236), .A(n10149), .B(n10148), .ZN(
        n10151) );
  AOI21_X1 U11050 ( .B1(n10152), .B2(n10241), .A(n10151), .ZN(n10154) );
  NAND2_X1 U11051 ( .A1(n10706), .A2(n10215), .ZN(n10153) );
  OAI211_X1 U11052 ( .C1(n10155), .C2(n10243), .A(n10154), .B(n10153), .ZN(
        P1_U3228) );
  NAND2_X1 U11053 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  XNOR2_X1 U11054 ( .A(n10159), .B(n10158), .ZN(n10164) );
  AOI22_X1 U11055 ( .A1(n10200), .A2(n10480), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10161) );
  NAND2_X1 U11056 ( .A1(n10241), .A2(n10508), .ZN(n10160) );
  OAI211_X1 U11057 ( .C1(n10668), .C2(n10169), .A(n10161), .B(n10160), .ZN(
        n10162) );
  AOI21_X1 U11058 ( .B1(n10654), .B2(n10215), .A(n10162), .ZN(n10163) );
  OAI21_X1 U11059 ( .B1(n10164), .B2(n10243), .A(n10163), .ZN(P1_U3229) );
  XOR2_X1 U11060 ( .A(n10165), .B(n10166), .Z(n10172) );
  AOI22_X1 U11061 ( .A1(n10200), .A2(n10577), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10168) );
  NAND2_X1 U11062 ( .A1(n10241), .A2(n10572), .ZN(n10167) );
  OAI211_X1 U11063 ( .C1(n10209), .C2(n10169), .A(n10168), .B(n10167), .ZN(
        n10170) );
  AOI21_X1 U11064 ( .B1(n10684), .B2(n10215), .A(n10170), .ZN(n10171) );
  OAI21_X1 U11065 ( .B1(n10172), .B2(n10243), .A(n10171), .ZN(P1_U3233) );
  AOI21_X1 U11066 ( .B1(n9185), .B2(n10175), .A(n10174), .ZN(n10176) );
  NAND2_X1 U11067 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10365)
         );
  INV_X1 U11068 ( .A(n10365), .ZN(n10177) );
  AOI21_X1 U11069 ( .B1(n10233), .B2(n10246), .A(n10177), .ZN(n10178) );
  OAI21_X1 U11070 ( .B1(n10179), .B2(n10236), .A(n10178), .ZN(n10180) );
  AOI21_X1 U11071 ( .B1(n10181), .B2(n10241), .A(n10180), .ZN(n10182) );
  OAI211_X1 U11072 ( .C1(n10184), .C2(n10237), .A(n10183), .B(n10182), .ZN(
        P1_U3234) );
  NAND2_X1 U11073 ( .A1(n10186), .A2(n10185), .ZN(n10187) );
  XOR2_X1 U11074 ( .A(n10188), .B(n10187), .Z(n10193) );
  AOI22_X1 U11075 ( .A1(n10233), .A2(n10577), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10190) );
  NAND2_X1 U11076 ( .A1(n10241), .A2(n10537), .ZN(n10189) );
  OAI211_X1 U11077 ( .C1(n10668), .C2(n10236), .A(n10190), .B(n10189), .ZN(
        n10191) );
  AOI21_X1 U11078 ( .B1(n10545), .B2(n10215), .A(n10191), .ZN(n10192) );
  OAI21_X1 U11079 ( .B1(n10193), .B2(n10243), .A(n10192), .ZN(P1_U3235) );
  OAI21_X1 U11080 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10197) );
  NAND2_X1 U11081 ( .A1(n10197), .A2(n10223), .ZN(n10203) );
  AOI22_X1 U11082 ( .A1(n10233), .A2(n5111), .B1(n10198), .B2(n10215), .ZN(
        n10202) );
  AOI22_X1 U11083 ( .A1(n10200), .A2(n10255), .B1(n10199), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10201) );
  NAND3_X1 U11084 ( .A1(n10203), .A2(n10202), .A3(n10201), .ZN(P1_U3237) );
  NAND2_X1 U11085 ( .A1(n10205), .A2(n10204), .ZN(n10207) );
  XNOR2_X1 U11086 ( .A(n10207), .B(n10206), .ZN(n10217) );
  OAI21_X1 U11087 ( .B1(n10236), .B2(n10209), .A(n10208), .ZN(n10210) );
  AOI21_X1 U11088 ( .B1(n10233), .B2(n10711), .A(n10210), .ZN(n10211) );
  OAI21_X1 U11089 ( .B1(n10213), .B2(n10212), .A(n10211), .ZN(n10214) );
  AOI21_X1 U11090 ( .B1(n10406), .B2(n10215), .A(n10214), .ZN(n10216) );
  OAI21_X1 U11091 ( .B1(n10217), .B2(n10243), .A(n10216), .ZN(P1_U3238) );
  INV_X1 U11092 ( .A(n10218), .ZN(n10221) );
  NAND3_X1 U11093 ( .A1(n10224), .A2(n10223), .A3(n10222), .ZN(n10228) );
  AOI22_X1 U11094 ( .A1(n10233), .A2(n10480), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10225) );
  OAI21_X1 U11095 ( .B1(n10633), .B2(n10236), .A(n10225), .ZN(n10226) );
  AOI21_X1 U11096 ( .B1(n10481), .B2(n10241), .A(n10226), .ZN(n10227) );
  OAI211_X1 U11097 ( .C1(n10758), .C2(n10237), .A(n10228), .B(n10227), .ZN(
        P1_U3240) );
  NAND2_X1 U11098 ( .A1(n10229), .A2(n10230), .ZN(n10232) );
  XNOR2_X1 U11099 ( .A(n10232), .B(n10231), .ZN(n10244) );
  NAND2_X1 U11100 ( .A1(n10233), .A2(n10720), .ZN(n10235) );
  OAI211_X1 U11101 ( .C1(n10703), .C2(n10236), .A(n10235), .B(n10234), .ZN(
        n10239) );
  NOR2_X1 U11102 ( .A1(n10723), .A2(n10237), .ZN(n10238) );
  AOI211_X1 U11103 ( .C1(n10241), .C2(n10240), .A(n10239), .B(n10238), .ZN(
        n10242) );
  OAI21_X1 U11104 ( .B1(n10244), .B2(n10243), .A(n10242), .ZN(P1_U3241) );
  MUX2_X1 U11105 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n10383), .S(P1_U3973), .Z(
        P1_U3585) );
  INV_X1 U11106 ( .A(n10245), .ZN(n10433) );
  MUX2_X1 U11107 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10433), .S(P1_U3973), .Z(
        P1_U3584) );
  INV_X1 U11108 ( .A(n10626), .ZN(n10427) );
  MUX2_X1 U11109 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10427), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U11110 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10425), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U11111 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10480), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U11112 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10659), .S(P1_U3973), .Z(
        P1_U3578) );
  INV_X1 U11113 ( .A(n10668), .ZN(n10416) );
  MUX2_X1 U11114 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10416), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U11115 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10658), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11116 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10577), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U11117 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10586), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U11118 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10694), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U11119 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10587), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U11120 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10711), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U11121 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10719), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U11122 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10730), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U11123 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n10720), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U11124 ( .A(n10733), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10278), .Z(
        P1_U3567) );
  MUX2_X1 U11125 ( .A(n10246), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10278), .Z(
        P1_U3566) );
  MUX2_X1 U11126 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10247), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U11127 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n10248), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U11128 ( .A(n10249), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10278), .Z(
        P1_U3563) );
  MUX2_X1 U11129 ( .A(n10250), .B(P1_DATAO_REG_8__SCAN_IN), .S(n10278), .Z(
        P1_U3562) );
  MUX2_X1 U11130 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n10251), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U11131 ( .A(n10252), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10278), .Z(
        P1_U3560) );
  MUX2_X1 U11132 ( .A(n10253), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10278), .Z(
        P1_U3559) );
  MUX2_X1 U11133 ( .A(n10254), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10278), .Z(
        P1_U3558) );
  MUX2_X1 U11134 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10255), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U11135 ( .A(n10256), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10278), .Z(
        P1_U3556) );
  MUX2_X1 U11136 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5111), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U11137 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10258), .S(P1_U3973), .Z(
        P1_U3554) );
  AND2_X1 U11138 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10260) );
  OAI211_X1 U11139 ( .C1(n10261), .C2(n10260), .A(n10354), .B(n10259), .ZN(
        n10270) );
  OAI211_X1 U11140 ( .C1(n10264), .C2(n10263), .A(n10372), .B(n10262), .ZN(
        n10269) );
  AOI22_X1 U11141 ( .A1(n10265), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10268) );
  NAND2_X1 U11142 ( .A1(n10369), .A2(n10266), .ZN(n10267) );
  NAND4_X1 U11143 ( .A1(n10270), .A2(n10269), .A3(n10268), .A4(n10267), .ZN(
        P1_U3244) );
  NOR3_X1 U11144 ( .A1(n10273), .A2(n10272), .A3(n10271), .ZN(n10279) );
  OAI22_X1 U11145 ( .A1(n10276), .A2(P1_IR_REG_0__SCAN_IN), .B1(n10275), .B2(
        n10274), .ZN(n10277) );
  OR3_X1 U11146 ( .A1(n10279), .A2(n10278), .A3(n10277), .ZN(n10319) );
  INV_X1 U11147 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10281) );
  INV_X1 U11148 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10280) );
  OAI22_X1 U11149 ( .A1(n10367), .A2(n10281), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10280), .ZN(n10282) );
  AOI21_X1 U11150 ( .B1(n10283), .B2(n10369), .A(n10282), .ZN(n10292) );
  OAI211_X1 U11151 ( .C1(n10286), .C2(n10285), .A(n10372), .B(n10284), .ZN(
        n10291) );
  OAI211_X1 U11152 ( .C1(n10289), .C2(n10288), .A(n10354), .B(n10287), .ZN(
        n10290) );
  NAND4_X1 U11153 ( .A1(n10319), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        P1_U3245) );
  INV_X1 U11154 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10294) );
  OAI21_X1 U11155 ( .B1(n10367), .B2(n10294), .A(n10293), .ZN(n10295) );
  AOI21_X1 U11156 ( .B1(n10296), .B2(n10369), .A(n10295), .ZN(n10305) );
  OAI211_X1 U11157 ( .C1(n10299), .C2(n10298), .A(n10372), .B(n10297), .ZN(
        n10304) );
  OAI211_X1 U11158 ( .C1(n10302), .C2(n10301), .A(n10354), .B(n10300), .ZN(
        n10303) );
  NAND3_X1 U11159 ( .A1(n10305), .A2(n10304), .A3(n10303), .ZN(P1_U3246) );
  INV_X1 U11160 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10307) );
  OAI21_X1 U11161 ( .B1(n10367), .B2(n10307), .A(n10306), .ZN(n10308) );
  AOI21_X1 U11162 ( .B1(n10309), .B2(n10369), .A(n10308), .ZN(n10318) );
  OAI211_X1 U11163 ( .C1(n10312), .C2(n10311), .A(n10354), .B(n10310), .ZN(
        n10317) );
  OAI211_X1 U11164 ( .C1(n10315), .C2(n10314), .A(n10372), .B(n10313), .ZN(
        n10316) );
  NAND4_X1 U11165 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        P1_U3247) );
  INV_X1 U11166 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10321) );
  OAI21_X1 U11167 ( .B1(n10367), .B2(n10321), .A(n10320), .ZN(n10322) );
  AOI21_X1 U11168 ( .B1(n10323), .B2(n10369), .A(n10322), .ZN(n10332) );
  OAI211_X1 U11169 ( .C1(n10326), .C2(n10325), .A(n10372), .B(n10324), .ZN(
        n10331) );
  OAI211_X1 U11170 ( .C1(n10329), .C2(n10328), .A(n10354), .B(n10327), .ZN(
        n10330) );
  NAND3_X1 U11171 ( .A1(n10332), .A2(n10331), .A3(n10330), .ZN(P1_U3248) );
  INV_X1 U11172 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10334) );
  OAI21_X1 U11173 ( .B1(n10367), .B2(n10334), .A(n10333), .ZN(n10335) );
  AOI21_X1 U11174 ( .B1(n10336), .B2(n10369), .A(n10335), .ZN(n10345) );
  OAI211_X1 U11175 ( .C1(n10339), .C2(n10338), .A(n10372), .B(n10337), .ZN(
        n10344) );
  OAI211_X1 U11176 ( .C1(n10342), .C2(n10341), .A(n10354), .B(n10340), .ZN(
        n10343) );
  NAND3_X1 U11177 ( .A1(n10345), .A2(n10344), .A3(n10343), .ZN(P1_U3249) );
  INV_X1 U11178 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10347) );
  OAI21_X1 U11179 ( .B1(n10367), .B2(n10347), .A(n10346), .ZN(n10348) );
  AOI21_X1 U11180 ( .B1(n10349), .B2(n10369), .A(n10348), .ZN(n10359) );
  OAI211_X1 U11181 ( .C1(n10352), .C2(n10351), .A(n10372), .B(n10350), .ZN(
        n10358) );
  OAI211_X1 U11182 ( .C1(n10356), .C2(n10355), .A(n10354), .B(n10353), .ZN(
        n10357) );
  NAND3_X1 U11183 ( .A1(n10359), .A2(n10358), .A3(n10357), .ZN(P1_U3250) );
  AOI211_X1 U11184 ( .C1(n10363), .C2(n10362), .A(n10361), .B(n10360), .ZN(
        n10364) );
  INV_X1 U11185 ( .A(n10364), .ZN(n10377) );
  INV_X1 U11186 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10366) );
  OAI21_X1 U11187 ( .B1(n10367), .B2(n10366), .A(n10365), .ZN(n10368) );
  AOI21_X1 U11188 ( .B1(n10370), .B2(n10369), .A(n10368), .ZN(n10376) );
  OAI211_X1 U11189 ( .C1(n10374), .C2(n10373), .A(n10372), .B(n10371), .ZN(
        n10375) );
  NAND3_X1 U11190 ( .A1(n10377), .A2(n10376), .A3(n10375), .ZN(P1_U3256) );
  NOR2_X2 U11191 ( .A1(n10592), .A2(n10593), .ZN(n10569) );
  NAND2_X1 U11192 ( .A1(n10510), .A2(n10505), .ZN(n10506) );
  NAND2_X1 U11193 ( .A1(n10747), .A2(n10431), .ZN(n10386) );
  XNOR2_X1 U11194 ( .A(n10386), .B(n10379), .ZN(n10380) );
  NOR2_X2 U11195 ( .A1(n10380), .A2(n10591), .ZN(n10606) );
  NAND2_X1 U11196 ( .A1(n10606), .A2(n10594), .ZN(n10385) );
  INV_X1 U11197 ( .A(P1_B_REG_SCAN_IN), .ZN(n10381) );
  NOR2_X1 U11198 ( .A1(n10795), .A2(n10381), .ZN(n10382) );
  NOR2_X1 U11199 ( .A1(n10667), .A2(n10382), .ZN(n10432) );
  AND2_X1 U11200 ( .A1(n10383), .A2(n10432), .ZN(n10605) );
  INV_X1 U11201 ( .A(n10605), .ZN(n10609) );
  NOR2_X1 U11202 ( .A1(n10596), .A2(n10609), .ZN(n10388) );
  AOI21_X1 U11203 ( .B1(n10596), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10388), 
        .ZN(n10384) );
  OAI211_X1 U11204 ( .C1(n10743), .C2(n10599), .A(n10385), .B(n10384), .ZN(
        P1_U3263) );
  OAI211_X1 U11205 ( .C1(n10747), .C2(n10431), .A(n10542), .B(n10386), .ZN(
        n10610) );
  NOR2_X1 U11206 ( .A1(n10747), .A2(n10599), .ZN(n10387) );
  AOI211_X1 U11207 ( .C1(n10596), .C2(P1_REG2_REG_30__SCAN_IN), .A(n10388), 
        .B(n10387), .ZN(n10389) );
  OAI21_X1 U11208 ( .B1(n10610), .B2(n11050), .A(n10389), .ZN(P1_U3264) );
  INV_X1 U11209 ( .A(n10390), .ZN(n10392) );
  NAND2_X1 U11210 ( .A1(n10396), .A2(n10395), .ZN(n10512) );
  NAND2_X1 U11211 ( .A1(n10490), .A2(n10399), .ZN(n10477) );
  NAND2_X1 U11212 ( .A1(n10477), .A2(n10479), .ZN(n10401) );
  NAND2_X1 U11213 ( .A1(n10401), .A2(n10400), .ZN(n10472) );
  NAND2_X1 U11214 ( .A1(n10470), .A2(n10402), .ZN(n10448) );
  INV_X1 U11215 ( .A(n10403), .ZN(n10404) );
  XOR2_X1 U11216 ( .A(n10405), .B(n10429), .Z(n10614) );
  NAND2_X1 U11217 ( .A1(n10406), .A2(n10587), .ZN(n10407) );
  NAND2_X1 U11218 ( .A1(n10408), .A2(n10407), .ZN(n10582) );
  OR2_X1 U11219 ( .A1(n10593), .A2(n10694), .ZN(n10409) );
  NAND2_X1 U11220 ( .A1(n10582), .A2(n10409), .ZN(n10411) );
  NAND2_X1 U11221 ( .A1(n10593), .A2(n10694), .ZN(n10410) );
  OR2_X1 U11222 ( .A1(n10684), .A2(n10586), .ZN(n10412) );
  OR2_X1 U11223 ( .A1(n10561), .A2(n10577), .ZN(n10413) );
  NAND2_X1 U11224 ( .A1(n10549), .A2(n10413), .ZN(n10534) );
  NAND2_X1 U11225 ( .A1(n10545), .A2(n10658), .ZN(n10415) );
  OR2_X1 U11226 ( .A1(n10529), .A2(n10416), .ZN(n10417) );
  NAND2_X1 U11227 ( .A1(n10654), .A2(n10659), .ZN(n10418) );
  OR2_X1 U11228 ( .A1(n10654), .A2(n10659), .ZN(n10419) );
  NAND2_X1 U11229 ( .A1(n10647), .A2(n10480), .ZN(n10421) );
  OR2_X1 U11230 ( .A1(n10487), .A2(n10464), .ZN(n10422) );
  NAND2_X1 U11231 ( .A1(n10487), .A2(n10464), .ZN(n10423) );
  NAND2_X1 U11232 ( .A1(n10424), .A2(n10423), .ZN(n10461) );
  OR2_X1 U11233 ( .A1(n10752), .A2(n10425), .ZN(n10426) );
  XNOR2_X1 U11234 ( .A(n10430), .B(n10429), .ZN(n10613) );
  NAND2_X1 U11235 ( .A1(n10613), .A2(n11053), .ZN(n10443) );
  AOI211_X1 U11236 ( .C1(n10618), .C2(n10454), .A(n10591), .B(n10431), .ZN(
        n10616) );
  NAND2_X1 U11237 ( .A1(n10618), .A2(n11047), .ZN(n10439) );
  NAND2_X1 U11238 ( .A1(n10433), .A2(n10432), .ZN(n10615) );
  INV_X1 U11239 ( .A(n10434), .ZN(n10436) );
  OAI22_X1 U11240 ( .A1(n10596), .A2(n10615), .B1(n10436), .B2(n10435), .ZN(
        n10437) );
  AOI21_X1 U11241 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n10596), .A(n10437), 
        .ZN(n10438) );
  OAI211_X1 U11242 ( .C1(n10626), .C2(n10440), .A(n10439), .B(n10438), .ZN(
        n10441) );
  AOI21_X1 U11243 ( .B1(n10616), .B2(n10594), .A(n10441), .ZN(n10442) );
  OAI211_X1 U11244 ( .C1(n10548), .C2(n10614), .A(n10443), .B(n10442), .ZN(
        P1_U3356) );
  AND2_X1 U11245 ( .A1(n10445), .A2(n10447), .ZN(n10446) );
  OR2_X2 U11246 ( .A1(n10444), .A2(n10446), .ZN(n10625) );
  XNOR2_X1 U11247 ( .A(n10448), .B(n10447), .ZN(n10449) );
  NAND2_X1 U11248 ( .A1(n10449), .A2(n10725), .ZN(n10453) );
  OAI22_X1 U11249 ( .A1(n10450), .A2(n10667), .B1(n10633), .B2(n10702), .ZN(
        n10451) );
  INV_X1 U11250 ( .A(n10451), .ZN(n10452) );
  NAND2_X1 U11251 ( .A1(n10453), .A2(n10452), .ZN(n10623) );
  AOI21_X1 U11252 ( .B1(n10620), .B2(n10462), .A(n10591), .ZN(n10455) );
  NAND2_X1 U11253 ( .A1(n10455), .A2(n10454), .ZN(n10621) );
  AOI22_X1 U11254 ( .A1(n10596), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n10456), 
        .B2(n11044), .ZN(n10458) );
  NAND2_X1 U11255 ( .A1(n10620), .A2(n11047), .ZN(n10457) );
  OAI211_X1 U11256 ( .C1(n10621), .C2(n11050), .A(n10458), .B(n10457), .ZN(
        n10459) );
  AOI21_X1 U11257 ( .B1(n10623), .B2(n10601), .A(n10459), .ZN(n10460) );
  OAI21_X1 U11258 ( .B1(n10625), .B2(n10603), .A(n10460), .ZN(P1_U3265) );
  AOI211_X1 U11259 ( .C1(n10752), .C2(n10484), .A(n10591), .B(n5114), .ZN(
        n10627) );
  INV_X1 U11260 ( .A(n10752), .ZN(n10463) );
  NOR2_X1 U11261 ( .A1(n10463), .A2(n10599), .ZN(n10469) );
  NAND2_X1 U11262 ( .A1(n10536), .A2(n10464), .ZN(n10467) );
  AOI22_X1 U11263 ( .A1(n10596), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10465), 
        .B2(n11044), .ZN(n10466) );
  OAI211_X1 U11264 ( .C1(n10626), .C2(n10540), .A(n10467), .B(n10466), .ZN(
        n10468) );
  AOI211_X1 U11265 ( .C1(n10627), .C2(n10594), .A(n10469), .B(n10468), .ZN(
        n10475) );
  OAI21_X1 U11266 ( .B1(n10472), .B2(n10471), .A(n10470), .ZN(n10629) );
  NAND2_X1 U11267 ( .A1(n10629), .A2(n10473), .ZN(n10474) );
  OAI211_X1 U11268 ( .C1(n10630), .C2(n10603), .A(n10475), .B(n10474), .ZN(
        P1_U3266) );
  XNOR2_X1 U11269 ( .A(n10477), .B(n10476), .ZN(n10638) );
  XNOR2_X1 U11270 ( .A(n10478), .B(n10479), .ZN(n10640) );
  NAND2_X1 U11271 ( .A1(n10640), .A2(n11053), .ZN(n10489) );
  NAND2_X1 U11272 ( .A1(n10536), .A2(n10480), .ZN(n10483) );
  AOI22_X1 U11273 ( .A1(n10596), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10481), 
        .B2(n11044), .ZN(n10482) );
  OAI211_X1 U11274 ( .C1(n10633), .C2(n10540), .A(n10483), .B(n10482), .ZN(
        n10486) );
  OAI211_X1 U11275 ( .C1(n10758), .C2(n10495), .A(n10542), .B(n10484), .ZN(
        n10636) );
  NOR2_X1 U11276 ( .A1(n10636), .A2(n11050), .ZN(n10485) );
  AOI211_X1 U11277 ( .C1(n11047), .C2(n10487), .A(n10486), .B(n10485), .ZN(
        n10488) );
  OAI211_X1 U11278 ( .C1(n10638), .C2(n10548), .A(n10489), .B(n10488), .ZN(
        P1_U3267) );
  OAI21_X1 U11279 ( .B1(n10491), .B2(n10493), .A(n10490), .ZN(n10492) );
  INV_X1 U11280 ( .A(n10492), .ZN(n10652) );
  NAND2_X1 U11281 ( .A1(n10494), .A2(n10493), .ZN(n10648) );
  NAND3_X1 U11282 ( .A1(n10649), .A2(n10648), .A3(n11053), .ZN(n10503) );
  AOI211_X1 U11283 ( .C1(n10647), .C2(n10506), .A(n10591), .B(n10495), .ZN(
        n10645) );
  NOR2_X1 U11284 ( .A1(n10496), .A2(n10599), .ZN(n10501) );
  NAND2_X1 U11285 ( .A1(n10536), .A2(n10659), .ZN(n10499) );
  AOI22_X1 U11286 ( .A1(n10596), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10497), 
        .B2(n11044), .ZN(n10498) );
  OAI211_X1 U11287 ( .C1(n10643), .C2(n10540), .A(n10499), .B(n10498), .ZN(
        n10500) );
  AOI211_X1 U11288 ( .C1(n10645), .C2(n10594), .A(n10501), .B(n10500), .ZN(
        n10502) );
  OAI211_X1 U11289 ( .C1(n10652), .C2(n10548), .A(n10503), .B(n10502), .ZN(
        P1_U3268) );
  XOR2_X1 U11290 ( .A(n10504), .B(n10511), .Z(n10657) );
  INV_X1 U11291 ( .A(n10505), .ZN(n10525) );
  INV_X1 U11292 ( .A(n10506), .ZN(n10507) );
  AOI211_X1 U11293 ( .C1(n10654), .C2(n10525), .A(n10591), .B(n10507), .ZN(
        n10653) );
  AOI22_X1 U11294 ( .A1(n10596), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n10508), 
        .B2(n11044), .ZN(n10509) );
  OAI21_X1 U11295 ( .B1(n10510), .B2(n10599), .A(n10509), .ZN(n10517) );
  AOI21_X1 U11296 ( .B1(n10512), .B2(n10511), .A(n11020), .ZN(n10515) );
  OAI22_X1 U11297 ( .A1(n10668), .A2(n10702), .B1(n10634), .B2(n10667), .ZN(
        n10513) );
  AOI21_X1 U11298 ( .B1(n10515), .B2(n10514), .A(n10513), .ZN(n10656) );
  NOR2_X1 U11299 ( .A1(n10656), .A2(n10596), .ZN(n10516) );
  AOI211_X1 U11300 ( .C1(n10653), .C2(n10594), .A(n10517), .B(n10516), .ZN(
        n10518) );
  OAI21_X1 U11301 ( .B1(n10657), .B2(n10603), .A(n10518), .ZN(P1_U3269) );
  XNOR2_X1 U11302 ( .A(n10519), .B(n10521), .ZN(n10662) );
  OAI21_X1 U11303 ( .B1(n5175), .B2(n10521), .A(n10520), .ZN(n10664) );
  NAND2_X1 U11304 ( .A1(n10664), .A2(n11053), .ZN(n10531) );
  NAND2_X1 U11305 ( .A1(n10536), .A2(n10658), .ZN(n10524) );
  AOI22_X1 U11306 ( .A1(n10596), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10522), 
        .B2(n11044), .ZN(n10523) );
  OAI211_X1 U11307 ( .C1(n10644), .C2(n10540), .A(n10524), .B(n10523), .ZN(
        n10528) );
  INV_X1 U11308 ( .A(n10541), .ZN(n10526) );
  OAI211_X1 U11309 ( .C1(n10764), .C2(n10526), .A(n10525), .B(n10542), .ZN(
        n10660) );
  NOR2_X1 U11310 ( .A1(n10660), .A2(n11050), .ZN(n10527) );
  AOI211_X1 U11311 ( .C1(n11047), .C2(n10529), .A(n10528), .B(n10527), .ZN(
        n10530) );
  OAI211_X1 U11312 ( .C1(n10662), .C2(n10548), .A(n10531), .B(n10530), .ZN(
        P1_U3270) );
  XNOR2_X1 U11313 ( .A(n10535), .B(n5142), .ZN(n10673) );
  INV_X1 U11314 ( .A(n10532), .ZN(n10533) );
  AOI21_X1 U11315 ( .B1(n10535), .B2(n10534), .A(n10533), .ZN(n10675) );
  NAND2_X1 U11316 ( .A1(n10675), .A2(n11053), .ZN(n10547) );
  NAND2_X1 U11317 ( .A1(n10536), .A2(n10577), .ZN(n10539) );
  AOI22_X1 U11318 ( .A1(n10596), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10537), 
        .B2(n11044), .ZN(n10538) );
  OAI211_X1 U11319 ( .C1(n10668), .C2(n10540), .A(n10539), .B(n10538), .ZN(
        n10544) );
  OAI211_X1 U11320 ( .C1(n10768), .C2(n10560), .A(n10542), .B(n10541), .ZN(
        n10671) );
  NOR2_X1 U11321 ( .A1(n10671), .A2(n11050), .ZN(n10543) );
  AOI211_X1 U11322 ( .C1(n11047), .C2(n10545), .A(n10544), .B(n10543), .ZN(
        n10546) );
  OAI211_X1 U11323 ( .C1(n10673), .C2(n10548), .A(n10547), .B(n10546), .ZN(
        P1_U3271) );
  OAI21_X1 U11324 ( .B1(n10550), .B2(n10555), .A(n10549), .ZN(n10680) );
  INV_X1 U11325 ( .A(n10680), .ZN(n10567) );
  INV_X1 U11326 ( .A(n10551), .ZN(n10552) );
  NOR2_X1 U11327 ( .A1(n10553), .A2(n10552), .ZN(n10575) );
  NAND2_X1 U11328 ( .A1(n10575), .A2(n10576), .ZN(n10574) );
  NAND2_X1 U11329 ( .A1(n10574), .A2(n10554), .ZN(n10556) );
  XNOR2_X1 U11330 ( .A(n10556), .B(n10555), .ZN(n10557) );
  OAI222_X1 U11331 ( .A1(n10667), .A2(n10559), .B1(n10702), .B2(n10558), .C1(
        n10557), .C2(n11020), .ZN(n10678) );
  AOI211_X1 U11332 ( .C1(n10561), .C2(n10570), .A(n10591), .B(n10560), .ZN(
        n10679) );
  NAND2_X1 U11333 ( .A1(n10679), .A2(n10594), .ZN(n10564) );
  AOI22_X1 U11334 ( .A1(n10596), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10562), 
        .B2(n11044), .ZN(n10563) );
  OAI211_X1 U11335 ( .C1(n10772), .C2(n10599), .A(n10564), .B(n10563), .ZN(
        n10565) );
  AOI21_X1 U11336 ( .B1(n10678), .B2(n10601), .A(n10565), .ZN(n10566) );
  OAI21_X1 U11337 ( .B1(n10567), .B2(n10603), .A(n10566), .ZN(P1_U3272) );
  XOR2_X1 U11338 ( .A(n10568), .B(n10576), .Z(n10687) );
  INV_X1 U11339 ( .A(n10569), .ZN(n10590) );
  INV_X1 U11340 ( .A(n10570), .ZN(n10571) );
  AOI211_X1 U11341 ( .C1(n10684), .C2(n10590), .A(n10591), .B(n10571), .ZN(
        n10683) );
  AOI22_X1 U11342 ( .A1(n10596), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10572), 
        .B2(n11044), .ZN(n10573) );
  OAI21_X1 U11343 ( .B1(n10378), .B2(n10599), .A(n10573), .ZN(n10580) );
  OAI21_X1 U11344 ( .B1(n10576), .B2(n10575), .A(n10574), .ZN(n10578) );
  AOI222_X1 U11345 ( .A1(n10725), .A2(n10578), .B1(n10694), .B2(n10732), .C1(
        n10577), .C2(n10731), .ZN(n10686) );
  NOR2_X1 U11346 ( .A1(n10686), .A2(n10596), .ZN(n10579) );
  AOI211_X1 U11347 ( .C1(n10683), .C2(n10594), .A(n10580), .B(n10579), .ZN(
        n10581) );
  OAI21_X1 U11348 ( .B1(n10603), .B2(n10687), .A(n10581), .ZN(P1_U3273) );
  XNOR2_X1 U11349 ( .A(n10582), .B(n10583), .ZN(n10690) );
  INV_X1 U11350 ( .A(n10690), .ZN(n10604) );
  XNOR2_X1 U11351 ( .A(n10584), .B(n10583), .ZN(n10585) );
  NAND2_X1 U11352 ( .A1(n10585), .A2(n10725), .ZN(n10589) );
  AOI22_X1 U11353 ( .A1(n10587), .A2(n10732), .B1(n10586), .B2(n10731), .ZN(
        n10588) );
  NAND2_X1 U11354 ( .A1(n10589), .A2(n10588), .ZN(n10688) );
  INV_X1 U11355 ( .A(n10593), .ZN(n10778) );
  AOI211_X1 U11356 ( .C1(n10593), .C2(n10592), .A(n10591), .B(n10569), .ZN(
        n10689) );
  NAND2_X1 U11357 ( .A1(n10689), .A2(n10594), .ZN(n10598) );
  AOI22_X1 U11358 ( .A1(n10596), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10595), 
        .B2(n11044), .ZN(n10597) );
  OAI211_X1 U11359 ( .C1(n10778), .C2(n10599), .A(n10598), .B(n10597), .ZN(
        n10600) );
  AOI21_X1 U11360 ( .B1(n10601), .B2(n10688), .A(n10600), .ZN(n10602) );
  OAI21_X1 U11361 ( .B1(n10604), .B2(n10603), .A(n10602), .ZN(P1_U3274) );
  NOR2_X1 U11362 ( .A1(n10606), .A2(n10605), .ZN(n10740) );
  MUX2_X1 U11363 ( .A(n10607), .B(n10740), .S(n11094), .Z(n10608) );
  OAI21_X1 U11364 ( .B1(n10743), .B2(n10693), .A(n10608), .ZN(P1_U3553) );
  INV_X1 U11365 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10611) );
  AND2_X1 U11366 ( .A1(n10610), .A2(n10609), .ZN(n10744) );
  MUX2_X1 U11367 ( .A(n10611), .B(n10744), .S(n11094), .Z(n10612) );
  OAI21_X1 U11368 ( .B1(n10747), .B2(n10693), .A(n10612), .ZN(P1_U3552) );
  NAND2_X1 U11369 ( .A1(n10613), .A2(n11091), .ZN(n10619) );
  OAI21_X1 U11370 ( .B1(n10626), .B2(n10702), .A(n10615), .ZN(n10617) );
  OAI21_X1 U11371 ( .B1(n5396), .B2(n11088), .A(n10621), .ZN(n10622) );
  NOR2_X1 U11372 ( .A1(n10623), .A2(n10622), .ZN(n10624) );
  MUX2_X1 U11373 ( .A(n10749), .B(P1_REG1_REG_28__SCAN_IN), .S(n11093), .Z(
        P1_U3550) );
  OAI22_X1 U11374 ( .A1(n10643), .A2(n10702), .B1(n10626), .B2(n10667), .ZN(
        n10628) );
  INV_X1 U11375 ( .A(n10632), .ZN(P1_U3549) );
  INV_X1 U11376 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10641) );
  OAI22_X1 U11377 ( .A1(n10634), .A2(n10702), .B1(n10633), .B2(n10667), .ZN(
        n10635) );
  INV_X1 U11378 ( .A(n10635), .ZN(n10637) );
  OAI211_X1 U11379 ( .C1(n10638), .C2(n11020), .A(n10637), .B(n10636), .ZN(
        n10639) );
  AOI21_X1 U11380 ( .B1(n10640), .B2(n11091), .A(n10639), .ZN(n10755) );
  MUX2_X1 U11381 ( .A(n10641), .B(n10755), .S(n11094), .Z(n10642) );
  OAI21_X1 U11382 ( .B1(n10758), .B2(n10693), .A(n10642), .ZN(P1_U3548) );
  OAI22_X1 U11383 ( .A1(n10644), .A2(n10702), .B1(n10643), .B2(n10667), .ZN(
        n10646) );
  AOI211_X1 U11384 ( .C1(n10707), .C2(n10647), .A(n10646), .B(n10645), .ZN(
        n10651) );
  NAND3_X1 U11385 ( .A1(n10649), .A2(n10648), .A3(n11091), .ZN(n10650) );
  OAI211_X1 U11386 ( .C1(n11020), .C2(n10652), .A(n10651), .B(n10650), .ZN(
        n10759) );
  MUX2_X1 U11387 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10759), .S(n11094), .Z(
        P1_U3547) );
  AOI21_X1 U11388 ( .B1(n10707), .B2(n10654), .A(n10653), .ZN(n10655) );
  OAI211_X1 U11389 ( .C1(n10657), .C2(n11021), .A(n10656), .B(n10655), .ZN(
        n10760) );
  MUX2_X1 U11390 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10760), .S(n11094), .Z(
        P1_U3546) );
  INV_X1 U11391 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U11392 ( .A1(n10659), .A2(n10731), .B1(n10732), .B2(n10658), .ZN(
        n10661) );
  OAI211_X1 U11393 ( .C1(n10662), .C2(n11020), .A(n10661), .B(n10660), .ZN(
        n10663) );
  AOI21_X1 U11394 ( .B1(n10664), .B2(n11091), .A(n10663), .ZN(n10761) );
  MUX2_X1 U11395 ( .A(n10665), .B(n10761), .S(n11094), .Z(n10666) );
  OAI21_X1 U11396 ( .B1(n10764), .B2(n10693), .A(n10666), .ZN(P1_U3545) );
  INV_X1 U11397 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10676) );
  OAI22_X1 U11398 ( .A1(n10669), .A2(n10702), .B1(n10668), .B2(n10667), .ZN(
        n10670) );
  INV_X1 U11399 ( .A(n10670), .ZN(n10672) );
  OAI211_X1 U11400 ( .C1(n10673), .C2(n11020), .A(n10672), .B(n10671), .ZN(
        n10674) );
  AOI21_X1 U11401 ( .B1(n10675), .B2(n11091), .A(n10674), .ZN(n10765) );
  MUX2_X1 U11402 ( .A(n10676), .B(n10765), .S(n11094), .Z(n10677) );
  OAI21_X1 U11403 ( .B1(n10768), .B2(n10693), .A(n10677), .ZN(P1_U3544) );
  INV_X1 U11404 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10681) );
  AOI211_X1 U11405 ( .C1(n10680), .C2(n11091), .A(n10679), .B(n10678), .ZN(
        n10769) );
  MUX2_X1 U11406 ( .A(n10681), .B(n10769), .S(n11094), .Z(n10682) );
  OAI21_X1 U11407 ( .B1(n10772), .B2(n10693), .A(n10682), .ZN(P1_U3543) );
  AOI21_X1 U11408 ( .B1(n10707), .B2(n10684), .A(n10683), .ZN(n10685) );
  OAI211_X1 U11409 ( .C1(n10687), .C2(n11021), .A(n10686), .B(n10685), .ZN(
        n10773) );
  MUX2_X1 U11410 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10773), .S(n11094), .Z(
        P1_U3542) );
  AOI211_X1 U11411 ( .C1(n10690), .C2(n11091), .A(n10689), .B(n10688), .ZN(
        n10774) );
  MUX2_X1 U11412 ( .A(n10691), .B(n10774), .S(n11094), .Z(n10692) );
  OAI21_X1 U11413 ( .B1(n10778), .B2(n10693), .A(n10692), .ZN(P1_U3541) );
  AOI22_X1 U11414 ( .A1(n10694), .A2(n10731), .B1(n10732), .B2(n10711), .ZN(
        n10695) );
  OAI211_X1 U11415 ( .C1(n10697), .C2(n11088), .A(n10696), .B(n10695), .ZN(
        n10698) );
  AOI21_X1 U11416 ( .B1(n10699), .B2(n10725), .A(n10698), .ZN(n10700) );
  OAI21_X1 U11417 ( .B1(n10701), .B2(n11021), .A(n10700), .ZN(n10779) );
  MUX2_X1 U11418 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10779), .S(n11094), .Z(
        P1_U3540) );
  NOR2_X1 U11419 ( .A1(n10703), .A2(n10702), .ZN(n10705) );
  AOI211_X1 U11420 ( .C1(n10707), .C2(n10706), .A(n10705), .B(n10704), .ZN(
        n10708) );
  OAI211_X1 U11421 ( .C1(n10710), .C2(n11021), .A(n10709), .B(n10708), .ZN(
        n10780) );
  MUX2_X1 U11422 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10780), .S(n11094), .Z(
        P1_U3539) );
  AOI22_X1 U11423 ( .A1(n10711), .A2(n10731), .B1(n10732), .B2(n10730), .ZN(
        n10712) );
  OAI211_X1 U11424 ( .C1(n10714), .C2(n11088), .A(n10713), .B(n10712), .ZN(
        n10715) );
  AOI21_X1 U11425 ( .B1(n10716), .B2(n10725), .A(n10715), .ZN(n10717) );
  OAI21_X1 U11426 ( .B1(n10718), .B2(n11021), .A(n10717), .ZN(n10781) );
  MUX2_X1 U11427 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10781), .S(n11094), .Z(
        P1_U3538) );
  AOI22_X1 U11428 ( .A1(n10720), .A2(n10732), .B1(n10731), .B2(n10719), .ZN(
        n10721) );
  OAI211_X1 U11429 ( .C1(n10723), .C2(n11088), .A(n10722), .B(n10721), .ZN(
        n10724) );
  AOI21_X1 U11430 ( .B1(n10726), .B2(n10725), .A(n10724), .ZN(n10727) );
  OAI21_X1 U11431 ( .B1(n10728), .B2(n11021), .A(n10727), .ZN(n10782) );
  MUX2_X1 U11432 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10782), .S(n11094), .Z(
        P1_U3537) );
  AOI22_X1 U11433 ( .A1(n10733), .A2(n10732), .B1(n10731), .B2(n10730), .ZN(
        n10734) );
  OAI211_X1 U11434 ( .C1(n5387), .C2(n11088), .A(n10735), .B(n10734), .ZN(
        n10736) );
  INV_X1 U11435 ( .A(n10736), .ZN(n10738) );
  OAI211_X1 U11436 ( .C1(n10739), .C2(n11021), .A(n10738), .B(n10737), .ZN(
        n10783) );
  MUX2_X1 U11437 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10783), .S(n11094), .Z(
        P1_U3536) );
  INV_X1 U11438 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10741) );
  INV_X2 U11439 ( .A(n11095), .ZN(n11079) );
  MUX2_X1 U11440 ( .A(n10741), .B(n10740), .S(n11079), .Z(n10742) );
  OAI21_X1 U11441 ( .B1(n10743), .B2(n10777), .A(n10742), .ZN(P1_U3521) );
  INV_X1 U11442 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10745) );
  MUX2_X1 U11443 ( .A(n10745), .B(n10744), .S(n11079), .Z(n10746) );
  OAI21_X1 U11444 ( .B1(n10747), .B2(n10777), .A(n10746), .ZN(P1_U3520) );
  MUX2_X1 U11445 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10748), .S(n11079), .Z(
        P1_U3519) );
  MUX2_X1 U11446 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10749), .S(n11079), .Z(
        P1_U3518) );
  INV_X1 U11447 ( .A(n10777), .ZN(n10753) );
  AOI21_X1 U11448 ( .B1(n10753), .B2(n10752), .A(n10751), .ZN(n10754) );
  INV_X1 U11449 ( .A(n10754), .ZN(P1_U3517) );
  INV_X1 U11450 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10756) );
  MUX2_X1 U11451 ( .A(n10756), .B(n10755), .S(n11079), .Z(n10757) );
  OAI21_X1 U11452 ( .B1(n10758), .B2(n10777), .A(n10757), .ZN(P1_U3516) );
  MUX2_X1 U11453 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10759), .S(n11079), .Z(
        P1_U3515) );
  MUX2_X1 U11454 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10760), .S(n11079), .Z(
        P1_U3514) );
  INV_X1 U11455 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10762) );
  MUX2_X1 U11456 ( .A(n10762), .B(n10761), .S(n11079), .Z(n10763) );
  OAI21_X1 U11457 ( .B1(n10764), .B2(n10777), .A(n10763), .ZN(P1_U3513) );
  INV_X1 U11458 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10766) );
  MUX2_X1 U11459 ( .A(n10766), .B(n10765), .S(n11079), .Z(n10767) );
  OAI21_X1 U11460 ( .B1(n10768), .B2(n10777), .A(n10767), .ZN(P1_U3512) );
  INV_X1 U11461 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10770) );
  MUX2_X1 U11462 ( .A(n10770), .B(n10769), .S(n11079), .Z(n10771) );
  OAI21_X1 U11463 ( .B1(n10772), .B2(n10777), .A(n10771), .ZN(P1_U3511) );
  MUX2_X1 U11464 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10773), .S(n11079), .Z(
        P1_U3510) );
  INV_X1 U11465 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10775) );
  MUX2_X1 U11466 ( .A(n10775), .B(n10774), .S(n11079), .Z(n10776) );
  OAI21_X1 U11467 ( .B1(n10778), .B2(n10777), .A(n10776), .ZN(P1_U3509) );
  MUX2_X1 U11468 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10779), .S(n11079), .Z(
        P1_U3507) );
  MUX2_X1 U11469 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10780), .S(n11079), .Z(
        P1_U3504) );
  MUX2_X1 U11470 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10781), .S(n11079), .Z(
        P1_U3501) );
  MUX2_X1 U11471 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10782), .S(n11079), .Z(
        P1_U3498) );
  MUX2_X1 U11472 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10783), .S(n11079), .Z(
        P1_U3495) );
  MUX2_X1 U11473 ( .A(P1_D_REG_1__SCAN_IN), .B(n10784), .S(n10803), .Z(
        P1_U3440) );
  MUX2_X1 U11474 ( .A(P1_D_REG_0__SCAN_IN), .B(n10785), .S(n10803), .Z(
        P1_U3439) );
  NOR4_X1 U11475 ( .A1(n6450), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n6447), .ZN(n10786) );
  AOI21_X1 U11476 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10796), .A(n10786), 
        .ZN(n10787) );
  OAI21_X1 U11477 ( .B1(n10788), .B2(n10799), .A(n10787), .ZN(P1_U3324) );
  INV_X1 U11478 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10789) );
  OAI222_X1 U11479 ( .A1(P1_U3086), .A2(n10791), .B1(n10799), .B2(n10790), 
        .C1(n10789), .C2(n10792), .ZN(P1_U3326) );
  INV_X1 U11480 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10793) );
  OAI222_X1 U11481 ( .A1(P1_U3086), .A2(n10795), .B1(n10799), .B2(n10794), 
        .C1(n10793), .C2(n10792), .ZN(P1_U3328) );
  AOI22_X1 U11482 ( .A1(n10797), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10796), .ZN(n10798) );
  OAI21_X1 U11483 ( .B1(n10800), .B2(n10799), .A(n10798), .ZN(P1_U3329) );
  INV_X1 U11484 ( .A(n10801), .ZN(n10802) );
  MUX2_X1 U11485 ( .A(n10802), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U11486 ( .A1(n10835), .A2(n10805), .ZN(P1_U3323) );
  NOR2_X1 U11487 ( .A1(n10835), .A2(n10806), .ZN(P1_U3322) );
  NOR2_X1 U11488 ( .A1(n10835), .A2(n10807), .ZN(P1_U3321) );
  NOR2_X1 U11489 ( .A1(n10835), .A2(n10808), .ZN(P1_U3320) );
  INV_X1 U11490 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10809) );
  NOR2_X1 U11491 ( .A1(n10835), .A2(n10809), .ZN(P1_U3319) );
  INV_X1 U11492 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10810) );
  NOR2_X1 U11493 ( .A1(n10835), .A2(n10810), .ZN(P1_U3318) );
  INV_X1 U11494 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10811) );
  NOR2_X1 U11495 ( .A1(n10835), .A2(n10811), .ZN(P1_U3317) );
  INV_X1 U11496 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10812) );
  NOR2_X1 U11497 ( .A1(n10835), .A2(n10812), .ZN(P1_U3316) );
  INV_X1 U11498 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10813) );
  NOR2_X1 U11499 ( .A1(n10835), .A2(n10813), .ZN(P1_U3315) );
  INV_X1 U11500 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10814) );
  NOR2_X1 U11501 ( .A1(n10835), .A2(n10814), .ZN(P1_U3314) );
  INV_X1 U11502 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10815) );
  NOR2_X1 U11503 ( .A1(n10835), .A2(n10815), .ZN(P1_U3313) );
  INV_X1 U11504 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10816) );
  NOR2_X1 U11505 ( .A1(n10835), .A2(n10816), .ZN(P1_U3312) );
  INV_X1 U11506 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10817) );
  NOR2_X1 U11507 ( .A1(n10835), .A2(n10817), .ZN(P1_U3311) );
  INV_X1 U11508 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10818) );
  NOR2_X1 U11509 ( .A1(n10835), .A2(n10818), .ZN(P1_U3310) );
  INV_X1 U11510 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10819) );
  NOR2_X1 U11511 ( .A1(n10835), .A2(n10819), .ZN(P1_U3309) );
  INV_X1 U11512 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10820) );
  NOR2_X1 U11513 ( .A1(n10835), .A2(n10820), .ZN(P1_U3308) );
  INV_X1 U11514 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10821) );
  NOR2_X1 U11515 ( .A1(n10835), .A2(n10821), .ZN(P1_U3307) );
  INV_X1 U11516 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10822) );
  NOR2_X1 U11517 ( .A1(n10835), .A2(n10822), .ZN(P1_U3306) );
  INV_X1 U11518 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10823) );
  NOR2_X1 U11519 ( .A1(n10835), .A2(n10823), .ZN(P1_U3305) );
  INV_X1 U11520 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10824) );
  NOR2_X1 U11521 ( .A1(n10835), .A2(n10824), .ZN(P1_U3304) );
  INV_X1 U11522 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10825) );
  NOR2_X1 U11523 ( .A1(n10835), .A2(n10825), .ZN(P1_U3303) );
  INV_X1 U11524 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10826) );
  NOR2_X1 U11525 ( .A1(n10835), .A2(n10826), .ZN(P1_U3302) );
  INV_X1 U11526 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10827) );
  NOR2_X1 U11527 ( .A1(n10835), .A2(n10827), .ZN(P1_U3301) );
  INV_X1 U11528 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10828) );
  NOR2_X1 U11529 ( .A1(n10835), .A2(n10828), .ZN(P1_U3300) );
  INV_X1 U11530 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10829) );
  NOR2_X1 U11531 ( .A1(n10835), .A2(n10829), .ZN(P1_U3299) );
  INV_X1 U11532 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10830) );
  NOR2_X1 U11533 ( .A1(n10835), .A2(n10830), .ZN(P1_U3298) );
  INV_X1 U11534 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U11535 ( .A1(n10835), .A2(n10831), .ZN(P1_U3297) );
  INV_X1 U11536 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10832) );
  NOR2_X1 U11537 ( .A1(n10835), .A2(n10832), .ZN(P1_U3296) );
  INV_X1 U11538 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10833) );
  NOR2_X1 U11539 ( .A1(n10835), .A2(n10833), .ZN(P1_U3295) );
  INV_X1 U11540 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10834) );
  NOR2_X1 U11541 ( .A1(n10835), .A2(n10834), .ZN(P1_U3294) );
  XOR2_X1 U11542 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11543 ( .A1(n10840), .A2(n10839), .B1(n10840), .B2(n10838), .C1(
        n10837), .C2(n10836), .ZN(ADD_1068_U5) );
  AOI21_X1 U11544 ( .B1(n10843), .B2(n10842), .A(n10841), .ZN(ADD_1068_U54) );
  AOI21_X1 U11545 ( .B1(n10846), .B2(n10845), .A(n10844), .ZN(ADD_1068_U53) );
  OAI21_X1 U11546 ( .B1(n10849), .B2(n10848), .A(n10847), .ZN(ADD_1068_U52) );
  OAI21_X1 U11547 ( .B1(n10852), .B2(n10851), .A(n10850), .ZN(ADD_1068_U51) );
  OAI21_X1 U11548 ( .B1(n10855), .B2(n10854), .A(n10853), .ZN(ADD_1068_U50) );
  OAI21_X1 U11549 ( .B1(n10858), .B2(n10857), .A(n10856), .ZN(ADD_1068_U49) );
  OAI21_X1 U11550 ( .B1(n10861), .B2(n10860), .A(n10859), .ZN(ADD_1068_U48) );
  OAI21_X1 U11551 ( .B1(n10864), .B2(n10863), .A(n10862), .ZN(ADD_1068_U47) );
  OAI21_X1 U11552 ( .B1(n10867), .B2(n10866), .A(n10865), .ZN(ADD_1068_U63) );
  OAI21_X1 U11553 ( .B1(n10870), .B2(n10869), .A(n10868), .ZN(ADD_1068_U62) );
  OAI21_X1 U11554 ( .B1(n10873), .B2(n10872), .A(n10871), .ZN(ADD_1068_U61) );
  OAI21_X1 U11555 ( .B1(n10876), .B2(n10875), .A(n10874), .ZN(ADD_1068_U60) );
  OAI21_X1 U11556 ( .B1(n10879), .B2(n10878), .A(n10877), .ZN(ADD_1068_U59) );
  OAI21_X1 U11557 ( .B1(n10882), .B2(n10881), .A(n10880), .ZN(ADD_1068_U58) );
  OAI21_X1 U11558 ( .B1(n10885), .B2(n10884), .A(n10883), .ZN(ADD_1068_U57) );
  OAI21_X1 U11559 ( .B1(n10888), .B2(n10887), .A(n10886), .ZN(ADD_1068_U56) );
  OAI21_X1 U11560 ( .B1(n10891), .B2(n10890), .A(n10889), .ZN(ADD_1068_U55) );
  AOI22_X1 U11561 ( .A1(n10976), .A2(P2_IR_REG_0__SCAN_IN), .B1(n10999), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10897) );
  OAI21_X1 U11562 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10893), .A(n10892), .ZN(
        n10894) );
  OAI21_X1 U11563 ( .B1(n10996), .B2(n10895), .A(n10894), .ZN(n10896) );
  OAI211_X1 U11564 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10898), .A(n10897), .B(
        n10896), .ZN(P2_U3182) );
  INV_X1 U11565 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10919) );
  OAI21_X1 U11566 ( .B1(n10901), .B2(n10900), .A(n10899), .ZN(n10904) );
  NOR2_X1 U11567 ( .A1(n10902), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10903) );
  AOI21_X1 U11568 ( .B1(n10983), .B2(n10904), .A(n10903), .ZN(n10911) );
  NOR2_X1 U11569 ( .A1(n10906), .A2(n10905), .ZN(n10908) );
  NOR2_X1 U11570 ( .A1(n10908), .A2(n10907), .ZN(n10909) );
  OR2_X1 U11571 ( .A1(n11011), .A2(n10909), .ZN(n10910) );
  OAI211_X1 U11572 ( .C1(n11000), .C2(n10912), .A(n10911), .B(n10910), .ZN(
        n10913) );
  INV_X1 U11573 ( .A(n10913), .ZN(n10918) );
  XOR2_X1 U11574 ( .A(n10915), .B(n10914), .Z(n10916) );
  NAND2_X1 U11575 ( .A1(n10916), .A2(n10996), .ZN(n10917) );
  OAI211_X1 U11576 ( .C1(n10919), .C2(n10940), .A(n10918), .B(n10917), .ZN(
        P2_U3184) );
  INV_X1 U11577 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10941) );
  INV_X1 U11578 ( .A(n10920), .ZN(n10923) );
  NAND2_X1 U11579 ( .A1(n10923), .A2(n10922), .ZN(n10924) );
  AND2_X1 U11580 ( .A1(n10925), .A2(n10924), .ZN(n10932) );
  XNOR2_X1 U11581 ( .A(n10927), .B(n10926), .ZN(n10928) );
  OR2_X1 U11582 ( .A1(n11008), .A2(n10928), .ZN(n10931) );
  INV_X1 U11583 ( .A(n10929), .ZN(n10930) );
  OAI211_X1 U11584 ( .C1(n10932), .C2(n11011), .A(n10931), .B(n10930), .ZN(
        n10933) );
  AOI21_X1 U11585 ( .B1(n10934), .B2(n10976), .A(n10933), .ZN(n10939) );
  OAI211_X1 U11586 ( .C1(n10937), .C2(n10936), .A(n10935), .B(n10996), .ZN(
        n10938) );
  OAI211_X1 U11587 ( .C1(n10941), .C2(n10940), .A(n10939), .B(n10938), .ZN(
        P2_U3186) );
  OAI21_X1 U11588 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n10943), .A(n10942), .ZN(
        n10945) );
  AOI22_X1 U11589 ( .A1(n10945), .A2(n10983), .B1(n10944), .B2(n10976), .ZN(
        n10956) );
  AOI21_X1 U11590 ( .B1(n10947), .B2(n5900), .A(n10946), .ZN(n10948) );
  NOR2_X1 U11591 ( .A1(n10948), .A2(n11011), .ZN(n10949) );
  AOI211_X1 U11592 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n10999), .A(n10950), .B(
        n10949), .ZN(n10955) );
  OAI211_X1 U11593 ( .C1(n10953), .C2(n10952), .A(n10951), .B(n10996), .ZN(
        n10954) );
  NAND3_X1 U11594 ( .A1(n10956), .A2(n10955), .A3(n10954), .ZN(P2_U3187) );
  AOI22_X1 U11595 ( .A1(n10976), .A2(n10957), .B1(n10999), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n10974) );
  INV_X1 U11596 ( .A(n10958), .ZN(n10960) );
  NAND2_X1 U11597 ( .A1(n10960), .A2(n10959), .ZN(n10961) );
  XNOR2_X1 U11598 ( .A(n10962), .B(n10961), .ZN(n10967) );
  OAI21_X1 U11599 ( .B1(n10965), .B2(n10964), .A(n10963), .ZN(n10966) );
  AOI22_X1 U11600 ( .A1(n10967), .A2(n10996), .B1(n10983), .B2(n10966), .ZN(
        n10973) );
  NAND2_X1 U11601 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3151), .ZN(n10972)
         );
  AOI21_X1 U11602 ( .B1(n5191), .B2(n10969), .A(n10968), .ZN(n10970) );
  OR2_X1 U11603 ( .A1(n10970), .A2(n11011), .ZN(n10971) );
  NAND4_X1 U11604 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        P2_U3192) );
  AOI22_X1 U11605 ( .A1(n10976), .A2(n10975), .B1(n10999), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n10991) );
  OAI21_X1 U11606 ( .B1(n10979), .B2(n10978), .A(n10977), .ZN(n10984) );
  OAI21_X1 U11607 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n10981), .A(n10980), 
        .ZN(n10982) );
  AOI22_X1 U11608 ( .A1(n10984), .A2(n10996), .B1(n10983), .B2(n10982), .ZN(
        n10990) );
  NAND2_X1 U11609 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3151), .ZN(n10989)
         );
  AOI21_X1 U11610 ( .B1(n10986), .B2(n6005), .A(n10985), .ZN(n10987) );
  OR2_X1 U11611 ( .A1(n11011), .A2(n10987), .ZN(n10988) );
  NAND4_X1 U11612 ( .A1(n10991), .A2(n10990), .A3(n10989), .A4(n10988), .ZN(
        P2_U3193) );
  INV_X1 U11613 ( .A(n10992), .ZN(n10994) );
  NAND2_X1 U11614 ( .A1(n10994), .A2(n10993), .ZN(n11002) );
  AND3_X1 U11615 ( .A1(n11002), .A2(n10996), .A3(n10995), .ZN(n10997) );
  AOI211_X1 U11616 ( .C1(n10999), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n10998), 
        .B(n10997), .ZN(n11018) );
  OAI21_X1 U11617 ( .B1(n11002), .B2(n11001), .A(n11000), .ZN(n11004) );
  NAND2_X1 U11618 ( .A1(n11004), .A2(n11003), .ZN(n11017) );
  AOI21_X1 U11619 ( .B1(n11007), .B2(n11006), .A(n11005), .ZN(n11009) );
  OR2_X1 U11620 ( .A1(n11009), .A2(n11008), .ZN(n11016) );
  AND2_X1 U11621 ( .A1(n5180), .A2(n11010), .ZN(n11014) );
  INV_X1 U11622 ( .A(n11011), .ZN(n11012) );
  OAI21_X1 U11623 ( .B1(n11014), .B2(n11013), .A(n11012), .ZN(n11015) );
  NAND4_X1 U11624 ( .A1(n11018), .A2(n11017), .A3(n11016), .A4(n11015), .ZN(
        P2_U3200) );
  XNOR2_X1 U11625 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11626 ( .B1(n11021), .B2(n11020), .A(n11019), .ZN(n11025) );
  INV_X1 U11627 ( .A(n11022), .ZN(n11023) );
  NOR3_X1 U11628 ( .A1(n11025), .A2(n11024), .A3(n11023), .ZN(n11028) );
  AOI22_X1 U11629 ( .A1(n11094), .A2(n11028), .B1(n11026), .B2(n11093), .ZN(
        P1_U3522) );
  INV_X1 U11630 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U11631 ( .A1(n11079), .A2(n11028), .B1(n11027), .B2(n11095), .ZN(
        P1_U3453) );
  INV_X1 U11632 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U11633 ( .A1(n11108), .A2(n11030), .B1(n11029), .B2(n11105), .ZN(
        P2_U3390) );
  INV_X1 U11634 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U11635 ( .A1(n11108), .A2(n11032), .B1(n11031), .B2(n11105), .ZN(
        P2_U3393) );
  MUX2_X1 U11636 ( .A(n11033), .B(P2_REG0_REG_2__SCAN_IN), .S(n11105), .Z(
        P2_U3396) );
  AOI22_X1 U11637 ( .A1(n11108), .A2(n11034), .B1(n5886), .B2(n11105), .ZN(
        P2_U3402) );
  OAI21_X1 U11638 ( .B1(n11036), .B2(n11088), .A(n11035), .ZN(n11038) );
  AOI211_X1 U11639 ( .C1(n11091), .C2(n11039), .A(n11038), .B(n11037), .ZN(
        n11041) );
  AOI22_X1 U11640 ( .A1(n11094), .A2(n11041), .B1(n7390), .B2(n11093), .ZN(
        P1_U3526) );
  INV_X1 U11641 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U11642 ( .A1(n11079), .A2(n11041), .B1(n11040), .B2(n11095), .ZN(
        P1_U3465) );
  INV_X1 U11643 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U11644 ( .A1(n11108), .A2(n11043), .B1(n11042), .B2(n11105), .ZN(
        P2_U3405) );
  AOI22_X1 U11645 ( .A1(n10596), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n11045), 
        .B2(n11044), .ZN(n11049) );
  NAND2_X1 U11646 ( .A1(n11047), .A2(n11046), .ZN(n11048) );
  OAI211_X1 U11647 ( .C1(n11051), .C2(n11050), .A(n11049), .B(n11048), .ZN(
        n11052) );
  AOI21_X1 U11648 ( .B1(n11054), .B2(n11053), .A(n11052), .ZN(n11055) );
  OAI21_X1 U11649 ( .B1(n10596), .B2(n11056), .A(n11055), .ZN(P1_U3288) );
  INV_X1 U11650 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U11651 ( .A1(n11108), .A2(n11058), .B1(n11057), .B2(n11105), .ZN(
        P2_U3408) );
  INV_X1 U11652 ( .A(n11059), .ZN(n11062) );
  OAI21_X1 U11653 ( .B1(n11062), .B2(n11061), .A(n11060), .ZN(n11068) );
  INV_X1 U11654 ( .A(n11063), .ZN(n11067) );
  AOI222_X1 U11655 ( .A1(n11069), .A2(n11068), .B1(n11067), .B2(n11066), .C1(
        n11065), .C2(n11064), .ZN(n11070) );
  OAI21_X1 U11656 ( .B1(n11071), .B2(n7771), .A(n11070), .ZN(P2_U3225) );
  OAI21_X1 U11657 ( .B1(n11073), .B2(n11088), .A(n11072), .ZN(n11075) );
  AOI211_X1 U11658 ( .C1(n11091), .C2(n11076), .A(n11075), .B(n11074), .ZN(
        n11078) );
  AOI22_X1 U11659 ( .A1(n11094), .A2(n11078), .B1(n7488), .B2(n11093), .ZN(
        P1_U3531) );
  INV_X1 U11660 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U11661 ( .A1(n11079), .A2(n11078), .B1(n11077), .B2(n11095), .ZN(
        P1_U3480) );
  INV_X1 U11662 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U11663 ( .A1(n11108), .A2(n11081), .B1(n11080), .B2(n11105), .ZN(
        P2_U3420) );
  INV_X1 U11664 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U11665 ( .A1(n11108), .A2(n11083), .B1(n11082), .B2(n11105), .ZN(
        P2_U3423) );
  INV_X1 U11666 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U11667 ( .A1(n11108), .A2(n11085), .B1(n11084), .B2(n11105), .ZN(
        P2_U3426) );
  OAI211_X1 U11668 ( .C1(n11089), .C2(n11088), .A(n11087), .B(n11086), .ZN(
        n11090) );
  AOI21_X1 U11669 ( .B1(n11092), .B2(n11091), .A(n11090), .ZN(n11097) );
  AOI22_X1 U11670 ( .A1(n11094), .A2(n11097), .B1(n7498), .B2(n11093), .ZN(
        P1_U3534) );
  INV_X1 U11671 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U11672 ( .A1(n11079), .A2(n11097), .B1(n11096), .B2(n11095), .ZN(
        P1_U3489) );
  INV_X1 U11673 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U11674 ( .A1(n11108), .A2(n11099), .B1(n11098), .B2(n11105), .ZN(
        P2_U3429) );
  INV_X1 U11675 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U11676 ( .A1(n11108), .A2(n11101), .B1(n11100), .B2(n11105), .ZN(
        P2_U3432) );
  INV_X1 U11677 ( .A(n11102), .ZN(n11104) );
  INV_X1 U11678 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11103) );
  AOI22_X1 U11679 ( .A1(n11108), .A2(n11104), .B1(n11103), .B2(n11105), .ZN(
        P2_U3435) );
  INV_X1 U11680 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U11681 ( .A1(n11108), .A2(n11107), .B1(n11106), .B2(n11105), .ZN(
        P2_U3438) );
  XNOR2_X1 U11682 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X2 U5180 ( .A(n6586), .ZN(n7262) );
  NAND2_X1 U5227 ( .A1(n9244), .A2(n5115), .ZN(n5491) );
  CLKBUF_X1 U5184 ( .A(n5879), .Z(n6127) );
  CLKBUF_X1 U5199 ( .A(n6586), .Z(n6764) );
  CLKBUF_X3 U5211 ( .A(n6519), .Z(n6576) );
  CLKBUF_X2 U5340 ( .A(n5397), .Z(n5114) );
  CLKBUF_X1 U7758 ( .A(n10257), .Z(n5111) );
endmodule

