

module b17_C_AntiSAT_k_128_8 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9631, n9632, n9633, n9634, n9635, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965;

  INV_X1 U11079 ( .A(n17527), .ZN(n17546) );
  INV_X2 U11080 ( .A(n17649), .ZN(n17570) );
  OAI211_X1 U11081 ( .C1(n19969), .C2(n9835), .A(n9834), .B(n13312), .ZN(
        n13311) );
  INV_X2 U11082 ( .A(n10476), .ZN(n10556) );
  INV_X2 U11083 ( .A(n18114), .ZN(n17197) );
  INV_X1 U11084 ( .A(n15462), .ZN(n13427) );
  INV_X4 U11085 ( .A(n13971), .ZN(n17066) );
  CLKBUF_X1 U11086 ( .A(n10729), .Z(n10854) );
  CLKBUF_X3 U11087 ( .A(n15521), .Z(n9633) );
  AND2_X1 U11088 ( .A1(n13220), .A2(n10588), .ZN(n12432) );
  AND2_X2 U11089 ( .A1(n12443), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10627) );
  INV_X1 U11091 ( .A(n12954), .ZN(n20756) );
  AND2_X2 U11092 ( .A1(n12575), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10647) );
  CLKBUF_X2 U11093 ( .A(n12554), .Z(n12548) );
  INV_X2 U11094 ( .A(n11205), .ZN(n11817) );
  BUF_X1 U11095 ( .A(n10564), .Z(n9647) );
  BUF_X1 U11096 ( .A(n10412), .Z(n12312) );
  OR2_X1 U11098 ( .A1(n10919), .A2(n10918), .ZN(n20022) );
  AND2_X1 U11099 ( .A1(n10903), .A2(n12928), .ZN(n11070) );
  CLKBUF_X2 U11100 ( .A(n10339), .Z(n9646) );
  INV_X2 U11101 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13075) );
  OR2_X1 U11105 ( .A1(n10464), .A2(n10456), .ZN(n10458) );
  CLKBUF_X3 U11106 ( .A(n10361), .Z(n12581) );
  AND2_X1 U11107 ( .A1(n10420), .A2(n10431), .ZN(n12593) );
  INV_X1 U11108 ( .A(n15537), .ZN(n16832) );
  INV_X1 U11109 ( .A(n9633), .ZN(n16903) );
  AOI22_X1 U11110 ( .A1(n20940), .A2(keyinput31), .B1(keyinput10), .B2(n20939), 
        .ZN(n20938) );
  BUF_X1 U11111 ( .A(n11032), .Z(n12929) );
  AND2_X2 U11112 ( .A1(n10929), .A2(n10243), .ZN(n11033) );
  NAND2_X1 U11113 ( .A1(n12991), .A2(n11126), .ZN(n11168) );
  OR2_X1 U11114 ( .A1(n10909), .A2(n10908), .ZN(n20018) );
  NOR2_X1 U11115 ( .A1(n10249), .A2(n10281), .ZN(n10247) );
  NAND2_X1 U11116 ( .A1(n12186), .A2(n12118), .ZN(n12113) );
  NOR2_X1 U11117 ( .A1(n12089), .A2(n12088), .ZN(n12100) );
  INV_X1 U11118 ( .A(n12270), .ZN(n12170) );
  INV_X1 U11119 ( .A(n15043), .ZN(n12025) );
  BUF_X1 U11120 ( .A(n11909), .Z(n9652) );
  AND2_X1 U11121 ( .A1(n10004), .A2(n11918), .ZN(n11965) );
  NOR2_X2 U11122 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13876) );
  OAI221_X1 U11123 ( .B1(n20940), .B2(keyinput31), .C1(n20939), .C2(keyinput10), .A(n20938), .ZN(n20953) );
  NAND2_X1 U11124 ( .A1(n20014), .A2(n20022), .ZN(n12870) );
  AND4_X1 U11125 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n12774) );
  XNOR2_X1 U11126 ( .A(n11168), .B(n19978), .ZN(n12988) );
  INV_X1 U11127 ( .A(n12312), .ZN(n12229) );
  INV_X1 U11128 ( .A(n10399), .ZN(n12617) );
  NAND2_X1 U11129 ( .A1(n12121), .A2(n15408), .ZN(n15188) );
  INV_X1 U11130 ( .A(n16764), .ZN(n16734) );
  NAND2_X1 U11131 ( .A1(n16292), .A2(n15567), .ZN(n17648) );
  INV_X1 U11132 ( .A(n18539), .ZN(n18552) );
  INV_X1 U11133 ( .A(n18085), .ZN(n18732) );
  INV_X1 U11134 ( .A(n19826), .ZN(n19837) );
  OAI21_X1 U11135 ( .B1(n11377), .B2(n11308), .A(n11123), .ZN(n12944) );
  INV_X1 U11137 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19731) );
  BUF_X1 U11138 ( .A(n10399), .Z(n13386) );
  INV_X1 U11139 ( .A(n19737), .ZN(n10635) );
  NOR2_X1 U11140 ( .A1(n18575), .A2(n16427), .ZN(n16778) );
  NAND2_X1 U11141 ( .A1(n17576), .A2(n17483), .ZN(n17737) );
  INV_X1 U11142 ( .A(n18045), .ZN(n18509) );
  INV_X1 U11143 ( .A(n13382), .ZN(n13380) );
  INV_X1 U11144 ( .A(n19797), .ZN(n15842) );
  INV_X2 U11145 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18702) );
  AND2_X1 U11146 ( .A1(n10146), .A2(n10145), .ZN(n9631) );
  NOR2_X2 U11147 ( .A1(n10258), .A2(n15115), .ZN(n10257) );
  AND2_X2 U11150 ( .A1(n10212), .A2(n10211), .ZN(n14104) );
  INV_X2 U11151 ( .A(n17745), .ZN(n17716) );
  OAI21_X2 U11152 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18726), .A(n16406), 
        .ZN(n17745) );
  NOR2_X2 U11153 ( .A1(n10410), .A2(n12047), .ZN(n13268) );
  INV_X2 U11154 ( .A(n12222), .ZN(n10410) );
  XNOR2_X2 U11155 ( .A(n12020), .B(n12024), .ZN(n12087) );
  AND2_X1 U11156 ( .A1(n10898), .A2(n10900), .ZN(n9632) );
  AND2_X1 U11157 ( .A1(n10898), .A2(n10900), .ZN(n11616) );
  NOR4_X4 U11158 ( .A1(n17189), .A2(n17319), .A3(n17317), .A4(n17114), .ZN(
        n17154) );
  NAND2_X2 U11159 ( .A1(n10299), .A2(n10298), .ZN(n10613) );
  AND2_X1 U11160 ( .A1(n11911), .A2(n11917), .ZN(n19464) );
  NOR2_X1 U11161 ( .A1(n18685), .A2(n13873), .ZN(n15521) );
  CLKBUF_X1 U11162 ( .A(n12443), .Z(n9634) );
  NAND2_X1 U11163 ( .A1(n14913), .A2(n14912), .ZN(n14911) );
  NOR2_X2 U11164 ( .A1(n15167), .A2(n15166), .ZN(n15385) );
  OR2_X1 U11166 ( .A1(n9842), .A2(n9635), .ZN(n9799) );
  NOR2_X1 U11167 ( .A1(n19475), .A2(n19474), .ZN(n19545) );
  NOR2_X1 U11168 ( .A1(n19435), .A2(n19208), .ZN(n19429) );
  INV_X2 U11169 ( .A(n19850), .ZN(n19833) );
  INV_X2 U11170 ( .A(n17737), .ZN(n17729) );
  INV_X2 U11171 ( .A(n14788), .ZN(n14628) );
  INV_X4 U11172 ( .A(n11289), .ZN(n14788) );
  NAND2_X1 U11173 ( .A1(n17231), .A2(n17734), .ZN(n17649) );
  AND2_X1 U11174 ( .A1(n11916), .A2(n11918), .ZN(n13447) );
  NOR2_X1 U11175 ( .A1(n12176), .A2(n12174), .ZN(n12179) );
  AND2_X1 U11176 ( .A1(n9651), .A2(n9877), .ZN(n11919) );
  AND2_X1 U11177 ( .A1(n17627), .A2(n9751), .ZN(n17547) );
  NAND2_X2 U11178 ( .A1(n18552), .A2(n18537), .ZN(n17972) );
  CLKBUF_X2 U11179 ( .A(n11377), .Z(n9650) );
  NOR2_X2 U11180 ( .A1(n15634), .A2(n18522), .ZN(n18530) );
  NOR2_X1 U11181 ( .A1(n11651), .A2(n20839), .ZN(n11671) );
  AOI21_X1 U11182 ( .B1(n14001), .B2(n18732), .A(n16421), .ZN(n18526) );
  NAND2_X1 U11183 ( .A1(n16752), .A2(n18114), .ZN(n13998) );
  NAND3_X1 U11184 ( .A1(n9686), .A2(n10665), .A3(n10077), .ZN(n11929) );
  AND2_X1 U11185 ( .A1(n20029), .A2(n13021), .ZN(n12780) );
  CLKBUF_X2 U11186 ( .A(n12774), .Z(n14122) );
  NOR2_X1 U11187 ( .A1(n20018), .A2(n20022), .ZN(n13277) );
  INV_X2 U11188 ( .A(n13021), .ZN(n11112) );
  NAND2_X1 U11189 ( .A1(n10269), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10266) );
  AND4_X2 U11190 ( .A1(n10948), .A2(n10946), .A3(n10947), .A4(n10225), .ZN(
        n13021) );
  INV_X4 U11191 ( .A(n16832), .ZN(n17068) );
  AND4_X1 U11192 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10948) );
  AND4_X1 U11193 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10947) );
  BUF_X2 U11194 ( .A(n12576), .Z(n12568) );
  CLKBUF_X3 U11195 ( .A(n10979), .Z(n11659) );
  CLKBUF_X3 U11196 ( .A(n14055), .Z(n9638) );
  AND2_X1 U11197 ( .A1(n9778), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10902) );
  AND2_X1 U11198 ( .A1(n15037), .A2(n19056), .ZN(n9661) );
  NAND2_X1 U11199 ( .A1(n15040), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15041) );
  OAI21_X1 U11200 ( .B1(n15134), .B2(n15112), .A(n15111), .ZN(n15123) );
  AND2_X1 U11201 ( .A1(n10206), .A2(n10205), .ZN(n15023) );
  NAND2_X1 U11202 ( .A1(n15147), .A2(n15144), .ZN(n15134) );
  XNOR2_X1 U11203 ( .A(n14556), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9953) );
  OR2_X1 U11204 ( .A1(n14106), .A2(n9663), .ZN(n14107) );
  NAND2_X1 U11205 ( .A1(n14911), .A2(n12520), .ZN(n9775) );
  NAND2_X1 U11206 ( .A1(n15186), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15389) );
  OR2_X1 U11207 ( .A1(n15046), .A2(n15045), .ZN(n10239) );
  NAND2_X1 U11208 ( .A1(n9769), .A2(n15176), .ZN(n15167) );
  AND2_X1 U11209 ( .A1(n14553), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14564) );
  NOR2_X1 U11210 ( .A1(n14293), .A2(n10119), .ZN(n14259) );
  NAND2_X1 U11211 ( .A1(n9770), .A2(n9724), .ZN(n9769) );
  NAND2_X1 U11212 ( .A1(n15187), .A2(n9767), .ZN(n9770) );
  NAND2_X1 U11213 ( .A1(n9997), .A2(n14788), .ZN(n14580) );
  AOI211_X1 U11214 ( .C1(n15204), .C2(n16200), .A(n15203), .B(n15202), .ZN(
        n15207) );
  NAND2_X1 U11215 ( .A1(n14595), .A2(n9753), .ZN(n9997) );
  NAND2_X1 U11216 ( .A1(n9801), .A2(n9684), .ZN(n13721) );
  NAND2_X1 U11217 ( .A1(n14414), .A2(n14413), .ZN(n14586) );
  NAND2_X1 U11218 ( .A1(n17386), .A2(n17385), .ZN(n17384) );
  OAI21_X1 U11219 ( .B1(n9845), .B2(n14223), .A(n9843), .ZN(n14619) );
  XNOR2_X1 U11220 ( .A(n12616), .B(n10857), .ZN(n18939) );
  NAND2_X1 U11221 ( .A1(n9772), .A2(n9828), .ZN(n9771) );
  AND2_X1 U11222 ( .A1(n14341), .A2(n14342), .ZN(n14414) );
  NAND2_X1 U11223 ( .A1(n14215), .A2(n14214), .ZN(n14964) );
  NAND2_X1 U11224 ( .A1(n13710), .A2(n10114), .ZN(n14620) );
  AND2_X1 U11225 ( .A1(n9852), .A2(n9851), .ZN(n16290) );
  NAND2_X1 U11226 ( .A1(n11999), .A2(n13690), .ZN(n10145) );
  NAND2_X1 U11227 ( .A1(n9849), .A2(n11272), .ZN(n13667) );
  INV_X1 U11228 ( .A(n12019), .ZN(n13687) );
  NAND2_X1 U11229 ( .A1(n11981), .A2(n13691), .ZN(n9905) );
  AND2_X1 U11230 ( .A1(n9813), .A2(n14628), .ZN(n9845) );
  AOI21_X1 U11231 ( .B1(n9894), .B2(n9823), .A(n9722), .ZN(n9822) );
  NAND2_X1 U11232 ( .A1(n14988), .A2(n14987), .ZN(n14990) );
  AOI21_X1 U11233 ( .B1(n15871), .B2(n14629), .A(n11299), .ZN(n14630) );
  NOR2_X1 U11234 ( .A1(n9895), .A2(n9657), .ZN(n9894) );
  NAND2_X1 U11235 ( .A1(n10151), .A2(n10150), .ZN(n15002) );
  NOR2_X1 U11236 ( .A1(n9807), .A2(n9796), .ZN(n14789) );
  AND3_X1 U11237 ( .A1(n9870), .A2(n17475), .A3(n9674), .ZN(n15616) );
  AND2_X1 U11238 ( .A1(n11980), .A2(n11979), .ZN(n12000) );
  INV_X1 U11239 ( .A(n15301), .ZN(n10151) );
  INV_X1 U11240 ( .A(n12960), .ZN(n12351) );
  NAND2_X1 U11241 ( .A1(n15298), .A2(n15299), .ZN(n15301) );
  INV_X1 U11242 ( .A(n9843), .ZN(n9635) );
  NAND2_X1 U11243 ( .A1(n16011), .A2(n12186), .ZN(n12191) );
  AND4_X1 U11244 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11927) );
  NOR2_X1 U11245 ( .A1(n13578), .A2(n11428), .ZN(n10111) );
  INV_X1 U11246 ( .A(n13834), .ZN(n15298) );
  OR2_X1 U11247 ( .A1(n13534), .A2(n13580), .ZN(n13578) );
  OAI21_X1 U11248 ( .B1(n17741), .B2(n17483), .A(n18427), .ZN(n17588) );
  AND2_X1 U11249 ( .A1(n15320), .A2(n15319), .ZN(n15322) );
  CLKBUF_X1 U11250 ( .A(n13715), .Z(n15865) );
  CLKBUF_X1 U11251 ( .A(n13714), .Z(n15866) );
  AOI21_X1 U11252 ( .B1(n17541), .B2(n17436), .A(n15610), .ZN(n15611) );
  OR2_X1 U11253 ( .A1(n12345), .A2(n12344), .ZN(n12346) );
  NOR2_X2 U11254 ( .A1(n11925), .A2(n11918), .ZN(n19433) );
  OR2_X1 U11255 ( .A1(n12159), .A2(n15335), .ZN(n15121) );
  AND2_X1 U11256 ( .A1(n11912), .A2(n11919), .ZN(n11959) );
  NAND2_X1 U11257 ( .A1(n9795), .A2(n19999), .ZN(n11285) );
  NAND2_X1 U11258 ( .A1(n12343), .A2(n12342), .ZN(n12345) );
  NOR2_X1 U11259 ( .A1(n20034), .A2(n20154), .ZN(n20552) );
  OR2_X1 U11260 ( .A1(n18798), .A2(n12025), .ZN(n12159) );
  NOR2_X1 U11261 ( .A1(n11202), .A2(n9728), .ZN(n9795) );
  INV_X1 U11262 ( .A(n11202), .ZN(n11203) );
  CLKBUF_X1 U11263 ( .A(n11364), .Z(n20292) );
  NOR2_X1 U11264 ( .A1(n20019), .A2(n20154), .ZN(n20532) );
  NOR2_X1 U11265 ( .A1(n20026), .A2(n20154), .ZN(n20542) );
  NOR2_X1 U11266 ( .A1(n20042), .A2(n20154), .ZN(n20558) );
  NOR2_X1 U11267 ( .A1(n20007), .A2(n20154), .ZN(n20513) );
  NOR2_X1 U11268 ( .A1(n20023), .A2(n20154), .ZN(n20537) );
  NOR2_X2 U11269 ( .A1(n19926), .A2(n13019), .ZN(n19916) );
  OR3_X1 U11270 ( .A1(n18803), .A2(n12025), .A3(n15349), .ZN(n15135) );
  XNOR2_X1 U11271 ( .A(n10001), .B(n11152), .ZN(n11171) );
  NAND2_X1 U11272 ( .A1(n13100), .A2(n13101), .ZN(n13467) );
  XNOR2_X1 U11273 ( .A(n12943), .B(n11124), .ZN(n12992) );
  NAND2_X1 U11274 ( .A1(n12944), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12943) );
  OAI21_X1 U11275 ( .B1(n11371), .B2(n11372), .A(n11162), .ZN(n11170) );
  OR2_X1 U11276 ( .A1(n11722), .A2(n14322), .ZN(n11764) );
  OR2_X1 U11277 ( .A1(n12146), .A2(n10876), .ZN(n12153) );
  NAND2_X1 U11278 ( .A1(n9808), .A2(n9811), .ZN(n20727) );
  NAND2_X1 U11279 ( .A1(n12329), .A2(n12328), .ZN(n15475) );
  NOR2_X1 U11280 ( .A1(n18795), .A2(n18796), .ZN(n18794) );
  OR2_X1 U11281 ( .A1(n11161), .A2(n11160), .ZN(n11162) );
  NAND2_X1 U11282 ( .A1(n9790), .A2(n10000), .ZN(n9999) );
  CLKBUF_X1 U11283 ( .A(n12927), .Z(n20433) );
  XNOR2_X1 U11284 ( .A(n11161), .B(n11160), .ZN(n11371) );
  NAND2_X1 U11285 ( .A1(n11154), .A2(n11153), .ZN(n11161) );
  NOR2_X1 U11286 ( .A1(n15012), .A2(n19469), .ZN(n19588) );
  NAND2_X1 U11287 ( .A1(n11140), .A2(n11139), .ZN(n9998) );
  NOR2_X1 U11288 ( .A1(n13837), .A2(n19469), .ZN(n19573) );
  NOR2_X1 U11289 ( .A1(n18993), .A2(n19469), .ZN(n19467) );
  NOR2_X1 U11290 ( .A1(n18982), .A2(n19469), .ZN(n19552) );
  NOR2_X1 U11291 ( .A1(n18975), .A2(n19469), .ZN(n19485) );
  NAND2_X1 U11292 ( .A1(n11060), .A2(n11061), .ZN(n20047) );
  NAND2_X1 U11293 ( .A1(n11120), .A2(n11119), .ZN(n11154) );
  NAND2_X1 U11294 ( .A1(n11111), .A2(n11110), .ZN(n11120) );
  XNOR2_X1 U11295 ( .A(n11127), .B(n9787), .ZN(n20110) );
  NAND2_X1 U11296 ( .A1(n9782), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11127) );
  AND2_X1 U11297 ( .A1(n11094), .A2(n11092), .ZN(n11062) );
  NAND2_X1 U11298 ( .A1(n10403), .A2(n10443), .ZN(n10470) );
  OR2_X1 U11299 ( .A1(n11136), .A2(n12918), .ZN(n11138) );
  NAND2_X2 U11300 ( .A1(n17305), .A2(n17304), .ZN(n17353) );
  AND3_X1 U11301 ( .A1(n10469), .A2(n10468), .A3(n10467), .ZN(n10473) );
  AND3_X1 U11302 ( .A1(n10446), .A2(n10445), .A3(n10444), .ZN(n10453) );
  NOR3_X1 U11303 ( .A1(n13017), .A2(n11058), .A3(n13022), .ZN(n11059) );
  INV_X1 U11304 ( .A(n12075), .ZN(n10099) );
  NOR2_X1 U11305 ( .A1(n12074), .A2(n12065), .ZN(n10096) );
  BUF_X2 U11306 ( .A(n10464), .Z(n10561) );
  OR2_X1 U11307 ( .A1(n12266), .A2(n12249), .ZN(n10443) );
  XNOR2_X1 U11308 ( .A(n10638), .B(n10619), .ZN(n13182) );
  AND2_X1 U11309 ( .A1(n13184), .A2(n13183), .ZN(n10638) );
  AND2_X1 U11310 ( .A1(n10250), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10251) );
  NAND2_X1 U11311 ( .A1(n10076), .A2(n10075), .ZN(n12043) );
  NAND2_X1 U11312 ( .A1(n10401), .A2(n9794), .ZN(n12313) );
  OR3_X2 U11313 ( .A1(n10255), .A2(n10020), .A3(n10019), .ZN(n9679) );
  NAND2_X1 U11314 ( .A1(n9805), .A2(n13713), .ZN(n11035) );
  AND2_X1 U11315 ( .A1(n10374), .A2(n10413), .ZN(n10376) );
  OR2_X2 U11316 ( .A1(n12597), .A2(n10614), .ZN(n10853) );
  OR2_X1 U11317 ( .A1(n11048), .A2(n11026), .ZN(n12889) );
  NOR2_X1 U11318 ( .A1(n11986), .A2(n12312), .ZN(n10862) );
  NOR2_X1 U11319 ( .A1(n17248), .A2(n15586), .ZN(n15568) );
  OR2_X1 U11320 ( .A1(n11040), .A2(n12870), .ZN(n13030) );
  XOR2_X1 U11321 ( .A(n15569), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17735) );
  NAND2_X1 U11322 ( .A1(n11025), .A2(n20039), .ZN(n11048) );
  NAND4_X2 U11323 ( .A1(n13895), .A2(n13894), .A3(n13893), .A4(n13892), .ZN(
        n18114) );
  AND2_X1 U11324 ( .A1(n11112), .A2(n20039), .ZN(n11027) );
  INV_X1 U11325 ( .A(n17115), .ZN(n18109) );
  NAND2_X1 U11326 ( .A1(n20033), .A2(n20039), .ZN(n13713) );
  AND2_X1 U11327 ( .A1(n13021), .A2(n11324), .ZN(n12874) );
  NAND4_X2 U11328 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n15043) );
  AND2_X1 U11329 ( .A1(n9793), .A2(n10373), .ZN(n10405) );
  INV_X1 U11330 ( .A(n12318), .ZN(n10373) );
  INV_X2 U11331 ( .A(U212), .ZN(n16360) );
  CLKBUF_X3 U11332 ( .A(n10587), .Z(n19737) );
  INV_X1 U11333 ( .A(n20029), .ZN(n11324) );
  INV_X2 U11334 ( .A(n20014), .ZN(n13019) );
  INV_X1 U11335 ( .A(n20039), .ZN(n14461) );
  CLKBUF_X1 U11336 ( .A(n12318), .Z(n13408) );
  OR2_X2 U11337 ( .A1(n16361), .A2(n16302), .ZN(n16363) );
  OR2_X2 U11338 ( .A1(n11002), .A2(n11001), .ZN(n20039) );
  NAND2_X1 U11339 ( .A1(n10325), .A2(n10324), .ZN(n12318) );
  NAND2_X1 U11340 ( .A1(n10336), .A2(n10335), .ZN(n10399) );
  AND4_X1 U11341 ( .A1(n10983), .A2(n10982), .A3(n10981), .A4(n10980), .ZN(
        n10990) );
  AND4_X1 U11342 ( .A1(n10973), .A2(n10972), .A3(n10971), .A4(n10970), .ZN(
        n10992) );
  NOR2_X1 U11343 ( .A1(n9696), .A2(n10226), .ZN(n10225) );
  AND4_X1 U11344 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10389) );
  AND4_X1 U11345 ( .A1(n10978), .A2(n10977), .A3(n10976), .A4(n10975), .ZN(
        n10991) );
  AND4_X1 U11346 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11020) );
  AND4_X1 U11347 ( .A1(n11015), .A2(n11014), .A3(n11013), .A4(n11012), .ZN(
        n11021) );
  AND4_X1 U11348 ( .A1(n10952), .A2(n10951), .A3(n10950), .A4(n10949), .ZN(
        n10968) );
  AND4_X1 U11349 ( .A1(n10956), .A2(n10955), .A3(n10954), .A4(n10953), .ZN(
        n10967) );
  AND4_X1 U11350 ( .A1(n10964), .A2(n10963), .A3(n10962), .A4(n10961), .ZN(
        n10965) );
  AND4_X1 U11351 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n10946) );
  AND2_X2 U11352 ( .A1(n12548), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10680) );
  AND4_X1 U11353 ( .A1(n10988), .A2(n10987), .A3(n10986), .A4(n10985), .ZN(
        n10989) );
  AND2_X1 U11354 ( .A1(n12443), .A2(n13075), .ZN(n10646) );
  AND4_X1 U11355 ( .A1(n11007), .A2(n11006), .A3(n11005), .A4(n11004), .ZN(
        n11023) );
  AND3_X1 U11356 ( .A1(n10320), .A2(n13075), .A3(n10319), .ZN(n10323) );
  AND4_X1 U11357 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10929) );
  AND2_X2 U11358 ( .A1(n12568), .A2(n13075), .ZN(n10662) );
  AND2_X1 U11359 ( .A1(n10307), .A2(n10306), .ZN(n10308) );
  AND3_X1 U11360 ( .A1(n10293), .A2(n10292), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10294) );
  BUF_X2 U11361 ( .A(n11095), .Z(n11848) );
  BUF_X2 U11362 ( .A(n11063), .Z(n11847) );
  NAND2_X2 U11363 ( .A1(n19744), .A2(n19619), .ZN(n19668) );
  NAND2_X2 U11364 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19744), .ZN(n19669) );
  BUF_X2 U11365 ( .A(n11068), .Z(n11841) );
  AND2_X2 U11366 ( .A1(n9645), .A2(n13075), .ZN(n10663) );
  NAND2_X2 U11368 ( .A1(n18669), .A2(n18609), .ZN(n18657) );
  AND2_X2 U11369 ( .A1(n9639), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10620) );
  INV_X2 U11370 ( .A(n16395), .ZN(U215) );
  BUF_X2 U11371 ( .A(n11070), .Z(n11751) );
  BUF_X2 U11372 ( .A(n10354), .Z(n12569) );
  CLKBUF_X3 U11373 ( .A(n15535), .Z(n16976) );
  BUF_X2 U11374 ( .A(n10339), .Z(n9645) );
  AND2_X2 U11375 ( .A1(n10902), .A2(n10903), .ZN(n11707) );
  INV_X2 U11377 ( .A(n16286), .ZN(n9637) );
  CLKBUF_X3 U11378 ( .A(n15531), .Z(n17067) );
  NAND2_X1 U11379 ( .A1(n18553), .A2(n9814), .ZN(n17043) );
  AND2_X2 U11380 ( .A1(n10901), .A2(n12928), .ZN(n11100) );
  NOR4_X2 U11381 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n18708), .ZN(n15535) );
  AND2_X1 U11382 ( .A1(n18708), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9814) );
  NOR2_X1 U11383 ( .A1(n16117), .A2(n10018), .ZN(n10017) );
  AND3_X1 U11384 ( .A1(n10021), .A2(n10275), .A3(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10274) );
  NAND2_X2 U11385 ( .A1(n20750), .A2(n20757), .ZN(n14113) );
  AND2_X1 U11386 ( .A1(n13221), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13219) );
  AND2_X1 U11387 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10903) );
  INV_X2 U11388 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18685) );
  INV_X2 U11389 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10892) );
  NAND2_X1 U11390 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10287) );
  AND2_X1 U11391 ( .A1(n13219), .A2(n10568), .ZN(n9639) );
  AND2_X2 U11392 ( .A1(n13219), .A2(n10568), .ZN(n12576) );
  NAND3_X1 U11393 ( .A1(n10396), .A2(n9658), .A3(n12280), .ZN(n12283) );
  AND2_X1 U11394 ( .A1(n12568), .A2(n13075), .ZN(n9640) );
  AND2_X1 U11395 ( .A1(n12568), .A2(n13075), .ZN(n9641) );
  NAND3_X2 U11396 ( .A1(n10221), .A2(n10222), .A3(n10219), .ZN(n14222) );
  AND2_X1 U11397 ( .A1(n11900), .A2(n11916), .ZN(n13511) );
  AND2_X4 U11398 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12050) );
  NAND2_X2 U11399 ( .A1(n12882), .A2(n11042), .ZN(n13017) );
  AND2_X2 U11400 ( .A1(n15068), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15040) );
  OAI21_X2 U11401 ( .B1(n12927), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11077), 
        .ZN(n11372) );
  NAND2_X2 U11402 ( .A1(n10428), .A2(n10427), .ZN(n11879) );
  AOI21_X2 U11403 ( .B1(n10470), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10409), .ZN(n10428) );
  NOR2_X2 U11404 ( .A1(n13640), .A2(n10180), .ZN(n13830) );
  NAND2_X2 U11405 ( .A1(n13627), .A2(n13641), .ZN(n13640) );
  AOI21_X2 U11406 ( .B1(n12029), .B2(n20776), .A(n9879), .ZN(n9878) );
  NAND2_X2 U11407 ( .A1(n12028), .A2(n12027), .ZN(n12029) );
  NAND2_X1 U11408 ( .A1(n10242), .A2(n13497), .ZN(n16143) );
  NOR2_X2 U11409 ( .A1(n14620), .A2(n14422), .ZN(n14341) );
  NAND2_X2 U11410 ( .A1(n12351), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13059) );
  AND2_X2 U11411 ( .A1(n9797), .A2(n11957), .ZN(n9680) );
  AOI21_X2 U11412 ( .B1(n15200), .B2(n15041), .A(n15025), .ZN(n15037) );
  BUF_X2 U11413 ( .A(n18908), .Z(n9642) );
  XNOR2_X2 U11414 ( .A(n11222), .B(n11201), .ZN(n19935) );
  NAND2_X2 U11415 ( .A1(n13311), .A2(n11200), .ZN(n11222) );
  NOR2_X1 U11417 ( .A1(n10287), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10339) );
  AND2_X4 U11418 ( .A1(n10899), .A2(n10898), .ZN(n9648) );
  AND2_X1 U11419 ( .A1(n10899), .A2(n10898), .ZN(n9649) );
  AND2_X1 U11420 ( .A1(n10899), .A2(n10898), .ZN(n11660) );
  OAI21_X1 U11421 ( .B1(n11120), .B2(n11119), .A(n11154), .ZN(n11377) );
  BUF_X1 U11422 ( .A(n11909), .Z(n9651) );
  BUF_X2 U11423 ( .A(n11909), .Z(n9653) );
  XNOR2_X1 U11424 ( .A(n11371), .B(n11372), .ZN(n14833) );
  AOI21_X1 U11425 ( .B1(n10455), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10459), .ZN(n10461) );
  AOI21_X1 U11426 ( .B1(n10470), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10454), .ZN(n10460) );
  INV_X1 U11427 ( .A(n13050), .ZN(n12493) );
  OR2_X1 U11428 ( .A1(n15074), .A2(n9889), .ZN(n15042) );
  NAND2_X1 U11429 ( .A1(n10183), .A2(n15067), .ZN(n9889) );
  INV_X1 U11430 ( .A(n15075), .ZN(n10183) );
  AND2_X1 U11431 ( .A1(n15591), .A2(n17235), .ZN(n15567) );
  AND4_X1 U11432 ( .A1(n10715), .A2(n10714), .A3(n10713), .A4(n10712), .ZN(
        n10726) );
  AND4_X1 U11433 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(
        n10724) );
  AND4_X1 U11434 ( .A1(n10711), .A2(n10710), .A3(n10709), .A4(n10708), .ZN(
        n10727) );
  AOI21_X1 U11435 ( .B1(n11958), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A(n9761), .ZN(n12005) );
  INV_X1 U11436 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n9762) );
  AND4_X1 U11437 ( .A1(n12012), .A2(n12011), .A3(n12010), .A4(n12009), .ZN(
        n12013) );
  INV_X1 U11438 ( .A(n14223), .ZN(n9842) );
  NOR2_X1 U11439 ( .A1(n9723), .A2(n11048), .ZN(n12901) );
  AND2_X2 U11440 ( .A1(n10891), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10901) );
  NOR2_X1 U11441 ( .A1(n14330), .A2(n14587), .ZN(n10118) );
  OR2_X1 U11442 ( .A1(n12929), .A2(n20759), .ZN(n11861) );
  XNOR2_X1 U11443 ( .A(n11285), .B(n11275), .ZN(n11448) );
  OAI21_X1 U11444 ( .B1(n11372), .B2(n13019), .A(n11091), .ZN(n11124) );
  NOR2_X2 U11445 ( .A1(n20033), .A2(n20750), .ZN(n11569) );
  NOR2_X1 U11446 ( .A1(n9844), .A2(n9702), .ZN(n9843) );
  NOR2_X1 U11447 ( .A1(n14628), .A2(n11295), .ZN(n9844) );
  NAND2_X1 U11448 ( .A1(n14165), .A2(n14161), .ZN(n14166) );
  NAND2_X1 U11449 ( .A1(n11032), .A2(n20022), .ZN(n11037) );
  INV_X1 U11450 ( .A(n14166), .ZN(n14155) );
  INV_X1 U11451 ( .A(n11088), .ZN(n11159) );
  NAND2_X1 U11452 ( .A1(n20110), .A2(n11062), .ZN(n11132) );
  OR2_X1 U11453 ( .A1(n15086), .A2(n9689), .ZN(n9895) );
  NOR2_X1 U11454 ( .A1(n10074), .A2(n13704), .ZN(n10073) );
  INV_X1 U11455 ( .A(n13661), .ZN(n10074) );
  NAND2_X1 U11456 ( .A1(n13688), .A2(n12019), .ZN(n12021) );
  MUX2_X1 U11457 ( .A(n10415), .B(n10634), .S(n10414), .Z(n10417) );
  NAND2_X1 U11458 ( .A1(n9777), .A2(n12322), .ZN(n12326) );
  NAND2_X1 U11459 ( .A1(n12493), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12332) );
  NAND2_X1 U11460 ( .A1(n10006), .A2(n10005), .ZN(n9886) );
  NAND2_X1 U11461 ( .A1(n9709), .A2(n11880), .ZN(n10006) );
  NAND2_X1 U11462 ( .A1(n10035), .A2(n10034), .ZN(n15723) );
  AND2_X1 U11463 ( .A1(n15670), .A2(n17760), .ZN(n10034) );
  INV_X1 U11464 ( .A(n15619), .ZN(n10035) );
  INV_X1 U11465 ( .A(n9874), .ZN(n9873) );
  NAND2_X1 U11466 ( .A1(n9659), .A2(n17981), .ZN(n9871) );
  OAI21_X1 U11467 ( .B1(n15602), .B2(n9872), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9874) );
  OAI21_X1 U11468 ( .B1(n17656), .B2(n17655), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15662) );
  AOI21_X1 U11469 ( .B1(n14007), .B2(n14006), .A(n14005), .ZN(n16222) );
  NAND2_X1 U11470 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  INV_X1 U11471 ( .A(n14261), .ZN(n10120) );
  NAND2_X1 U11472 ( .A1(n10124), .A2(n10121), .ZN(n14260) );
  NAND2_X1 U11473 ( .A1(n20727), .A2(n20759), .ZN(n11192) );
  OR2_X1 U11474 ( .A1(n11351), .A2(n11318), .ZN(n11363) );
  NAND2_X1 U11475 ( .A1(n10572), .A2(n10574), .ZN(n12248) );
  OR2_X1 U11476 ( .A1(n10575), .A2(n10571), .ZN(n10572) );
  AND2_X1 U11477 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15738), .ZN(
        n10571) );
  AND2_X1 U11478 ( .A1(n10405), .A2(n12270), .ZN(n9794) );
  NAND2_X1 U11479 ( .A1(n10102), .A2(n10101), .ZN(n12171) );
  INV_X1 U11480 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10101) );
  NAND2_X1 U11481 ( .A1(n12356), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10176) );
  AND2_X1 U11482 ( .A1(n13562), .A2(n13415), .ZN(n12356) );
  AND2_X1 U11483 ( .A1(n10635), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12323) );
  OR2_X1 U11484 ( .A1(n18983), .A2(n12620), .ZN(n12815) );
  INV_X1 U11485 ( .A(n10405), .ZN(n12620) );
  NOR2_X1 U11486 ( .A1(n9752), .A2(n15227), .ZN(n10147) );
  NAND2_X1 U11487 ( .A1(n9687), .A2(n10207), .ZN(n10204) );
  NOR2_X1 U11488 ( .A1(n10200), .A2(n15409), .ZN(n10199) );
  INV_X1 U11489 ( .A(n9828), .ZN(n9773) );
  OR2_X1 U11490 ( .A1(n18786), .A2(n12158), .ZN(n15105) );
  NAND2_X1 U11491 ( .A1(n15373), .A2(n9915), .ZN(n15139) );
  NOR2_X1 U11492 ( .A1(n15358), .A2(n9918), .ZN(n9915) );
  NAND2_X1 U11493 ( .A1(n11998), .A2(n13475), .ZN(n10146) );
  AOI21_X1 U11494 ( .B1(n15462), .B2(n12337), .A(n12331), .ZN(n12767) );
  XNOR2_X1 U11495 ( .A(n15475), .B(n12332), .ZN(n12769) );
  AND2_X1 U11496 ( .A1(n13371), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12337) );
  INV_X1 U11497 ( .A(n19516), .ZN(n19469) );
  AND2_X1 U11498 ( .A1(n9920), .A2(n9736), .ZN(n16522) );
  OR2_X1 U11499 ( .A1(n16764), .A2(n16539), .ZN(n9921) );
  INV_X1 U11500 ( .A(n18104), .ZN(n17118) );
  NAND2_X1 U11501 ( .A1(n17602), .A2(n17915), .ZN(n17917) );
  INV_X1 U11502 ( .A(n9857), .ZN(n9856) );
  NAND2_X1 U11503 ( .A1(n9860), .A2(n15593), .ZN(n9859) );
  OR2_X1 U11504 ( .A1(n20029), .A2(n11033), .ZN(n11025) );
  AND2_X1 U11505 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n9980)
         );
  CLKBUF_X1 U11506 ( .A(n11707), .Z(n11822) );
  OR2_X1 U11508 ( .A1(n11108), .A2(n11107), .ZN(n11291) );
  OR2_X1 U11509 ( .A1(n11150), .A2(n11149), .ZN(n11151) );
  INV_X1 U11510 ( .A(n11151), .ZN(n11193) );
  INV_X1 U11511 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U11512 ( .A1(n12000), .A2(n9887), .ZN(n12024) );
  INV_X1 U11513 ( .A(n12020), .ZN(n12023) );
  NAND2_X1 U11514 ( .A1(n12261), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10408) );
  NOR2_X1 U11515 ( .A1(n17240), .A2(n15589), .ZN(n15591) );
  OR3_X1 U11516 ( .A1(n11319), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n19995), .ZN(n12738) );
  NOR2_X1 U11517 ( .A1(n14271), .A2(n14285), .ZN(n10122) );
  INV_X1 U11518 ( .A(n11861), .ZN(n11829) );
  AND2_X1 U11519 ( .A1(n14317), .A2(n10118), .ZN(n10117) );
  AND2_X1 U11520 ( .A1(n11577), .A2(n14429), .ZN(n13711) );
  AOI21_X1 U11521 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n9993), .ZN(n11471) );
  AND2_X1 U11522 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n9993)
         );
  AND2_X1 U11523 ( .A1(n9743), .A2(n10133), .ZN(n10132) );
  INV_X1 U11524 ( .A(n14415), .ZN(n10133) );
  INV_X1 U11525 ( .A(n9962), .ZN(n9961) );
  NOR2_X1 U11526 ( .A1(n14619), .A2(n11302), .ZN(n14595) );
  INV_X1 U11527 ( .A(n9964), .ZN(n9963) );
  OAI211_X1 U11528 ( .C1(n9800), .C2(n9635), .A(n9799), .B(n14618), .ZN(n14593) );
  INV_X1 U11529 ( .A(n9845), .ZN(n9800) );
  AND2_X1 U11530 ( .A1(n15872), .A2(n15876), .ZN(n14629) );
  NAND2_X1 U11531 ( .A1(n14789), .A2(n11297), .ZN(n15871) );
  OR2_X1 U11532 ( .A1(n11289), .A2(n15936), .ZN(n15876) );
  AND2_X1 U11533 ( .A1(n9719), .A2(n10144), .ZN(n10143) );
  INV_X1 U11534 ( .A(n14441), .ZN(n10144) );
  INV_X1 U11535 ( .A(n9960), .ZN(n9959) );
  NAND2_X1 U11536 ( .A1(n10003), .A2(n10002), .ZN(n10224) );
  NAND2_X1 U11537 ( .A1(n13547), .A2(n10137), .ZN(n10138) );
  INV_X1 U11538 ( .A(n10139), .ZN(n10137) );
  INV_X1 U11539 ( .A(n15916), .ZN(n10214) );
  NAND2_X1 U11540 ( .A1(n19969), .A2(n11169), .ZN(n11199) );
  INV_X1 U11541 ( .A(n9958), .ZN(n9957) );
  NAND2_X1 U11542 ( .A1(n10141), .A2(n10140), .ZN(n10139) );
  INV_X1 U11543 ( .A(n19816), .ZN(n10140) );
  INV_X1 U11544 ( .A(n13096), .ZN(n10141) );
  AND2_X1 U11545 ( .A1(n12987), .A2(n13088), .ZN(n9837) );
  INV_X1 U11546 ( .A(n11169), .ZN(n9841) );
  NOR2_X2 U11547 ( .A1(n14168), .A2(n14161), .ZN(n14163) );
  AND2_X1 U11548 ( .A1(n12890), .A2(n12897), .ZN(n13010) );
  NAND2_X2 U11549 ( .A1(n9956), .A2(n9955), .ZN(n9968) );
  INV_X1 U11550 ( .A(n20022), .ZN(n9955) );
  OR2_X1 U11551 ( .A1(n11087), .A2(n11086), .ZN(n11121) );
  NOR2_X1 U11552 ( .A1(n14122), .A2(n20759), .ZN(n11113) );
  NAND2_X1 U11553 ( .A1(n10217), .A2(n10215), .ZN(n11094) );
  NOR2_X1 U11554 ( .A1(n12914), .A2(n9786), .ZN(n10218) );
  NAND2_X1 U11555 ( .A1(n13021), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11178) );
  NAND2_X1 U11556 ( .A1(n11178), .A2(n11177), .ZN(n11331) );
  INV_X1 U11557 ( .A(n11356), .ZN(n11354) );
  OR2_X1 U11558 ( .A1(n11040), .A2(n9956), .ZN(n11041) );
  NAND2_X1 U11559 ( .A1(n11043), .A2(n9785), .ZN(n9784) );
  INV_X1 U11560 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20351) );
  AND3_X1 U11561 ( .A1(n13383), .A2(n10375), .A3(n10414), .ZN(n10401) );
  NAND2_X1 U11562 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10020) );
  AOI211_X1 U11563 ( .C1(n12535), .C2(n12533), .A(n13050), .B(n14898), .ZN(
        n12534) );
  OR2_X1 U11564 ( .A1(n10172), .A2(n10170), .ZN(n10169) );
  INV_X1 U11565 ( .A(n12650), .ZN(n10170) );
  INV_X1 U11566 ( .A(n13324), .ZN(n10154) );
  AND4_X1 U11567 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n10725) );
  NAND2_X1 U11568 ( .A1(n10051), .A2(n14853), .ZN(n10050) );
  INV_X1 U11569 ( .A(n14211), .ZN(n10051) );
  NAND2_X1 U11570 ( .A1(n9888), .A2(n12194), .ZN(n12198) );
  NAND2_X1 U11571 ( .A1(n15042), .A2(n15227), .ZN(n9888) );
  INV_X1 U11572 ( .A(n9826), .ZN(n9823) );
  NAND2_X1 U11573 ( .A1(n10068), .A2(n14930), .ZN(n10067) );
  INV_X1 U11574 ( .A(n14939), .ZN(n10068) );
  INV_X1 U11575 ( .A(n13773), .ZN(n10072) );
  NAND2_X1 U11576 ( .A1(n10173), .A2(n12660), .ZN(n10172) );
  INV_X1 U11577 ( .A(n13617), .ZN(n10173) );
  INV_X1 U11578 ( .A(n13466), .ZN(n10171) );
  OR2_X1 U11579 ( .A1(n13465), .A2(n12025), .ZN(n12120) );
  OR2_X1 U11580 ( .A1(n16126), .A2(n9910), .ZN(n9909) );
  NAND2_X1 U11581 ( .A1(n9792), .A2(n9791), .ZN(n9907) );
  AND2_X1 U11582 ( .A1(n12029), .A2(n12033), .ZN(n9791) );
  NAND2_X1 U11583 ( .A1(n10060), .A2(n13364), .ZN(n10059) );
  INV_X1 U11584 ( .A(n10061), .ZN(n10060) );
  INV_X1 U11585 ( .A(n16126), .ZN(n9879) );
  OR2_X1 U11586 ( .A1(n10614), .A2(n12170), .ZN(n10831) );
  AOI21_X1 U11587 ( .B1(n12813), .B2(n9677), .A(n10165), .ZN(n10164) );
  INV_X1 U11588 ( .A(n12818), .ZN(n10165) );
  INV_X1 U11589 ( .A(n10185), .ZN(n10184) );
  OAI21_X1 U11590 ( .B1(n13490), .B2(n10188), .A(n10186), .ZN(n10185) );
  AOI21_X1 U11591 ( .B1(n10192), .B2(n10187), .A(n9731), .ZN(n10186) );
  INV_X1 U11592 ( .A(n10192), .ZN(n10188) );
  OR2_X1 U11593 ( .A1(n10598), .A2(n10597), .ZN(n10868) );
  NAND2_X1 U11594 ( .A1(n13687), .A2(n12023), .ZN(n9803) );
  NAND2_X1 U11595 ( .A1(n10097), .A2(n10099), .ZN(n12083) );
  INV_X1 U11596 ( .A(n12000), .ZN(n10195) );
  NAND2_X1 U11597 ( .A1(n10472), .A2(n10471), .ZN(n10475) );
  INV_X1 U11598 ( .A(n13383), .ZN(n12252) );
  INV_X1 U11599 ( .A(n10831), .ZN(n10818) );
  NAND2_X1 U11600 ( .A1(n10462), .A2(n10463), .ZN(n11880) );
  INV_X1 U11601 ( .A(n12247), .ZN(n12253) );
  INV_X1 U11602 ( .A(n10399), .ZN(n9793) );
  NAND2_X1 U11603 ( .A1(n10004), .A2(n11900), .ZN(n11949) );
  OR2_X1 U11604 ( .A1(n11911), .A2(n13427), .ZN(n11914) );
  NAND2_X1 U11605 ( .A1(n13868), .A2(n13876), .ZN(n13971) );
  NOR3_X1 U11606 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18685), .A3(
        n18523), .ZN(n14055) );
  INV_X1 U11607 ( .A(n18099), .ZN(n14013) );
  NOR2_X1 U11608 ( .A1(n18109), .A2(n13995), .ZN(n13999) );
  AND2_X1 U11609 ( .A1(n17605), .A2(n9671), .ZN(n17535) );
  NAND4_X1 U11610 ( .A1(n9919), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16698) );
  NAND2_X1 U11611 ( .A1(n15618), .A2(n15617), .ZN(n9853) );
  OAI21_X1 U11612 ( .B1(n17568), .B2(n9750), .A(n17648), .ZN(n15608) );
  CLKBUF_X1 U11613 ( .A(n12736), .Z(n12737) );
  NAND2_X1 U11614 ( .A1(n19827), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14173) );
  AOI21_X1 U11615 ( .B1(n14389), .B2(n14165), .A(n13041), .ZN(n13093) );
  INV_X1 U11616 ( .A(n14381), .ZN(n12968) );
  AND2_X1 U11617 ( .A1(n12887), .A2(n12886), .ZN(n12971) );
  OR2_X1 U11618 ( .A1(n11870), .A2(n14264), .ZN(n11871) );
  NAND2_X1 U11619 ( .A1(n11810), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11834) );
  INV_X1 U11620 ( .A(n14294), .ZN(n11770) );
  INV_X1 U11621 ( .A(n14292), .ZN(n11771) );
  NAND2_X1 U11622 ( .A1(n11765), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11808) );
  CLKBUF_X1 U11623 ( .A(n14292), .Z(n14303) );
  OR2_X1 U11624 ( .A1(n14588), .A2(n14113), .ZN(n11674) );
  XNOR2_X1 U11625 ( .A(n14628), .B(n13747), .ZN(n9807) );
  INV_X1 U11626 ( .A(n13590), .ZN(n11414) );
  INV_X1 U11627 ( .A(n12981), .ZN(n11385) );
  AND2_X1 U11628 ( .A1(n14720), .A2(n14333), .ZN(n14331) );
  NAND2_X1 U11629 ( .A1(n14149), .A2(n9965), .ZN(n14150) );
  INV_X1 U11630 ( .A(n9966), .ZN(n9965) );
  NOR2_X1 U11631 ( .A1(n14434), .A2(n13761), .ZN(n14771) );
  OR2_X1 U11632 ( .A1(n15885), .A2(n15884), .ZN(n15887) );
  INV_X1 U11633 ( .A(n10003), .ZN(n11293) );
  INV_X1 U11634 ( .A(n10224), .ZN(n13783) );
  NOR2_X1 U11635 ( .A1(n13585), .A2(n13586), .ZN(n13603) );
  NAND2_X1 U11636 ( .A1(n19935), .A2(n19934), .ZN(n19933) );
  NAND2_X1 U11637 ( .A1(n9836), .A2(n9840), .ZN(n9835) );
  NAND2_X1 U11638 ( .A1(n19969), .A2(n9838), .ZN(n9832) );
  INV_X1 U11639 ( .A(n9839), .ZN(n9838) );
  OR2_X1 U11640 ( .A1(n11136), .A2(n10890), .ZN(n11176) );
  INV_X1 U11641 ( .A(n19750), .ZN(n13012) );
  NAND2_X1 U11642 ( .A1(n20292), .A2(n20151), .ZN(n20259) );
  AND2_X1 U11643 ( .A1(n20293), .A2(n20730), .ZN(n20726) );
  NOR2_X1 U11644 ( .A1(n20001), .A2(n20154), .ZN(n20356) );
  INV_X1 U11645 ( .A(n20294), .ZN(n20429) );
  AOI21_X1 U11646 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20464), .A(n20154), 
        .ZN(n20472) );
  NAND2_X1 U11647 ( .A1(n20759), .A2(n20000), .ZN(n20154) );
  AND2_X1 U11648 ( .A1(n20571), .A2(n20350), .ZN(n20462) );
  OAI22_X1 U11649 ( .A1(n19721), .A2(n12260), .B1(n19718), .B2(n12054), .ZN(
        n12226) );
  NAND2_X1 U11650 ( .A1(n12191), .A2(n16014), .ZN(n16012) );
  AND2_X1 U11651 ( .A1(n12179), .A2(n14932), .ZN(n12188) );
  NAND2_X1 U11652 ( .A1(n12096), .A2(n10109), .ZN(n12108) );
  NOR2_X1 U11653 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13266) );
  AND2_X1 U11654 ( .A1(n13566), .A2(n12647), .ZN(n13662) );
  AND2_X1 U11655 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13415) );
  INV_X1 U11656 ( .A(n10853), .ZN(n10855) );
  AOI21_X1 U11657 ( .B1(n14905), .B2(n14900), .A(n12562), .ZN(n14894) );
  INV_X1 U11658 ( .A(n10177), .ZN(n12460) );
  NAND2_X1 U11659 ( .A1(n9664), .A2(n14954), .ZN(n10180) );
  NOR2_X1 U11660 ( .A1(n10171), .A2(n10169), .ZN(n13643) );
  NAND2_X1 U11661 ( .A1(n10043), .A2(n12318), .ZN(n12596) );
  AND2_X1 U11662 ( .A1(n13248), .A2(n10635), .ZN(n12790) );
  NOR2_X1 U11663 ( .A1(n9676), .A2(n14939), .ZN(n14940) );
  AND3_X1 U11664 ( .A1(n10523), .A2(n10522), .A3(n10521), .ZN(n13862) );
  NAND2_X1 U11665 ( .A1(n13662), .A2(n13661), .ZN(n13705) );
  INV_X1 U11666 ( .A(n10049), .ZN(n10047) );
  NAND2_X1 U11667 ( .A1(n10204), .A2(n10093), .ZN(n9892) );
  AND2_X1 U11668 ( .A1(n15020), .A2(n10095), .ZN(n10093) );
  OR2_X1 U11669 ( .A1(n14852), .A2(n12025), .ZN(n15047) );
  NOR2_X1 U11670 ( .A1(n14917), .A2(n14908), .ZN(n14907) );
  OR2_X1 U11671 ( .A1(n14915), .A2(n14914), .ZN(n14917) );
  AND2_X1 U11672 ( .A1(n9884), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9883) );
  NOR2_X1 U11673 ( .A1(n9899), .A2(n9827), .ZN(n9826) );
  NAND2_X1 U11674 ( .A1(n15097), .A2(n9900), .ZN(n9899) );
  INV_X1 U11675 ( .A(n10196), .ZN(n9900) );
  NOR2_X1 U11676 ( .A1(n9657), .A2(n9689), .ZN(n9893) );
  NOR2_X1 U11677 ( .A1(n9685), .A2(n9904), .ZN(n9903) );
  INV_X1 U11678 ( .A(n15292), .ZN(n9904) );
  NAND2_X1 U11679 ( .A1(n15124), .A2(n15310), .ZN(n15126) );
  NAND2_X1 U11680 ( .A1(n13662), .A2(n10073), .ZN(n13774) );
  INV_X1 U11681 ( .A(n16158), .ZN(n10010) );
  NOR2_X1 U11682 ( .A1(n10172), .A2(n10171), .ZN(n13615) );
  NOR2_X1 U11683 ( .A1(n9704), .A2(n9829), .ZN(n9828) );
  INV_X1 U11684 ( .A(n12106), .ZN(n9829) );
  INV_X1 U11685 ( .A(n15427), .ZN(n10203) );
  NOR2_X1 U11686 ( .A1(n13353), .A2(n13354), .ZN(n13355) );
  NAND2_X1 U11687 ( .A1(n10162), .A2(n10164), .ZN(n13111) );
  AND2_X1 U11688 ( .A1(n10191), .A2(n9720), .ZN(n13681) );
  NAND2_X1 U11689 ( .A1(n10193), .A2(n10192), .ZN(n10191) );
  NAND2_X1 U11690 ( .A1(n11982), .A2(n9680), .ZN(n11996) );
  NOR2_X1 U11691 ( .A1(n10056), .A2(n10053), .ZN(n13057) );
  INV_X1 U11692 ( .A(n10055), .ZN(n10053) );
  NAND2_X1 U11693 ( .A1(n13490), .A2(n12080), .ZN(n10193) );
  AND2_X1 U11694 ( .A1(n12292), .A2(n12291), .ZN(n13725) );
  NAND2_X1 U11695 ( .A1(n11886), .A2(n11887), .ZN(n11885) );
  NOR2_X1 U11696 ( .A1(n10659), .A2(n10156), .ZN(n10155) );
  OR2_X1 U11697 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  AOI21_X1 U11698 ( .B1(n12769), .B2(n12767), .A(n12334), .ZN(n12940) );
  NAND2_X1 U11699 ( .A1(n13045), .A2(n13046), .ZN(n13064) );
  NOR2_X1 U11700 ( .A1(n19697), .A2(n19076), .ZN(n19361) );
  OR2_X1 U11701 ( .A1(n11911), .A2(n11895), .ZN(n11892) );
  INV_X1 U11702 ( .A(n11915), .ZN(n9755) );
  OR2_X1 U11703 ( .A1(n13451), .A2(n19708), .ZN(n19302) );
  NOR2_X2 U11704 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19682) );
  NAND2_X1 U11705 ( .A1(n13451), .A2(n18989), .ZN(n19475) );
  NAND2_X1 U11706 ( .A1(n13451), .A2(n19708), .ZN(n19435) );
  NAND2_X1 U11707 ( .A1(n16215), .A2(n13371), .ZN(n13375) );
  OR2_X1 U11708 ( .A1(n16546), .A2(n9733), .ZN(n9920) );
  OR2_X1 U11709 ( .A1(n16546), .A2(n16547), .ZN(n9922) );
  INV_X1 U11710 ( .A(n18536), .ZN(n15742) );
  NAND2_X1 U11711 ( .A1(n16264), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16236) );
  AND2_X1 U11712 ( .A1(n17495), .A2(n9947), .ZN(n17374) );
  AND2_X1 U11713 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  INV_X1 U11714 ( .A(n16429), .ZN(n9948) );
  INV_X1 U11715 ( .A(n17506), .ZN(n17495) );
  NAND2_X1 U11716 ( .A1(n15599), .A2(n17976), .ZN(n15601) );
  OR2_X1 U11717 ( .A1(n15619), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9851) );
  NAND2_X1 U11718 ( .A1(n15619), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16284) );
  AND2_X1 U11719 ( .A1(n15612), .A2(n9869), .ZN(n9868) );
  NAND2_X1 U11720 ( .A1(n17443), .A2(n17474), .ZN(n17475) );
  NAND2_X1 U11721 ( .A1(n17942), .A2(n17834), .ZN(n9818) );
  NAND2_X1 U11722 ( .A1(n17869), .A2(n9819), .ZN(n17832) );
  AND2_X1 U11723 ( .A1(n17808), .A2(n17809), .ZN(n9819) );
  INV_X1 U11724 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U11725 ( .A1(n17640), .A2(n15664), .ZN(n17602) );
  INV_X1 U11726 ( .A(n15662), .ZN(n15660) );
  NAND2_X1 U11727 ( .A1(n15600), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17937) );
  INV_X1 U11728 ( .A(n15599), .ZN(n15600) );
  NAND2_X1 U11729 ( .A1(n10032), .A2(n9690), .ZN(n9855) );
  AND3_X1 U11730 ( .A1(n9855), .A2(n9856), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17662) );
  OAI21_X1 U11731 ( .B1(n15590), .B2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n17682), .ZN(n17673) );
  OR2_X1 U11732 ( .A1(n17673), .A2(n17672), .ZN(n10032) );
  NOR2_X1 U11733 ( .A1(n17695), .A2(n15588), .ZN(n17683) );
  AND2_X1 U11734 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15587), .ZN(
        n15588) );
  INV_X1 U11735 ( .A(n18041), .ZN(n18515) );
  NOR2_X1 U11736 ( .A1(n12745), .A2(n19750), .ZN(n12746) );
  NAND2_X1 U11737 ( .A1(n14242), .A2(n14243), .ZN(n20752) );
  INV_X1 U11738 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20757) );
  INV_X1 U11739 ( .A(n15909), .ZN(n19943) );
  NAND2_X1 U11740 ( .A1(n12988), .A2(n12987), .ZN(n19969) );
  INV_X1 U11741 ( .A(n19938), .ZN(n19998) );
  AND2_X1 U11742 ( .A1(n15914), .A2(n12945), .ZN(n15909) );
  INV_X1 U11743 ( .A(n19939), .ZN(n15902) );
  INV_X1 U11744 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20464) );
  NAND2_X1 U11745 ( .A1(n9999), .A2(n9998), .ZN(n12915) );
  INV_X1 U11746 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20737) );
  NAND2_X1 U11747 ( .A1(n12124), .A2(n12123), .ZN(n18786) );
  INV_X1 U11748 ( .A(n19697), .ZN(n13554) );
  AND2_X1 U11749 ( .A1(n18966), .A2(n12598), .ZN(n16065) );
  NAND2_X1 U11750 ( .A1(n12595), .A2(n16213), .ZN(n18983) );
  INV_X1 U11751 ( .A(n15389), .ZN(n9788) );
  AND2_X1 U11752 ( .A1(n16151), .A2(n12057), .ZN(n16137) );
  XNOR2_X1 U11753 ( .A(n14210), .B(n9688), .ZN(n15039) );
  INV_X1 U11754 ( .A(n10204), .ZN(n14210) );
  NAND2_X1 U11755 ( .A1(n12314), .A2(n12264), .ZN(n16188) );
  AND2_X1 U11756 ( .A1(n12314), .A2(n19719), .ZN(n19065) );
  INV_X1 U11757 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19705) );
  INV_X1 U11758 ( .A(n13451), .ZN(n19683) );
  INV_X1 U11759 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12703) );
  NOR2_X1 U11760 ( .A1(n18512), .A2(n17303), .ZN(n18746) );
  INV_X1 U11761 ( .A(n16794), .ZN(n9938) );
  NAND2_X1 U11762 ( .A1(n9934), .A2(n9931), .ZN(n9930) );
  INV_X1 U11763 ( .A(n16445), .ZN(n9934) );
  NOR2_X1 U11764 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  INV_X1 U11765 ( .A(n16809), .ZN(n16792) );
  AND2_X1 U11766 ( .A1(n17257), .A2(n15569), .ZN(n10030) );
  NOR2_X1 U11767 ( .A1(n18536), .A2(n17259), .ZN(n17257) );
  NOR2_X1 U11768 ( .A1(n17239), .A2(n15742), .ZN(n17258) );
  NAND2_X1 U11769 ( .A1(n9943), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9941) );
  OR2_X1 U11770 ( .A1(n16264), .A2(n16447), .ZN(n9940) );
  INV_X1 U11771 ( .A(n9851), .ZN(n17391) );
  AOI21_X2 U11772 ( .B1(n15633), .B2(n15632), .A(n18581), .ZN(n18019) );
  AOI21_X1 U11773 ( .B1(n11958), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A(n9759), .ZN(n11964) );
  INV_X1 U11774 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U11775 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n9974) );
  NAND2_X1 U11776 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n9975) );
  NAND2_X1 U11777 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U11778 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n9972) );
  AOI21_X1 U11779 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A(n9996), .ZN(n11753) );
  AND2_X1 U11780 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n9996)
         );
  AOI21_X1 U11781 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A(n9995), .ZN(n11733) );
  AND2_X1 U11782 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n9995)
         );
  AOI21_X1 U11783 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A(n9994), .ZN(n11712) );
  AND2_X1 U11784 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n9994)
         );
  AOI21_X1 U11785 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A(n9990), .ZN(n11682) );
  AND2_X1 U11786 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n9990)
         );
  AOI21_X1 U11787 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n9991), .ZN(n11688) );
  AND2_X1 U11788 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n9991)
         );
  AOI21_X1 U11789 ( .B1(n12569), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n10082), .ZN(n12453) );
  AND2_X1 U11790 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10082) );
  AND2_X1 U11791 ( .A1(n12017), .A2(n12016), .ZN(n12020) );
  AOI22_X1 U11792 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n13447), .B1(
        n11931), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U11793 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11936), .B1(
        n12006), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11906) );
  OR2_X1 U11794 ( .A1(n11949), .A2(n11901), .ZN(n11905) );
  NAND2_X1 U11795 ( .A1(n12229), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10430) );
  NOR2_X1 U11796 ( .A1(n10420), .A2(n12273), .ZN(n10447) );
  AND2_X1 U11797 ( .A1(n9977), .A2(n9976), .ZN(n11842) );
  NAND2_X1 U11798 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n9976) );
  NAND2_X1 U11799 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n9977) );
  AND2_X1 U11800 ( .A1(n9975), .A2(n9974), .ZN(n11823) );
  AND2_X1 U11801 ( .A1(n9973), .A2(n9972), .ZN(n11796) );
  AOI21_X1 U11802 ( .B1(n13274), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n9981), .ZN(n11600) );
  AND2_X1 U11803 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n9981)
         );
  AOI21_X1 U11804 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n9992), .ZN(n11583) );
  AND2_X1 U11805 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n9992)
         );
  AOI21_X1 U11806 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n9988), .ZN(n11498) );
  AND2_X1 U11807 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n9988)
         );
  AOI21_X1 U11808 ( .B1(n13274), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A(n9978), .ZN(n11517) );
  AND2_X1 U11809 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n9978)
         );
  AOI21_X1 U11810 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n9985), .ZN(n11536) );
  AND2_X1 U11811 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n9985)
         );
  AOI21_X1 U11812 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n9987), .ZN(n11565) );
  AND2_X1 U11813 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n9987)
         );
  AOI21_X1 U11814 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n9986), .ZN(n11551) );
  AND2_X1 U11815 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n9986)
         );
  AOI21_X1 U11816 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n9989), .ZN(n11456) );
  AND2_X1 U11817 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n9989)
         );
  AOI21_X1 U11818 ( .B1(n11751), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A(n9982), .ZN(n11419) );
  AND2_X1 U11819 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n9982)
         );
  AOI21_X1 U11820 ( .B1(n13274), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A(n9979), .ZN(n11429) );
  AND2_X1 U11821 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n9979)
         );
  INV_X1 U11822 ( .A(n11027), .ZN(n9805) );
  OR2_X1 U11823 ( .A1(n11236), .A2(n11235), .ZN(n11277) );
  AOI21_X1 U11824 ( .B1(n11752), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n9984), .ZN(n11210) );
  AND2_X1 U11825 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n9984)
         );
  AOI21_X1 U11826 ( .B1(n11840), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n9983), .ZN(n11083) );
  AND2_X1 U11827 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n9983) );
  INV_X1 U11828 ( .A(n11045), .ZN(n10216) );
  NOR2_X1 U11829 ( .A1(n10892), .A2(n9786), .ZN(n9785) );
  CLKBUF_X3 U11830 ( .A(n10979), .Z(n11839) );
  NAND2_X1 U11831 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10986) );
  AND2_X1 U11832 ( .A1(n10573), .A2(n10566), .ZN(n10576) );
  OR2_X1 U11833 ( .A1(n12230), .A2(n12038), .ZN(n10573) );
  INV_X1 U11834 ( .A(n10868), .ZN(n12015) );
  AOI21_X1 U11835 ( .B1(n12568), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n10092), .ZN(n12558) );
  AND2_X1 U11836 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10092) );
  AOI21_X1 U11837 ( .B1(n10354), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n10091), .ZN(n12552) );
  AND2_X1 U11838 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10091) );
  AOI21_X1 U11839 ( .B1(n12569), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n10090), .ZN(n12544) );
  AND2_X1 U11840 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10090) );
  AOI21_X1 U11841 ( .B1(n12569), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n10089), .ZN(n12539) );
  AND2_X1 U11842 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10089) );
  AND2_X1 U11843 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10081) );
  AOI21_X1 U11844 ( .B1(n10354), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n10088), .ZN(n12529) );
  AND2_X1 U11845 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10088) );
  AND2_X1 U11846 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10086) );
  AOI21_X1 U11847 ( .B1(n12569), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n10087), .ZN(n12510) );
  AND2_X1 U11848 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10087) );
  AOI21_X1 U11849 ( .B1(n12577), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n10080), .ZN(n12489) );
  AND2_X1 U11850 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10080) );
  AOI21_X1 U11851 ( .B1(n12569), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n10085), .ZN(n12484) );
  AND2_X1 U11852 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10085) );
  AND2_X1 U11853 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10084) );
  AOI21_X1 U11854 ( .B1(n12577), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n10083), .ZN(n12472) );
  AND2_X1 U11855 ( .A1(n12575), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10083) );
  NAND2_X1 U11856 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10284) );
  NAND2_X1 U11857 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10285) );
  OR2_X1 U11858 ( .A1(n13621), .A2(n12025), .ZN(n12160) );
  INV_X1 U11859 ( .A(n12080), .ZN(n10187) );
  NAND2_X1 U11860 ( .A1(n18902), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10190) );
  NAND2_X1 U11861 ( .A1(n11929), .A2(n19737), .ZN(n11930) );
  AOI21_X1 U11862 ( .B1(n11958), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A(n9756), .ZN(n11923) );
  NOR3_X1 U11863 ( .A1(n11915), .A2(n11913), .A3(n9757), .ZN(n9756) );
  INV_X1 U11864 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U11865 ( .A1(n10667), .A2(n10664), .ZN(n10078) );
  NAND2_X1 U11867 ( .A1(n9776), .A2(n12617), .ZN(n12218) );
  INV_X1 U11868 ( .A(n10376), .ZN(n9776) );
  NOR2_X1 U11869 ( .A1(n11889), .A2(n11891), .ZN(n11902) );
  NAND2_X1 U11870 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10307) );
  AOI22_X1 U11871 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U11872 ( .A1(n18708), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13874) );
  NAND2_X1 U11873 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18685), .ZN(
        n13875) );
  OR2_X1 U11874 ( .A1(n9876), .A2(n17858), .ZN(n9872) );
  AOI21_X1 U11875 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18541), .A(
        n13959), .ZN(n13964) );
  AND2_X1 U11876 ( .A1(n15569), .A2(n17744), .ZN(n15649) );
  NOR2_X1 U11877 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18708), .ZN(
        n14003) );
  OR2_X1 U11878 ( .A1(n18562), .A2(n13965), .ZN(n13966) );
  AND2_X1 U11879 ( .A1(n10122), .A2(n14106), .ZN(n10121) );
  AND2_X1 U11880 ( .A1(n11809), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11810) );
  NOR2_X1 U11881 ( .A1(n11764), .A2(n14309), .ZN(n11765) );
  AND2_X1 U11882 ( .A1(n10117), .A2(n14304), .ZN(n10116) );
  AOI21_X1 U11883 ( .B1(n13274), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n9980), .ZN(n11655) );
  AND2_X1 U11884 ( .A1(n13712), .A2(n13711), .ZN(n11578) );
  AND2_X1 U11885 ( .A1(n11576), .A2(n13799), .ZN(n14429) );
  AND2_X1 U11886 ( .A1(n13716), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11392) );
  NAND2_X1 U11887 ( .A1(n14532), .A2(n14543), .ZN(n9806) );
  INV_X1 U11888 ( .A(n14295), .ZN(n10128) );
  NOR2_X1 U11889 ( .A1(n14305), .A2(n10130), .ZN(n10129) );
  INV_X1 U11890 ( .A(n14319), .ZN(n10130) );
  NAND2_X1 U11891 ( .A1(n14630), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9813) );
  OR2_X1 U11892 ( .A1(n11289), .A2(n11298), .ZN(n15872) );
  OR2_X1 U11893 ( .A1(n11289), .A2(n11301), .ZN(n15873) );
  INV_X1 U11894 ( .A(n12780), .ZN(n11040) );
  OR2_X1 U11895 ( .A1(n11260), .A2(n11259), .ZN(n11276) );
  INV_X1 U11896 ( .A(n19934), .ZN(n9848) );
  NAND2_X1 U11897 ( .A1(n11203), .A2(n19999), .ZN(n11225) );
  NAND2_X1 U11898 ( .A1(n11169), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9839) );
  NAND3_X1 U11899 ( .A1(n10936), .A2(n10935), .A3(n10937), .ZN(n10226) );
  AND3_X1 U11900 ( .A1(n12901), .A2(n11029), .A3(n11307), .ZN(n12888) );
  OAI211_X1 U11901 ( .C1(n11159), .C2(n11177), .A(n11158), .B(n11157), .ZN(
        n11160) );
  NAND2_X1 U11902 ( .A1(n20750), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11867) );
  AND2_X1 U11903 ( .A1(n11173), .A2(n20638), .ZN(n20004) );
  INV_X1 U11904 ( .A(n12973), .ZN(n11028) );
  AND2_X1 U11905 ( .A1(n11317), .A2(n11316), .ZN(n12744) );
  OR2_X1 U11906 ( .A1(n11319), .A2(n11315), .ZN(n11317) );
  AOI21_X1 U11907 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20759), .A(
        n11359), .ZN(n11360) );
  OR3_X1 U11908 ( .A1(n11356), .A2(n11355), .A3(n12738), .ZN(n11357) );
  OR2_X1 U11909 ( .A1(n11356), .A2(n11308), .ZN(n11351) );
  AOI22_X1 U11910 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_7__2__SCAN_IN), .B2(n11100), .ZN(n10893) );
  NAND2_X1 U11911 ( .A1(n12312), .A2(n12240), .ZN(n10075) );
  NAND2_X1 U11912 ( .A1(n11929), .A2(n12229), .ZN(n10076) );
  OR2_X1 U11913 ( .A1(n12189), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16011) );
  NOR2_X1 U11914 ( .A1(n10104), .A2(n10873), .ZN(n10103) );
  AND2_X1 U11915 ( .A1(n13389), .A2(n10872), .ZN(n10873) );
  INV_X1 U11916 ( .A(n10105), .ZN(n10104) );
  NOR2_X1 U11917 ( .A1(n12140), .A2(n10106), .ZN(n10105) );
  INV_X1 U11918 ( .A(n10870), .ZN(n10106) );
  NOR2_X1 U11919 ( .A1(n10108), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10107) );
  INV_X1 U11920 ( .A(n10109), .ZN(n10108) );
  NOR2_X1 U11921 ( .A1(n10110), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10109) );
  INV_X1 U11922 ( .A(n12095), .ZN(n10110) );
  MUX2_X1 U11923 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n12040), .S(n12270), .Z(
        n12070) );
  NOR2_X1 U11924 ( .A1(n14858), .A2(n14213), .ZN(n12612) );
  NOR2_X1 U11925 ( .A1(n14990), .A2(n14977), .ZN(n10167) );
  AOI21_X1 U11926 ( .B1(n12577), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n10081), .ZN(n12524) );
  AOI21_X1 U11927 ( .B1(n12577), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n10086), .ZN(n12505) );
  NAND2_X1 U11928 ( .A1(n9738), .A2(n14926), .ZN(n10178) );
  NAND2_X1 U11929 ( .A1(n12431), .A2(n12430), .ZN(n12458) );
  NAND2_X1 U11930 ( .A1(n13830), .A2(n13832), .ZN(n13831) );
  INV_X1 U11931 ( .A(n13791), .ZN(n10181) );
  INV_X1 U11932 ( .A(n13640), .ZN(n10182) );
  NAND2_X1 U11933 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U11934 ( .A1(n10024), .A2(n10233), .ZN(n10023) );
  INV_X1 U11935 ( .A(n10025), .ZN(n10024) );
  OR2_X1 U11936 ( .A1(n10026), .A2(n10263), .ZN(n10025) );
  NAND2_X1 U11937 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10026) );
  INV_X1 U11938 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10018) );
  OR2_X1 U11939 ( .A1(n12024), .A2(n12023), .ZN(n12031) );
  NAND2_X1 U11940 ( .A1(n10063), .A2(n10062), .ZN(n10061) );
  INV_X1 U11941 ( .A(n13106), .ZN(n10062) );
  INV_X1 U11942 ( .A(n13124), .ZN(n10063) );
  OR2_X1 U11943 ( .A1(n12200), .A2(n12201), .ZN(n12203) );
  INV_X1 U11944 ( .A(n14209), .ZN(n10095) );
  OR3_X1 U11945 ( .A1(n12195), .A2(n12025), .A3(n15252), .ZN(n15065) );
  INV_X1 U11946 ( .A(n12117), .ZN(n10200) );
  AND2_X1 U11947 ( .A1(n9747), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9884) );
  INV_X1 U11948 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U11949 ( .A1(n10161), .A2(n10742), .ZN(n10160) );
  INV_X1 U11950 ( .A(n10164), .ZN(n10161) );
  NAND2_X1 U11951 ( .A1(n9890), .A2(n18886), .ZN(n12093) );
  NAND2_X1 U11952 ( .A1(n12087), .A2(n12025), .ZN(n9890) );
  NOR2_X1 U11953 ( .A1(n12079), .A2(n9742), .ZN(n10192) );
  INV_X1 U11954 ( .A(n9798), .ZN(n11982) );
  NOR2_X2 U11955 ( .A1(n9798), .A2(n9763), .ZN(n9887) );
  NOR2_X1 U11956 ( .A1(n9765), .A2(n11995), .ZN(n9764) );
  OAI211_X1 U11957 ( .C1(n10853), .C2(n18919), .A(n10617), .B(n10616), .ZN(
        n13183) );
  INV_X1 U11958 ( .A(n11925), .ZN(n11950) );
  NAND3_X1 U11959 ( .A1(n19682), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19516), 
        .ZN(n13381) );
  NAND2_X1 U11960 ( .A1(n10330), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10336) );
  AND4_X1 U11961 ( .A1(n10329), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        n10330) );
  NAND3_X1 U11962 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18702), .ZN(n13873) );
  NAND2_X1 U11963 ( .A1(n13876), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13877) );
  NOR2_X1 U11964 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13873), .ZN(
        n14087) );
  NOR3_X1 U11965 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n13874), .ZN(n14076) );
  NOR2_X1 U11966 ( .A1(n13875), .A2(n16791), .ZN(n15572) );
  NOR3_X1 U11967 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18523), .ZN(n15531) );
  NOR2_X1 U11968 ( .A1(n17741), .A2(n9945), .ZN(n9944) );
  NOR2_X1 U11969 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  NAND2_X1 U11970 ( .A1(n9668), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9950) );
  INV_X1 U11971 ( .A(n17461), .ZN(n9951) );
  AND2_X1 U11972 ( .A1(n9876), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10033) );
  NOR2_X1 U11973 ( .A1(n17883), .A2(n16283), .ZN(n16254) );
  INV_X1 U11974 ( .A(n18096), .ZN(n13989) );
  AND2_X1 U11975 ( .A1(n9749), .A2(n17614), .ZN(n10041) );
  AND2_X1 U11976 ( .A1(n10032), .A2(n10031), .ZN(n15595) );
  INV_X1 U11977 ( .A(n15594), .ZN(n9860) );
  XNOR2_X1 U11978 ( .A(n15649), .B(n9815), .ZN(n15650) );
  XNOR2_X1 U11979 ( .A(n17252), .B(n15569), .ZN(n15584) );
  NAND2_X1 U11980 ( .A1(n17302), .A2(n14008), .ZN(n16421) );
  AOI221_X1 U11981 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18688), .C1(n18742), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n18703), .ZN(n18080) );
  NAND2_X1 U11982 ( .A1(n14122), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11177) );
  NOR2_X1 U11983 ( .A1(n11449), .A2(n19774), .ZN(n11479) );
  NAND2_X1 U11984 ( .A1(n12996), .A2(n10232), .ZN(n13041) );
  INV_X1 U11985 ( .A(n19827), .ZN(n19836) );
  NAND2_X1 U11986 ( .A1(n14385), .A2(n14123), .ZN(n19826) );
  INV_X1 U11987 ( .A(n11867), .ZN(n11864) );
  OR2_X1 U11988 ( .A1(n11814), .A2(n11813), .ZN(n14271) );
  NAND2_X1 U11989 ( .A1(n10124), .A2(n10123), .ZN(n14283) );
  OR2_X1 U11990 ( .A1(n11769), .A2(n11768), .ZN(n14294) );
  OR2_X1 U11991 ( .A1(n11721), .A2(n14575), .ZN(n11722) );
  NAND2_X1 U11992 ( .A1(n11671), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11721) );
  NAND2_X1 U11993 ( .A1(n11677), .A2(n11676), .ZN(n14584) );
  AND2_X1 U11994 ( .A1(n11654), .A2(n11653), .ZN(n14413) );
  AND2_X1 U11995 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n11632), .ZN(
        n11633) );
  NAND2_X1 U11996 ( .A1(n11633), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11651) );
  NAND2_X1 U11997 ( .A1(n11596), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11631) );
  NOR2_X1 U11998 ( .A1(n11593), .A2(n15786), .ZN(n11596) );
  NOR2_X1 U11999 ( .A1(n10115), .A2(n14623), .ZN(n10114) );
  INV_X1 U12000 ( .A(n11578), .ZN(n10115) );
  NAND2_X1 U12001 ( .A1(n13710), .A2(n11578), .ZN(n14622) );
  NAND2_X1 U12002 ( .A1(n11531), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11515) );
  INV_X1 U12003 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20939) );
  NOR2_X1 U12004 ( .A1(n20939), .A2(n11515), .ZN(n11514) );
  NOR2_X1 U12005 ( .A1(n11572), .A2(n14644), .ZN(n11531) );
  OR2_X1 U12006 ( .A1(n14357), .A2(n13801), .ZN(n14438) );
  OR2_X1 U12007 ( .A1(n11557), .A2(n15820), .ZN(n11572) );
  AND2_X1 U12008 ( .A1(n11479), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11480) );
  AND2_X1 U12009 ( .A1(n11569), .A2(n11477), .ZN(n14354) );
  INV_X1 U12010 ( .A(n13653), .ZN(n11466) );
  NAND2_X1 U12011 ( .A1(n11443), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11449) );
  NAND2_X1 U12012 ( .A1(n11409), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11442) );
  NOR2_X1 U12013 ( .A1(n11401), .A2(n19809), .ZN(n11409) );
  NOR2_X1 U12014 ( .A1(n13333), .A2(n13334), .ZN(n13337) );
  NAND2_X1 U12015 ( .A1(n13337), .A2(n13336), .ZN(n13589) );
  NAND2_X1 U12016 ( .A1(n11394), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11401) );
  NOR2_X1 U12017 ( .A1(n11387), .A2(n13315), .ZN(n11394) );
  NAND2_X1 U12018 ( .A1(n12992), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12991) );
  AND2_X1 U12019 ( .A1(n11289), .A2(n10238), .ZN(n11305) );
  NAND2_X1 U12020 ( .A1(n9806), .A2(n14193), .ZN(n14510) );
  NOR2_X1 U12021 ( .A1(n14628), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10210) );
  NAND2_X1 U12022 ( .A1(n14510), .A2(n11289), .ZN(n10211) );
  NOR2_X1 U12023 ( .A1(n14281), .A2(n14273), .ZN(n14272) );
  NAND2_X1 U12024 ( .A1(n9969), .A2(n9967), .ZN(n14164) );
  NAND2_X1 U12025 ( .A1(n14169), .A2(n9970), .ZN(n9969) );
  NAND2_X1 U12026 ( .A1(n14331), .A2(n10127), .ZN(n14281) );
  AND2_X1 U12027 ( .A1(n9673), .A2(n14282), .ZN(n10127) );
  OAI21_X1 U12028 ( .B1(n14517), .B2(n14519), .A(n14788), .ZN(n14543) );
  NAND2_X1 U12029 ( .A1(n14331), .A2(n10129), .ZN(n14307) );
  NAND2_X1 U12030 ( .A1(n14331), .A2(n14319), .ZN(n14321) );
  AND2_X1 U12031 ( .A1(n14769), .A2(n9745), .ZN(n14720) );
  INV_X1 U12032 ( .A(n14722), .ZN(n10131) );
  OAI21_X1 U12033 ( .B1(n14593), .B2(n9754), .A(n14628), .ZN(n14579) );
  NAND2_X1 U12034 ( .A1(n14579), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14581) );
  NAND2_X1 U12035 ( .A1(n14769), .A2(n10132), .ZN(n14721) );
  AND2_X1 U12036 ( .A1(n14145), .A2(n14144), .ZN(n14344) );
  NAND2_X1 U12037 ( .A1(n14143), .A2(n9961), .ZN(n14144) );
  NAND2_X1 U12038 ( .A1(n14769), .A2(n9743), .ZN(n14416) );
  AND2_X1 U12039 ( .A1(n14769), .A2(n14423), .ZN(n14425) );
  AND2_X1 U12040 ( .A1(n14139), .A2(n14138), .ZN(n14772) );
  NAND2_X1 U12041 ( .A1(n14137), .A2(n9963), .ZN(n14138) );
  AND2_X1 U12042 ( .A1(n14771), .A2(n14772), .ZN(n14769) );
  NAND2_X1 U12043 ( .A1(n14455), .A2(n9725), .ZN(n14434) );
  INV_X1 U12044 ( .A(n14432), .ZN(n10142) );
  AND2_X1 U12045 ( .A1(n13755), .A2(n13754), .ZN(n14441) );
  NAND2_X1 U12046 ( .A1(n14455), .A2(n10143), .ZN(n14444) );
  AND2_X1 U12047 ( .A1(n14455), .A2(n14360), .ZN(n14362) );
  NAND2_X1 U12048 ( .A1(n14455), .A2(n9719), .ZN(n14442) );
  NAND2_X1 U12049 ( .A1(n14641), .A2(n14639), .ZN(n9796) );
  NAND2_X1 U12050 ( .A1(n13744), .A2(n9959), .ZN(n13745) );
  NOR2_X1 U12051 ( .A1(n14456), .A2(n14457), .ZN(n14455) );
  OR2_X1 U12052 ( .A1(n13769), .A2(n13768), .ZN(n14456) );
  NAND2_X1 U12053 ( .A1(n20720), .A2(n20759), .ZN(n11872) );
  AND2_X1 U12054 ( .A1(n13781), .A2(n9710), .ZN(n10219) );
  AND2_X1 U12055 ( .A1(n13603), .A2(n13602), .ZN(n13659) );
  NAND2_X1 U12056 ( .A1(n10136), .A2(n10134), .ZN(n13585) );
  NOR2_X1 U12057 ( .A1(n10138), .A2(n10135), .ZN(n10134) );
  INV_X1 U12058 ( .A(n9748), .ZN(n10135) );
  OR2_X1 U12059 ( .A1(n13667), .A2(n13666), .ZN(n13669) );
  NAND2_X1 U12060 ( .A1(n13537), .A2(n9957), .ZN(n13538) );
  NOR2_X1 U12061 ( .A1(n13095), .A2(n10139), .ZN(n19814) );
  OR2_X1 U12062 ( .A1(n13095), .A2(n13096), .ZN(n19815) );
  NAND2_X1 U12063 ( .A1(n13013), .A2(n13012), .ZN(n13025) );
  AND2_X1 U12064 ( .A1(n15938), .A2(n15943), .ZN(n14805) );
  NAND2_X1 U12065 ( .A1(n13033), .A2(n13284), .ZN(n15943) );
  NAND2_X1 U12066 ( .A1(n13033), .A2(n13032), .ZN(n14767) );
  NAND2_X1 U12067 ( .A1(n13020), .A2(n20014), .ZN(n11042) );
  NAND2_X1 U12068 ( .A1(n11118), .A2(n11117), .ZN(n11119) );
  NAND2_X1 U12069 ( .A1(n20047), .A2(n11132), .ZN(n12927) );
  INV_X1 U12070 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12918) );
  NAND2_X1 U12071 ( .A1(n12895), .A2(n12894), .ZN(n15688) );
  NOR2_X1 U12072 ( .A1(n20115), .A2(n9650), .ZN(n20108) );
  NOR2_X1 U12073 ( .A1(n20259), .A2(n9650), .ZN(n20262) );
  AND3_X1 U12074 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20759), .A3(n20000), 
        .ZN(n20040) );
  AND2_X1 U12075 ( .A1(n20292), .A2(n19999), .ZN(n20571) );
  NOR2_X1 U12076 ( .A1(n20750), .A2(n14128), .ZN(n13298) );
  AND2_X1 U12077 ( .A1(n13243), .A2(n13241), .ZN(n13252) );
  NAND2_X1 U12078 ( .A1(n10167), .A2(n10166), .ZN(n14858) );
  INV_X1 U12079 ( .A(n14856), .ZN(n10166) );
  OR2_X1 U12080 ( .A1(n16012), .A2(n12192), .ZN(n12200) );
  OR2_X1 U12081 ( .A1(n16021), .A2(n16022), .ZN(n10022) );
  NAND2_X1 U12082 ( .A1(n12188), .A2(n14923), .ZN(n12189) );
  NOR3_X1 U12083 ( .A1(n10255), .A2(n10020), .A3(n15081), .ZN(n10254) );
  AOI21_X1 U12084 ( .B1(n18782), .B2(n16078), .A(n18891), .ZN(n14876) );
  OR2_X1 U12085 ( .A1(n18782), .A2(n18891), .ZN(n10027) );
  NAND2_X1 U12086 ( .A1(n12122), .A2(n10877), .ZN(n12176) );
  NAND2_X1 U12087 ( .A1(n12171), .A2(n12186), .ZN(n12122) );
  INV_X1 U12088 ( .A(n10102), .ZN(n12155) );
  OR2_X1 U12089 ( .A1(n13849), .A2(n10280), .ZN(n10029) );
  AND2_X1 U12090 ( .A1(n12113), .A2(n10103), .ZN(n12135) );
  NAND2_X1 U12091 ( .A1(n12113), .A2(n10105), .ZN(n12143) );
  AND2_X1 U12092 ( .A1(n13389), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U12093 ( .A1(n12113), .A2(n10870), .ZN(n12141) );
  NAND2_X1 U12094 ( .A1(n13355), .A2(n13345), .ZN(n13344) );
  NAND2_X1 U12095 ( .A1(n12612), .A2(n12613), .ZN(n12616) );
  INV_X1 U12096 ( .A(n10167), .ZN(n14978) );
  NAND2_X1 U12097 ( .A1(n14911), .A2(n9697), .ZN(n10174) );
  INV_X1 U12098 ( .A(n12534), .ZN(n9774) );
  XNOR2_X1 U12099 ( .A(n12497), .B(n12499), .ZN(n14922) );
  NAND2_X1 U12100 ( .A1(n14922), .A2(n14921), .ZN(n14920) );
  INV_X1 U12101 ( .A(n12458), .ZN(n14942) );
  CLKBUF_X1 U12102 ( .A(n13831), .Z(n14943) );
  NOR2_X1 U12103 ( .A1(n10169), .A2(n9727), .ZN(n10168) );
  OR2_X1 U12104 ( .A1(n12376), .A2(n12375), .ZN(n13641) );
  INV_X1 U12105 ( .A(n13629), .ZN(n10175) );
  NOR2_X1 U12106 ( .A1(n16175), .A2(n16176), .ZN(n13100) );
  NAND2_X1 U12107 ( .A1(n10162), .A2(n10157), .ZN(n16175) );
  NOR2_X1 U12108 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  INV_X1 U12109 ( .A(n12951), .ZN(n10158) );
  INV_X1 U12110 ( .A(n10160), .ZN(n10159) );
  NAND2_X1 U12111 ( .A1(n10153), .A2(n9700), .ZN(n10152) );
  INV_X1 U12112 ( .A(n10659), .ZN(n10153) );
  INV_X1 U12113 ( .A(n12608), .ZN(n13382) );
  AND3_X1 U12114 ( .A1(n10552), .A2(n10551), .A3(n10550), .ZN(n14211) );
  AND3_X1 U12115 ( .A1(n10532), .A2(n10531), .A3(n10530), .ZN(n14939) );
  INV_X1 U12116 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15115) );
  AND2_X1 U12117 ( .A1(n13662), .A2(n9735), .ZN(n14958) );
  INV_X1 U12118 ( .A(n13862), .ZN(n10071) );
  INV_X1 U12119 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10263) );
  NOR2_X1 U12120 ( .A1(n10266), .A2(n10025), .ZN(n10264) );
  NOR2_X1 U12121 ( .A1(n13344), .A2(n12659), .ZN(n13565) );
  AND2_X1 U12122 ( .A1(n13565), .A2(n13564), .ZN(n13566) );
  NAND2_X1 U12123 ( .A1(n10014), .A2(n10017), .ZN(n10279) );
  NOR2_X1 U12124 ( .A1(n13125), .A2(n10059), .ZN(n13502) );
  NOR2_X1 U12125 ( .A1(n13125), .A2(n10061), .ZN(n13365) );
  OR2_X1 U12126 ( .A1(n13125), .A2(n13124), .ZN(n13127) );
  NAND2_X1 U12127 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10276) );
  NOR2_X1 U12128 ( .A1(n10050), .A2(n10052), .ZN(n10049) );
  INV_X1 U12129 ( .A(n10050), .ZN(n10048) );
  NAND2_X1 U12130 ( .A1(n10204), .A2(n10095), .ZN(n10206) );
  OAI211_X1 U12131 ( .C1(n14964), .C2(n19070), .A(n14216), .B(n10229), .ZN(
        n14217) );
  AND2_X1 U12132 ( .A1(n15249), .A2(n12295), .ZN(n15214) );
  AND3_X1 U12133 ( .A1(n10546), .A2(n10545), .A3(n10544), .ZN(n14908) );
  NAND2_X1 U12134 ( .A1(n10066), .A2(n10065), .ZN(n10064) );
  NOR2_X1 U12135 ( .A1(n10070), .A2(n14862), .ZN(n10065) );
  INV_X1 U12136 ( .A(n10067), .ZN(n10066) );
  NAND2_X1 U12137 ( .A1(n9824), .A2(n9822), .ZN(n15074) );
  OR2_X1 U12138 ( .A1(n9825), .A2(n12121), .ZN(n9824) );
  INV_X1 U12139 ( .A(n9894), .ZN(n9825) );
  NOR3_X1 U12140 ( .A1(n9676), .A2(n10070), .A3(n14939), .ZN(n14931) );
  AND3_X1 U12141 ( .A1(n10529), .A2(n10528), .A3(n10527), .ZN(n14949) );
  INV_X1 U12142 ( .A(n9916), .ZN(n9914) );
  AND2_X1 U12143 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n9917), .ZN(
        n9916) );
  NOR2_X1 U12144 ( .A1(n15349), .A2(n9918), .ZN(n9917) );
  AND3_X1 U12145 ( .A1(n10520), .A2(n10519), .A3(n10518), .ZN(n13773) );
  NAND2_X1 U12146 ( .A1(n13662), .A2(n9718), .ZN(n13863) );
  OR3_X1 U12147 ( .A1(n13853), .A2(n12025), .A3(n15358), .ZN(n15144) );
  OR2_X1 U12148 ( .A1(n18827), .A2(n12131), .ZN(n15156) );
  AND2_X1 U12149 ( .A1(n9660), .A2(n16170), .ZN(n9906) );
  NOR2_X1 U12150 ( .A1(n16081), .A2(n9768), .ZN(n9767) );
  INV_X1 U12151 ( .A(n15191), .ZN(n9768) );
  NAND2_X1 U12152 ( .A1(n13466), .A2(n12660), .ZN(n13616) );
  NAND2_X1 U12153 ( .A1(n9907), .A2(n9660), .ZN(n15423) );
  NAND2_X1 U12154 ( .A1(n10202), .A2(n12111), .ZN(n15426) );
  INV_X1 U12155 ( .A(n15448), .ZN(n10202) );
  AND3_X1 U12156 ( .A1(n10503), .A2(n10502), .A3(n10501), .ZN(n13354) );
  NAND2_X1 U12157 ( .A1(n10058), .A2(n13501), .ZN(n10057) );
  INV_X1 U12158 ( .A(n10059), .ZN(n10058) );
  AND2_X1 U12159 ( .A1(n12110), .A2(n12109), .ZN(n16104) );
  INV_X1 U12160 ( .A(n12029), .ZN(n9880) );
  OR2_X1 U12161 ( .A1(n12116), .A2(n15455), .ZN(n16101) );
  NAND2_X1 U12162 ( .A1(n10486), .A2(n10240), .ZN(n13125) );
  OAI21_X1 U12163 ( .B1(n12085), .B2(n13691), .A(n10184), .ZN(n10189) );
  XNOR2_X1 U12164 ( .A(n12093), .B(n13729), .ZN(n12091) );
  NAND2_X1 U12165 ( .A1(n13688), .A2(n9802), .ZN(n9801) );
  NOR2_X1 U12166 ( .A1(n13687), .A2(n12018), .ZN(n9802) );
  OR2_X1 U12167 ( .A1(n11887), .A2(n11886), .ZN(n11890) );
  OAI21_X1 U12168 ( .B1(n13408), .B2(n13371), .A(n19731), .ZN(n12341) );
  AND2_X1 U12169 ( .A1(n11881), .A2(n11880), .ZN(n11882) );
  NAND2_X1 U12170 ( .A1(n12250), .A2(n12793), .ZN(n12251) );
  INV_X1 U12171 ( .A(n19361), .ZN(n19367) );
  NOR2_X1 U12172 ( .A1(n13382), .A2(n13381), .ZN(n13405) );
  NOR2_X1 U12173 ( .A1(n13380), .A2(n13381), .ZN(n13406) );
  INV_X1 U12174 ( .A(n13407), .ZN(n13398) );
  NAND2_X2 U12175 ( .A1(n10391), .A2(n10390), .ZN(n13383) );
  INV_X1 U12176 ( .A(n19303), .ZN(n19266) );
  INV_X1 U12177 ( .A(n13405), .ZN(n13402) );
  INV_X1 U12178 ( .A(n13406), .ZN(n13403) );
  OR2_X1 U12179 ( .A1(n19475), .A2(n19266), .ZN(n19078) );
  NAND2_X1 U12180 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19516), .ZN(n13407) );
  NOR2_X1 U12181 ( .A1(n19683), .A2(n19736), .ZN(n19471) );
  NOR2_X1 U12182 ( .A1(n13511), .A2(n13510), .ZN(n13516) );
  INV_X1 U12183 ( .A(n16446), .ZN(n9933) );
  NOR2_X1 U12184 ( .A1(n16447), .A2(n16793), .ZN(n9932) );
  INV_X1 U12185 ( .A(n17439), .ZN(n9928) );
  NAND2_X1 U12186 ( .A1(n16764), .A2(n9927), .ZN(n9926) );
  NAND2_X1 U12187 ( .A1(n16734), .A2(n9928), .ZN(n9927) );
  NOR3_X1 U12188 ( .A1(n17036), .A2(n17056), .A3(n17075), .ZN(n17034) );
  INV_X1 U12189 ( .A(n13885), .ZN(n15558) );
  OAI21_X1 U12190 ( .B1(n13997), .B2(n13969), .A(n14020), .ZN(n15739) );
  NOR2_X1 U12191 ( .A1(n13905), .A2(n13904), .ZN(n16752) );
  OAI211_X1 U12192 ( .C1(n18530), .C2(n14019), .A(n18513), .B(n18733), .ZN(
        n15741) );
  NOR2_X1 U12193 ( .A1(n17303), .A2(n17266), .ZN(n17284) );
  NAND2_X1 U12194 ( .A1(n17495), .A2(n9949), .ZN(n17419) );
  INV_X1 U12195 ( .A(n17520), .ZN(n16604) );
  NOR3_X1 U12196 ( .A1(n16698), .A2(n17643), .A3(n16233), .ZN(n17605) );
  INV_X1 U12197 ( .A(n9875), .ZN(n17647) );
  AND3_X1 U12198 ( .A1(n9919), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17658) );
  NOR2_X1 U12199 ( .A1(n15569), .A2(n18689), .ZN(n15582) );
  XNOR2_X1 U12200 ( .A(n15584), .B(n15583), .ZN(n17723) );
  XNOR2_X1 U12201 ( .A(n15650), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17727) );
  NOR2_X1 U12202 ( .A1(n15569), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15651) );
  NAND2_X1 U12203 ( .A1(n17726), .A2(n17727), .ZN(n17725) );
  AOI22_X1 U12204 ( .A1(n18510), .A2(n18509), .B1(n18514), .B2(n18041), .ZN(
        n16232) );
  NAND2_X1 U12205 ( .A1(n17574), .A2(n17745), .ZN(n17483) );
  NOR2_X1 U12206 ( .A1(n17755), .A2(n16272), .ZN(n16255) );
  OR2_X1 U12207 ( .A1(n16295), .A2(n17913), .ZN(n9864) );
  NAND2_X1 U12208 ( .A1(n17384), .A2(n9866), .ZN(n9865) );
  AND2_X1 U12209 ( .A1(n16293), .A2(n9867), .ZN(n9866) );
  AND2_X1 U12210 ( .A1(n18041), .A2(n16292), .ZN(n9867) );
  NOR2_X1 U12211 ( .A1(n17402), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17401) );
  NOR2_X1 U12212 ( .A1(n15616), .A2(n17648), .ZN(n17427) );
  NOR2_X1 U12213 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n9876), .ZN(
        n17513) );
  INV_X1 U12214 ( .A(n15608), .ZN(n15606) );
  NAND2_X1 U12215 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17567), .ZN(
        n17806) );
  NOR2_X1 U12216 ( .A1(n17118), .A2(n18089), .ZN(n15629) );
  INV_X1 U12217 ( .A(n16222), .ZN(n18513) );
  NAND2_X1 U12218 ( .A1(n9875), .A2(n9659), .ZN(n15607) );
  NOR2_X1 U12219 ( .A1(n17560), .A2(n15597), .ZN(n17555) );
  NOR2_X1 U12220 ( .A1(n17937), .A2(n17885), .ZN(n17567) );
  NOR2_X1 U12221 ( .A1(n17917), .A2(n10040), .ZN(n17561) );
  NAND2_X1 U12222 ( .A1(n17561), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17560) );
  INV_X1 U12223 ( .A(n17937), .ZN(n17914) );
  NAND2_X1 U12224 ( .A1(n17627), .A2(n10041), .ZN(n17592) );
  NAND2_X1 U12225 ( .A1(n17668), .A2(n15659), .ZN(n17656) );
  NAND2_X1 U12226 ( .A1(n10037), .A2(n10036), .ZN(n17696) );
  NAND2_X1 U12227 ( .A1(n17713), .A2(n10039), .ZN(n10036) );
  NOR2_X1 U12228 ( .A1(n15630), .A2(n15621), .ZN(n18041) );
  NAND2_X1 U12229 ( .A1(n17744), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17743) );
  INV_X1 U12230 ( .A(n13876), .ZN(n16791) );
  NAND2_X1 U12231 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18523) );
  INV_X1 U12232 ( .A(n18526), .ZN(n18522) );
  INV_X1 U12233 ( .A(n18039), .ZN(n18548) );
  AND2_X1 U12234 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18553) );
  NAND2_X1 U12235 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18553), .ZN(
        n18556) );
  INV_X1 U12236 ( .A(n16752), .ZN(n18082) );
  NAND3_X1 U12237 ( .A1(n13980), .A2(n13979), .A3(n13978), .ZN(n18085) );
  AOI22_X1 U12238 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16976), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13979) );
  AOI22_X1 U12239 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13980) );
  AOI211_X1 U12240 ( .C1(n9638), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n13977), .B(n13976), .ZN(n13978) );
  INV_X1 U12241 ( .A(n18374), .ZN(n18426) );
  INV_X1 U12242 ( .A(n16232), .ZN(n18570) );
  NOR2_X1 U12243 ( .A1(n16423), .A2(n18742), .ZN(n18727) );
  INV_X1 U12244 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n20899) );
  OR2_X1 U12245 ( .A1(n12772), .A2(n19750), .ZN(n14242) );
  AND2_X1 U12246 ( .A1(n19827), .A2(n14116), .ZN(n19797) );
  AND2_X1 U12247 ( .A1(n14129), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14116) );
  INV_X1 U12248 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19809) );
  INV_X1 U12249 ( .A(n19849), .ZN(n19847) );
  AND2_X1 U12250 ( .A1(n19827), .A2(n14130), .ZN(n19850) );
  NOR2_X2 U12251 ( .A1(n14173), .A2(n14172), .ZN(n19834) );
  INV_X1 U12252 ( .A(n19834), .ZN(n19865) );
  INV_X1 U12253 ( .A(n19830), .ZN(n19858) );
  AND2_X2 U12254 ( .A1(n12877), .A2(n13012), .ZN(n19873) );
  OR2_X1 U12255 ( .A1(n12998), .A2(n12969), .ZN(n12875) );
  INV_X1 U12256 ( .A(n15870), .ZN(n14493) );
  NOR2_X1 U12257 ( .A1(n15863), .A2(n12974), .ZN(n15867) );
  NAND2_X1 U12258 ( .A1(n12971), .A2(n12970), .ZN(n12972) );
  OR2_X1 U12259 ( .A1(n12969), .A2(n12968), .ZN(n12970) );
  INV_X1 U12260 ( .A(n15863), .ZN(n14505) );
  NAND2_X1 U12261 ( .A1(n14505), .A2(n12974), .ZN(n14504) );
  AND2_X1 U12262 ( .A1(n12843), .A2(n14121), .ZN(n19877) );
  INV_X2 U12263 ( .A(n13140), .ZN(n19929) );
  OR2_X1 U12264 ( .A1(n9707), .A2(n14318), .ZN(n14571) );
  XNOR2_X1 U12265 ( .A(n14642), .B(n9807), .ZN(n15942) );
  AND2_X1 U12266 ( .A1(n13579), .A2(n13535), .ZN(n19790) );
  INV_X1 U12267 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U12268 ( .A1(n11370), .A2(n11386), .ZN(n12982) );
  XNOR2_X1 U12269 ( .A(n9779), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14682) );
  NAND2_X1 U12270 ( .A1(n9781), .A2(n9780), .ZN(n9779) );
  NAND2_X1 U12271 ( .A1(n14534), .A2(n11289), .ZN(n9780) );
  NAND2_X1 U12272 ( .A1(n14533), .A2(n14788), .ZN(n9781) );
  OR2_X1 U12273 ( .A1(n14773), .A2(n14190), .ZN(n14715) );
  AND2_X1 U12274 ( .A1(n15887), .A2(n15886), .ZN(n15931) );
  OR2_X1 U12275 ( .A1(n11872), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15922) );
  AND2_X1 U12276 ( .A1(n10222), .A2(n13781), .ZN(n10220) );
  NAND2_X1 U12277 ( .A1(n15917), .A2(n15916), .ZN(n15915) );
  NAND2_X1 U12278 ( .A1(n19933), .A2(n11223), .ZN(n15917) );
  NAND2_X1 U12279 ( .A1(n9833), .A2(n9832), .ZN(n13313) );
  INV_X1 U12280 ( .A(n9835), .ZN(n9833) );
  INV_X1 U12281 ( .A(n14805), .ZN(n19961) );
  INV_X1 U12282 ( .A(n14832), .ZN(n19988) );
  INV_X1 U12283 ( .A(n20576), .ZN(n20573) );
  NAND2_X1 U12284 ( .A1(n10000), .A2(n20148), .ZN(n9811) );
  INV_X1 U12285 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19995) );
  OAI21_X1 U12286 ( .B1(n13299), .B2(n15998), .A(n20154), .ZN(n20738) );
  INV_X1 U12287 ( .A(n20719), .ZN(n15714) );
  NOR2_X1 U12288 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20720) );
  OAI211_X1 U12289 ( .C1(n20041), .C2(n20301), .A(n20356), .B(n20006), .ZN(
        n20044) );
  INV_X1 U12290 ( .A(n20215), .ZN(n20187) );
  INV_X1 U12291 ( .A(n20261), .ZN(n20288) );
  OAI211_X1 U12292 ( .C1(n20317), .C2(n20301), .A(n20356), .B(n20300), .ZN(
        n20319) );
  OAI21_X1 U12293 ( .B1(n20398), .B2(n20397), .A(n20472), .ZN(n20425) );
  INV_X1 U12294 ( .A(n20582), .ZN(n20514) );
  INV_X1 U12295 ( .A(n20589), .ZN(n20528) );
  INV_X1 U12296 ( .A(n20597), .ZN(n20533) );
  INV_X1 U12297 ( .A(n20605), .ZN(n20538) );
  INV_X1 U12298 ( .A(n20613), .ZN(n20543) );
  INV_X1 U12299 ( .A(n20621), .ZN(n20548) );
  INV_X1 U12300 ( .A(n20629), .ZN(n20553) );
  OAI211_X1 U12301 ( .C1(n20559), .C2(n20523), .A(n20522), .B(n20521), .ZN(
        n20561) );
  INV_X1 U12302 ( .A(n20639), .ZN(n20560) );
  NAND2_X1 U12303 ( .A1(n20462), .A2(n20461), .ZN(n20564) );
  AND2_X1 U12304 ( .A1(n20462), .A2(n9654), .ZN(n20644) );
  OR2_X1 U12305 ( .A1(n20649), .A2(n20759), .ZN(n19750) );
  NAND2_X1 U12306 ( .A1(n14128), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20649) );
  INV_X2 U12307 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20750) );
  NAND2_X1 U12308 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20661) );
  OR2_X1 U12309 ( .A1(n10882), .A2(n12665), .ZN(n12670) );
  OR2_X1 U12310 ( .A1(n18891), .A2(n14842), .ZN(n16001) );
  NOR2_X1 U12311 ( .A1(n16031), .A2(n18891), .ZN(n16021) );
  INV_X1 U12312 ( .A(n10022), .ZN(n16020) );
  AOI21_X1 U12313 ( .B1(n13849), .B2(n10028), .A(n10280), .ZN(n18795) );
  AND2_X1 U12314 ( .A1(n10029), .A2(n10028), .ZN(n18807) );
  AND2_X1 U12315 ( .A1(n18751), .A2(n10858), .ZN(n18922) );
  OR2_X1 U12316 ( .A1(n18751), .A2(n10861), .ZN(n18918) );
  INV_X1 U12317 ( .A(n18922), .ZN(n18916) );
  INV_X1 U12318 ( .A(n18878), .ZN(n18927) );
  OR2_X1 U12319 ( .A1(n10815), .A2(n10814), .ZN(n13562) );
  OR2_X1 U12320 ( .A1(n10803), .A2(n10802), .ZN(n13416) );
  OR2_X1 U12321 ( .A1(n10778), .A2(n10777), .ZN(n13352) );
  INV_X1 U12322 ( .A(n14961), .ZN(n14945) );
  NOR2_X1 U12323 ( .A1(n14934), .A2(n12460), .ZN(n14927) );
  INV_X1 U12324 ( .A(n13643), .ZN(n12649) );
  CLKBUF_X1 U12325 ( .A(n12960), .Z(n13051) );
  OR2_X1 U12326 ( .A1(n16065), .A2(n12816), .ZN(n18958) );
  NOR2_X1 U12327 ( .A1(n15475), .A2(n12762), .ZN(n18989) );
  AND4_X1 U12328 ( .A1(n13408), .A2(n12761), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19731), .ZN(n12762) );
  INV_X1 U12329 ( .A(n18958), .ZN(n18992) );
  INV_X2 U12330 ( .A(n18998), .ZN(n19028) );
  INV_X2 U12331 ( .A(n12869), .ZN(n19035) );
  AOI21_X1 U12332 ( .B1(n9903), .B2(n10196), .A(n9901), .ZN(n9898) );
  NAND2_X1 U12333 ( .A1(n15188), .A2(n9903), .ZN(n9897) );
  AND2_X1 U12334 ( .A1(n13774), .A2(n13706), .ZN(n18823) );
  NAND2_X1 U12335 ( .A1(n15187), .A2(n15191), .ZN(n16084) );
  NAND2_X1 U12336 ( .A1(n9792), .A2(n12029), .ZN(n16127) );
  OR2_X1 U12337 ( .A1(n18757), .A2(n10635), .ZN(n16133) );
  INV_X1 U12338 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16152) );
  NAND2_X1 U12339 ( .A1(n18757), .A2(n12056), .ZN(n16151) );
  INV_X1 U12340 ( .A(n16142), .ZN(n19052) );
  INV_X1 U12341 ( .A(n16151), .ZN(n19039) );
  INV_X1 U12342 ( .A(n16133), .ZN(n19042) );
  NAND3_X1 U12343 ( .A1(n10045), .A2(n10044), .A3(n10046), .ZN(n14889) );
  NAND2_X1 U12344 ( .A1(n10047), .A2(n10563), .ZN(n10046) );
  OR2_X1 U12345 ( .A1(n14907), .A2(n10562), .ZN(n10045) );
  XNOR2_X1 U12346 ( .A(n9891), .B(n9691), .ZN(n12315) );
  NAND2_X1 U12347 ( .A1(n9892), .A2(n10094), .ZN(n9891) );
  NOR2_X1 U12348 ( .A1(n9752), .A2(n10149), .ZN(n10148) );
  NAND2_X1 U12349 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10149) );
  NAND2_X1 U12350 ( .A1(n15225), .A2(n10239), .ZN(n15049) );
  NAND2_X1 U12351 ( .A1(n9896), .A2(n9893), .ZN(n15088) );
  NAND2_X1 U12352 ( .A1(n12121), .A2(n9826), .ZN(n9896) );
  OR2_X1 U12353 ( .A1(n15188), .A2(n10196), .ZN(n9902) );
  XNOR2_X1 U12354 ( .A(n9766), .B(n9721), .ZN(n15317) );
  OAI21_X1 U12355 ( .B1(n15123), .B2(n15113), .A(n15121), .ZN(n9766) );
  NAND2_X1 U12356 ( .A1(n9912), .A2(n9911), .ZN(n15338) );
  OR2_X1 U12357 ( .A1(n15127), .A2(n15335), .ZN(n9911) );
  NOR2_X1 U12358 ( .A1(n15127), .A2(n9914), .ZN(n9913) );
  INV_X1 U12359 ( .A(n15139), .ZN(n15148) );
  NAND2_X1 U12360 ( .A1(n16189), .A2(n19075), .ZN(n10011) );
  NAND2_X1 U12361 ( .A1(n10010), .A2(n10009), .ZN(n10008) );
  NAND2_X1 U12362 ( .A1(n15371), .A2(n15370), .ZN(n10009) );
  INV_X1 U12363 ( .A(n13635), .ZN(n16159) );
  NAND2_X1 U12364 ( .A1(n10201), .A2(n12117), .ZN(n15411) );
  NAND2_X1 U12365 ( .A1(n9830), .A2(n9828), .ZN(n10201) );
  NOR2_X1 U12366 ( .A1(n13725), .A2(n12293), .ZN(n16194) );
  NAND2_X1 U12367 ( .A1(n10163), .A2(n9677), .ZN(n12819) );
  OR2_X1 U12368 ( .A1(n12814), .A2(n12813), .ZN(n10163) );
  NAND2_X1 U12369 ( .A1(n12085), .A2(n12066), .ZN(n13683) );
  INV_X1 U12370 ( .A(n9905), .ZN(n13685) );
  AND2_X1 U12371 ( .A1(n10055), .A2(n10241), .ZN(n13055) );
  AND2_X1 U12372 ( .A1(n10193), .A2(n10194), .ZN(n13478) );
  INV_X1 U12373 ( .A(n16188), .ZN(n19067) );
  INV_X1 U12374 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19714) );
  INV_X1 U12375 ( .A(n18989), .ZN(n19708) );
  XNOR2_X1 U12376 ( .A(n12769), .B(n12768), .ZN(n19699) );
  NOR2_X1 U12377 ( .A1(n13178), .A2(n10659), .ZN(n13196) );
  INV_X1 U12378 ( .A(n19699), .ZN(n19076) );
  XNOR2_X1 U12379 ( .A(n12939), .B(n12941), .ZN(n19697) );
  AND2_X1 U12380 ( .A1(n13065), .A2(n13064), .ZN(n13451) );
  AND2_X1 U12381 ( .A1(n13248), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16215) );
  INV_X1 U12382 ( .A(n10396), .ZN(n9885) );
  INV_X1 U12383 ( .A(n19147), .ZN(n19156) );
  OR2_X1 U12384 ( .A1(n19207), .A2(n19469), .ZN(n19225) );
  NOR2_X2 U12385 ( .A1(n19302), .A2(n19208), .ZN(n19259) );
  NAND2_X1 U12386 ( .A1(n9758), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19264) );
  OR2_X1 U12387 ( .A1(n19367), .A2(n19435), .ZN(n19354) );
  INV_X1 U12388 ( .A(n19345), .ZN(n19349) );
  OAI21_X1 U12389 ( .B1(n19458), .B2(n19731), .A(n19441), .ZN(n19461) );
  NOR2_X1 U12390 ( .A1(n19475), .A2(n19208), .ZN(n19460) );
  INV_X1 U12391 ( .A(n19501), .ZN(n19494) );
  OAI22_X1 U12392 ( .A1(n16311), .A2(n13403), .B1(n20933), .B2(n13402), .ZN(
        n19530) );
  AND2_X1 U12393 ( .A1(n10414), .A2(n13398), .ZN(n19529) );
  AND2_X1 U12394 ( .A1(n10635), .A2(n13398), .ZN(n19551) );
  INV_X1 U12395 ( .A(n19528), .ZN(n19559) );
  INV_X1 U12396 ( .A(n19452), .ZN(n19567) );
  INV_X1 U12397 ( .A(n19491), .ZN(n19568) );
  INV_X1 U12398 ( .A(n19537), .ZN(n19566) );
  INV_X1 U12399 ( .A(n19543), .ZN(n19580) );
  NOR2_X2 U12400 ( .A1(n19435), .A2(n19266), .ZN(n19593) );
  INV_X1 U12401 ( .A(n19078), .ZN(n19591) );
  AND2_X1 U12402 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10584), .ZN(n16213) );
  AND2_X1 U12403 ( .A1(n13270), .A2(n13269), .ZN(n16214) );
  NAND2_X1 U12404 ( .A1(n18727), .A2(n18513), .ZN(n17303) );
  INV_X1 U12405 ( .A(n16450), .ZN(n9937) );
  NOR2_X1 U12406 ( .A1(n16515), .A2(n17439), .ZN(n16514) );
  NOR2_X1 U12407 ( .A1(n16521), .A2(n16734), .ZN(n16515) );
  NOR2_X1 U12408 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16550), .ZN(n16536) );
  INV_X1 U12409 ( .A(n16778), .ZN(n16799) );
  AND2_X1 U12410 ( .A1(n9922), .A2(n16764), .ZN(n16538) );
  INV_X1 U12411 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16671) );
  NOR2_X1 U12412 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16673), .ZN(n16672) );
  INV_X1 U12413 ( .A(n16784), .ZN(n16793) );
  INV_X1 U12414 ( .A(n16569), .ZN(n16798) );
  INV_X1 U12415 ( .A(n16798), .ZN(n16807) );
  OAI211_X1 U12416 ( .C1(n16423), .C2(n18451), .A(n16422), .B(n18725), .ZN(
        n16809) );
  NOR2_X1 U12417 ( .A1(n16508), .A2(n16860), .ZN(n16864) );
  NOR2_X1 U12418 ( .A1(n16529), .A2(n16870), .ZN(n16875) );
  NOR4_X1 U12419 ( .A1(n16583), .A2(n16593), .A3(n14023), .A4(n16929), .ZN(
        n16941) );
  INV_X2 U12420 ( .A(n17105), .ZN(n17101) );
  AND2_X1 U12421 ( .A1(n17107), .A2(n18114), .ZN(n17105) );
  INV_X1 U12422 ( .A(n17124), .ZN(n17120) );
  NOR2_X1 U12423 ( .A1(n17327), .A2(n17143), .ZN(n17138) );
  INV_X1 U12424 ( .A(n17149), .ZN(n17144) );
  NAND2_X1 U12425 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17144), .ZN(n17143) );
  INV_X1 U12426 ( .A(n17168), .ZN(n17163) );
  INV_X1 U12427 ( .A(n17182), .ZN(n17178) );
  INV_X1 U12428 ( .A(n17171), .ZN(n17188) );
  NOR2_X1 U12429 ( .A1(n17259), .A2(n17197), .ZN(n17212) );
  NOR2_X1 U12430 ( .A1(n15508), .A2(n15507), .ZN(n17240) );
  INV_X1 U12431 ( .A(n17258), .ZN(n17256) );
  INV_X1 U12432 ( .A(n17257), .ZN(n17253) );
  CLKBUF_X2 U12433 ( .A(n17330), .Z(n17368) );
  NOR2_X1 U12434 ( .A1(n17372), .A2(n16234), .ZN(n16264) );
  NAND2_X1 U12436 ( .A1(n17495), .A2(n9666), .ZN(n17485) );
  NAND2_X1 U12437 ( .A1(n16604), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17506) );
  NAND2_X1 U12438 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17742), .ZN(n17576) );
  INV_X1 U12439 ( .A(n17806), .ZN(n17884) );
  NAND2_X1 U12440 ( .A1(n17605), .A2(n9665), .ZN(n17564) );
  INV_X1 U12441 ( .A(n17917), .ZN(n17583) );
  NAND2_X1 U12442 ( .A1(n9919), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17680) );
  NOR2_X1 U12443 ( .A1(n18085), .A2(n16406), .ZN(n17738) );
  NOR2_X1 U12444 ( .A1(n17716), .A2(n17532), .ZN(n17742) );
  INV_X1 U12445 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17741) );
  INV_X1 U12446 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18688) );
  INV_X1 U12447 ( .A(n17734), .ZN(n17748) );
  XNOR2_X1 U12448 ( .A(n15725), .B(n15724), .ZN(n16252) );
  NAND2_X1 U12449 ( .A1(n16284), .A2(n9876), .ZN(n9852) );
  NAND2_X1 U12450 ( .A1(n9862), .A2(n9861), .ZN(n16296) );
  NOR2_X1 U12451 ( .A1(n18017), .A2(n15670), .ZN(n9861) );
  NAND2_X1 U12452 ( .A1(n9865), .A2(n9863), .ZN(n9862) );
  AND2_X1 U12453 ( .A1(n16294), .A2(n9864), .ZN(n9863) );
  INV_X1 U12454 ( .A(n16284), .ZN(n17390) );
  NAND2_X1 U12455 ( .A1(n17443), .A2(n15612), .ZN(n17435) );
  NAND2_X1 U12456 ( .A1(n17475), .A2(n15614), .ZN(n17444) );
  INV_X1 U12457 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18742) );
  NOR2_X1 U12458 ( .A1(n17832), .A2(n9816), .ZN(n17835) );
  NAND2_X1 U12459 ( .A1(n9818), .A2(n9817), .ZN(n9816) );
  INV_X1 U12460 ( .A(n17833), .ZN(n9817) );
  AND2_X1 U12461 ( .A1(n9821), .A2(n9820), .ZN(n17869) );
  NAND2_X1 U12462 ( .A1(n17806), .A2(n17938), .ZN(n9820) );
  OR2_X1 U12463 ( .A1(n17555), .A2(n18045), .ZN(n9821) );
  INV_X1 U12464 ( .A(n17555), .ZN(n17883) );
  INV_X1 U12465 ( .A(n17967), .ZN(n17982) );
  OAI21_X2 U12466 ( .B1(n18520), .B2(n18522), .A(n18519), .ZN(n18524) );
  AND2_X1 U12467 ( .A1(n17627), .A2(n9749), .ZN(n17609) );
  NAND2_X1 U12468 ( .A1(n17627), .A2(n17962), .ZN(n17618) );
  INV_X1 U12469 ( .A(n17602), .ZN(n17939) );
  NAND2_X1 U12470 ( .A1(n9855), .A2(n9856), .ZN(n17663) );
  INV_X1 U12471 ( .A(n10032), .ZN(n17671) );
  INV_X1 U12472 ( .A(n18019), .ZN(n18065) );
  INV_X1 U12473 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18541) );
  INV_X1 U12474 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18561) );
  INV_X1 U12475 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18563) );
  INV_X1 U12476 ( .A(n16757), .ZN(n18585) );
  AND2_X1 U12477 ( .A1(n12635), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19996)
         );
  AND2_X1 U12479 ( .A1(n14462), .A2(n19938), .ZN(n11876) );
  AOI211_X1 U12480 ( .C1(n15909), .C2(n14131), .A(n14109), .B(n14108), .ZN(
        n14110) );
  NAND2_X1 U12481 ( .A1(n9953), .A2(n19939), .ZN(n14561) );
  OAI211_X1 U12482 ( .C1(n14656), .C2(n14832), .A(n10126), .B(n10125), .ZN(
        P1_U3001) );
  OR2_X1 U12483 ( .A1(n14652), .A2(n19981), .ZN(n10125) );
  AOI21_X1 U12484 ( .B1(n14655), .B2(n14654), .A(n14653), .ZN(n10126) );
  AND2_X1 U12485 ( .A1(n12622), .A2(n12621), .ZN(n12623) );
  OAI21_X1 U12486 ( .B1(n15039), .B2(n16204), .A(n9831), .ZN(P2_U3017) );
  NOR2_X1 U12487 ( .A1(n9701), .A2(n9661), .ZN(n9831) );
  OR2_X1 U12488 ( .A1(n16449), .A2(n9936), .ZN(n9935) );
  AOI21_X1 U12489 ( .B1(n16454), .B2(n16818), .A(n9930), .ZN(n9929) );
  NAND2_X1 U12490 ( .A1(n9938), .A2(n9937), .ZN(n9936) );
  AOI21_X1 U12491 ( .B1(n17258), .B2(BUF2_REG_1__SCAN_IN), .A(n10030), .ZN(
        n17264) );
  NOR2_X2 U12492 ( .A1(n18523), .A2(n13875), .ZN(n13937) );
  AND2_X1 U12493 ( .A1(n10182), .A2(n9664), .ZN(n9655) );
  NAND2_X1 U12494 ( .A1(n10017), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10016) );
  AND2_X1 U12495 ( .A1(n12575), .A2(n13075), .ZN(n10641) );
  CLKBUF_X3 U12496 ( .A(n10354), .Z(n12577) );
  AND2_X1 U12497 ( .A1(n15124), .A2(n9747), .ZN(n9656) );
  NOR2_X1 U12498 ( .A1(n10266), .A2(n15180), .ZN(n10267) );
  NAND2_X1 U12499 ( .A1(n11889), .A2(n11899), .ZN(n15462) );
  NOR2_X1 U12500 ( .A1(n9903), .A2(n9901), .ZN(n9657) );
  OR2_X1 U12501 ( .A1(n10394), .A2(n10395), .ZN(n9658) );
  AND2_X1 U12502 ( .A1(n15601), .A2(n16282), .ZN(n9659) );
  AND2_X1 U12503 ( .A1(n9909), .A2(n15125), .ZN(n9660) );
  OR3_X1 U12504 ( .A1(n9676), .A2(n10067), .A3(n10070), .ZN(n9662) );
  AND2_X1 U12505 ( .A1(n10124), .A2(n10122), .ZN(n9663) );
  INV_X1 U12506 ( .A(n15373), .ZN(n10012) );
  AND2_X1 U12507 ( .A1(n11885), .A2(n11890), .ZN(n18928) );
  INV_X1 U12508 ( .A(n18928), .ZN(n9877) );
  INV_X1 U12509 ( .A(n10016), .ZN(n10015) );
  OR2_X1 U12510 ( .A1(n13019), .A2(n12774), .ZN(n12998) );
  NAND2_X1 U12512 ( .A1(n10182), .A2(n12387), .ZN(n13776) );
  OR2_X1 U12513 ( .A1(n13059), .A2(n10176), .ZN(n13561) );
  AND2_X1 U12514 ( .A1(n12387), .A2(n10181), .ZN(n9664) );
  AND2_X1 U12515 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9665) );
  AND2_X1 U12516 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9666) );
  AND2_X1 U12517 ( .A1(n10210), .A2(n11304), .ZN(n9667) );
  AND2_X1 U12518 ( .A1(n9666), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9668) );
  AND2_X1 U12519 ( .A1(n11224), .A2(n11248), .ZN(n9669) );
  AND2_X1 U12520 ( .A1(n10027), .A2(n16078), .ZN(n9670) );
  AND2_X1 U12521 ( .A1(n9665), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9671) );
  AND2_X1 U12522 ( .A1(n9667), .A2(n14650), .ZN(n9672) );
  NAND2_X1 U12523 ( .A1(n13179), .A2(n10155), .ZN(n13197) );
  NAND3_X1 U12524 ( .A1(n9940), .A2(n9939), .A3(n9941), .ZN(n16764) );
  NAND2_X1 U12525 ( .A1(n11910), .A2(n9755), .ZN(n19270) );
  AND2_X1 U12526 ( .A1(n10129), .A2(n10128), .ZN(n9673) );
  AND2_X1 U12527 ( .A1(n15614), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9674) );
  AND2_X1 U12528 ( .A1(n15310), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9675) );
  INV_X4 U12529 ( .A(n13939), .ZN(n15536) );
  OR2_X1 U12530 ( .A1(n14956), .A2(n14949), .ZN(n9676) );
  NOR2_X2 U12531 ( .A1(n13874), .A2(n13875), .ZN(n13884) );
  NAND2_X1 U12532 ( .A1(n11192), .A2(n11191), .ZN(n19999) );
  OR2_X1 U12533 ( .A1(n12025), .A2(n10831), .ZN(n9677) );
  INV_X1 U12534 ( .A(n15534), .ZN(n15487) );
  INV_X1 U12535 ( .A(n17648), .ZN(n9876) );
  OR2_X1 U12536 ( .A1(n18685), .A2(n9854), .ZN(n9678) );
  XNOR2_X1 U12537 ( .A(n10247), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12060) );
  INV_X2 U12538 ( .A(n12774), .ZN(n9956) );
  INV_X1 U12539 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13371) );
  INV_X1 U12540 ( .A(n10418), .ZN(n10431) );
  NAND2_X1 U12541 ( .A1(n12096), .A2(n12095), .ZN(n12094) );
  NAND2_X1 U12542 ( .A1(n9898), .A2(n9897), .ZN(n15098) );
  NAND2_X1 U12543 ( .A1(n15124), .A2(n9884), .ZN(n15089) );
  NAND2_X1 U12544 ( .A1(n10021), .A2(n10275), .ZN(n10273) );
  AND2_X1 U12545 ( .A1(n15124), .A2(n9675), .ZN(n15114) );
  AND2_X1 U12546 ( .A1(n11917), .A2(n11918), .ZN(n11931) );
  NOR2_X1 U12547 ( .A1(n17647), .A2(n15602), .ZN(n9681) );
  NOR2_X1 U12548 ( .A1(n10271), .A2(n16117), .ZN(n10272) );
  AND2_X1 U12549 ( .A1(n15065), .A2(n12197), .ZN(n9682) );
  INV_X1 U12550 ( .A(n9870), .ZN(n17434) );
  NAND2_X1 U12551 ( .A1(n9868), .A2(n17443), .ZN(n9870) );
  NAND2_X1 U12552 ( .A1(n11896), .A2(n11900), .ZN(n11968) );
  OR2_X1 U12553 ( .A1(n10176), .A2(n13636), .ZN(n9683) );
  AND2_X1 U12554 ( .A1(n9804), .A2(n9803), .ZN(n9684) );
  NOR2_X1 U12555 ( .A1(n10198), .A2(n12168), .ZN(n9685) );
  AND4_X1 U12556 ( .A1(n10672), .A2(n10671), .A3(n10670), .A4(n10669), .ZN(
        n9686) );
  OAI211_X1 U12557 ( .C1(n20008), .C2(n11872), .A(n11138), .B(n11137), .ZN(
        n11139) );
  INV_X1 U12558 ( .A(n11139), .ZN(n10000) );
  AND2_X1 U12559 ( .A1(n12198), .A2(n9682), .ZN(n9687) );
  AND3_X1 U12560 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10275) );
  INV_X1 U12561 ( .A(n10414), .ZN(n10404) );
  OR2_X1 U12562 ( .A1(n15018), .A2(n14209), .ZN(n9688) );
  NOR2_X1 U12563 ( .A1(n12177), .A2(n15283), .ZN(n9689) );
  NOR2_X1 U12564 ( .A1(n11478), .A2(n11466), .ZN(n13652) );
  AND2_X1 U12565 ( .A1(n15594), .A2(n10031), .ZN(n9690) );
  XOR2_X1 U12566 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12207), .Z(
        n9691) );
  AND4_X1 U12567 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n13075), .ZN(
        n9692) );
  NAND2_X1 U12568 ( .A1(n10338), .A2(n10337), .ZN(n10394) );
  NAND2_X1 U12569 ( .A1(n9902), .A2(n9903), .ZN(n15096) );
  INV_X1 U12570 ( .A(n10613), .ZN(n10043) );
  AND4_X1 U12571 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n9693) );
  AND4_X1 U12572 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n9694) );
  NAND2_X1 U12573 ( .A1(n13764), .A2(n11484), .ZN(n13710) );
  INV_X1 U12574 ( .A(n13195), .ZN(n10156) );
  NAND2_X1 U12575 ( .A1(n12092), .A2(n12091), .ZN(n13822) );
  INV_X1 U12576 ( .A(n9887), .ZN(n11994) );
  AND2_X1 U12577 ( .A1(n15373), .A2(n9916), .ZN(n9695) );
  AND2_X1 U12578 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n9696) );
  AND2_X1 U12579 ( .A1(n12520), .A2(n9774), .ZN(n9697) );
  NAND2_X1 U12580 ( .A1(n14907), .A2(n10048), .ZN(n9698) );
  AND2_X1 U12581 ( .A1(n12327), .A2(n12335), .ZN(n12939) );
  NAND2_X1 U12582 ( .A1(n11771), .A2(n11770), .ZN(n14293) );
  AND2_X1 U12583 ( .A1(n11926), .A2(n11930), .ZN(n9699) );
  AND2_X1 U12584 ( .A1(n10154), .A2(n13195), .ZN(n9700) );
  NAND2_X1 U12585 ( .A1(n14221), .A2(n10230), .ZN(n9701) );
  INV_X1 U12586 ( .A(n15097), .ZN(n9901) );
  INV_X1 U12587 ( .A(n15593), .ZN(n10031) );
  AND2_X1 U12588 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15592), .ZN(
        n15593) );
  NAND2_X1 U12589 ( .A1(n14629), .A2(n15873), .ZN(n9702) );
  AND2_X1 U12590 ( .A1(n10586), .A2(n10585), .ZN(n9703) );
  NAND2_X1 U12591 ( .A1(n10146), .A2(n10145), .ZN(n13684) );
  NAND2_X1 U12592 ( .A1(n10203), .A2(n12111), .ZN(n9704) );
  NAND2_X1 U12593 ( .A1(n11900), .A2(n15462), .ZN(n11913) );
  NAND3_X1 U12594 ( .A1(n11203), .A2(n19999), .A3(n9669), .ZN(n9705) );
  OAI21_X1 U12595 ( .B1(n10179), .B2(n14934), .A(n10178), .ZN(n12497) );
  OR2_X1 U12596 ( .A1(n9683), .A2(n10175), .ZN(n9706) );
  AND2_X1 U12597 ( .A1(n11677), .A2(n10117), .ZN(n9707) );
  NAND2_X1 U12598 ( .A1(n9830), .A2(n12106), .ZN(n15448) );
  AND2_X1 U12599 ( .A1(n11677), .A2(n10118), .ZN(n9708) );
  NAND2_X1 U12600 ( .A1(n11881), .A2(n11879), .ZN(n9709) );
  INV_X1 U12601 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15180) );
  OR2_X1 U12602 ( .A1(n14628), .A2(n15957), .ZN(n9710) );
  AND2_X1 U12603 ( .A1(n11967), .A2(n11966), .ZN(n9711) );
  INV_X1 U12604 ( .A(n12033), .ZN(n9910) );
  NOR2_X1 U12605 ( .A1(n14927), .A2(n14926), .ZN(n9712) );
  AND2_X1 U12606 ( .A1(n10107), .A2(n10500), .ZN(n9713) );
  NAND2_X1 U12607 ( .A1(n12096), .A2(n10107), .ZN(n9714) );
  AND2_X1 U12608 ( .A1(n10174), .A2(n14900), .ZN(n9715) );
  INV_X1 U12609 ( .A(n12081), .ZN(n10098) );
  INV_X1 U12610 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10283) );
  INV_X1 U12611 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13825) );
  BUF_X1 U12612 ( .A(n12870), .Z(n14161) );
  NOR2_X1 U12613 ( .A1(n13059), .A2(n12352), .ZN(n13123) );
  NAND2_X1 U12614 ( .A1(n12814), .A2(n9677), .ZN(n10162) );
  AND2_X1 U12615 ( .A1(n17495), .A2(n9668), .ZN(n9716) );
  NOR2_X1 U12616 ( .A1(n13059), .A2(n9683), .ZN(n13626) );
  INV_X1 U12617 ( .A(n11380), .ZN(n20111) );
  NAND2_X1 U12618 ( .A1(n18732), .A2(n18020), .ZN(n18045) );
  NOR2_X1 U12619 ( .A1(n10268), .A2(n15193), .ZN(n10269) );
  INV_X1 U12620 ( .A(n10455), .ZN(n10476) );
  NOR2_X1 U12621 ( .A1(n10016), .A2(n10271), .ZN(n10270) );
  XNOR2_X1 U12622 ( .A(n14258), .B(n14257), .ZN(n14652) );
  AND2_X1 U12623 ( .A1(n14331), .A2(n9673), .ZN(n9717) );
  AND2_X1 U12624 ( .A1(n10073), .A2(n10072), .ZN(n9718) );
  AND2_X1 U12625 ( .A1(n10162), .A2(n10160), .ZN(n12950) );
  INV_X1 U12626 ( .A(n12065), .ZN(n10100) );
  AND2_X1 U12627 ( .A1(n13803), .A2(n14360), .ZN(n9719) );
  NAND2_X1 U12628 ( .A1(n10220), .A2(n10221), .ZN(n13807) );
  INV_X1 U12629 ( .A(n12091), .ZN(n13722) );
  OR2_X1 U12630 ( .A1(n13328), .A2(n13690), .ZN(n9720) );
  AND2_X1 U12631 ( .A1(n15106), .A2(n15105), .ZN(n9721) );
  AND2_X1 U12632 ( .A1(n12183), .A2(n15262), .ZN(n9722) );
  NOR2_X1 U12633 ( .A1(n12973), .A2(n11112), .ZN(n9723) );
  INV_X1 U12634 ( .A(n11478), .ZN(n13654) );
  AND2_X1 U12635 ( .A1(n15173), .A2(n15175), .ZN(n9724) );
  NAND2_X1 U12636 ( .A1(n11414), .A2(n10113), .ZN(n13588) );
  INV_X1 U12637 ( .A(n13588), .ZN(n10112) );
  AND2_X1 U12638 ( .A1(n10143), .A2(n10142), .ZN(n9725) );
  NOR2_X1 U12639 ( .A1(n9676), .A2(n10064), .ZN(n10069) );
  AND2_X1 U12640 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9726) );
  INV_X1 U12641 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17486) );
  NAND2_X1 U12642 ( .A1(n13644), .A2(n13642), .ZN(n9727) );
  INV_X1 U12643 ( .A(n14285), .ZN(n10123) );
  INV_X1 U12644 ( .A(n14587), .ZN(n11676) );
  NAND2_X1 U12645 ( .A1(n9669), .A2(n11263), .ZN(n9728) );
  AND3_X1 U12646 ( .A1(n11292), .A2(n20756), .A3(n11291), .ZN(n9729) );
  OR2_X1 U12647 ( .A1(n10266), .A2(n10026), .ZN(n9730) );
  INV_X1 U12648 ( .A(n10867), .ZN(n11995) );
  OR2_X1 U12649 ( .A1(n10687), .A2(n10686), .ZN(n10867) );
  NAND2_X1 U12650 ( .A1(n9720), .A2(n10190), .ZN(n9731) );
  AND2_X1 U12651 ( .A1(n10103), .A2(n13663), .ZN(n9732) );
  OR2_X1 U12652 ( .A1(n16539), .A2(n16547), .ZN(n9733) );
  OR2_X1 U12653 ( .A1(n11193), .A2(n11178), .ZN(n9734) );
  AND2_X1 U12654 ( .A1(n9718), .A2(n10071), .ZN(n9735) );
  AND2_X1 U12655 ( .A1(n9921), .A2(n16764), .ZN(n9736) );
  AND2_X1 U12656 ( .A1(n9671), .A2(n9726), .ZN(n9737) );
  INV_X2 U12657 ( .A(n12444), .ZN(n13067) );
  NAND2_X1 U12658 ( .A1(n12765), .A2(n16213), .ZN(n12964) );
  OR3_X1 U12659 ( .A1(n12479), .A2(n12478), .A3(n14929), .ZN(n9738) );
  OR2_X1 U12660 ( .A1(n10255), .A2(n10020), .ZN(n9739) );
  OR2_X1 U12661 ( .A1(n13125), .A2(n10057), .ZN(n13353) );
  NOR2_X1 U12662 ( .A1(n13095), .A2(n10138), .ZN(n9740) );
  NOR2_X1 U12663 ( .A1(n20003), .A2(n20727), .ZN(n9741) );
  NAND2_X1 U12664 ( .A1(n11176), .A2(n11175), .ZN(n20148) );
  INV_X1 U12665 ( .A(n20148), .ZN(n9812) );
  AND2_X1 U12666 ( .A1(n12593), .A2(n12229), .ZN(n12288) );
  XOR2_X1 U12667 ( .A(n13328), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n9742) );
  AND2_X1 U12668 ( .A1(n14344), .A2(n14423), .ZN(n9743) );
  BUF_X1 U12669 ( .A(n10280), .Z(n18891) );
  OAI22_X1 U12670 ( .A1(n13371), .A2(n10248), .B1(n12060), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n18908) );
  AND2_X1 U12671 ( .A1(n12314), .A2(n19720), .ZN(n19056) );
  INV_X1 U12672 ( .A(n19056), .ZN(n16189) );
  INV_X1 U12673 ( .A(n12961), .ZN(n10486) );
  INV_X1 U12674 ( .A(n15408), .ZN(n9827) );
  INV_X1 U12675 ( .A(n17858), .ZN(n16282) );
  INV_X1 U12676 ( .A(n9943), .ZN(n9942) );
  NAND2_X1 U12677 ( .A1(n9944), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9943) );
  AND2_X1 U12678 ( .A1(n10049), .A2(n10562), .ZN(n9744) );
  AND2_X1 U12679 ( .A1(n10132), .A2(n10131), .ZN(n9745) );
  INV_X1 U12680 ( .A(n12079), .ZN(n10194) );
  INV_X1 U12681 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9952) );
  INV_X1 U12682 ( .A(n16134), .ZN(n19040) );
  AND2_X1 U12683 ( .A1(n16264), .A2(n9944), .ZN(n9746) );
  INV_X1 U12684 ( .A(n14236), .ZN(n10052) );
  AND2_X1 U12685 ( .A1(n9675), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9747) );
  NAND2_X1 U12686 ( .A1(n10251), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10249) );
  OR2_X1 U12687 ( .A1(n13550), .A2(n13549), .ZN(n9748) );
  AND2_X1 U12688 ( .A1(n17962), .A2(n10042), .ZN(n9749) );
  NOR2_X1 U12689 ( .A1(n9679), .A2(n15060), .ZN(n10250) );
  NAND2_X1 U12690 ( .A1(n15598), .A2(n15597), .ZN(n9750) );
  AND2_X1 U12691 ( .A1(n10041), .A2(n10040), .ZN(n9751) );
  INV_X1 U12692 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10040) );
  INV_X1 U12693 ( .A(n17252), .ZN(n9815) );
  OR2_X1 U12694 ( .A1(n15200), .A2(n15213), .ZN(n9752) );
  INV_X1 U12695 ( .A(n16745), .ZN(n9919) );
  AND2_X1 U12696 ( .A1(n14737), .A2(n14744), .ZN(n9753) );
  NAND2_X1 U12697 ( .A1(n14729), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9754) );
  INV_X1 U12698 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9946) );
  INV_X1 U12699 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9945) );
  INV_X1 U12700 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n9970) );
  INV_X1 U12701 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9869) );
  INV_X1 U12702 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10002) );
  NOR2_X1 U12703 ( .A1(n18427), .A2(n18100), .ZN(n18481) );
  INV_X1 U12704 ( .A(n16235), .ZN(n18427) );
  AOI22_X2 U12705 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20037), .B1(DATAI_28_), 
        .B2(n20038), .ZN(n20546) );
  AOI22_X2 U12706 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20037), .B1(DATAI_26_), 
        .B2(n20038), .ZN(n20536) );
  AOI22_X2 U12707 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20037), .B1(DATAI_27_), 
        .B2(n20038), .ZN(n20541) );
  NOR2_X2 U12708 ( .A1(n19998), .A2(n19997), .ZN(n20037) );
  NOR2_X2 U12709 ( .A1(n19996), .A2(n19998), .ZN(n20038) );
  NOR3_X2 U12710 ( .A1(n18571), .A2(n18372), .A3(n18347), .ZN(n18342) );
  NAND2_X1 U12711 ( .A1(n19270), .A2(n19269), .ZN(n9758) );
  NOR2_X1 U12712 ( .A1(n19270), .A2(n9760), .ZN(n9759) );
  NOR2_X1 U12713 ( .A1(n19270), .A2(n9762), .ZN(n9761) );
  NAND2_X1 U12714 ( .A1(n9797), .A2(n9764), .ZN(n9763) );
  INV_X1 U12715 ( .A(n11957), .ZN(n9765) );
  INV_X1 U12716 ( .A(n9770), .ZN(n15174) );
  OAI211_X2 U12717 ( .C1(n13822), .C2(n9773), .A(n9771), .B(n10199), .ZN(
        n12121) );
  INV_X1 U12718 ( .A(n12101), .ZN(n9772) );
  NAND2_X1 U12719 ( .A1(n13822), .A2(n12101), .ZN(n9830) );
  NAND2_X2 U12720 ( .A1(n9775), .A2(n12534), .ZN(n14900) );
  NAND3_X1 U12721 ( .A1(n10174), .A2(n14906), .A3(n14900), .ZN(n14905) );
  NOR2_X2 U12722 ( .A1(n13059), .A2(n9706), .ZN(n13627) );
  NAND2_X2 U12723 ( .A1(n14920), .A2(n12501), .ZN(n12517) );
  NAND2_X1 U12724 ( .A1(n14942), .A2(n12459), .ZN(n10177) );
  NAND2_X1 U12725 ( .A1(n11911), .A2(n12337), .ZN(n9777) );
  INV_X2 U12726 ( .A(n9806), .ZN(n14533) );
  INV_X1 U12727 ( .A(n11059), .ZN(n9782) );
  OAI21_X1 U12728 ( .B1(n11043), .B2(n13017), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11136) );
  NAND3_X1 U12729 ( .A1(n9784), .A2(n11056), .A3(n9783), .ZN(n9787) );
  NAND2_X1 U12730 ( .A1(n13017), .A2(n9785), .ZN(n9783) );
  INV_X1 U12731 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9786) );
  AND2_X2 U12732 ( .A1(n9788), .A2(n15372), .ZN(n15373) );
  NAND2_X1 U12733 ( .A1(n9789), .A2(n9734), .ZN(n10001) );
  NAND3_X1 U12734 ( .A1(n9999), .A2(n9786), .A3(n9998), .ZN(n9789) );
  INV_X1 U12735 ( .A(n11140), .ZN(n9790) );
  OR2_X2 U12737 ( .A1(n9653), .A2(n18928), .ZN(n11915) );
  XNOR2_X2 U12738 ( .A(n9886), .B(n11878), .ZN(n11909) );
  NAND2_X1 U12739 ( .A1(n13821), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9792) );
  XNOR2_X2 U12740 ( .A(n12028), .B(n12026), .ZN(n13821) );
  NAND2_X2 U12741 ( .A1(n11285), .A2(n11288), .ZN(n11289) );
  NAND2_X2 U12742 ( .A1(n9881), .A2(n9882), .ZN(n9798) );
  XNOR2_X2 U12743 ( .A(n9798), .B(n9680), .ZN(n10242) );
  NAND3_X1 U12744 ( .A1(n11955), .A2(n11953), .A3(n11954), .ZN(n9797) );
  NAND2_X1 U12745 ( .A1(n9631), .A2(n9905), .ZN(n13688) );
  NAND3_X1 U12746 ( .A1(n9631), .A2(n9905), .A3(n12018), .ZN(n9804) );
  NAND2_X1 U12747 ( .A1(n9812), .A2(n11139), .ZN(n9810) );
  OAI21_X1 U12748 ( .B1(n20148), .B2(n11140), .A(n9809), .ZN(n9808) );
  NAND2_X1 U12749 ( .A1(n9810), .A2(n11140), .ZN(n9809) );
  NOR2_X1 U12750 ( .A1(n9998), .A2(n9812), .ZN(n13293) );
  INV_X2 U12751 ( .A(n17043), .ZN(n13910) );
  AOI22_X1 U12752 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n19433), .ZN(n11951) );
  NAND4_X1 U12753 ( .A1(n10431), .A2(n12592), .A3(n12170), .A4(n10405), .ZN(
        n10406) );
  NAND3_X1 U12754 ( .A1(n9836), .A2(n9839), .A3(n9840), .ZN(n9834) );
  NAND2_X1 U12755 ( .A1(n9837), .A2(n12988), .ZN(n9836) );
  NAND2_X1 U12756 ( .A1(n9841), .A2(n13088), .ZN(n9840) );
  NAND2_X1 U12757 ( .A1(n19935), .A2(n9847), .ZN(n9846) );
  NAND2_X1 U12758 ( .A1(n9850), .A2(n9846), .ZN(n13606) );
  NOR2_X1 U12759 ( .A1(n10214), .A2(n9848), .ZN(n9847) );
  NAND2_X1 U12760 ( .A1(n13606), .A2(n11271), .ZN(n9849) );
  INV_X1 U12761 ( .A(n10213), .ZN(n9850) );
  NOR2_X2 U12762 ( .A1(n17401), .A2(n9853), .ZN(n15619) );
  NAND3_X1 U12763 ( .A1(n18708), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n18695), .ZN(n9854) );
  INV_X2 U12764 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18708) );
  OAI21_X1 U12765 ( .B1(n17673), .B2(n9858), .A(n9859), .ZN(n9857) );
  OR2_X1 U12766 ( .A1(n17672), .A2(n15594), .ZN(n9858) );
  NAND2_X1 U12767 ( .A1(n9871), .A2(n9873), .ZN(n15604) );
  OR2_X1 U12768 ( .A1(n17981), .A2(n17648), .ZN(n9875) );
  XNOR2_X2 U12769 ( .A(n10473), .B(n10475), .ZN(n11878) );
  OAI21_X1 U12770 ( .B1(n9880), .B2(n13821), .A(n9878), .ZN(n9908) );
  NAND3_X1 U12771 ( .A1(n9699), .A2(n11928), .A3(n11927), .ZN(n9881) );
  NAND2_X1 U12772 ( .A1(n11930), .A2(n19737), .ZN(n9882) );
  NAND2_X2 U12773 ( .A1(n15124), .A2(n9883), .ZN(n15083) );
  NAND4_X1 U12774 ( .A1(n10405), .A2(n10392), .A3(n10393), .A4(n12280), .ZN(
        n10564) );
  NAND3_X1 U12775 ( .A1(n10392), .A2(n10393), .A3(n10405), .ZN(n10396) );
  NAND2_X1 U12776 ( .A1(n9885), .A2(n12701), .ZN(n13254) );
  NAND2_X1 U12777 ( .A1(n11878), .A2(n9886), .ZN(n10055) );
  XNOR2_X1 U12778 ( .A(n10195), .B(n9887), .ZN(n12064) );
  AND2_X2 U12779 ( .A1(n9907), .A2(n9906), .ZN(n15186) );
  NAND2_X2 U12780 ( .A1(n9908), .A2(n12033), .ZN(n15124) );
  NAND2_X1 U12781 ( .A1(n15373), .A2(n9913), .ZN(n9912) );
  NAND2_X1 U12782 ( .A1(n15373), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15162) );
  NAND2_X1 U12783 ( .A1(n17605), .A2(n9737), .ZN(n17520) );
  NAND2_X1 U12784 ( .A1(n9920), .A2(n9921), .ZN(n16537) );
  INV_X1 U12785 ( .A(n9922), .ZN(n16545) );
  AOI21_X1 U12786 ( .B1(n16521), .B2(n9928), .A(n9926), .ZN(n9925) );
  INV_X1 U12787 ( .A(n9923), .ZN(n16501) );
  AOI22_X1 U12788 ( .A1(n16521), .A2(n9924), .B1(n9926), .B2(n17421), .ZN(
        n9923) );
  AND2_X1 U12789 ( .A1(n17421), .A2(n9928), .ZN(n9924) );
  NAND2_X1 U12790 ( .A1(n9935), .A2(n9929), .ZN(P3_U2640) );
  NOR2_X1 U12791 ( .A1(n16457), .A2(n16734), .ZN(n16449) );
  NAND3_X1 U12792 ( .A1(n16264), .A2(n16447), .A3(n9942), .ZN(n9939) );
  NAND2_X1 U12793 ( .A1(n9953), .A2(n19988), .ZN(n14700) );
  CLKBUF_X1 U12794 ( .A(n9968), .Z(n9954) );
  INV_X1 U12795 ( .A(n9968), .ZN(n14158) );
  NAND2_X4 U12796 ( .A1(n9968), .A2(n12870), .ZN(n14180) );
  NAND2_X1 U12797 ( .A1(n9954), .A2(n13088), .ZN(n13089) );
  NAND2_X1 U12798 ( .A1(n9954), .A2(n13747), .ZN(n13748) );
  NAND2_X1 U12799 ( .A1(n9954), .A2(n15936), .ZN(n13753) );
  NAND2_X1 U12800 ( .A1(n9954), .A2(n14751), .ZN(n14140) );
  NAND2_X1 U12801 ( .A1(n9954), .A2(n14737), .ZN(n14146) );
  NAND2_X1 U12802 ( .A1(n9954), .A2(n14705), .ZN(n14152) );
  OAI22_X1 U12803 ( .A1(n14161), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n12871), .B2(
        n9968), .ZN(n12997) );
  OAI211_X1 U12804 ( .C1(n14168), .C2(P1_EBX_REG_6__SCAN_IN), .A(n13544), .B(
        n9954), .ZN(n13545) );
  OAI211_X1 U12805 ( .C1(n14168), .C2(P1_EBX_REG_8__SCAN_IN), .A(n13582), .B(
        n9954), .ZN(n13583) );
  OAI21_X1 U12806 ( .B1(n14168), .B2(P1_EBX_REG_4__SCAN_IN), .A(n9968), .ZN(
        n9958) );
  OAI21_X1 U12807 ( .B1(n14168), .B2(P1_EBX_REG_12__SCAN_IN), .A(n9954), .ZN(
        n9960) );
  OAI21_X1 U12808 ( .B1(n14168), .B2(P1_EBX_REG_20__SCAN_IN), .A(n9954), .ZN(
        n9962) );
  OAI21_X1 U12809 ( .B1(n14168), .B2(P1_EBX_REG_18__SCAN_IN), .A(n9954), .ZN(
        n9964) );
  OAI21_X1 U12810 ( .B1(n12998), .B2(P1_EBX_REG_22__SCAN_IN), .A(n9954), .ZN(
        n9966) );
  NAND2_X1 U12811 ( .A1(n9954), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n9967) );
  CLKBUF_X1 U12812 ( .A(n11616), .Z(n9971) );
  NOR2_X1 U12813 ( .A1(n14788), .A2(n9729), .ZN(n10003) );
  NAND3_X1 U12814 ( .A1(n11203), .A2(n19999), .A3(n11224), .ZN(n11249) );
  NAND2_X1 U12815 ( .A1(n10461), .A2(n10460), .ZN(n11881) );
  NAND2_X2 U12816 ( .A1(n10007), .A2(n11885), .ZN(n11889) );
  NAND3_X1 U12817 ( .A1(n10007), .A2(n11885), .A3(n11880), .ZN(n10005) );
  INV_X1 U12818 ( .A(n11884), .ZN(n10007) );
  AOI21_X2 U12819 ( .B1(n10012), .B2(n10011), .A(n10008), .ZN(n15394) );
  NAND2_X2 U12820 ( .A1(n10013), .A2(n12022), .ZN(n12028) );
  NAND2_X1 U12821 ( .A1(n13721), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10013) );
  INV_X1 U12822 ( .A(n10271), .ZN(n10014) );
  NAND3_X1 U12823 ( .A1(n10015), .A2(n10014), .A3(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10268) );
  NOR2_X1 U12824 ( .A1(n10255), .A2(n10246), .ZN(n10256) );
  AND3_X1 U12825 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10021) );
  NOR2_X2 U12826 ( .A1(n14849), .A2(n15053), .ZN(n14848) );
  AND2_X2 U12827 ( .A1(n10022), .A2(n9642), .ZN(n14849) );
  OR2_X2 U12828 ( .A1(n10266), .A2(n10023), .ZN(n10258) );
  INV_X1 U12829 ( .A(n10027), .ZN(n15679) );
  NOR2_X2 U12830 ( .A1(n14876), .A2(n15100), .ZN(n14875) );
  INV_X1 U12831 ( .A(n10029), .ZN(n18809) );
  INV_X1 U12832 ( .A(n18808), .ZN(n10028) );
  NAND2_X1 U12833 ( .A1(n15619), .A2(n10033), .ZN(n16293) );
  AOI21_X2 U12834 ( .B1(n15723), .B2(n16293), .A(n16285), .ZN(n15620) );
  NAND2_X1 U12835 ( .A1(n17712), .A2(n17713), .ZN(n17711) );
  NAND2_X1 U12836 ( .A1(n17712), .A2(n10038), .ZN(n10037) );
  OR2_X1 U12837 ( .A1(n17713), .A2(n10039), .ZN(n10038) );
  NOR2_X1 U12838 ( .A1(n17696), .A2(n17697), .ZN(n17695) );
  INV_X1 U12839 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10039) );
  INV_X2 U12840 ( .A(n12596), .ZN(n10634) );
  NAND2_X1 U12841 ( .A1(n14907), .A2(n10049), .ZN(n14238) );
  NAND2_X1 U12842 ( .A1(n14907), .A2(n9744), .ZN(n10044) );
  NAND2_X1 U12843 ( .A1(n14907), .A2(n14853), .ZN(n14855) );
  INV_X1 U12844 ( .A(n10056), .ZN(n10054) );
  NAND2_X1 U12845 ( .A1(n10241), .A2(n13054), .ZN(n10056) );
  NAND3_X1 U12846 ( .A1(n10054), .A2(n10055), .A3(n12962), .ZN(n12961) );
  INV_X1 U12847 ( .A(n10069), .ZN(n14915) );
  INV_X1 U12848 ( .A(n14879), .ZN(n10070) );
  INV_X1 U12849 ( .A(n12043), .ZN(n10866) );
  NOR2_X1 U12850 ( .A1(n10079), .A2(n10078), .ZN(n10077) );
  INV_X1 U12851 ( .A(n10666), .ZN(n10079) );
  AOI21_X1 U12852 ( .B1(n12577), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n10084), .ZN(n12467) );
  NOR2_X1 U12853 ( .A1(n15018), .A2(n15019), .ZN(n10094) );
  NOR2_X1 U12854 ( .A1(n10098), .A2(n12074), .ZN(n10097) );
  NAND3_X1 U12855 ( .A1(n12081), .A2(n10099), .A3(n10096), .ZN(n12089) );
  NOR2_X1 U12856 ( .A1(n12075), .A2(n12074), .ZN(n12076) );
  NOR2_X2 U12857 ( .A1(n12153), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10102) );
  NAND2_X1 U12858 ( .A1(n12113), .A2(n9732), .ZN(n12130) );
  NAND2_X1 U12859 ( .A1(n12096), .A2(n9713), .ZN(n12118) );
  NAND2_X1 U12860 ( .A1(n10112), .A2(n10111), .ZN(n11478) );
  AOI21_X1 U12861 ( .B1(n11448), .B2(n11569), .A(n11447), .ZN(n13534) );
  INV_X1 U12862 ( .A(n13589), .ZN(n10113) );
  NAND2_X1 U12863 ( .A1(n11677), .A2(n10116), .ZN(n14292) );
  NAND3_X1 U12864 ( .A1(n11370), .A2(n11385), .A3(n11386), .ZN(n12984) );
  NAND2_X1 U12865 ( .A1(n12984), .A2(n11386), .ZN(n13086) );
  INV_X1 U12866 ( .A(n14293), .ZN(n10124) );
  INV_X1 U12867 ( .A(n13095), .ZN(n10136) );
  NAND2_X2 U12868 ( .A1(n16143), .A2(n11993), .ZN(n13477) );
  AND2_X1 U12869 ( .A1(n15068), .A2(n10147), .ZN(n15025) );
  NAND2_X1 U12870 ( .A1(n15068), .A2(n10148), .ZN(n12037) );
  NOR2_X2 U12871 ( .A1(n15002), .A2(n15003), .ZN(n15001) );
  INV_X1 U12872 ( .A(n14881), .ZN(n10150) );
  NOR2_X2 U12873 ( .A1(n13178), .A2(n10152), .ZN(n13697) );
  NOR2_X1 U12874 ( .A1(n13177), .A2(n13176), .ZN(n13178) );
  NAND2_X1 U12875 ( .A1(n13466), .A2(n10168), .ZN(n13855) );
  NAND2_X1 U12876 ( .A1(n10177), .A2(n9738), .ZN(n10179) );
  NOR2_X1 U12877 ( .A1(n15074), .A2(n15075), .ZN(n15064) );
  NAND2_X1 U12878 ( .A1(n12086), .A2(n10189), .ZN(n13723) );
  NAND2_X1 U12879 ( .A1(n10197), .A2(n15291), .ZN(n10196) );
  INV_X1 U12880 ( .A(n12169), .ZN(n10197) );
  INV_X1 U12881 ( .A(n15291), .ZN(n10198) );
  OAI21_X1 U12882 ( .B1(n15188), .B2(n12169), .A(n12168), .ZN(n15293) );
  INV_X1 U12883 ( .A(n15018), .ZN(n10205) );
  NAND2_X1 U12884 ( .A1(n12199), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10207) );
  NAND2_X1 U12885 ( .A1(n14533), .A2(n9667), .ZN(n14508) );
  NAND2_X1 U12886 ( .A1(n10209), .A2(n10208), .ZN(n11306) );
  NAND2_X1 U12887 ( .A1(n14533), .A2(n9672), .ZN(n10208) );
  NAND3_X1 U12888 ( .A1(n10211), .A2(n10212), .A3(n11305), .ZN(n10209) );
  NAND2_X1 U12889 ( .A1(n14533), .A2(n11304), .ZN(n10212) );
  OAI21_X1 U12890 ( .B1(n10214), .B2(n11223), .A(n11247), .ZN(n10213) );
  NAND2_X1 U12891 ( .A1(n11043), .A2(n10218), .ZN(n10217) );
  AOI21_X1 U12892 ( .B1(n13017), .B2(n10218), .A(n10216), .ZN(n10215) );
  NAND3_X1 U12893 ( .A1(n13667), .A2(n10224), .A3(n11284), .ZN(n10221) );
  OR2_X1 U12894 ( .A1(n13783), .A2(n10223), .ZN(n10222) );
  NAND2_X1 U12895 ( .A1(n13666), .A2(n11284), .ZN(n10223) );
  NAND2_X1 U12896 ( .A1(n13669), .A2(n11284), .ZN(n13785) );
  OR2_X1 U12897 ( .A1(n15057), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15226) );
  NAND2_X1 U12898 ( .A1(n15057), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15225) );
  INV_X1 U12899 ( .A(n13831), .ZN(n12431) );
  OR3_X1 U12900 ( .A1(n11331), .A2(n13019), .A3(n11325), .ZN(n11355) );
  NAND2_X1 U12901 ( .A1(n12346), .A2(n13048), .ZN(n13062) );
  NOR2_X1 U12902 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  AND2_X2 U12903 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12928) );
  INV_X1 U12904 ( .A(n11931), .ZN(n19360) );
  NAND2_X1 U12905 ( .A1(n11910), .A2(n11919), .ZN(n11943) );
  INV_X1 U12906 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U12907 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10320) );
  NOR2_X4 U12908 ( .A1(n13467), .A2(n13468), .ZN(n13466) );
  CLKBUF_X1 U12909 ( .A(n12882), .Z(n15984) );
  NAND2_X1 U12910 ( .A1(n18939), .A2(n18922), .ZN(n10889) );
  AND2_X2 U12911 ( .A1(n11950), .A2(n11918), .ZN(n11960) );
  NAND2_X1 U12912 ( .A1(n12336), .A2(n12335), .ZN(n13045) );
  XNOR2_X1 U12913 ( .A(n10658), .B(n10657), .ZN(n13177) );
  NAND2_X1 U12914 ( .A1(n11172), .A2(n11171), .ZN(n11202) );
  XNOR2_X1 U12915 ( .A(n11171), .B(n11170), .ZN(n11364) );
  AND2_X4 U12916 ( .A1(n10900), .A2(n10903), .ZN(n10930) );
  INV_X2 U12917 ( .A(n10613), .ZN(n12270) );
  AND2_X1 U12918 ( .A1(n12349), .A2(n12348), .ZN(n10227) );
  AND2_X1 U12919 ( .A1(n10889), .A2(n10888), .ZN(n10228) );
  NAND2_X1 U12920 ( .A1(n19873), .A2(n14461), .ZN(n14448) );
  NOR2_X1 U12921 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13877), .ZN(
        n15534) );
  CLKBUF_X3 U12922 ( .A(n14076), .Z(n17041) );
  INV_X1 U12923 ( .A(n10466), .ZN(n10506) );
  NAND2_X2 U12924 ( .A1(n12288), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10464) );
  OR2_X1 U12925 ( .A1(n15201), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10229) );
  OR2_X1 U12926 ( .A1(n15035), .A2(n16188), .ZN(n10230) );
  AND2_X1 U12927 ( .A1(n12314), .A2(n12269), .ZN(n16200) );
  OR2_X1 U12928 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20750), .ZN(n10231) );
  INV_X2 U12929 ( .A(n18740), .ZN(n18669) );
  OR2_X1 U12930 ( .A1(n14180), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10232) );
  AND2_X1 U12931 ( .A1(n10245), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10233) );
  OR2_X1 U12932 ( .A1(n10440), .A2(n19705), .ZN(n10234) );
  AND2_X1 U12933 ( .A1(n12617), .A2(n10416), .ZN(n10235) );
  AND3_X1 U12934 ( .A1(n10332), .A2(n10331), .A3(n13075), .ZN(n10236) );
  OR2_X1 U12935 ( .A1(n12354), .A2(n13342), .ZN(n10237) );
  INV_X1 U12936 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n18920) );
  AND2_X1 U12937 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10238) );
  OR2_X1 U12938 ( .A1(n19601), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19745) );
  INV_X1 U12939 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15193) );
  INV_X1 U12940 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19774) );
  INV_X1 U12941 ( .A(n9642), .ZN(n10280) );
  INV_X1 U12942 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12319) );
  INV_X1 U12943 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11003) );
  NOR2_X1 U12944 ( .A1(n18685), .A2(n18556), .ZN(n13885) );
  NAND2_X1 U12945 ( .A1(n19682), .A2(n13266), .ZN(n18900) );
  NOR3_X1 U12946 ( .A1(n18683), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n16286) );
  INV_X1 U12947 ( .A(n9637), .ZN(n18032) );
  INV_X1 U12948 ( .A(n9637), .ZN(n18017) );
  INV_X1 U12949 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13528) );
  NAND3_X1 U12950 ( .A1(n10485), .A2(n10484), .A3(n10483), .ZN(n10240) );
  OR2_X1 U12951 ( .A1(n10475), .A2(n10474), .ZN(n10241) );
  INV_X1 U12952 ( .A(n11885), .ZN(n11898) );
  AND2_X2 U12953 ( .A1(n10899), .A2(n10901), .ZN(n11095) );
  AND4_X1 U12954 ( .A1(n11051), .A2(n12906), .A3(n11031), .A4(n12778), .ZN(
        n10244) );
  AOI22_X1 U12955 ( .A1(n11958), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11959), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11942) );
  INV_X1 U12956 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10890) );
  AND2_X1 U12957 ( .A1(n20464), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11328) );
  BUF_X2 U12958 ( .A(n10984), .Z(n11840) );
  OR2_X1 U12959 ( .A1(n11215), .A2(n11214), .ZN(n11239) );
  AND4_X1 U12960 ( .A1(n11051), .A2(n13028), .A3(n11050), .A4(n11049), .ZN(
        n11054) );
  OR2_X1 U12961 ( .A1(n11076), .A2(n11075), .ZN(n11088) );
  NAND2_X1 U12962 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10293) );
  INV_X1 U12963 ( .A(n10430), .ZN(n10432) );
  NAND2_X1 U12964 ( .A1(n10404), .A2(n13383), .ZN(n10418) );
  INV_X1 U12965 ( .A(n11902), .ZN(n11895) );
  OR2_X1 U12966 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19995), .ZN(
        n11316) );
  INV_X1 U12967 ( .A(n13594), .ZN(n11428) );
  NAND2_X1 U12968 ( .A1(n11262), .A2(n11261), .ZN(n11263) );
  NOR2_X1 U12969 ( .A1(n11115), .A2(n20759), .ZN(n11287) );
  NAND2_X1 U12970 ( .A1(n11113), .A2(n11112), .ZN(n11356) );
  OR2_X1 U12971 ( .A1(n11190), .A2(n11189), .ZN(n11240) );
  INV_X1 U12972 ( .A(n12518), .ZN(n12519) );
  AND3_X1 U12973 ( .A1(n10285), .A2(n10284), .A3(n13075), .ZN(n10291) );
  NAND2_X1 U12974 ( .A1(n10421), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10444) );
  AND2_X1 U12975 ( .A1(n10301), .A2(n10300), .ZN(n10302) );
  AOI21_X1 U12976 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18561), .A(
        n13960), .ZN(n13961) );
  NAND2_X1 U12977 ( .A1(n11028), .A2(n11027), .ZN(n11032) );
  INV_X1 U12978 ( .A(n11631), .ZN(n11632) );
  NOR2_X1 U12979 ( .A1(n12907), .A2(n13713), .ZN(n13022) );
  AND3_X1 U12980 ( .A1(n12905), .A2(n12904), .A3(n12903), .ZN(n13029) );
  OR2_X1 U12981 ( .A1(n11159), .A2(n11178), .ZN(n11077) );
  OR2_X1 U12982 ( .A1(n11356), .A2(n11114), .ZN(n11118) );
  INV_X1 U12983 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10246) );
  NAND2_X1 U12984 ( .A1(n12517), .A2(n12519), .ZN(n12520) );
  INV_X1 U12985 ( .A(n12498), .ZN(n12499) );
  INV_X1 U12986 ( .A(n12570), .ZN(n12578) );
  AND2_X1 U12987 ( .A1(n10314), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10318) );
  INV_X1 U12988 ( .A(n15047), .ZN(n12194) );
  AND2_X1 U12989 ( .A1(n12132), .A2(n15156), .ZN(n15108) );
  OR2_X1 U12990 ( .A1(n12658), .A2(n12025), .ZN(n12163) );
  INV_X1 U12991 ( .A(n16104), .ZN(n12111) );
  INV_X1 U12992 ( .A(n10451), .ZN(n10452) );
  NOR2_X1 U12993 ( .A1(n13961), .A2(n18685), .ZN(n13965) );
  INV_X1 U12994 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n20929) );
  INV_X1 U12995 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20848) );
  INV_X1 U12996 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n20943) );
  INV_X1 U12997 ( .A(n13020), .ZN(n12745) );
  INV_X1 U12998 ( .A(n14173), .ZN(n14385) );
  INV_X1 U12999 ( .A(n11805), .ZN(n11865) );
  XNOR2_X1 U13000 ( .A(n11871), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14129) );
  INV_X1 U13001 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14309) );
  OR2_X1 U13002 ( .A1(n13652), .A2(n13765), .ZN(n13766) );
  INV_X1 U13003 ( .A(n14113), .ZN(n11858) );
  AND2_X1 U13004 ( .A1(n14148), .A2(n14147), .ZN(n14415) );
  AND2_X1 U13005 ( .A1(n12898), .A2(n13007), .ZN(n13032) );
  AND2_X1 U13006 ( .A1(n12737), .A2(n20014), .ZN(n13284) );
  INV_X1 U13007 ( .A(n20389), .ZN(n20567) );
  AND2_X1 U13008 ( .A1(n20388), .A2(n11135), .ZN(n20008) );
  INV_X1 U13009 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20428) );
  NOR2_X1 U13010 ( .A1(n18918), .A2(n19671), .ZN(n10886) );
  AND2_X1 U13011 ( .A1(n13389), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12174) );
  NAND2_X2 U13012 ( .A1(n12096), .A2(n12270), .ZN(n12186) );
  AND3_X1 U13013 ( .A1(n10489), .A2(n10488), .A3(n10487), .ZN(n13124) );
  NAND2_X1 U13014 ( .A1(n12500), .A2(n12499), .ZN(n12501) );
  AND3_X1 U13015 ( .A1(n10517), .A2(n10516), .A3(n10515), .ZN(n13704) );
  AND3_X1 U13016 ( .A1(n10493), .A2(n10492), .A3(n10491), .ZN(n13106) );
  AND2_X1 U13017 ( .A1(n15273), .A2(n12294), .ZN(n15249) );
  INV_X1 U13018 ( .A(n15108), .ZN(n15166) );
  NOR2_X1 U13019 ( .A1(n13451), .A2(n19736), .ZN(n19298) );
  AND2_X1 U13020 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19296), .ZN(
        n12338) );
  AOI22_X1 U13021 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18563), .B1(
        n13967), .B2(n13966), .ZN(n14006) );
  INV_X1 U13022 ( .A(n15487), .ZN(n15502) );
  OR2_X1 U13023 ( .A1(n14009), .A2(n18520), .ZN(n13997) );
  INV_X1 U13024 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15583) );
  NOR2_X1 U13025 ( .A1(n15585), .A2(n17722), .ZN(n17712) );
  NAND4_X1 U13026 ( .A1(n15635), .A2(n17118), .A3(n13999), .A4(n18082), .ZN(
        n17302) );
  INV_X1 U13027 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15820) );
  NOR2_X1 U13028 ( .A1(n20945), .A2(n11442), .ZN(n11443) );
  INV_X1 U13029 ( .A(n19853), .ZN(n19819) );
  AND2_X1 U13030 ( .A1(n11635), .A2(n11634), .ZN(n14342) );
  NAND2_X1 U13031 ( .A1(n11033), .A2(n20029), .ZN(n12973) );
  INV_X1 U13032 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20839) );
  INV_X1 U13033 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15786) );
  INV_X1 U13034 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14644) );
  AND3_X1 U13035 ( .A1(n11441), .A2(n11440), .A3(n11439), .ZN(n13580) );
  AND2_X1 U13036 ( .A1(n12888), .A2(n12780), .ZN(n15700) );
  NAND2_X1 U13037 ( .A1(n19961), .A2(n19985), .ZN(n19965) );
  OAI21_X1 U13038 ( .B1(n20765), .B2(n13298), .A(n15714), .ZN(n20000) );
  AND2_X1 U13039 ( .A1(n11363), .A2(n11362), .ZN(n13008) );
  AND2_X1 U13040 ( .A1(n20181), .A2(n20180), .ZN(n20208) );
  INV_X1 U13041 ( .A(n19999), .ZN(n20151) );
  AND2_X1 U13042 ( .A1(n20393), .A2(n20392), .ZN(n20421) );
  NOR2_X1 U13043 ( .A1(n20155), .A2(n20154), .ZN(n20522) );
  AND2_X1 U13044 ( .A1(n20580), .A2(n20579), .ZN(n20637) );
  OR2_X1 U13045 ( .A1(n13292), .A2(n13291), .ZN(n15699) );
  OR2_X1 U13046 ( .A1(n14889), .A2(n18878), .ZN(n10585) );
  AND2_X1 U13047 ( .A1(n12248), .A2(n10583), .ZN(n13241) );
  NAND2_X1 U13048 ( .A1(n12323), .A2(n13408), .ZN(n13050) );
  OAI21_X1 U13049 ( .B1(n12607), .B2(n12606), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12608) );
  INV_X1 U13050 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15081) );
  AND2_X1 U13051 ( .A1(n12302), .A2(n12301), .ZN(n15452) );
  INV_X1 U13052 ( .A(n16200), .ZN(n19070) );
  INV_X1 U13053 ( .A(n15397), .ZN(n18885) );
  AND2_X1 U13054 ( .A1(n13180), .A2(n13179), .ZN(n19692) );
  NAND2_X1 U13055 ( .A1(n18928), .A2(n12337), .ZN(n12329) );
  NAND2_X1 U13056 ( .A1(n12253), .A2(n12251), .ZN(n13248) );
  OR2_X1 U13057 ( .A1(n19120), .A2(n19117), .ZN(n19154) );
  INV_X1 U13058 ( .A(n19077), .ZN(n19265) );
  NAND2_X1 U13059 ( .A1(n13554), .A2(n19076), .ZN(n19208) );
  AND2_X1 U13060 ( .A1(n19697), .A2(n19699), .ZN(n19472) );
  INV_X1 U13061 ( .A(n19472), .ZN(n19474) );
  INV_X2 U13062 ( .A(n12270), .ZN(n13389) );
  NOR2_X1 U13063 ( .A1(n18732), .A2(n18082), .ZN(n15640) );
  NOR2_X1 U13064 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16592), .ZN(n16577) );
  NOR2_X1 U13065 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16619), .ZN(n16600) );
  NOR2_X1 U13066 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16663), .ZN(n16647) );
  INV_X1 U13067 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16741) );
  NAND2_X1 U13068 ( .A1(n18746), .A2(n18082), .ZN(n16427) );
  INV_X1 U13069 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17036) );
  AOI211_X1 U13070 ( .C1(n13910), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n15494), .B(n15493), .ZN(n15495) );
  INV_X1 U13071 ( .A(n17110), .ZN(n17259) );
  INV_X1 U13072 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17422) );
  INV_X1 U13073 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17563) );
  INV_X1 U13074 ( .A(n16254), .ZN(n17755) );
  NOR2_X1 U13075 ( .A1(n16283), .A2(n17806), .ZN(n17759) );
  INV_X1 U13076 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17446) );
  INV_X2 U13077 ( .A(n18524), .ZN(n18537) );
  INV_X1 U13078 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17664) );
  NOR2_X1 U13079 ( .A1(n17972), .A2(n18548), .ZN(n18020) );
  NAND2_X1 U13080 ( .A1(n18744), .A2(n15641), .ZN(n18039) );
  NOR2_X1 U13081 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18080), .ZN(n18374) );
  NOR2_X1 U13082 ( .A1(n13916), .A2(n13915), .ZN(n17115) );
  INV_X1 U13083 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18572) );
  INV_X1 U13084 ( .A(n13008), .ZN(n13001) );
  AND2_X1 U13085 ( .A1(n20759), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20754) );
  AND2_X1 U13086 ( .A1(n19827), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19853) );
  OR2_X1 U13087 ( .A1(n20752), .A2(n14115), .ZN(n19827) );
  NOR2_X1 U13088 ( .A1(n19753), .A2(n19836), .ZN(n19776) );
  INV_X1 U13089 ( .A(n14448), .ZN(n19869) );
  INV_X1 U13090 ( .A(n14504), .ZN(n14234) );
  NAND2_X2 U13091 ( .A1(n12972), .A2(n13012), .ZN(n15863) );
  INV_X2 U13092 ( .A(n19875), .ZN(n19901) );
  NAND2_X1 U13093 ( .A1(n11514), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11593) );
  AND2_X1 U13094 ( .A1(n14440), .A2(n14439), .ZN(n15889) );
  NAND2_X1 U13095 ( .A1(n11480), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11557) );
  INV_X1 U13096 ( .A(n15914), .ZN(n19932) );
  AND3_X1 U13097 ( .A1(n15700), .A2(n13012), .A3(n13001), .ZN(n19939) );
  AND2_X1 U13098 ( .A1(n20725), .A2(n20754), .ZN(n19938) );
  AND2_X1 U13099 ( .A1(n14703), .A2(n14188), .ZN(n14773) );
  INV_X1 U13100 ( .A(n15922), .ZN(n19944) );
  NOR2_X2 U13101 ( .A1(n13025), .A2(n13024), .ZN(n19974) );
  INV_X1 U13102 ( .A(n13025), .ZN(n13033) );
  NOR2_X1 U13103 ( .A1(n20301), .A2(n13008), .ZN(n20719) );
  OAI22_X1 U13104 ( .A1(n20011), .A2(n20010), .B1(n20358), .B2(n20150), .ZN(
        n20043) );
  INV_X1 U13105 ( .A(n20107), .ZN(n20065) );
  OAI22_X1 U13106 ( .A1(n20080), .A2(n20079), .B1(n20358), .B2(n20221), .ZN(
        n20103) );
  OR2_X1 U13107 ( .A1(n20730), .A2(n20292), .ZN(n20115) );
  OAI21_X1 U13108 ( .B1(n20173), .B2(n20156), .A(n20522), .ZN(n20174) );
  INV_X1 U13109 ( .A(n20250), .ZN(n20211) );
  OR2_X1 U13110 ( .A1(n9654), .A2(n20350), .ZN(n20294) );
  OAI22_X1 U13111 ( .A1(n20223), .A2(n20222), .B1(n20512), .B2(n20221), .ZN(
        n20246) );
  INV_X1 U13112 ( .A(n20284), .ZN(n20318) );
  INV_X1 U13113 ( .A(n20387), .ZN(n20345) );
  OAI22_X1 U13114 ( .A1(n20360), .A2(n20359), .B1(n20511), .B2(n20358), .ZN(
        n20383) );
  INV_X1 U13115 ( .A(n9650), .ZN(n20350) );
  OAI22_X1 U13116 ( .A1(n20440), .A2(n20439), .B1(n20512), .B2(n20438), .ZN(
        n20456) );
  AND2_X1 U13117 ( .A1(n20571), .A2(n20429), .ZN(n20505) );
  NOR2_X1 U13118 ( .A1(n20015), .A2(n20154), .ZN(n20527) );
  NOR2_X1 U13119 ( .A1(n20030), .A2(n20154), .ZN(n20547) );
  INV_X1 U13120 ( .A(n9654), .ZN(n20461) );
  AND2_X1 U13121 ( .A1(n20571), .A2(n20516), .ZN(n20642) );
  INV_X1 U13122 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n14128) );
  INV_X1 U13123 ( .A(n20661), .ZN(n20751) );
  INV_X1 U13124 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20659) );
  INV_X1 U13125 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19733) );
  INV_X1 U13126 ( .A(n18925), .ZN(n18901) );
  INV_X1 U13127 ( .A(n18918), .ZN(n18829) );
  OR2_X1 U13128 ( .A1(n12644), .A2(n10560), .ZN(n18925) );
  INV_X1 U13129 ( .A(n18883), .ZN(n18912) );
  OR2_X1 U13130 ( .A1(n10791), .A2(n10790), .ZN(n13343) );
  OR2_X1 U13131 ( .A1(n13307), .A2(n13306), .ZN(n13361) );
  INV_X1 U13132 ( .A(n12588), .ZN(n12589) );
  OR2_X1 U13133 ( .A1(n18983), .A2(n12617), .ZN(n18967) );
  INV_X1 U13134 ( .A(n18967), .ZN(n18984) );
  AND2_X1 U13135 ( .A1(n13357), .A2(n13356), .ZN(n18844) );
  AND2_X1 U13136 ( .A1(n16151), .A2(n12679), .ZN(n16142) );
  AND2_X1 U13137 ( .A1(n15329), .A2(n16169), .ZN(n16153) );
  AND2_X1 U13138 ( .A1(n12259), .A2(n16213), .ZN(n12314) );
  INV_X1 U13139 ( .A(n19680), .ZN(n13574) );
  INV_X1 U13140 ( .A(n19107), .ZN(n19112) );
  NOR2_X1 U13141 ( .A1(n13451), .A2(n18989), .ZN(n19077) );
  NOR2_X2 U13142 ( .A1(n19367), .A2(n19302), .ZN(n19189) );
  NOR2_X2 U13143 ( .A1(n19265), .A2(n19208), .ZN(n19224) );
  NOR2_X2 U13144 ( .A1(n19265), .A2(n19474), .ZN(n19251) );
  NOR2_X2 U13145 ( .A1(n19302), .A2(n19474), .ZN(n19290) );
  NOR2_X1 U13146 ( .A1(n19266), .A2(n19265), .ZN(n19321) );
  AND2_X1 U13147 ( .A1(n19697), .A2(n19076), .ZN(n19303) );
  INV_X1 U13148 ( .A(n19354), .ZN(n19382) );
  NOR2_X2 U13149 ( .A1(n19475), .A2(n19367), .ZN(n19412) );
  OR3_X1 U13150 ( .A1(n13450), .A2(n13454), .A3(n13449), .ZN(n19430) );
  NOR2_X1 U13151 ( .A1(n19435), .A2(n19474), .ZN(n19501) );
  NAND2_X1 U13152 ( .A1(n13375), .A2(n13374), .ZN(n19516) );
  NOR2_X1 U13153 ( .A1(n13528), .A2(n19733), .ZN(n19711) );
  INV_X1 U13154 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19619) );
  INV_X1 U13155 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19601) );
  NOR2_X1 U13156 ( .A1(n18530), .A2(n16421), .ZN(n18512) );
  NOR2_X1 U13157 ( .A1(n16799), .A2(n16440), .ZN(n16469) );
  NOR2_X1 U13158 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16528), .ZN(n16513) );
  NOR2_X1 U13159 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16565), .ZN(n16555) );
  NOR2_X1 U13160 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16636), .ZN(n16626) );
  INV_X1 U13161 ( .A(n16701), .ZN(n16730) );
  NOR2_X2 U13162 ( .A1(n18679), .A2(n16792), .ZN(n16784) );
  NAND2_X1 U13163 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16916), .ZN(n16900) );
  NOR2_X1 U13164 ( .A1(n16671), .A2(n17020), .ZN(n17007) );
  INV_X1 U13165 ( .A(n15739), .ZN(n13981) );
  NAND2_X1 U13166 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17138), .ZN(n17133) );
  NOR2_X1 U13167 ( .A1(n18114), .A2(n17153), .ZN(n17150) );
  NOR2_X1 U13168 ( .A1(n17313), .A2(n17177), .ZN(n17172) );
  NAND2_X1 U13169 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17193), .ZN(n17189) );
  NAND3_X1 U13170 ( .A1(n15497), .A2(n15496), .A3(n15495), .ZN(n16292) );
  INV_X1 U13171 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17472) );
  NOR2_X1 U13172 ( .A1(n17858), .A2(n17639), .ZN(n17527) );
  INV_X1 U13173 ( .A(n17576), .ZN(n17597) );
  NOR2_X2 U13174 ( .A1(n17748), .A2(n17231), .ZN(n17636) );
  NOR2_X1 U13175 ( .A1(n18426), .A2(n18324), .ZN(n16235) );
  INV_X1 U13176 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15724) );
  INV_X1 U13177 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20898) );
  NOR2_X1 U13178 ( .A1(n18019), .A2(n18017), .ZN(n18058) );
  INV_X1 U13179 ( .A(n18558), .ZN(n18535) );
  NOR2_X1 U13180 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18679), .ZN(
        n18703) );
  INV_X1 U13181 ( .A(n18508), .ZN(n18159) );
  INV_X1 U13182 ( .A(n18153), .ZN(n18181) );
  INV_X1 U13183 ( .A(n18185), .ZN(n18249) );
  INV_X1 U13184 ( .A(n18229), .ZN(n18255) );
  INV_X1 U13185 ( .A(n18266), .ZN(n18298) );
  INV_X1 U13186 ( .A(n18276), .ZN(n18343) );
  INV_X1 U13187 ( .A(n18335), .ZN(n18365) );
  INV_X1 U13188 ( .A(n18347), .ZN(n18369) );
  INV_X1 U13189 ( .A(n18383), .ZN(n18419) );
  INV_X1 U13190 ( .A(n18412), .ZN(n18446) );
  INV_X1 U13191 ( .A(n18733), .ZN(n18599) );
  NOR2_X1 U13192 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12638), .ZN(n16387)
         );
  NAND2_X1 U13193 ( .A1(n12746), .A2(n13001), .ZN(n14243) );
  INV_X1 U13194 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20759) );
  INV_X1 U13195 ( .A(n19776), .ZN(n19817) );
  OR2_X1 U13196 ( .A1(n14414), .A2(n14343), .ZN(n14603) );
  OR2_X1 U13197 ( .A1(n15863), .A2(n13717), .ZN(n15870) );
  OR2_X1 U13198 ( .A1(n14454), .A2(n14453), .ZN(n15897) );
  INV_X1 U13199 ( .A(n15867), .ZN(n14489) );
  INV_X1 U13200 ( .A(n15867), .ZN(n14507) );
  NAND2_X1 U13201 ( .A1(n19877), .A2(n9956), .ZN(n13139) );
  INV_X1 U13202 ( .A(n19877), .ZN(n19903) );
  INV_X1 U13203 ( .A(n19926), .ZN(n13141) );
  OR2_X1 U13204 ( .A1(n13652), .A2(n13655), .ZN(n15843) );
  OR2_X1 U13205 ( .A1(n19939), .A2(n11868), .ZN(n15914) );
  INV_X1 U13206 ( .A(n19974), .ZN(n19981) );
  OR2_X1 U13207 ( .A1(n14773), .A2(n14791), .ZN(n15937) );
  AND2_X1 U13208 ( .A1(n13672), .A2(n13671), .ZN(n19977) );
  NAND2_X1 U13209 ( .A1(n13033), .A2(n13018), .ZN(n14832) );
  INV_X1 U13210 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12914) );
  OR2_X1 U13211 ( .A1(n20115), .A2(n20294), .ZN(n20068) );
  NAND2_X1 U13212 ( .A1(n20108), .A2(n20461), .ZN(n20107) );
  OR2_X1 U13213 ( .A1(n20115), .A2(n20515), .ZN(n20147) );
  NAND2_X1 U13214 ( .A1(n20108), .A2(n9654), .ZN(n20177) );
  OR2_X1 U13215 ( .A1(n20259), .A2(n20294), .ZN(n20215) );
  NAND2_X1 U13216 ( .A1(n20262), .A2(n20461), .ZN(n20250) );
  OR2_X1 U13217 ( .A1(n20259), .A2(n20515), .ZN(n20291) );
  NAND2_X1 U13218 ( .A1(n20726), .A2(n20429), .ZN(n20349) );
  NAND2_X1 U13219 ( .A1(n20726), .A2(n20328), .ZN(n20387) );
  OR2_X1 U13220 ( .A1(n20396), .A2(n20350), .ZN(n20417) );
  OR2_X1 U13221 ( .A1(n20396), .A2(n9650), .ZN(n20460) );
  INV_X1 U13222 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20301) );
  INV_X1 U13223 ( .A(n20717), .ZN(n20651) );
  AND2_X1 U13224 ( .A1(n20659), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20749) );
  INV_X1 U13225 ( .A(n20706), .ZN(n20704) );
  AND2_X1 U13226 ( .A1(n13252), .A2(n16213), .ZN(n18751) );
  NAND2_X1 U13227 ( .A1(n12226), .A2(n12055), .ZN(n18757) );
  OR2_X1 U13228 ( .A1(n10881), .A2(n10880), .ZN(n18878) );
  INV_X1 U13229 ( .A(n14890), .ZN(n14946) );
  INV_X1 U13230 ( .A(n12964), .ZN(n14890) );
  OR2_X1 U13231 ( .A1(n14946), .A2(n13386), .ZN(n14961) );
  INV_X1 U13232 ( .A(n18983), .ZN(n18966) );
  OR2_X1 U13233 ( .A1(n18983), .A2(n12596), .ZN(n18978) );
  NAND2_X1 U13234 ( .A1(n19030), .A2(n19728), .ZN(n18998) );
  NAND2_X1 U13235 ( .A1(n12794), .A2(n12793), .ZN(n18995) );
  OR2_X1 U13236 ( .A1(n12792), .A2(n19735), .ZN(n19030) );
  OR2_X1 U13237 ( .A1(n12670), .A2(n10635), .ZN(n12869) );
  OR2_X1 U13238 ( .A1(n18757), .A2(n19737), .ZN(n16134) );
  INV_X1 U13239 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20946) );
  INV_X1 U13240 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16140) );
  INV_X1 U13241 ( .A(n16137), .ZN(n19047) );
  INV_X1 U13242 ( .A(n19065), .ZN(n16204) );
  INV_X1 U13243 ( .A(n15468), .ZN(n16209) );
  AOI21_X1 U13244 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13371), .A(n12697), 
        .ZN(n15477) );
  AND2_X1 U13245 ( .A1(n19087), .A2(n19516), .ZN(n19107) );
  NAND2_X1 U13246 ( .A1(n19361), .A2(n19077), .ZN(n19147) );
  AOI21_X1 U13247 ( .B1(n19165), .B2(n19682), .A(n19164), .ZN(n19193) );
  NOR2_X1 U13248 ( .A1(n19200), .A2(n19199), .ZN(n19228) );
  INV_X1 U13249 ( .A(n19259), .ZN(n19254) );
  INV_X1 U13250 ( .A(n19321), .ZN(n19317) );
  NAND2_X1 U13251 ( .A1(n19304), .A2(n19303), .ZN(n19345) );
  INV_X1 U13252 ( .A(n19412), .ZN(n19407) );
  INV_X1 U13253 ( .A(n19429), .ZN(n19424) );
  INV_X1 U13254 ( .A(n19460), .ZN(n19455) );
  INV_X1 U13255 ( .A(n19530), .ZN(n19488) );
  INV_X1 U13256 ( .A(n19545), .ZN(n19506) );
  AOI21_X1 U13257 ( .B1(n19513), .B2(n19517), .A(n19510), .ZN(n19550) );
  INV_X1 U13258 ( .A(n19678), .ZN(n19599) );
  INV_X1 U13259 ( .A(n16760), .ZN(n18747) );
  NAND2_X1 U13260 ( .A1(n18727), .A2(n18570), .ZN(n16406) );
  INV_X1 U13261 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17432) );
  INV_X1 U13262 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17462) );
  INV_X1 U13263 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17056) );
  NAND2_X1 U13264 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18590), .ZN(n16757) );
  INV_X1 U13265 ( .A(n16806), .ZN(n16805) );
  NAND2_X1 U13266 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16864), .ZN(n16858) );
  AND2_X1 U13267 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16902), .ZN(n16916) );
  INV_X1 U13268 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17084) );
  INV_X1 U13269 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17091) );
  INV_X1 U13270 ( .A(n16292), .ZN(n17231) );
  NOR2_X1 U13271 ( .A1(n15519), .A2(n15518), .ZN(n17248) );
  AOI21_X1 U13272 ( .B1(n15741), .B2(n15740), .A(n18581), .ZN(n17110) );
  NAND2_X1 U13273 ( .A1(n17284), .A2(n18082), .ZN(n17283) );
  INV_X1 U13274 ( .A(n17284), .ZN(n17301) );
  INV_X1 U13275 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17845) );
  INV_X1 U13276 ( .A(n17636), .ZN(n17650) );
  INV_X1 U13277 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17962) );
  INV_X1 U13278 ( .A(n17738), .ZN(n17750) );
  INV_X1 U13279 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17820) );
  INV_X1 U13280 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17933) );
  INV_X1 U13281 ( .A(n18058), .ZN(n18035) );
  NAND2_X1 U13282 ( .A1(n18019), .A2(n18509), .ZN(n18068) );
  INV_X1 U13283 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18562) );
  INV_X1 U13284 ( .A(n18319), .ZN(n18291) );
  INV_X1 U13285 ( .A(n18453), .ZN(n18400) );
  INV_X1 U13286 ( .A(n18430), .ZN(n18450) );
  INV_X1 U13287 ( .A(n18727), .ZN(n18581) );
  INV_X1 U13288 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18679) );
  INV_X1 U13289 ( .A(n18676), .ZN(n18591) );
  INV_X1 U13290 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18607) );
  NAND2_X1 U13291 ( .A1(n18607), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18740) );
  INV_X1 U13292 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n18999) );
  INV_X1 U13293 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19624) );
  CLKBUF_X1 U13294 ( .A(n16398), .Z(n20962) );
  OR4_X1 U13295 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        P2_U2840) );
  INV_X1 U13296 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10248) );
  NAND2_X1 U13297 ( .A1(n10274), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10271) );
  INV_X1 U13298 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16117) );
  AND2_X1 U13299 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U13300 ( .A1(n10257), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10255) );
  INV_X1 U13301 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15060) );
  INV_X1 U13302 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15050) );
  INV_X1 U13303 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10281) );
  OAI21_X1 U13304 ( .B1(n10251), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n10249), .ZN(n15031) );
  INV_X1 U13305 ( .A(n15031), .ZN(n14844) );
  INV_X1 U13306 ( .A(n10250), .ZN(n10252) );
  AOI21_X1 U13307 ( .B1(n15050), .B2(n10252), .A(n10251), .ZN(n15053) );
  AOI21_X1 U13308 ( .B1(n15060), .B2(n9679), .A(n10250), .ZN(n16022) );
  OR2_X1 U13309 ( .A1(n10254), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10253) );
  NAND2_X1 U13310 ( .A1(n9679), .A2(n10253), .ZN(n15069) );
  INV_X1 U13311 ( .A(n15069), .ZN(n16033) );
  AOI21_X1 U13312 ( .B1(n15081), .B2(n9739), .A(n10254), .ZN(n15079) );
  OAI21_X1 U13313 ( .B1(n10256), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n9739), .ZN(n15091) );
  INV_X1 U13314 ( .A(n15091), .ZN(n16041) );
  AOI21_X1 U13315 ( .B1(n10246), .B2(n10255), .A(n10256), .ZN(n15100) );
  OAI21_X1 U13316 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10257), .A(
        n10255), .ZN(n16078) );
  INV_X1 U13317 ( .A(n16078), .ZN(n15680) );
  AOI21_X1 U13318 ( .B1(n15115), .B2(n10258), .A(n10257), .ZN(n18784) );
  AND2_X1 U13319 ( .A1(n10264), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10262) );
  AND2_X1 U13320 ( .A1(n10262), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10260) );
  OAI21_X1 U13321 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10260), .A(
        n10258), .ZN(n15129) );
  INV_X1 U13322 ( .A(n15129), .ZN(n18796) );
  NOR2_X1 U13323 ( .A1(n10262), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10259) );
  NOR2_X1 U13324 ( .A1(n10260), .A2(n10259), .ZN(n18808) );
  NOR2_X1 U13325 ( .A1(n10264), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10261) );
  NOR2_X1 U13326 ( .A1(n10262), .A2(n10261), .ZN(n15149) );
  AND2_X1 U13327 ( .A1(n9730), .A2(n10263), .ZN(n10265) );
  OR2_X1 U13328 ( .A1(n10265), .A2(n10264), .ZN(n18826) );
  INV_X1 U13329 ( .A(n18826), .ZN(n18817) );
  AOI21_X1 U13330 ( .B1(n15180), .B2(n10266), .A(n10267), .ZN(n12645) );
  AOI21_X1 U13331 ( .B1(n15193), .B2(n10268), .A(n10269), .ZN(n12657) );
  AOI21_X1 U13332 ( .B1(n20946), .B2(n10279), .A(n10270), .ZN(n18840) );
  AOI21_X1 U13333 ( .B1(n16117), .B2(n10271), .A(n10272), .ZN(n18862) );
  AOI21_X1 U13334 ( .B1(n13825), .B2(n10273), .A(n10274), .ZN(n18873) );
  NAND2_X1 U13335 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10275), .ZN(
        n10277) );
  NOR2_X1 U13336 ( .A1(n16140), .A2(n10277), .ZN(n10278) );
  AOI21_X1 U13337 ( .B1(n16140), .B2(n10277), .A(n10278), .ZN(n18910) );
  AOI21_X1 U13338 ( .B1(n16152), .B2(n10276), .A(n10275), .ZN(n16141) );
  OAI22_X1 U13339 ( .A1(n13371), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n18937) );
  INV_X1 U13340 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13422) );
  OAI22_X1 U13341 ( .A1(n13371), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13422), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13429) );
  AND2_X1 U13342 ( .A1(n18937), .A2(n13429), .ZN(n13428) );
  OAI21_X1 U13343 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n10276), .ZN(n13434) );
  NAND2_X1 U13344 ( .A1(n13428), .A2(n13434), .ZN(n13193) );
  NOR2_X1 U13345 ( .A1(n16141), .A2(n13193), .ZN(n13319) );
  OAI21_X1 U13346 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10275), .A(
        n10277), .ZN(n19051) );
  NAND2_X1 U13347 ( .A1(n13319), .A2(n19051), .ZN(n18907) );
  NOR2_X1 U13348 ( .A1(n18910), .A2(n18907), .ZN(n18890) );
  OAI21_X1 U13349 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10278), .A(
        n10273), .ZN(n18892) );
  NAND2_X1 U13350 ( .A1(n18890), .A2(n18892), .ZN(n18872) );
  NOR2_X1 U13351 ( .A1(n18873), .A2(n18872), .ZN(n13108) );
  OAI21_X1 U13352 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10274), .A(
        n10271), .ZN(n16131) );
  NAND2_X1 U13353 ( .A1(n13108), .A2(n16131), .ZN(n18861) );
  NOR2_X1 U13354 ( .A1(n18862), .A2(n18861), .ZN(n18854) );
  OAI21_X1 U13355 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10272), .A(
        n10279), .ZN(n18855) );
  NAND2_X1 U13356 ( .A1(n18854), .A2(n18855), .ZN(n18839) );
  NOR2_X1 U13357 ( .A1(n18840), .A2(n18839), .ZN(n13462) );
  OAI21_X1 U13358 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10270), .A(
        n10268), .ZN(n16093) );
  NAND2_X1 U13359 ( .A1(n13462), .A2(n16093), .ZN(n12655) );
  NOR2_X1 U13360 ( .A1(n12657), .A2(n12655), .ZN(n13612) );
  OAI21_X1 U13361 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10269), .A(
        n10266), .ZN(n16087) );
  NAND2_X1 U13362 ( .A1(n13612), .A2(n16087), .ZN(n12639) );
  NOR2_X1 U13363 ( .A1(n12645), .A2(n12639), .ZN(n18830) );
  OAI21_X1 U13364 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10267), .A(
        n9730), .ZN(n18832) );
  NAND2_X1 U13365 ( .A1(n18830), .A2(n18832), .ZN(n18816) );
  NOR2_X1 U13366 ( .A1(n18817), .A2(n18816), .ZN(n18815) );
  NOR2_X1 U13367 ( .A1(n12060), .A2(n18815), .ZN(n13850) );
  NOR2_X1 U13368 ( .A1(n15149), .A2(n13850), .ZN(n13849) );
  NOR2_X1 U13369 ( .A1(n18891), .A2(n18794), .ZN(n18783) );
  NOR2_X1 U13370 ( .A1(n18784), .A2(n18783), .ZN(n18782) );
  NOR2_X1 U13371 ( .A1(n18891), .A2(n14875), .ZN(n16040) );
  NOR2_X1 U13372 ( .A1(n16041), .A2(n16040), .ZN(n16039) );
  NOR2_X1 U13373 ( .A1(n18891), .A2(n16039), .ZN(n14870) );
  NOR2_X2 U13374 ( .A1(n15079), .A2(n14870), .ZN(n14869) );
  NOR2_X1 U13375 ( .A1(n12060), .A2(n14869), .ZN(n16032) );
  NOR2_X1 U13376 ( .A1(n16033), .A2(n16032), .ZN(n16031) );
  NOR2_X1 U13377 ( .A1(n18891), .A2(n14848), .ZN(n14843) );
  NOR2_X1 U13378 ( .A1(n14844), .A2(n14843), .ZN(n14842) );
  NOR3_X1 U13379 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15736) );
  NAND2_X1 U13380 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15736), .ZN(n18883) );
  NAND2_X1 U13381 ( .A1(n18912), .A2(n9642), .ZN(n18936) );
  INV_X1 U13382 ( .A(n18936), .ZN(n10282) );
  XNOR2_X1 U13383 ( .A(n10249), .B(n10281), .ZN(n16000) );
  NAND3_X1 U13384 ( .A1(n16001), .A2(n10282), .A3(n16000), .ZN(n10586) );
  AND2_X4 U13385 ( .A1(n12050), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10384) );
  AND2_X4 U13386 ( .A1(n12050), .A2(n10283), .ZN(n10361) );
  AND2_X2 U13387 ( .A1(n10283), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13220) );
  INV_X2 U13388 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10568) );
  AND2_X4 U13389 ( .A1(n13220), .A2(n10568), .ZN(n12443) );
  AND2_X2 U13390 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13069) );
  AND2_X4 U13391 ( .A1(n13069), .A2(n10568), .ZN(n12554) );
  AOI22_X1 U13392 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10290) );
  NOR2_X4 U13393 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10286) );
  AND2_X4 U13394 ( .A1(n10286), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10354) );
  AND2_X4 U13395 ( .A1(n10286), .A2(n10568), .ZN(n12575) );
  AOI22_X1 U13396 ( .A1(n12577), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13397 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10288) );
  NAND4_X1 U13398 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10299) );
  AOI22_X1 U13399 ( .A1(n12577), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U13400 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13401 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10295) );
  NAND2_X1 U13402 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10292) );
  NAND4_X1 U13403 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  AOI22_X1 U13404 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13405 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13406 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U13407 ( .A1(n10361), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10301) );
  NAND2_X1 U13408 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10300) );
  NAND4_X1 U13409 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10313) );
  AOI22_X1 U13410 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13411 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13412 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10309) );
  NAND2_X1 U13413 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10306) );
  NAND4_X1 U13414 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10312) );
  MUX2_X2 U13415 ( .A(n10313), .B(n10312), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10416) );
  AOI22_X1 U13416 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13417 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13418 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13419 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10315) );
  NAND4_X1 U13420 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10325) );
  AOI22_X1 U13421 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13422 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10321) );
  NAND3_X1 U13423 ( .A1(n10323), .A2(n10322), .A3(n10321), .ZN(n10324) );
  MUX2_X1 U13424 ( .A(n10613), .B(n10416), .S(n12318), .Z(n10338) );
  AOI22_X1 U13425 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13426 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13427 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13428 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13429 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10384), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13430 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13431 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13432 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10331) );
  NAND3_X1 U13433 ( .A1(n10334), .A2(n10333), .A3(n10236), .ZN(n10335) );
  NAND2_X1 U13434 ( .A1(n10399), .A2(n10416), .ZN(n10337) );
  NOR2_X2 U13435 ( .A1(n10394), .A2(n12617), .ZN(n10420) );
  AOI22_X1 U13436 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13437 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13438 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13439 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10340) );
  NAND4_X1 U13440 ( .A1(n10343), .A2(n10342), .A3(n10341), .A4(n10340), .ZN(
        n10349) );
  AOI22_X1 U13441 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13442 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13443 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13444 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U13445 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10348) );
  MUX2_X2 U13446 ( .A(n10349), .B(n10348), .S(n13075), .Z(n10615) );
  NAND2_X1 U13448 ( .A1(n12596), .A2(n19737), .ZN(n12273) );
  AOI22_X1 U13449 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10354), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13450 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13451 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13452 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10350) );
  NAND4_X1 U13453 ( .A1(n10353), .A2(n10352), .A3(n10351), .A4(n10350), .ZN(
        n10360) );
  AOI22_X1 U13454 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9644), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13455 ( .A1(n10354), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13456 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13457 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10361), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10355) );
  NAND4_X1 U13458 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10359) );
  MUX2_X2 U13459 ( .A(n10360), .B(n10359), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13399) );
  INV_X1 U13460 ( .A(n10420), .ZN(n10372) );
  AOI22_X1 U13461 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13462 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12577), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13463 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10363) );
  BUF_X2 U13464 ( .A(n10361), .Z(n10383) );
  AOI22_X1 U13465 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10362) );
  NAND4_X1 U13466 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10371) );
  AOI22_X1 U13467 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13468 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13469 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10367) );
  INV_X1 U13470 ( .A(n10384), .ZN(n12444) );
  AOI22_X1 U13471 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10366) );
  NAND4_X1 U13472 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10370) );
  MUX2_X2 U13473 ( .A(n10371), .B(n10370), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10414) );
  NAND2_X1 U13474 ( .A1(n10372), .A2(n10404), .ZN(n10378) );
  NAND2_X1 U13475 ( .A1(n12318), .A2(n10613), .ZN(n10413) );
  NAND2_X1 U13476 ( .A1(n10373), .A2(n10043), .ZN(n10374) );
  INV_X2 U13477 ( .A(n10416), .ZN(n10375) );
  NAND2_X1 U13478 ( .A1(n10376), .A2(n10375), .ZN(n12212) );
  NAND2_X1 U13479 ( .A1(n12596), .A2(n10416), .ZN(n12210) );
  NAND3_X1 U13480 ( .A1(n12212), .A2(n12210), .A3(n12617), .ZN(n12278) );
  NAND2_X1 U13481 ( .A1(n12278), .A2(n10414), .ZN(n10377) );
  NAND2_X1 U13482 ( .A1(n10378), .A2(n10377), .ZN(n10449) );
  NAND2_X1 U13483 ( .A1(n10615), .A2(n13399), .ZN(n10412) );
  NAND2_X1 U13484 ( .A1(n10449), .A2(n12229), .ZN(n10397) );
  AOI22_X1 U13485 ( .A1(n9639), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9644), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13486 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13487 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13488 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10379) );
  NAND2_X1 U13489 ( .A1(n10382), .A2(n9692), .ZN(n10391) );
  AOI22_X1 U13490 ( .A1(n12576), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13491 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13492 ( .A1(n12443), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13493 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10385) );
  NAND2_X1 U13494 ( .A1(n10389), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10390) );
  NOR2_X1 U13495 ( .A1(n13383), .A2(n10613), .ZN(n10393) );
  NOR2_X1 U13496 ( .A1(n10416), .A2(n10414), .ZN(n10392) );
  OAI21_X1 U13497 ( .B1(n10634), .B2(n10404), .A(n13383), .ZN(n10395) );
  INV_X4 U13498 ( .A(n13399), .ZN(n12280) );
  OAI211_X1 U13499 ( .C1(n10447), .C2(n13399), .A(n10397), .B(n12283), .ZN(
        n10398) );
  NAND2_X1 U13500 ( .A1(n10398), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10403) );
  NOR2_X1 U13501 ( .A1(n10413), .A2(n13386), .ZN(n10400) );
  AND2_X2 U13502 ( .A1(n10401), .A2(n10400), .ZN(n12222) );
  NAND3_X1 U13503 ( .A1(n12313), .A2(n13383), .A3(n10615), .ZN(n10402) );
  NAND2_X1 U13504 ( .A1(n10410), .A2(n10402), .ZN(n12266) );
  NAND2_X1 U13505 ( .A1(n13399), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12249) );
  NAND2_X2 U13506 ( .A1(n12280), .A2(n10587), .ZN(n12700) );
  INV_X1 U13507 ( .A(n12700), .ZN(n12592) );
  NAND2_X1 U13508 ( .A1(n9647), .A2(n10406), .ZN(n10411) );
  INV_X1 U13509 ( .A(n10411), .ZN(n10407) );
  NAND2_X1 U13510 ( .A1(n12222), .A2(n13399), .ZN(n10882) );
  NAND2_X1 U13511 ( .A1(n10407), .A2(n10882), .ZN(n12261) );
  INV_X1 U13512 ( .A(n13266), .ZN(n10440) );
  NAND2_X1 U13513 ( .A1(n10408), .A2(n10234), .ZN(n10409) );
  INV_X1 U13514 ( .A(n10428), .ZN(n10426) );
  NAND2_X1 U13515 ( .A1(n19737), .A2(n13399), .ZN(n12047) );
  OAI21_X1 U13516 ( .B1(n13268), .B2(n10411), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10419) );
  NAND2_X2 U13517 ( .A1(n12700), .A2(n10412), .ZN(n12275) );
  NOR2_X1 U13518 ( .A1(n10413), .A2(n10615), .ZN(n10415) );
  NAND3_X2 U13519 ( .A1(n12275), .A2(n10417), .A3(n10235), .ZN(n12265) );
  NOR2_X2 U13520 ( .A1(n12265), .A2(n10418), .ZN(n13066) );
  NAND2_X1 U13521 ( .A1(n13066), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10436) );
  NAND2_X1 U13522 ( .A1(n10419), .A2(n10436), .ZN(n10455) );
  NAND2_X1 U13523 ( .A1(n10455), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10424) );
  INV_X1 U13524 ( .A(n10464), .ZN(n10421) );
  NAND2_X1 U13525 ( .A1(n10421), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10423) );
  NOR2_X2 U13526 ( .A1(n10430), .A2(n10410), .ZN(n10466) );
  AOI22_X1 U13527 ( .A1(n10466), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10422) );
  AND3_X2 U13528 ( .A1(n10424), .A2(n10423), .A3(n10422), .ZN(n10427) );
  INV_X1 U13529 ( .A(n10427), .ZN(n10425) );
  NAND2_X1 U13530 ( .A1(n10426), .A2(n10425), .ZN(n10429) );
  NAND2_X1 U13531 ( .A1(n10429), .A2(n11879), .ZN(n11884) );
  AND2_X1 U13532 ( .A1(n10432), .A2(n10431), .ZN(n10434) );
  INV_X2 U13533 ( .A(n10464), .ZN(n10433) );
  OAI22_X1 U13534 ( .A1(n10470), .A2(n10434), .B1(n10433), .B2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U13535 ( .A1(n13266), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10435) );
  AND2_X1 U13536 ( .A1(n10436), .A2(n10435), .ZN(n10437) );
  NAND2_X1 U13537 ( .A1(n10438), .A2(n10437), .ZN(n11887) );
  NAND2_X1 U13538 ( .A1(n10455), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10446) );
  NAND2_X1 U13539 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10439) );
  NAND2_X1 U13540 ( .A1(n10440), .A2(n10439), .ZN(n10441) );
  AOI21_X1 U13541 ( .B1(n10466), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10441), .ZN(
        n10442) );
  AND2_X1 U13542 ( .A1(n10443), .A2(n10442), .ZN(n10445) );
  INV_X1 U13543 ( .A(n10447), .ZN(n10448) );
  OAI21_X1 U13544 ( .B1(n10449), .B2(n12280), .A(n10448), .ZN(n10450) );
  AOI21_X1 U13545 ( .B1(n10450), .B2(n12283), .A(n13371), .ZN(n10451) );
  NAND2_X1 U13546 ( .A1(n10453), .A2(n10452), .ZN(n11886) );
  OAI21_X1 U13547 ( .B1(n12319), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13528), 
        .ZN(n10454) );
  INV_X1 U13548 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13549 ( .A1(n10466), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10457) );
  NAND2_X1 U13550 ( .A1(n10458), .A2(n10457), .ZN(n10459) );
  INV_X1 U13551 ( .A(n10460), .ZN(n10463) );
  INV_X1 U13552 ( .A(n10461), .ZN(n10462) );
  NAND2_X1 U13553 ( .A1(n10455), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10469) );
  INV_X1 U13554 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10465) );
  OR2_X1 U13555 ( .A1(n10561), .A2(n10465), .ZN(n10468) );
  AOI22_X1 U13556 ( .A1(n10466), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10467) );
  NAND2_X1 U13557 ( .A1(n10470), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10472) );
  NAND2_X1 U13558 ( .A1(n13266), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10471) );
  INV_X1 U13559 ( .A(n10473), .ZN(n10474) );
  INV_X1 U13560 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13561 ( .A1(n10557), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10478) );
  NAND2_X1 U13562 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10477) );
  OAI211_X1 U13563 ( .C1(n10561), .C2(n10479), .A(n10478), .B(n10477), .ZN(
        n13054) );
  INV_X1 U13564 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U13565 ( .A1(n10557), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10481) );
  NAND2_X1 U13566 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10480) );
  OAI211_X1 U13567 ( .C1(n10561), .C2(n12967), .A(n10481), .B(n10480), .ZN(
        n12962) );
  NAND2_X1 U13568 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10485) );
  INV_X1 U13569 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10482) );
  OR2_X1 U13570 ( .A1(n10561), .A2(n10482), .ZN(n10484) );
  INV_X2 U13571 ( .A(n10506), .ZN(n10557) );
  AOI22_X1 U13572 ( .A1(n10557), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10483) );
  NAND2_X1 U13573 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10489) );
  INV_X1 U13574 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10869) );
  OR2_X1 U13575 ( .A1(n10561), .A2(n10869), .ZN(n10488) );
  AOI22_X1 U13576 ( .A1(n10557), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10487) );
  NAND2_X1 U13577 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10493) );
  INV_X1 U13578 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10490) );
  OR2_X1 U13579 ( .A1(n10561), .A2(n10490), .ZN(n10492) );
  AOI22_X1 U13580 ( .A1(n10557), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10491) );
  INV_X1 U13581 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13582 ( .A1(n10557), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10495) );
  NAND2_X1 U13583 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10494) );
  OAI211_X1 U13584 ( .C1(n10561), .C2(n10496), .A(n10495), .B(n10494), .ZN(
        n13364) );
  INV_X1 U13585 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13586 ( .A1(n10557), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10498) );
  NAND2_X1 U13587 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10497) );
  OAI211_X1 U13588 ( .C1(n10561), .C2(n10499), .A(n10498), .B(n10497), .ZN(
        n13501) );
  NAND2_X1 U13589 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10503) );
  INV_X1 U13590 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10500) );
  OR2_X1 U13591 ( .A1(n10561), .A2(n10500), .ZN(n10502) );
  AOI22_X1 U13592 ( .A1(n10557), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10501) );
  INV_X1 U13593 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15418) );
  AOI22_X1 U13594 ( .A1(n10557), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10505) );
  NAND2_X1 U13595 ( .A1(n10433), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10504) );
  OAI211_X1 U13596 ( .C1(n10476), .C2(n15418), .A(n10505), .B(n10504), .ZN(
        n13345) );
  INV_X1 U13597 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20932) );
  OAI22_X1 U13598 ( .A1(n10506), .A2(n20932), .B1(n13528), .B2(n15193), .ZN(
        n10508) );
  INV_X1 U13599 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15395) );
  NOR2_X1 U13600 ( .A1(n10476), .A2(n15395), .ZN(n10507) );
  AOI211_X1 U13601 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n10433), .A(n10508), .B(
        n10507), .ZN(n12659) );
  INV_X1 U13602 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13571) );
  AOI22_X1 U13603 ( .A1(n10557), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10510) );
  NAND2_X1 U13604 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10509) );
  OAI211_X1 U13605 ( .C1(n10561), .C2(n13571), .A(n10510), .B(n10509), .ZN(
        n13564) );
  INV_X1 U13606 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13607 ( .A1(n10557), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10512) );
  NAND2_X1 U13608 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10511) );
  OAI211_X1 U13609 ( .C1(n10561), .C2(n10871), .A(n10512), .B(n10511), .ZN(
        n12647) );
  INV_X1 U13610 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U13611 ( .A1(n10557), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10514) );
  NAND2_X1 U13612 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10513) );
  OAI211_X1 U13613 ( .C1(n10561), .C2(n13663), .A(n10514), .B(n10513), .ZN(
        n13661) );
  NAND2_X1 U13614 ( .A1(n10433), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10517) );
  NAND2_X1 U13615 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10516) );
  AOI22_X1 U13616 ( .A1(n10557), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10515) );
  NAND2_X1 U13617 ( .A1(n10433), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U13618 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10519) );
  AOI22_X1 U13619 ( .A1(n10557), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10518) );
  NAND2_X1 U13620 ( .A1(n10433), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10523) );
  NAND2_X1 U13621 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10522) );
  AOI22_X1 U13622 ( .A1(n10557), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10521) );
  INV_X1 U13623 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13624 ( .A1(n10557), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10525) );
  NAND2_X1 U13625 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10524) );
  OAI211_X1 U13626 ( .C1(n10561), .C2(n10526), .A(n10525), .B(n10524), .ZN(
        n14957) );
  NAND2_X1 U13627 ( .A1(n14958), .A2(n14957), .ZN(n14956) );
  NAND2_X1 U13628 ( .A1(n10433), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10529) );
  NAND2_X1 U13629 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10528) );
  AOI22_X1 U13630 ( .A1(n10557), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10527) );
  NAND2_X1 U13631 ( .A1(n10433), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10532) );
  NAND2_X1 U13632 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10531) );
  AOI22_X1 U13633 ( .A1(n10557), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10530) );
  INV_X1 U13634 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13635 ( .A1(n10557), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10534) );
  NAND2_X1 U13636 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10533) );
  OAI211_X1 U13637 ( .C1(n10561), .C2(n10535), .A(n10534), .B(n10533), .ZN(
        n14879) );
  INV_X1 U13638 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14932) );
  AOI22_X1 U13639 ( .A1(n10557), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10537) );
  NAND2_X1 U13640 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10536) );
  OAI211_X1 U13641 ( .C1(n10561), .C2(n14932), .A(n10537), .B(n10536), .ZN(
        n14930) );
  NAND2_X1 U13642 ( .A1(n10433), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U13643 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10539) );
  AOI22_X1 U13644 ( .A1(n10557), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10538) );
  AND3_X1 U13645 ( .A1(n10540), .A2(n10539), .A3(n10538), .ZN(n14862) );
  NAND2_X1 U13646 ( .A1(n10433), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10543) );
  NAND2_X1 U13647 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10542) );
  AOI22_X1 U13648 ( .A1(n10557), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10541) );
  AND3_X1 U13649 ( .A1(n10543), .A2(n10542), .A3(n10541), .ZN(n14914) );
  NAND2_X1 U13650 ( .A1(n10433), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10546) );
  NAND2_X1 U13651 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10545) );
  AOI22_X1 U13652 ( .A1(n10557), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10544) );
  INV_X1 U13653 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13654 ( .A1(n10557), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10548) );
  NAND2_X1 U13655 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10547) );
  OAI211_X1 U13656 ( .C1(n10561), .C2(n10549), .A(n10548), .B(n10547), .ZN(
        n14853) );
  NAND2_X1 U13657 ( .A1(n10433), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10552) );
  NAND2_X1 U13658 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10551) );
  AOI22_X1 U13659 ( .A1(n10557), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10550) );
  INV_X1 U13660 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10555) );
  AOI22_X1 U13661 ( .A1(n10557), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10554) );
  NAND2_X1 U13662 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10553) );
  OAI211_X1 U13663 ( .C1(n10561), .C2(n10555), .A(n10554), .B(n10553), .ZN(
        n14236) );
  INV_X1 U13664 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13665 ( .A1(n10556), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10559) );
  AOI22_X1 U13666 ( .A1(n10557), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10558) );
  OAI211_X1 U13667 ( .C1(n10561), .C2(n10560), .A(n10559), .B(n10558), .ZN(
        n10562) );
  INV_X1 U13668 ( .A(n10562), .ZN(n10563) );
  NAND2_X1 U13669 ( .A1(n10882), .A2(n9647), .ZN(n13243) );
  NAND2_X1 U13670 ( .A1(n19705), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10566) );
  NAND2_X1 U13671 ( .A1(n13221), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10565) );
  NAND2_X1 U13672 ( .A1(n10566), .A2(n10565), .ZN(n12230) );
  NAND2_X1 U13673 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19714), .ZN(
        n12038) );
  NAND2_X1 U13674 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12319), .ZN(
        n10567) );
  NAND2_X1 U13675 ( .A1(n10576), .A2(n10567), .ZN(n10570) );
  NAND2_X1 U13676 ( .A1(n13070), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10569) );
  NAND2_X1 U13677 ( .A1(n10570), .A2(n10569), .ZN(n10581) );
  XNOR2_X1 U13678 ( .A(n13075), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10579) );
  OAI22_X1 U13679 ( .A1(n10581), .A2(n10579), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13075), .ZN(n10575) );
  INV_X1 U13680 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15738) );
  NAND2_X1 U13681 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12703), .ZN(
        n10574) );
  NAND2_X1 U13682 ( .A1(n12230), .A2(n12038), .ZN(n12039) );
  AND2_X1 U13683 ( .A1(n10573), .A2(n12039), .ZN(n12232) );
  OR2_X1 U13684 ( .A1(n10575), .A2(n10574), .ZN(n12242) );
  MUX2_X1 U13685 ( .A(n12319), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10577) );
  INV_X1 U13686 ( .A(n10577), .ZN(n10578) );
  MUX2_X1 U13687 ( .A(n10578), .B(n10577), .S(n10576), .Z(n12228) );
  INV_X1 U13688 ( .A(n10579), .ZN(n10580) );
  XNOR2_X1 U13689 ( .A(n10581), .B(n10580), .ZN(n12240) );
  NAND3_X1 U13690 ( .A1(n12242), .A2(n12228), .A3(n12240), .ZN(n12048) );
  INV_X1 U13691 ( .A(n12048), .ZN(n10582) );
  NAND2_X1 U13692 ( .A1(n12232), .A2(n10582), .ZN(n10583) );
  NAND2_X1 U13693 ( .A1(n13528), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10859) );
  INV_X1 U13694 ( .A(n10859), .ZN(n10584) );
  NAND2_X1 U13695 ( .A1(n18751), .A2(n12229), .ZN(n10881) );
  NAND2_X1 U13696 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19600) );
  INV_X1 U13697 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19736) );
  NAND2_X1 U13698 ( .A1(n19600), .A2(n19736), .ZN(n10880) );
  NAND2_X1 U13699 ( .A1(n10587), .A2(n19731), .ZN(n10614) );
  AND2_X2 U13700 ( .A1(n9646), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10692) );
  AOI22_X1 U13701 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13702 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10591) );
  AND2_X2 U13703 ( .A1(n12577), .A2(n13075), .ZN(n10681) );
  AOI22_X1 U13704 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10681), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10590) );
  AND2_X2 U13705 ( .A1(n12577), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10599) );
  AND2_X1 U13706 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13707 ( .A1(n10599), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10589) );
  NAND4_X1 U13708 ( .A1(n10592), .A2(n10591), .A3(n10590), .A4(n10589), .ZN(
        n10598) );
  AND2_X2 U13709 ( .A1(n12548), .A2(n13075), .ZN(n10668) );
  AOI22_X1 U13710 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n10668), .ZN(n10596) );
  AOI22_X1 U13711 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10595) );
  AND2_X2 U13712 ( .A1(n13067), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10626) );
  AOI22_X1 U13713 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10594) );
  AND2_X2 U13714 ( .A1(n12581), .A2(n13075), .ZN(n10621) );
  AND2_X2 U13715 ( .A1(n10384), .A2(n13075), .ZN(n13078) );
  AOI22_X1 U13716 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10621), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10593) );
  NAND4_X1 U13717 ( .A1(n10596), .A2(n10595), .A3(n10594), .A4(n10593), .ZN(
        n10597) );
  AOI22_X1 U13718 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13719 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13720 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13721 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10600) );
  NAND4_X1 U13722 ( .A1(n10603), .A2(n10602), .A3(n10601), .A4(n10600), .ZN(
        n10609) );
  AOI22_X1 U13723 ( .A1(n10641), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13724 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13725 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10681), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13726 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10604) );
  NAND4_X1 U13727 ( .A1(n10607), .A2(n10606), .A3(n10605), .A4(n10604), .ZN(
        n10608) );
  NOR2_X1 U13728 ( .A1(n10609), .A2(n10608), .ZN(n12676) );
  OR2_X1 U13729 ( .A1(n12676), .A2(n10831), .ZN(n10612) );
  MUX2_X1 U13730 ( .A(n12617), .B(n19714), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10610) );
  AND2_X1 U13731 ( .A1(n10615), .A2(n19731), .ZN(n10729) );
  NAND2_X1 U13732 ( .A1(n10634), .A2(n10729), .ZN(n10654) );
  AND2_X1 U13733 ( .A1(n10610), .A2(n10654), .ZN(n10611) );
  NAND2_X1 U13734 ( .A1(n10612), .A2(n10611), .ZN(n13184) );
  NAND2_X1 U13735 ( .A1(n12617), .A2(n10613), .ZN(n12597) );
  INV_X1 U13736 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18919) );
  AOI21_X1 U13737 ( .B1(n10615), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13738 ( .A1(n13386), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10616) );
  INV_X1 U13739 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19620) );
  AND2_X2 U13740 ( .A1(n13386), .A2(n19731), .ZN(n10728) );
  INV_X1 U13741 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U13742 ( .A1(n10728), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10729), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10618) );
  OAI21_X1 U13743 ( .B1(n10853), .B2(n19620), .A(n10618), .ZN(n10637) );
  INV_X1 U13744 ( .A(n10637), .ZN(n10619) );
  AOI22_X1 U13745 ( .A1(n10599), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13746 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13747 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13748 ( .A1(n9641), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10681), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10622) );
  NAND4_X1 U13749 ( .A1(n10625), .A2(n10624), .A3(n10623), .A4(n10622), .ZN(
        n10633) );
  AOI22_X1 U13750 ( .A1(n10641), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12432), .ZN(n10631) );
  AOI22_X1 U13751 ( .A1(n10646), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10630) );
  AOI22_X1 U13752 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13753 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10692), .B1(
        n10627), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10628) );
  NAND4_X1 U13754 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .ZN(
        n10632) );
  NOR2_X1 U13755 ( .A1(n10633), .A2(n10632), .ZN(n11983) );
  OR2_X1 U13756 ( .A1(n11983), .A2(n12170), .ZN(n10864) );
  OAI22_X1 U13757 ( .A1(n10864), .A2(n10635), .B1(n13386), .B2(n10634), .ZN(
        n10636) );
  MUX2_X1 U13758 ( .A(n10636), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_3__SCAN_IN), .Z(n13181) );
  INV_X1 U13759 ( .A(n13181), .ZN(n10640) );
  NOR2_X1 U13760 ( .A1(n10638), .A2(n10637), .ZN(n10639) );
  AOI21_X2 U13761 ( .B1(n13182), .B2(n10640), .A(n10639), .ZN(n10658) );
  AOI22_X1 U13762 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10663), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13763 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n12432), .ZN(n10644) );
  AOI22_X1 U13764 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U13765 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10642) );
  NAND4_X1 U13766 ( .A1(n10645), .A2(n10644), .A3(n10643), .A4(n10642), .ZN(
        n10653) );
  AOI22_X1 U13767 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n10680), .ZN(n10651) );
  AOI22_X1 U13768 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13769 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13770 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10621), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10648) );
  NAND4_X1 U13771 ( .A1(n10651), .A2(n10650), .A3(n10649), .A4(n10648), .ZN(
        n10652) );
  NOR2_X1 U13772 ( .A1(n10653), .A2(n10652), .ZN(n11986) );
  NAND2_X1 U13773 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10655) );
  OAI211_X1 U13774 ( .C1(n10831), .C2(n11986), .A(n10655), .B(n10654), .ZN(
        n10657) );
  INV_X1 U13775 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19622) );
  AOI22_X1 U13776 ( .A1(n10728), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10854), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10656) );
  OAI21_X1 U13777 ( .B1(n10853), .B2(n19622), .A(n10656), .ZN(n13176) );
  NOR2_X1 U13778 ( .A1(n10658), .A2(n10657), .ZN(n10659) );
  INV_X1 U13779 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13780 ( .A1(n10854), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10661) );
  NAND2_X1 U13781 ( .A1(n10728), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10660) );
  AND2_X1 U13782 ( .A1(n10661), .A2(n10660), .ZN(n10674) );
  AOI22_X1 U13783 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10662), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13784 ( .A1(n10641), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n12432), .ZN(n10666) );
  AOI22_X1 U13785 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13786 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13787 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n10680), .ZN(n10672) );
  AOI22_X1 U13788 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13789 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10670) );
  AOI22_X1 U13790 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10621), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10669) );
  NAND2_X1 U13791 ( .A1(n10818), .A2(n11929), .ZN(n10673) );
  OAI211_X1 U13792 ( .C1(n10853), .C2(n10675), .A(n10674), .B(n10673), .ZN(
        n13195) );
  AOI22_X1 U13793 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10662), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13794 ( .A1(n10641), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n12432), .ZN(n10678) );
  AOI22_X1 U13795 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13796 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10676) );
  NAND4_X1 U13797 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(
        n10687) );
  AOI22_X1 U13798 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n10680), .ZN(n10685) );
  AOI22_X1 U13799 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13800 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13801 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10626), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10682) );
  NAND4_X1 U13802 ( .A1(n10685), .A2(n10684), .A3(n10683), .A4(n10682), .ZN(
        n10686) );
  AOI22_X1 U13803 ( .A1(n10728), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10854), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10688) );
  OAI21_X1 U13804 ( .B1(n11995), .B2(n10831), .A(n10688), .ZN(n10689) );
  INV_X1 U13805 ( .A(n10689), .ZN(n10691) );
  NAND2_X1 U13806 ( .A1(n10855), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10690) );
  AND2_X1 U13807 ( .A1(n10691), .A2(n10690), .ZN(n13324) );
  INV_X1 U13808 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13809 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13810 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13811 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13812 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10693) );
  NAND4_X1 U13813 ( .A1(n10696), .A2(n10695), .A3(n10694), .A4(n10693), .ZN(
        n10702) );
  AOI22_X1 U13814 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13815 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13816 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13817 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10697) );
  NAND4_X1 U13818 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10701) );
  NOR2_X1 U13819 ( .A1(n10702), .A2(n10701), .ZN(n11978) );
  OAI22_X1 U13820 ( .A1(n10853), .A2(n10703), .B1(n10831), .B2(n11978), .ZN(
        n10704) );
  INV_X1 U13821 ( .A(n10704), .ZN(n10706) );
  AOI22_X1 U13822 ( .A1(n10728), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10854), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U13823 ( .A1(n10706), .A2(n10705), .ZN(n13696) );
  NAND2_X1 U13824 ( .A1(n13697), .A2(n13696), .ZN(n13695) );
  INV_X1 U13825 ( .A(n13695), .ZN(n10707) );
  AOI21_X1 U13826 ( .B1(n10818), .B2(n10868), .A(n10707), .ZN(n12814) );
  AOI222_X1 U13827 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n10855), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n10728), .ZN(n12813) );
  NAND2_X1 U13828 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U13829 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10710) );
  NAND2_X1 U13830 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10709) );
  NAND2_X1 U13831 ( .A1(n10641), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10708) );
  NAND2_X1 U13832 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10715) );
  NAND2_X1 U13833 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10714) );
  NAND2_X1 U13834 ( .A1(n10599), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10713) );
  NAND2_X1 U13835 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10712) );
  NAND2_X1 U13836 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10719) );
  NAND2_X1 U13837 ( .A1(n10668), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10718) );
  NAND2_X1 U13838 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10717) );
  NAND2_X1 U13839 ( .A1(n10680), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10716) );
  NAND2_X1 U13840 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10723) );
  NAND2_X1 U13841 ( .A1(n13078), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10722) );
  NAND2_X1 U13842 ( .A1(n10626), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10721) );
  NAND2_X1 U13843 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10720) );
  INV_X1 U13844 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20776) );
  INV_X1 U13845 ( .A(n10729), .ZN(n10849) );
  INV_X1 U13846 ( .A(n10728), .ZN(n10850) );
  INV_X1 U13847 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19015) );
  INV_X1 U13848 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19630) );
  OAI222_X1 U13849 ( .A1(n20776), .A2(n10849), .B1(n10850), .B2(n19015), .C1(
        n10853), .C2(n19630), .ZN(n12818) );
  INV_X1 U13850 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U13851 ( .A1(n10728), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10854), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U13852 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13853 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13854 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13855 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10730) );
  NAND4_X1 U13856 ( .A1(n10733), .A2(n10732), .A3(n10731), .A4(n10730), .ZN(
        n10739) );
  AOI22_X1 U13857 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13858 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13859 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U13860 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10734) );
  NAND4_X1 U13861 ( .A1(n10737), .A2(n10736), .A3(n10735), .A4(n10734), .ZN(
        n10738) );
  NOR2_X1 U13862 ( .A1(n10739), .A2(n10738), .ZN(n13306) );
  INV_X1 U13863 ( .A(n13306), .ZN(n13308) );
  NAND2_X1 U13864 ( .A1(n10818), .A2(n13308), .ZN(n10740) );
  OAI211_X1 U13865 ( .C1(n10853), .C2(n13116), .A(n10741), .B(n10740), .ZN(
        n13113) );
  INV_X1 U13866 ( .A(n13113), .ZN(n10742) );
  INV_X1 U13867 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13868 ( .A1(n10728), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10854), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13869 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10662), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13870 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12432), .ZN(n10745) );
  AOI22_X1 U13871 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13872 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10743) );
  NAND4_X1 U13873 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10752) );
  AOI22_X1 U13874 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n10680), .ZN(n10750) );
  AOI22_X1 U13875 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13876 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13877 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10621), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10747) );
  NAND4_X1 U13878 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10751) );
  NOR2_X1 U13879 ( .A1(n10752), .A2(n10751), .ZN(n13360) );
  INV_X1 U13880 ( .A(n13360), .ZN(n13362) );
  NAND2_X1 U13881 ( .A1(n10818), .A2(n13362), .ZN(n10753) );
  OAI211_X1 U13882 ( .C1(n10853), .C2(n10755), .A(n10754), .B(n10753), .ZN(
        n12951) );
  AOI22_X1 U13883 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13884 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13885 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10681), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13886 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12432), .ZN(n10756) );
  NAND4_X1 U13887 ( .A1(n10759), .A2(n10758), .A3(n10757), .A4(n10756), .ZN(
        n10765) );
  AOI22_X1 U13888 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n10680), .ZN(n10763) );
  AOI22_X1 U13889 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13890 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13891 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10626), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10760) );
  NAND4_X1 U13892 ( .A1(n10763), .A2(n10762), .A3(n10761), .A4(n10760), .ZN(
        n10764) );
  NOR2_X1 U13893 ( .A1(n10765), .A2(n10764), .ZN(n13506) );
  NOR2_X1 U13894 ( .A1(n10831), .A2(n13506), .ZN(n10768) );
  INV_X1 U13895 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n10766) );
  INV_X1 U13896 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12109) );
  OAI22_X1 U13897 ( .A1(n10850), .A2(n10766), .B1(n10849), .B2(n12109), .ZN(
        n10767) );
  AOI211_X1 U13898 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n10855), .A(n10768), 
        .B(n10767), .ZN(n16176) );
  INV_X1 U13899 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U13900 ( .A1(n10728), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13901 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10662), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13902 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12432), .ZN(n10771) );
  AOI22_X1 U13903 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13904 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10769) );
  NAND4_X1 U13905 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10778) );
  AOI22_X1 U13906 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .B2(n10680), .ZN(n10776) );
  AOI22_X1 U13907 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13908 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13909 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10621), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10773) );
  NAND4_X1 U13910 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        n10777) );
  NAND2_X1 U13911 ( .A1(n10818), .A2(n13352), .ZN(n10779) );
  OAI211_X1 U13912 ( .C1(n10853), .C2(n10781), .A(n10780), .B(n10779), .ZN(
        n13101) );
  AOI22_X1 U13913 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10662), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10785) );
  AOI22_X1 U13914 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12432), .ZN(n10784) );
  AOI22_X1 U13915 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13916 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10782) );
  NAND4_X1 U13917 ( .A1(n10785), .A2(n10784), .A3(n10783), .A4(n10782), .ZN(
        n10791) );
  AOI22_X1 U13918 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(n10680), .ZN(n10789) );
  INV_X1 U13919 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n20925) );
  AOI22_X1 U13920 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13921 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13922 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10621), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10786) );
  NAND4_X1 U13923 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10790) );
  INV_X1 U13924 ( .A(n13343), .ZN(n12354) );
  AOI22_X1 U13925 ( .A1(n10728), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10792) );
  OAI21_X1 U13926 ( .B1(n12354), .B2(n10831), .A(n10792), .ZN(n10793) );
  AOI21_X1 U13927 ( .B1(n10855), .B2(P2_REIP_REG_12__SCAN_IN), .A(n10793), 
        .ZN(n13468) );
  AOI22_X1 U13928 ( .A1(n10728), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13929 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U13930 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13931 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13932 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10794) );
  NAND4_X1 U13933 ( .A1(n10797), .A2(n10796), .A3(n10795), .A4(n10794), .ZN(
        n10803) );
  AOI22_X1 U13934 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13935 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U13936 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13937 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10798) );
  NAND4_X1 U13938 ( .A1(n10801), .A2(n10800), .A3(n10799), .A4(n10798), .ZN(
        n10802) );
  NAND2_X1 U13939 ( .A1(n10818), .A2(n13416), .ZN(n10804) );
  OAI211_X1 U13940 ( .C1(n10853), .C2(n20932), .A(n10805), .B(n10804), .ZN(
        n12660) );
  AOI22_X1 U13941 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10662), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13942 ( .A1(n10599), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12432), .ZN(n10808) );
  AOI22_X1 U13943 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13944 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10681), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10806) );
  NAND4_X1 U13945 ( .A1(n10809), .A2(n10808), .A3(n10807), .A4(n10806), .ZN(
        n10815) );
  AOI22_X1 U13946 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(n10680), .ZN(n10813) );
  AOI22_X1 U13947 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13948 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U13949 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n13078), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10810) );
  NAND4_X1 U13950 ( .A1(n10813), .A2(n10812), .A3(n10811), .A4(n10810), .ZN(
        n10814) );
  INV_X1 U13951 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n13619) );
  AOI22_X1 U13952 ( .A1(n10728), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10816) );
  OAI21_X1 U13953 ( .B1(n10853), .B2(n13619), .A(n10816), .ZN(n10817) );
  AOI21_X1 U13954 ( .B1(n10818), .B2(n13562), .A(n10817), .ZN(n13617) );
  AOI22_X1 U13955 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10662), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13956 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12432), .ZN(n10821) );
  AOI22_X1 U13957 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13958 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U13959 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10828) );
  AOI22_X1 U13960 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n10680), .ZN(n10826) );
  AOI22_X1 U13961 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13962 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13963 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10621), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10823) );
  NAND4_X1 U13964 ( .A1(n10826), .A2(n10825), .A3(n10824), .A4(n10823), .ZN(
        n10827) );
  NOR2_X1 U13965 ( .A1(n10828), .A2(n10827), .ZN(n13636) );
  NAND2_X1 U13966 ( .A1(n10855), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13967 ( .A1(n10728), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10829) );
  OAI211_X1 U13968 ( .C1(n13636), .C2(n10831), .A(n10830), .B(n10829), .ZN(
        n12650) );
  INV_X1 U13969 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13970 ( .A1(n10728), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10832) );
  OAI21_X1 U13971 ( .B1(n10853), .B2(n10833), .A(n10832), .ZN(n13644) );
  INV_X1 U13972 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19644) );
  AOI22_X1 U13973 ( .A1(n10728), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10834) );
  OAI21_X1 U13974 ( .B1(n10853), .B2(n19644), .A(n10834), .ZN(n13642) );
  INV_X1 U13975 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19646) );
  AOI22_X1 U13976 ( .A1(n10728), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10835) );
  OAI21_X1 U13977 ( .B1(n10853), .B2(n19646), .A(n10835), .ZN(n10836) );
  INV_X1 U13978 ( .A(n10836), .ZN(n13854) );
  OR2_X2 U13979 ( .A1(n13855), .A2(n13854), .ZN(n13857) );
  INV_X1 U13980 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19648) );
  AOI22_X1 U13981 ( .A1(n10728), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10837) );
  OAI21_X1 U13982 ( .B1(n10853), .B2(n19648), .A(n10837), .ZN(n10838) );
  INV_X1 U13983 ( .A(n10838), .ZN(n13793) );
  NOR2_X2 U13984 ( .A1(n13857), .A2(n13793), .ZN(n15320) );
  INV_X1 U13985 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U13986 ( .A1(n10728), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10839) );
  OAI21_X1 U13987 ( .B1(n10853), .B2(n15128), .A(n10839), .ZN(n15319) );
  INV_X1 U13988 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19651) );
  AOI22_X1 U13989 ( .A1(n10728), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10840) );
  OAI21_X1 U13990 ( .B1(n10853), .B2(n19651), .A(n10840), .ZN(n13833) );
  NAND2_X1 U13991 ( .A1(n15322), .A2(n13833), .ZN(n13834) );
  INV_X1 U13992 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13993 ( .A1(n10728), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10841) );
  OAI21_X1 U13994 ( .B1(n10853), .B2(n10842), .A(n10841), .ZN(n15299) );
  INV_X1 U13995 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15011) );
  INV_X1 U13996 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15283) );
  OAI22_X1 U13997 ( .A1(n10850), .A2(n15011), .B1(n10849), .B2(n15283), .ZN(
        n10843) );
  AOI21_X1 U13998 ( .B1(n10855), .B2(P2_REIP_REG_23__SCAN_IN), .A(n10843), 
        .ZN(n14881) );
  INV_X1 U13999 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15004) );
  INV_X1 U14000 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15262) );
  OAI22_X1 U14001 ( .A1(n10850), .A2(n15004), .B1(n10849), .B2(n15262), .ZN(
        n10844) );
  AOI21_X1 U14002 ( .B1(n10855), .B2(P2_REIP_REG_24__SCAN_IN), .A(n10844), 
        .ZN(n15003) );
  INV_X1 U14003 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19658) );
  AOI22_X1 U14004 ( .A1(n10728), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10845) );
  OAI21_X1 U14005 ( .B1(n10853), .B2(n19658), .A(n10845), .ZN(n14863) );
  AND2_X2 U14006 ( .A1(n15001), .A2(n14863), .ZN(n14988) );
  INV_X1 U14007 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19660) );
  AOI22_X1 U14008 ( .A1(n10728), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10846) );
  OAI21_X1 U14009 ( .B1(n10853), .B2(n19660), .A(n10846), .ZN(n14987) );
  INV_X1 U14010 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14981) );
  INV_X1 U14011 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15227) );
  OAI22_X1 U14012 ( .A1(n10850), .A2(n14981), .B1(n10849), .B2(n15227), .ZN(
        n10847) );
  AOI21_X1 U14013 ( .B1(n10855), .B2(P2_REIP_REG_27__SCAN_IN), .A(n10847), 
        .ZN(n14977) );
  INV_X1 U14014 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14970) );
  INV_X1 U14015 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15213) );
  OAI22_X1 U14016 ( .A1(n10850), .A2(n14970), .B1(n10849), .B2(n15213), .ZN(
        n10848) );
  AOI21_X1 U14017 ( .B1(n10855), .B2(P2_REIP_REG_28__SCAN_IN), .A(n10848), 
        .ZN(n14856) );
  INV_X1 U14018 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14963) );
  INV_X1 U14019 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15200) );
  OAI22_X1 U14020 ( .A1(n10850), .A2(n14963), .B1(n10849), .B2(n15200), .ZN(
        n10851) );
  AOI21_X1 U14021 ( .B1(n10855), .B2(P2_REIP_REG_29__SCAN_IN), .A(n10851), 
        .ZN(n14213) );
  INV_X1 U14022 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n15026) );
  AOI22_X1 U14023 ( .A1(n10728), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10852) );
  OAI21_X1 U14024 ( .B1(n10853), .B2(n15026), .A(n10852), .ZN(n12613) );
  AOI222_X1 U14025 ( .A1(n10855), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10854), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n10728), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n10856) );
  INV_X1 U14026 ( .A(n10856), .ZN(n10857) );
  NOR2_X1 U14027 ( .A1(n19601), .A2(n19619), .ZN(n19610) );
  NOR2_X1 U14028 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19612) );
  NOR3_X1 U14029 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19610), .A3(n19612), 
        .ZN(n12791) );
  NAND2_X1 U14030 ( .A1(n19600), .A2(n12791), .ZN(n12691) );
  INV_X1 U14031 ( .A(n12691), .ZN(n13249) );
  NAND2_X1 U14032 ( .A1(n19736), .A2(n13249), .ZN(n13265) );
  NOR2_X1 U14033 ( .A1(n12047), .A2(n13265), .ZN(n10858) );
  INV_X1 U14034 ( .A(n18900), .ZN(n15397) );
  NOR3_X1 U14035 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10859), .A3(n19731), 
        .ZN(n16211) );
  NOR2_X1 U14036 ( .A1(n16211), .A2(n18912), .ZN(n10860) );
  NAND2_X1 U14037 ( .A1(n18885), .A2(n10860), .ZN(n10861) );
  NAND2_X1 U14038 ( .A1(n18918), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18931) );
  INV_X2 U14039 ( .A(n18931), .ZN(n18906) );
  AND2_X1 U14040 ( .A1(n12312), .A2(n12228), .ZN(n12238) );
  NOR2_X1 U14041 ( .A1(n10862), .A2(n12238), .ZN(n12040) );
  INV_X1 U14042 ( .A(n12070), .ZN(n10865) );
  INV_X1 U14043 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13421) );
  NAND3_X1 U14044 ( .A1(n12170), .A2(n13421), .A3(n18920), .ZN(n10863) );
  NAND2_X1 U14045 ( .A1(n10864), .A2(n10863), .ZN(n12071) );
  NAND2_X1 U14046 ( .A1(n10865), .A2(n12071), .ZN(n12075) );
  MUX2_X1 U14047 ( .A(n10866), .B(P2_EBX_REG_3__SCAN_IN), .S(n12170), .Z(
        n12074) );
  MUX2_X1 U14048 ( .A(n10867), .B(n12242), .S(n12312), .Z(n12042) );
  MUX2_X1 U14049 ( .A(n12042), .B(n10479), .S(n13389), .Z(n12081) );
  MUX2_X1 U14050 ( .A(n11978), .B(P2_EBX_REG_5__SCAN_IN), .S(n13389), .Z(
        n12065) );
  MUX2_X1 U14051 ( .A(n12015), .B(P2_EBX_REG_6__SCAN_IN), .S(n13389), .Z(
        n12088) );
  MUX2_X1 U14052 ( .A(n15043), .B(n10869), .S(n13389), .Z(n12098) );
  AND2_X2 U14053 ( .A1(n12100), .A2(n12098), .ZN(n12096) );
  NAND2_X1 U14054 ( .A1(n13389), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12095) );
  NAND2_X1 U14055 ( .A1(n12170), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10870) );
  NAND2_X1 U14056 ( .A1(n10871), .A2(n13571), .ZN(n10872) );
  NAND2_X1 U14057 ( .A1(n12186), .A2(n12130), .ZN(n12128) );
  NAND2_X1 U14058 ( .A1(n12170), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12126) );
  NAND2_X1 U14059 ( .A1(n12128), .A2(n12126), .ZN(n12146) );
  INV_X1 U14060 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n13865) );
  INV_X1 U14061 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U14062 ( .A1(n13865), .A2(n10874), .ZN(n10875) );
  AND2_X1 U14063 ( .A1(n13389), .A2(n10875), .ZN(n10876) );
  NAND2_X1 U14064 ( .A1(n13389), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10877) );
  INV_X1 U14065 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14923) );
  INV_X1 U14066 ( .A(n12191), .ZN(n10879) );
  NAND2_X1 U14067 ( .A1(n12170), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16014) );
  AND2_X1 U14068 ( .A1(n12170), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12192) );
  AND2_X1 U14069 ( .A1(n13389), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12201) );
  NOR2_X1 U14070 ( .A1(n12203), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10878) );
  MUX2_X1 U14071 ( .A(n10879), .B(n10878), .S(n13389), .Z(n12206) );
  INV_X1 U14072 ( .A(n12206), .ZN(n10883) );
  INV_X1 U14073 ( .A(n10880), .ZN(n12640) );
  OR2_X1 U14074 ( .A1(n10881), .A2(n12640), .ZN(n12644) );
  NAND2_X1 U14075 ( .A1(n13241), .A2(n16213), .ZN(n12665) );
  NAND2_X1 U14076 ( .A1(n19035), .A2(n13265), .ZN(n12642) );
  OAI21_X1 U14077 ( .B1(n10883), .B2(n12644), .A(n12642), .ZN(n10884) );
  AOI22_X1 U14078 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18906), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n10884), .ZN(n10885) );
  INV_X1 U14079 ( .A(n10885), .ZN(n10887) );
  INV_X1 U14080 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19671) );
  NOR2_X1 U14081 ( .A1(n10887), .A2(n10886), .ZN(n10888) );
  NAND2_X1 U14082 ( .A1(n9703), .A2(n10228), .ZN(P2_U2824) );
  NOR2_X2 U14083 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n10890), .ZN(
        n10897) );
  AND2_X2 U14084 ( .A1(n10897), .A2(n12928), .ZN(n11063) );
  INV_X1 U14085 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10891) );
  NOR2_X4 U14086 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10900) );
  AND2_X2 U14087 ( .A1(n10901), .A2(n10900), .ZN(n11068) );
  AOI22_X1 U14088 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10896) );
  NOR2_X4 U14089 ( .A1(n10892), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10899) );
  AND2_X2 U14090 ( .A1(n10897), .A2(n10899), .ZN(n10984) );
  NOR2_X4 U14091 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10898) );
  AND2_X2 U14092 ( .A1(n10902), .A2(n10898), .ZN(n11101) );
  AOI22_X1 U14093 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11101), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10895) );
  AND2_X2 U14094 ( .A1(n10897), .A2(n10900), .ZN(n10969) );
  AOI22_X1 U14095 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10894) );
  NAND4_X1 U14096 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n10909) );
  AND2_X2 U14097 ( .A1(n10902), .A2(n10897), .ZN(n10974) );
  AOI22_X1 U14098 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10907) );
  AND2_X2 U14099 ( .A1(n10898), .A2(n12928), .ZN(n11069) );
  AOI22_X1 U14100 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10906) );
  AND2_X2 U14101 ( .A1(n10899), .A2(n10903), .ZN(n11102) );
  AOI22_X1 U14102 ( .A1(n11102), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10905) );
  AND2_X2 U14103 ( .A1(n10902), .A2(n10901), .ZN(n10979) );
  BUF_X2 U14104 ( .A(n10979), .Z(n11641) );
  AOI22_X1 U14105 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11070), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10904) );
  NAND4_X1 U14106 ( .A1(n10907), .A2(n10906), .A3(n10905), .A4(n10904), .ZN(
        n10908) );
  INV_X1 U14107 ( .A(n20018), .ZN(n10920) );
  AOI22_X1 U14108 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U14109 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11095), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U14110 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U14111 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10910) );
  NAND4_X1 U14112 ( .A1(n10913), .A2(n10912), .A3(n10911), .A4(n10910), .ZN(
        n10919) );
  AOI22_X1 U14113 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U14114 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11102), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U14115 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11070), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U14116 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10914) );
  NAND4_X1 U14117 ( .A1(n10917), .A2(n10916), .A3(n10915), .A4(n10914), .ZN(
        n10918) );
  AND2_X2 U14118 ( .A1(n10920), .A2(n20022), .ZN(n11029) );
  AOI22_X1 U14119 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11063), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U14120 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11101), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U14121 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9649), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U14122 ( .A1(n11102), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11070), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U14123 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U14124 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U14125 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U14126 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10925) );
  NAND2_X1 U14127 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10934) );
  NAND2_X1 U14128 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10933) );
  NAND2_X1 U14129 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10932) );
  NAND2_X1 U14130 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10931) );
  NAND2_X1 U14131 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10937) );
  NAND2_X1 U14132 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10936) );
  NAND2_X1 U14133 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10935) );
  NAND2_X1 U14134 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10941) );
  NAND2_X1 U14135 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10940) );
  NAND2_X1 U14136 ( .A1(n11102), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10939) );
  NAND2_X1 U14137 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10938) );
  NAND2_X1 U14138 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10945) );
  NAND2_X1 U14139 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10944) );
  NAND2_X1 U14140 ( .A1(n10979), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10943) );
  NAND2_X1 U14141 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10942) );
  NAND2_X1 U14142 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10952) );
  NAND2_X1 U14143 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10951) );
  NAND2_X1 U14144 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10950) );
  NAND2_X1 U14145 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10949) );
  NAND2_X1 U14146 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10956) );
  NAND2_X1 U14147 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10955) );
  NAND2_X1 U14148 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10954) );
  NAND2_X1 U14149 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10953) );
  NAND2_X1 U14150 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10960) );
  NAND2_X1 U14151 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10959) );
  NAND2_X1 U14152 ( .A1(n11102), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10958) );
  NAND2_X1 U14153 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10957) );
  AND4_X2 U14154 ( .A1(n10960), .A2(n10959), .A3(n10958), .A4(n10957), .ZN(
        n10966) );
  NAND2_X1 U14155 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10964) );
  NAND2_X1 U14156 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10963) );
  NAND2_X1 U14157 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10962) );
  NAND2_X1 U14158 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10961) );
  NAND4_X4 U14159 ( .A1(n10968), .A2(n10967), .A3(n10966), .A4(n10965), .ZN(
        n20029) );
  AND3_X2 U14160 ( .A1(n11029), .A2(n11033), .A3(n12874), .ZN(n12892) );
  NAND2_X1 U14161 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10973) );
  NAND2_X1 U14162 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10972) );
  NAND2_X1 U14163 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10971) );
  NAND2_X1 U14164 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10970) );
  NAND2_X1 U14165 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10978) );
  NAND2_X1 U14166 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10977) );
  NAND2_X1 U14167 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10976) );
  NAND2_X1 U14168 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10975) );
  NAND2_X1 U14169 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10983) );
  NAND2_X1 U14170 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10982) );
  NAND2_X1 U14171 ( .A1(n11102), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10981) );
  NAND2_X1 U14172 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10980) );
  NAND2_X1 U14173 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U14174 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10987) );
  NAND2_X1 U14175 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10985) );
  NAND2_X2 U14176 ( .A1(n12892), .A2(n9956), .ZN(n12782) );
  AOI22_X1 U14177 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U14178 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11095), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U14179 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14180 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10993) );
  NAND4_X1 U14181 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n11002) );
  AOI22_X1 U14182 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14183 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11102), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14184 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11070), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14185 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10997) );
  NAND4_X1 U14186 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11001) );
  NOR2_X4 U14187 ( .A1(n12782), .A2(n14461), .ZN(n13020) );
  XNOR2_X1 U14188 ( .A(n11003), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n12773) );
  NAND2_X1 U14189 ( .A1(n13020), .A2(n12773), .ZN(n11057) );
  NAND2_X1 U14190 ( .A1(n11063), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11007) );
  NAND2_X1 U14191 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11006) );
  NAND2_X1 U14192 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11005) );
  NAND2_X1 U14193 ( .A1(n11102), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11004) );
  NAND2_X1 U14194 ( .A1(n10969), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U14195 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U14196 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U14197 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11008) );
  AND4_X2 U14198 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n11022) );
  NAND2_X1 U14199 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11015) );
  NAND2_X1 U14200 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11014) );
  NAND2_X1 U14201 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U14202 ( .A1(n11069), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11012) );
  NAND2_X1 U14203 ( .A1(n11101), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U14204 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11018) );
  NAND2_X1 U14205 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U14206 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11016) );
  NAND4_X4 U14207 ( .A1(n11023), .A2(n11022), .A3(n11021), .A4(n11020), .ZN(
        n20014) );
  OR2_X1 U14208 ( .A1(n12774), .A2(n20014), .ZN(n12954) );
  OAI21_X1 U14209 ( .B1(n12954), .B2(n13021), .A(n13030), .ZN(n11024) );
  INV_X1 U14210 ( .A(n11024), .ZN(n11051) );
  NAND2_X1 U14211 ( .A1(n9956), .A2(n20018), .ZN(n12906) );
  NAND2_X1 U14212 ( .A1(n12973), .A2(n13021), .ZN(n11026) );
  NAND2_X1 U14213 ( .A1(n12889), .A2(n12929), .ZN(n11031) );
  INV_X1 U14214 ( .A(n11029), .ZN(n11030) );
  NAND2_X1 U14215 ( .A1(n14180), .A2(n11030), .ZN(n12778) );
  INV_X2 U14216 ( .A(n11033), .ZN(n20033) );
  NAND2_X1 U14217 ( .A1(n20029), .A2(n20033), .ZN(n11034) );
  MUX2_X1 U14218 ( .A(n11034), .B(n12780), .S(n20018), .Z(n11036) );
  NAND3_X2 U14219 ( .A1(n11037), .A2(n11036), .A3(n11035), .ZN(n12899) );
  INV_X1 U14220 ( .A(n13277), .ZN(n12900) );
  NAND2_X1 U14221 ( .A1(n12900), .A2(n13019), .ZN(n11038) );
  OAI21_X1 U14222 ( .B1(n12899), .B2(n11038), .A(n14122), .ZN(n11039) );
  NAND3_X1 U14223 ( .A1(n11057), .A2(n10244), .A3(n11039), .ZN(n11043) );
  NOR2_X1 U14224 ( .A1(n12899), .A2(n11041), .ZN(n12736) );
  NAND2_X1 U14225 ( .A1(n12736), .A2(n13019), .ZN(n12882) );
  INV_X1 U14226 ( .A(n20649), .ZN(n11044) );
  MUX2_X1 U14227 ( .A(n11044), .B(n11872), .S(n20464), .Z(n11045) );
  NAND2_X1 U14228 ( .A1(n13277), .A2(n11033), .ZN(n11046) );
  AND2_X1 U14229 ( .A1(n11046), .A2(n12906), .ZN(n13028) );
  NAND2_X1 U14230 ( .A1(n14122), .A2(n20014), .ZN(n14383) );
  NAND3_X1 U14231 ( .A1(n14383), .A2(n20720), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11047) );
  AOI21_X1 U14232 ( .B1(n20756), .B2(n11048), .A(n11047), .ZN(n11050) );
  NAND3_X1 U14233 ( .A1(n12889), .A2(n20014), .A3(n12929), .ZN(n11049) );
  AND2_X2 U14234 ( .A1(n14122), .A2(n13019), .ZN(n14381) );
  NAND3_X1 U14235 ( .A1(n12968), .A2(n12973), .A3(n20022), .ZN(n11052) );
  NAND2_X1 U14236 ( .A1(n12899), .A2(n11052), .ZN(n11053) );
  NAND2_X1 U14237 ( .A1(n11054), .A2(n11053), .ZN(n11092) );
  INV_X1 U14238 ( .A(n11062), .ZN(n11061) );
  NAND2_X1 U14239 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11134) );
  OAI21_X1 U14240 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11134), .ZN(n20354) );
  NAND2_X1 U14241 ( .A1(n20649), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11128) );
  OAI21_X1 U14242 ( .B1(n11872), .B2(n20354), .A(n11128), .ZN(n11055) );
  INV_X1 U14243 ( .A(n11055), .ZN(n11056) );
  INV_X1 U14244 ( .A(n11057), .ZN(n11058) );
  NAND3_X1 U14245 ( .A1(n14381), .A2(n11324), .A3(n13277), .ZN(n12907) );
  INV_X1 U14246 ( .A(n20110), .ZN(n11060) );
  AOI22_X1 U14247 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11067) );
  BUF_X2 U14248 ( .A(n11101), .Z(n11838) );
  AOI22_X1 U14249 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14250 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U14251 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11064) );
  NAND4_X1 U14252 ( .A1(n11067), .A2(n11066), .A3(n11065), .A4(n11064), .ZN(
        n11076) );
  AOI22_X1 U14253 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11074) );
  INV_X1 U14254 ( .A(n11100), .ZN(n11184) );
  AOI22_X1 U14255 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11073) );
  BUF_X1 U14256 ( .A(n11069), .Z(n11636) );
  AOI22_X1 U14257 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11072) );
  BUF_X2 U14258 ( .A(n11102), .Z(n11849) );
  AOI22_X1 U14259 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11071) );
  NAND4_X1 U14260 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11075) );
  AOI22_X1 U14261 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U14262 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14263 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14264 ( .A1(n11100), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11078) );
  NAND4_X1 U14265 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11087) );
  AOI22_X1 U14266 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14267 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14268 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11082) );
  NAND4_X1 U14269 ( .A1(n11085), .A2(n11084), .A3(n11083), .A4(n11082), .ZN(
        n11086) );
  NAND2_X1 U14270 ( .A1(n11088), .A2(n11121), .ZN(n11194) );
  OAI21_X1 U14271 ( .B1(n11088), .B2(n11121), .A(n11194), .ZN(n11089) );
  OAI211_X1 U14272 ( .C1(n11089), .C2(n12954), .A(n11029), .B(n20029), .ZN(
        n11090) );
  INV_X1 U14273 ( .A(n11090), .ZN(n11091) );
  INV_X1 U14274 ( .A(n11092), .ZN(n11093) );
  XNOR2_X1 U14275 ( .A(n11094), .B(n11093), .ZN(n11379) );
  NAND2_X1 U14276 ( .A1(n11379), .A2(n20759), .ZN(n11111) );
  AOI22_X1 U14277 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14278 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14279 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14280 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11096) );
  NAND4_X1 U14281 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11108) );
  AOI22_X1 U14282 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11100), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14283 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14284 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14285 ( .A1(n9632), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11103) );
  NAND4_X1 U14286 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n11107) );
  NAND2_X1 U14287 ( .A1(n13021), .A2(n11291), .ZN(n11115) );
  NOR2_X1 U14288 ( .A1(n11178), .A2(n11291), .ZN(n11156) );
  MUX2_X1 U14289 ( .A(n11287), .B(n11156), .S(n11121), .Z(n11109) );
  INV_X1 U14290 ( .A(n11109), .ZN(n11110) );
  INV_X1 U14291 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11114) );
  AOI21_X1 U14292 ( .B1(n14122), .B2(n11121), .A(n20759), .ZN(n11116) );
  AND2_X1 U14293 ( .A1(n11116), .A2(n11115), .ZN(n11117) );
  NAND2_X1 U14294 ( .A1(n20014), .A2(n20029), .ZN(n11308) );
  NAND2_X1 U14295 ( .A1(n14122), .A2(n20022), .ZN(n11163) );
  OAI21_X1 U14296 ( .B1(n12954), .B2(n11121), .A(n11163), .ZN(n11122) );
  INV_X1 U14297 ( .A(n11122), .ZN(n11123) );
  INV_X1 U14298 ( .A(n11124), .ZN(n11125) );
  OR2_X1 U14299 ( .A1(n12943), .A2(n11125), .ZN(n11126) );
  INV_X1 U14300 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19978) );
  INV_X1 U14301 ( .A(n11127), .ZN(n11130) );
  NAND2_X1 U14302 ( .A1(n11128), .A2(n10892), .ZN(n11129) );
  NAND2_X1 U14303 ( .A1(n11130), .A2(n11129), .ZN(n11131) );
  NAND2_X2 U14304 ( .A1(n11132), .A2(n11131), .ZN(n11140) );
  INV_X1 U14305 ( .A(n11134), .ZN(n11133) );
  NAND2_X1 U14306 ( .A1(n11133), .A2(n20428), .ZN(n20388) );
  NAND2_X1 U14307 ( .A1(n11134), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11135) );
  NAND2_X1 U14308 ( .A1(n20649), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11137) );
  AOI22_X1 U14309 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14310 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14311 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14312 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11141) );
  NAND4_X1 U14313 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11150) );
  AOI22_X1 U14314 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14315 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14316 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11146) );
  AOI22_X1 U14317 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11145) );
  NAND4_X1 U14318 ( .A1(n11148), .A2(n11147), .A3(n11146), .A4(n11145), .ZN(
        n11149) );
  INV_X1 U14319 ( .A(n11177), .ZN(n20763) );
  AOI22_X1 U14320 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n20763), .B2(n11151), .ZN(n11152) );
  INV_X1 U14321 ( .A(n11287), .ZN(n11153) );
  INV_X1 U14322 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11155) );
  OR2_X1 U14323 ( .A1(n11356), .A2(n11155), .ZN(n11158) );
  INV_X1 U14324 ( .A(n11156), .ZN(n11157) );
  INV_X1 U14325 ( .A(n11308), .ZN(n11286) );
  NAND2_X1 U14326 ( .A1(n11364), .A2(n11286), .ZN(n11167) );
  XNOR2_X1 U14327 ( .A(n11194), .B(n11193), .ZN(n11165) );
  INV_X1 U14328 ( .A(n11163), .ZN(n11164) );
  AOI21_X1 U14329 ( .B1(n11165), .B2(n20756), .A(n11164), .ZN(n11166) );
  NAND2_X1 U14330 ( .A1(n11167), .A2(n11166), .ZN(n12987) );
  NAND2_X1 U14331 ( .A1(n11168), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11169) );
  INV_X1 U14332 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13088) );
  INV_X1 U14333 ( .A(n11170), .ZN(n11172) );
  INV_X1 U14334 ( .A(n11872), .ZN(n11174) );
  NAND3_X1 U14335 ( .A1(n20737), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20260) );
  INV_X1 U14336 ( .A(n20260), .ZN(n20254) );
  NAND2_X1 U14337 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20254), .ZN(
        n20286) );
  NAND2_X1 U14338 ( .A1(n20737), .A2(n20286), .ZN(n11173) );
  NAND3_X1 U14339 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20574) );
  INV_X1 U14340 ( .A(n20574), .ZN(n20578) );
  NAND2_X1 U14341 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20578), .ZN(
        n20638) );
  AOI22_X1 U14342 ( .A1(n11174), .A2(n20004), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20649), .ZN(n11175) );
  INV_X1 U14343 ( .A(n10974), .ZN(n11179) );
  INV_X2 U14344 ( .A(n11179), .ZN(n11846) );
  AOI22_X1 U14345 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14346 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14347 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11181) );
  AOI22_X1 U14348 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11180) );
  NAND4_X1 U14349 ( .A1(n11183), .A2(n11182), .A3(n11181), .A4(n11180), .ZN(
        n11190) );
  INV_X2 U14350 ( .A(n11184), .ZN(n13274) );
  AOI22_X1 U14351 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14352 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14353 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14354 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11185) );
  NAND4_X1 U14355 ( .A1(n11188), .A2(n11187), .A3(n11186), .A4(n11185), .ZN(
        n11189) );
  AOI22_X1 U14356 ( .A1(n11354), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11331), .B2(n11240), .ZN(n11191) );
  XNOR2_X2 U14357 ( .A(n11202), .B(n19999), .ZN(n20730) );
  NAND2_X1 U14358 ( .A1(n20730), .A2(n11286), .ZN(n11198) );
  NAND2_X1 U14359 ( .A1(n11194), .A2(n11193), .ZN(n11242) );
  INV_X1 U14360 ( .A(n11240), .ZN(n11195) );
  XNOR2_X1 U14361 ( .A(n11242), .B(n11195), .ZN(n11196) );
  NAND2_X1 U14362 ( .A1(n11196), .A2(n20756), .ZN(n11197) );
  NAND2_X1 U14363 ( .A1(n11198), .A2(n11197), .ZN(n13312) );
  NAND2_X1 U14364 ( .A1(n11199), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11200) );
  INV_X1 U14365 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11201) );
  INV_X1 U14366 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11204) );
  OR2_X1 U14367 ( .A1(n11356), .A2(n11204), .ZN(n11217) );
  AOI22_X1 U14368 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11846), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11209) );
  INV_X1 U14369 ( .A(n10969), .ZN(n11205) );
  AOI22_X1 U14370 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11817), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14371 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11847), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14372 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11206) );
  NAND4_X1 U14373 ( .A1(n11209), .A2(n11208), .A3(n11207), .A4(n11206), .ZN(
        n11215) );
  AOI22_X1 U14374 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14375 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11838), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14376 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11211) );
  INV_X1 U14377 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20913) );
  NAND4_X1 U14378 ( .A1(n11213), .A2(n11212), .A3(n11211), .A4(n11210), .ZN(
        n11214) );
  NAND2_X1 U14379 ( .A1(n11331), .A2(n11239), .ZN(n11216) );
  NAND2_X1 U14380 ( .A1(n11217), .A2(n11216), .ZN(n11224) );
  XNOR2_X1 U14381 ( .A(n11225), .B(n11224), .ZN(n11399) );
  NAND2_X1 U14382 ( .A1(n11399), .A2(n11286), .ZN(n11221) );
  NAND2_X1 U14383 ( .A1(n11242), .A2(n11240), .ZN(n11218) );
  XNOR2_X1 U14384 ( .A(n11218), .B(n11239), .ZN(n11219) );
  NAND2_X1 U14385 ( .A1(n11219), .A2(n20756), .ZN(n11220) );
  NAND2_X1 U14386 ( .A1(n11221), .A2(n11220), .ZN(n19934) );
  NAND2_X1 U14387 ( .A1(n11222), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11223) );
  INV_X1 U14388 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11226) );
  OR2_X1 U14389 ( .A1(n11356), .A2(n11226), .ZN(n11238) );
  AOI22_X1 U14390 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14391 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14392 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14393 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11227) );
  NAND4_X1 U14394 ( .A1(n11230), .A2(n11229), .A3(n11228), .A4(n11227), .ZN(
        n11236) );
  AOI22_X1 U14395 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14396 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11233) );
  AOI22_X1 U14397 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11232) );
  AOI22_X1 U14398 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11231) );
  NAND4_X1 U14399 ( .A1(n11234), .A2(n11233), .A3(n11232), .A4(n11231), .ZN(
        n11235) );
  NAND2_X1 U14400 ( .A1(n11331), .A2(n11277), .ZN(n11237) );
  NAND2_X1 U14401 ( .A1(n11238), .A2(n11237), .ZN(n11248) );
  XNOR2_X1 U14402 ( .A(n11249), .B(n11248), .ZN(n11400) );
  NAND2_X1 U14403 ( .A1(n11400), .A2(n11286), .ZN(n11245) );
  AND2_X1 U14404 ( .A1(n11240), .A2(n11239), .ZN(n11241) );
  NAND2_X1 U14405 ( .A1(n11242), .A2(n11241), .ZN(n11279) );
  XNOR2_X1 U14406 ( .A(n11279), .B(n11277), .ZN(n11243) );
  NAND2_X1 U14407 ( .A1(n11243), .A2(n20756), .ZN(n11244) );
  NAND2_X1 U14408 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  INV_X1 U14409 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15982) );
  XNOR2_X1 U14410 ( .A(n11246), .B(n15982), .ZN(n15916) );
  NAND2_X1 U14411 ( .A1(n11246), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11247) );
  INV_X1 U14412 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11250) );
  OR2_X1 U14413 ( .A1(n11356), .A2(n11250), .ZN(n11262) );
  AOI22_X1 U14414 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14415 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14416 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14417 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11251) );
  NAND4_X1 U14418 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11260) );
  AOI22_X1 U14419 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14420 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14421 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14422 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11255) );
  NAND4_X1 U14423 ( .A1(n11258), .A2(n11257), .A3(n11256), .A4(n11255), .ZN(
        n11259) );
  NAND2_X1 U14424 ( .A1(n11331), .A2(n11276), .ZN(n11261) );
  INV_X1 U14425 ( .A(n11263), .ZN(n11264) );
  NAND2_X1 U14426 ( .A1(n9705), .A2(n11264), .ZN(n11265) );
  AND2_X1 U14427 ( .A1(n11285), .A2(n11265), .ZN(n11413) );
  NAND2_X1 U14428 ( .A1(n11413), .A2(n11286), .ZN(n11270) );
  INV_X1 U14429 ( .A(n11279), .ZN(n11266) );
  NAND2_X1 U14430 ( .A1(n11266), .A2(n11277), .ZN(n11267) );
  XNOR2_X1 U14431 ( .A(n11267), .B(n11276), .ZN(n11268) );
  NAND2_X1 U14432 ( .A1(n11268), .A2(n20756), .ZN(n11269) );
  NAND2_X1 U14433 ( .A1(n11270), .A2(n11269), .ZN(n13607) );
  OR2_X1 U14434 ( .A1(n13607), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11271) );
  NAND2_X1 U14435 ( .A1(n13607), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11272) );
  INV_X1 U14436 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11274) );
  NAND2_X1 U14437 ( .A1(n11331), .A2(n11291), .ZN(n11273) );
  OAI21_X1 U14438 ( .B1(n11356), .B2(n11274), .A(n11273), .ZN(n11275) );
  NAND2_X1 U14439 ( .A1(n11448), .A2(n11286), .ZN(n11282) );
  NAND2_X1 U14440 ( .A1(n11277), .A2(n11276), .ZN(n11278) );
  OR2_X1 U14441 ( .A1(n11279), .A2(n11278), .ZN(n11290) );
  XNOR2_X1 U14442 ( .A(n11290), .B(n11291), .ZN(n11280) );
  NAND2_X1 U14443 ( .A1(n11280), .A2(n20756), .ZN(n11281) );
  NAND2_X1 U14444 ( .A1(n11282), .A2(n11281), .ZN(n11283) );
  XNOR2_X1 U14445 ( .A(n11283), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13666) );
  OR2_X1 U14446 ( .A1(n11283), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11284) );
  AND2_X1 U14447 ( .A1(n11287), .A2(n11286), .ZN(n11288) );
  INV_X1 U14448 ( .A(n11290), .ZN(n11292) );
  NAND2_X1 U14449 ( .A1(n11293), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13781) );
  INV_X1 U14450 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15957) );
  NAND2_X1 U14451 ( .A1(n11289), .A2(n15957), .ZN(n11294) );
  NAND2_X2 U14452 ( .A1(n14222), .A2(n11294), .ZN(n14223) );
  NOR2_X1 U14453 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11295) );
  INV_X1 U14454 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14813) );
  NAND2_X1 U14455 ( .A1(n14628), .A2(n14813), .ZN(n14641) );
  NAND2_X1 U14456 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U14457 ( .A1(n14628), .A2(n11296), .ZN(n14639) );
  INV_X1 U14458 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14791) );
  NAND2_X1 U14459 ( .A1(n11289), .A2(n14791), .ZN(n11297) );
  NOR2_X1 U14460 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11298) );
  INV_X1 U14461 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15936) );
  XNOR2_X1 U14462 ( .A(n14628), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15878) );
  NAND2_X1 U14463 ( .A1(n11289), .A2(n15936), .ZN(n15877) );
  NAND2_X1 U14464 ( .A1(n15878), .A2(n15877), .ZN(n11299) );
  INV_X1 U14465 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11300) );
  INV_X1 U14466 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U14467 ( .A1(n11300), .A2(n14226), .ZN(n14638) );
  NOR2_X1 U14468 ( .A1(n14638), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11301) );
  XNOR2_X1 U14469 ( .A(n14628), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14618) );
  AND2_X1 U14470 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14729) );
  INV_X1 U14471 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14610) );
  INV_X1 U14472 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14751) );
  NAND2_X1 U14473 ( .A1(n14610), .A2(n14751), .ZN(n11302) );
  INV_X1 U14474 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14737) );
  INV_X1 U14475 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14744) );
  NAND2_X2 U14476 ( .A1(n14581), .A2(n14580), .ZN(n14517) );
  AND2_X1 U14477 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14687) );
  NAND2_X1 U14478 ( .A1(n14687), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14518) );
  NAND2_X1 U14479 ( .A1(n14517), .A2(n14518), .ZN(n11303) );
  NAND2_X1 U14480 ( .A1(n14581), .A2(n14628), .ZN(n14553) );
  NAND3_X1 U14481 ( .A1(n11303), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14553), .ZN(n14532) );
  INV_X1 U14482 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14705) );
  INV_X1 U14483 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14686) );
  INV_X1 U14484 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14565) );
  NAND3_X1 U14485 ( .A1(n14705), .A2(n14686), .A3(n14565), .ZN(n14519) );
  NOR2_X1 U14486 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11304) );
  INV_X1 U14487 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14658) );
  AND2_X1 U14488 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14193) );
  XNOR2_X1 U14489 ( .A(n11306), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14208) );
  NAND2_X1 U14490 ( .A1(n12929), .A2(n14122), .ZN(n11307) );
  XNOR2_X1 U14491 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11323) );
  NAND2_X1 U14492 ( .A1(n11328), .A2(n11323), .ZN(n11310) );
  NAND2_X1 U14493 ( .A1(n20351), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11309) );
  NAND2_X1 U14494 ( .A1(n11310), .A2(n11309), .ZN(n11343) );
  XNOR2_X1 U14495 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14496 ( .A1(n11343), .A2(n11342), .ZN(n11312) );
  NAND2_X1 U14497 ( .A1(n20428), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14498 ( .A1(n11312), .A2(n11311), .ZN(n11321) );
  XNOR2_X1 U14499 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U14500 ( .A1(n11321), .A2(n11320), .ZN(n11314) );
  NAND2_X1 U14501 ( .A1(n20737), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11313) );
  NAND2_X1 U14502 ( .A1(n11314), .A2(n11313), .ZN(n11319) );
  INV_X1 U14503 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15988) );
  NOR2_X1 U14504 ( .A1(n15988), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11315) );
  INV_X1 U14505 ( .A(n12744), .ZN(n11318) );
  NAND2_X1 U14506 ( .A1(n12744), .A2(n11331), .ZN(n11361) );
  XNOR2_X1 U14507 ( .A(n11321), .B(n11320), .ZN(n12741) );
  INV_X1 U14508 ( .A(n12741), .ZN(n11352) );
  OR2_X1 U14509 ( .A1(n14122), .A2(n20029), .ZN(n11322) );
  NAND2_X1 U14510 ( .A1(n11322), .A2(n13019), .ZN(n11347) );
  XNOR2_X1 U14511 ( .A(n11323), .B(n11328), .ZN(n12740) );
  NAND2_X1 U14512 ( .A1(n11324), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11326) );
  INV_X1 U14513 ( .A(n11326), .ZN(n11325) );
  INV_X1 U14514 ( .A(n11331), .ZN(n11344) );
  OAI21_X1 U14515 ( .B1(n11344), .B2(n13019), .A(n11326), .ZN(n11327) );
  AOI21_X1 U14516 ( .B1(n11354), .B2(n12740), .A(n11327), .ZN(n11337) );
  AOI21_X1 U14517 ( .B1(n12740), .B2(n11355), .A(n11337), .ZN(n11341) );
  INV_X1 U14518 ( .A(n11328), .ZN(n11330) );
  NAND2_X1 U14519 ( .A1(n12914), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11329) );
  NAND2_X1 U14520 ( .A1(n11330), .A2(n11329), .ZN(n11334) );
  INV_X1 U14521 ( .A(n11334), .ZN(n11332) );
  NAND2_X1 U14522 ( .A1(n11332), .A2(n11331), .ZN(n11336) );
  INV_X1 U14523 ( .A(n12874), .ZN(n11333) );
  OAI211_X1 U14524 ( .C1(n13021), .C2(n11334), .A(n11333), .B(n9956), .ZN(
        n11335) );
  AOI22_X1 U14525 ( .A1(n11351), .A2(n11336), .B1(n11347), .B2(n11335), .ZN(
        n11340) );
  INV_X1 U14526 ( .A(n12740), .ZN(n11339) );
  INV_X1 U14527 ( .A(n11337), .ZN(n11338) );
  OAI22_X1 U14528 ( .A1(n11341), .A2(n11340), .B1(n11339), .B2(n11338), .ZN(
        n11345) );
  XNOR2_X1 U14529 ( .A(n11343), .B(n11342), .ZN(n12739) );
  AOI211_X1 U14530 ( .C1(n11347), .C2(n11345), .A(n11344), .B(n12739), .ZN(
        n11349) );
  NAND2_X1 U14531 ( .A1(n11354), .A2(n12739), .ZN(n11346) );
  AOI21_X1 U14532 ( .B1(n11347), .B2(n11346), .A(n11345), .ZN(n11348) );
  OAI22_X1 U14533 ( .A1(n11354), .A2(n11352), .B1(n11349), .B2(n11348), .ZN(
        n11350) );
  OAI21_X1 U14534 ( .B1(n11352), .B2(n11351), .A(n11350), .ZN(n11353) );
  OAI21_X1 U14535 ( .B1(n11354), .B2(n12738), .A(n11353), .ZN(n11358) );
  NAND2_X1 U14536 ( .A1(n11358), .A2(n11357), .ZN(n11359) );
  NAND2_X1 U14537 ( .A1(n11361), .A2(n11360), .ZN(n11362) );
  NAND2_X1 U14538 ( .A1(n11364), .A2(n11569), .ZN(n11369) );
  INV_X1 U14539 ( .A(n13713), .ZN(n13716) );
  NAND2_X1 U14540 ( .A1(n11392), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11367) );
  NOR2_X2 U14541 ( .A1(n20039), .A2(n20750), .ZN(n11408) );
  INV_X1 U14542 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12985) );
  XNOR2_X1 U14543 ( .A(n12985), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19851) );
  OAI21_X1 U14544 ( .B1(n19851), .B2(n14113), .A(n11867), .ZN(n11365) );
  AOI21_X1 U14545 ( .B1(n11408), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11365), .ZN(
        n11366) );
  AND2_X1 U14546 ( .A1(n11367), .A2(n11366), .ZN(n11368) );
  NAND2_X1 U14547 ( .A1(n11369), .A2(n11368), .ZN(n11370) );
  NAND2_X1 U14548 ( .A1(n11864), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11386) );
  NAND2_X1 U14549 ( .A1(n14833), .A2(n11569), .ZN(n11376) );
  AOI22_X1 U14550 ( .A1(n11865), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20750), .ZN(n11374) );
  NAND2_X1 U14551 ( .A1(n11392), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11373) );
  AND2_X1 U14552 ( .A1(n11374), .A2(n11373), .ZN(n11375) );
  NAND2_X1 U14553 ( .A1(n11376), .A2(n11375), .ZN(n12978) );
  NAND2_X1 U14554 ( .A1(n9650), .A2(n11033), .ZN(n11378) );
  NAND2_X1 U14555 ( .A1(n11378), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12880) );
  INV_X1 U14556 ( .A(n11379), .ZN(n11380) );
  INV_X1 U14557 ( .A(n11392), .ZN(n11391) );
  NAND2_X1 U14558 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11382) );
  NAND2_X1 U14559 ( .A1(n11865), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11381) );
  OAI211_X1 U14560 ( .C1(n11391), .C2(n12914), .A(n11382), .B(n11381), .ZN(
        n11383) );
  AOI21_X1 U14561 ( .B1(n20111), .B2(n11569), .A(n11383), .ZN(n12881) );
  OR2_X1 U14562 ( .A1(n12880), .A2(n12881), .ZN(n12878) );
  NAND2_X1 U14563 ( .A1(n12881), .A2(n11858), .ZN(n11384) );
  NAND2_X1 U14564 ( .A1(n12878), .A2(n11384), .ZN(n12977) );
  NAND2_X1 U14565 ( .A1(n12978), .A2(n12977), .ZN(n12981) );
  NAND2_X1 U14566 ( .A1(n20730), .A2(n11569), .ZN(n11390) );
  NAND2_X1 U14567 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11387) );
  AOI21_X1 U14568 ( .B1(n13315), .B2(n11387), .A(n11394), .ZN(n19835) );
  OAI22_X1 U14569 ( .A1(n19835), .A2(n14113), .B1(n11867), .B2(n13315), .ZN(
        n11388) );
  AOI21_X1 U14570 ( .B1(n11408), .B2(P1_EAX_REG_3__SCAN_IN), .A(n11388), .ZN(
        n11389) );
  OAI211_X1 U14571 ( .C1(n11391), .C2(n10890), .A(n11390), .B(n11389), .ZN(
        n13085) );
  NAND2_X1 U14572 ( .A1(n13086), .A2(n13085), .ZN(n13333) );
  NAND2_X1 U14573 ( .A1(n11392), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11397) );
  INV_X1 U14574 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19818) );
  AOI21_X1 U14575 ( .B1(n19818), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11393) );
  AOI21_X1 U14576 ( .B1(n11408), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11393), .ZN(
        n11396) );
  OAI21_X1 U14577 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11394), .A(
        n11401), .ZN(n19942) );
  NOR2_X1 U14578 ( .A1(n19942), .A2(n14113), .ZN(n11395) );
  AOI21_X1 U14579 ( .B1(n11397), .B2(n11396), .A(n11395), .ZN(n11398) );
  AOI21_X1 U14580 ( .B1(n11399), .B2(n11569), .A(n11398), .ZN(n13334) );
  NAND2_X1 U14581 ( .A1(n11400), .A2(n11569), .ZN(n11407) );
  INV_X1 U14582 ( .A(n11401), .ZN(n11403) );
  INV_X1 U14583 ( .A(n11409), .ZN(n11402) );
  OAI21_X1 U14584 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11403), .A(
        n11402), .ZN(n19813) );
  NAND2_X1 U14585 ( .A1(n19813), .A2(n11858), .ZN(n11404) );
  OAI21_X1 U14586 ( .B1(n19809), .B2(n11867), .A(n11404), .ZN(n11405) );
  AOI21_X1 U14587 ( .B1(n11408), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11405), .ZN(
        n11406) );
  NAND2_X1 U14588 ( .A1(n11407), .A2(n11406), .ZN(n13336) );
  INV_X1 U14589 ( .A(n11408), .ZN(n11805) );
  INV_X1 U14590 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11411) );
  OAI21_X1 U14591 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11409), .A(
        n11442), .ZN(n19805) );
  AOI22_X1 U14592 ( .A1(n11858), .A2(n19805), .B1(n11864), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11410) );
  OAI21_X1 U14593 ( .B1(n11805), .B2(n11411), .A(n11410), .ZN(n11412) );
  AOI21_X1 U14594 ( .B1(n11413), .B2(n11569), .A(n11412), .ZN(n13590) );
  INV_X1 U14595 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20945) );
  XOR2_X1 U14596 ( .A(n19774), .B(n11449), .Z(n19778) );
  AOI22_X1 U14597 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11817), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14598 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14599 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14600 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11415) );
  NAND4_X1 U14601 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(
        n11424) );
  AOI22_X1 U14602 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14603 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14604 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11420) );
  NAND4_X1 U14605 ( .A1(n11422), .A2(n11421), .A3(n11420), .A4(n11419), .ZN(
        n11423) );
  OR2_X1 U14606 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  AOI22_X1 U14607 ( .A1(n11569), .A2(n11425), .B1(n11864), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11427) );
  NAND2_X1 U14608 ( .A1(n11865), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11426) );
  OAI211_X1 U14609 ( .C1(n19778), .C2(n14113), .A(n11427), .B(n11426), .ZN(
        n13594) );
  AOI22_X1 U14610 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14611 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14612 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11430) );
  NAND4_X1 U14613 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n11438) );
  AOI22_X1 U14614 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14615 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14616 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14617 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U14618 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11437) );
  OAI21_X1 U14619 ( .B1(n11438), .B2(n11437), .A(n11569), .ZN(n11441) );
  XNOR2_X1 U14620 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11443), .ZN(
        n14373) );
  AOI22_X1 U14621 ( .A1(n11858), .A2(n14373), .B1(n11864), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U14622 ( .A1(n11865), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11439) );
  INV_X1 U14623 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13536) );
  INV_X1 U14624 ( .A(n11442), .ZN(n11445) );
  INV_X1 U14625 ( .A(n11443), .ZN(n11444) );
  OAI21_X1 U14626 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11445), .A(
        n11444), .ZN(n19793) );
  AOI22_X1 U14627 ( .A1(n11858), .A2(n19793), .B1(n11864), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11446) );
  OAI21_X1 U14628 ( .B1(n11805), .B2(n13536), .A(n11446), .ZN(n11447) );
  INV_X1 U14629 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11450) );
  XNOR2_X1 U14630 ( .A(n11479), .B(n11450), .ZN(n15846) );
  OR2_X1 U14631 ( .A1(n15846), .A2(n14113), .ZN(n11465) );
  AOI22_X1 U14632 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14633 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14634 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14635 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11451) );
  NAND4_X1 U14636 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11460) );
  AOI22_X1 U14637 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14638 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14639 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11455) );
  NAND4_X1 U14640 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(
        n11459) );
  OAI21_X1 U14641 ( .B1(n11460), .B2(n11459), .A(n11569), .ZN(n11463) );
  NAND2_X1 U14642 ( .A1(n11865), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U14643 ( .A1(n11864), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11461) );
  AND3_X1 U14644 ( .A1(n11463), .A2(n11462), .A3(n11461), .ZN(n11464) );
  NAND2_X1 U14645 ( .A1(n11465), .A2(n11464), .ZN(n13653) );
  AOI22_X1 U14646 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14647 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14648 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14649 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11467) );
  NAND4_X1 U14650 ( .A1(n11470), .A2(n11469), .A3(n11468), .A4(n11467), .ZN(
        n11476) );
  AOI22_X1 U14651 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14652 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14653 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11472) );
  NAND4_X1 U14654 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n11475) );
  OR2_X1 U14655 ( .A1(n11476), .A2(n11475), .ZN(n11477) );
  NAND2_X1 U14656 ( .A1(n13652), .A2(n14354), .ZN(n11484) );
  NAND2_X1 U14657 ( .A1(n11865), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11482) );
  OAI21_X1 U14658 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11480), .A(
        n11557), .ZN(n15908) );
  AOI22_X1 U14659 ( .A1(n11858), .A2(n15908), .B1(n11864), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11481) );
  NAND2_X1 U14660 ( .A1(n11482), .A2(n11481), .ZN(n13765) );
  AND2_X1 U14661 ( .A1(n13765), .A2(n13653), .ZN(n11483) );
  NAND2_X1 U14662 ( .A1(n13654), .A2(n11483), .ZN(n13764) );
  AOI22_X1 U14663 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14664 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14665 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14666 ( .A1(n13274), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11485) );
  NAND4_X1 U14667 ( .A1(n11488), .A2(n11487), .A3(n11486), .A4(n11485), .ZN(
        n11494) );
  AOI22_X1 U14668 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14669 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14670 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9971), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14671 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11489) );
  NAND4_X1 U14672 ( .A1(n11492), .A2(n11491), .A3(n11490), .A4(n11489), .ZN(
        n11493) );
  NOR2_X1 U14673 ( .A1(n11494), .A2(n11493), .ZN(n11497) );
  XNOR2_X1 U14674 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11593), .ZN(
        n15784) );
  OAI22_X1 U14675 ( .A1(n15784), .A2(n14113), .B1(n11867), .B2(n15786), .ZN(
        n11495) );
  AOI21_X1 U14676 ( .B1(n11408), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11495), .ZN(
        n11496) );
  OAI21_X1 U14677 ( .B1(n11861), .B2(n11497), .A(n11496), .ZN(n13712) );
  AOI22_X1 U14678 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14679 ( .A1(n11841), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14680 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11499) );
  NAND4_X1 U14681 ( .A1(n11501), .A2(n11500), .A3(n11499), .A4(n11498), .ZN(
        n11507) );
  AOI22_X1 U14682 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14683 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14684 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14685 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11502) );
  NAND4_X1 U14686 ( .A1(n11505), .A2(n11504), .A3(n11503), .A4(n11502), .ZN(
        n11506) );
  NOR2_X1 U14687 ( .A1(n11507), .A2(n11506), .ZN(n11511) );
  NAND2_X1 U14688 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14689 ( .A1(n14113), .A2(n11508), .ZN(n11509) );
  AOI21_X1 U14690 ( .B1(n11408), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11509), .ZN(
        n11510) );
  OAI21_X1 U14691 ( .B1(n11861), .B2(n11511), .A(n11510), .ZN(n11513) );
  OAI21_X1 U14692 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11514), .A(
        n11593), .ZN(n15883) );
  OR2_X1 U14693 ( .A1(n14113), .A2(n15883), .ZN(n11512) );
  NAND2_X1 U14694 ( .A1(n11513), .A2(n11512), .ZN(n14431) );
  INV_X1 U14695 ( .A(n14431), .ZN(n11577) );
  AOI21_X1 U14696 ( .B1(n11515), .B2(n20939), .A(n11514), .ZN(n15888) );
  OR2_X1 U14697 ( .A1(n15888), .A2(n14113), .ZN(n11530) );
  AOI22_X1 U14698 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14699 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14700 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11516) );
  NAND4_X1 U14701 ( .A1(n11519), .A2(n11518), .A3(n11517), .A4(n11516), .ZN(
        n11525) );
  AOI22_X1 U14702 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14703 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14704 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14705 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11520) );
  NAND4_X1 U14706 ( .A1(n11523), .A2(n11522), .A3(n11521), .A4(n11520), .ZN(
        n11524) );
  OAI21_X1 U14707 ( .B1(n11525), .B2(n11524), .A(n11569), .ZN(n11528) );
  NAND2_X1 U14708 ( .A1(n11865), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U14709 ( .A1(n11864), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11526) );
  AND3_X1 U14710 ( .A1(n11528), .A2(n11527), .A3(n11526), .ZN(n11529) );
  AND2_X1 U14711 ( .A1(n11530), .A2(n11529), .ZN(n14437) );
  INV_X1 U14712 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15813) );
  XNOR2_X1 U14713 ( .A(n15813), .B(n11531), .ZN(n15892) );
  INV_X1 U14714 ( .A(n15892), .ZN(n11546) );
  AOI22_X1 U14715 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14716 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14717 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14718 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11532) );
  NAND4_X1 U14719 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n11541) );
  AOI22_X1 U14720 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14721 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14722 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11537) );
  NAND4_X1 U14723 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n11540) );
  OAI21_X1 U14724 ( .B1(n11541), .B2(n11540), .A(n11569), .ZN(n11544) );
  NAND2_X1 U14725 ( .A1(n11865), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11543) );
  NAND2_X1 U14726 ( .A1(n11864), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11542) );
  NAND3_X1 U14727 ( .A1(n11544), .A2(n11543), .A3(n11542), .ZN(n11545) );
  AOI21_X1 U14728 ( .B1(n11546), .B2(n11858), .A(n11545), .ZN(n13801) );
  NOR2_X1 U14729 ( .A1(n14437), .A2(n13801), .ZN(n11576) );
  INV_X1 U14730 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U14731 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11847), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14732 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14733 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14734 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11547) );
  NAND4_X1 U14735 ( .A1(n11550), .A2(n11549), .A3(n11548), .A4(n11547), .ZN(
        n11556) );
  AOI22_X1 U14736 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11817), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14737 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14738 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11552) );
  NAND4_X1 U14739 ( .A1(n11554), .A2(n11553), .A3(n11552), .A4(n11551), .ZN(
        n11555) );
  OAI21_X1 U14740 ( .B1(n11556), .B2(n11555), .A(n11569), .ZN(n11560) );
  XNOR2_X1 U14741 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11557), .ZN(
        n15899) );
  OAI22_X1 U14742 ( .A1(n15899), .A2(n14113), .B1(n11867), .B2(n15820), .ZN(
        n11558) );
  INV_X1 U14743 ( .A(n11558), .ZN(n11559) );
  OAI211_X1 U14744 ( .C1(n11805), .C2(n14506), .A(n11560), .B(n11559), .ZN(
        n14451) );
  INV_X1 U14745 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14501) );
  AOI22_X1 U14746 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14747 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14748 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14749 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11561) );
  NAND4_X1 U14750 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11571) );
  AOI22_X1 U14751 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14752 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14753 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11566) );
  NAND4_X1 U14754 ( .A1(n11568), .A2(n11567), .A3(n11566), .A4(n11565), .ZN(
        n11570) );
  OAI21_X1 U14755 ( .B1(n11571), .B2(n11570), .A(n11569), .ZN(n11575) );
  XNOR2_X1 U14756 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11572), .ZN(
        n14648) );
  OAI22_X1 U14757 ( .A1(n14648), .A2(n14113), .B1(n11867), .B2(n14644), .ZN(
        n11573) );
  INV_X1 U14758 ( .A(n11573), .ZN(n11574) );
  OAI211_X1 U14759 ( .C1(n11805), .C2(n14501), .A(n11575), .B(n11574), .ZN(
        n14358) );
  AND2_X1 U14760 ( .A1(n14451), .A2(n14358), .ZN(n13799) );
  AOI22_X1 U14761 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14762 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14763 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9649), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14764 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11579) );
  NAND4_X1 U14765 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11588) );
  AOI22_X1 U14766 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14767 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14768 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11584) );
  NAND4_X1 U14769 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n11587) );
  NOR2_X1 U14770 ( .A1(n11588), .A2(n11587), .ZN(n11592) );
  NAND2_X1 U14771 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11589) );
  NAND2_X1 U14772 ( .A1(n14113), .A2(n11589), .ZN(n11590) );
  AOI21_X1 U14773 ( .B1(n11408), .B2(P1_EAX_REG_18__SCAN_IN), .A(n11590), .ZN(
        n11591) );
  OAI21_X1 U14774 ( .B1(n11861), .B2(n11592), .A(n11591), .ZN(n11599) );
  INV_X1 U14775 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11595) );
  INV_X1 U14776 ( .A(n11596), .ZN(n11594) );
  NAND2_X1 U14777 ( .A1(n11595), .A2(n11594), .ZN(n11597) );
  AND2_X1 U14778 ( .A1(n11597), .A2(n11631), .ZN(n15776) );
  NAND2_X1 U14779 ( .A1(n15776), .A2(n11858), .ZN(n11598) );
  NAND2_X1 U14780 ( .A1(n11599), .A2(n11598), .ZN(n14623) );
  AOI22_X1 U14781 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14782 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14783 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11601) );
  NAND4_X1 U14784 ( .A1(n11603), .A2(n11602), .A3(n11601), .A4(n11600), .ZN(
        n11609) );
  AOI22_X1 U14785 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14786 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U14787 ( .A1(n9649), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14788 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11604) );
  NAND4_X1 U14789 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n11608) );
  NOR2_X1 U14790 ( .A1(n11609), .A2(n11608), .ZN(n11613) );
  NAND2_X1 U14791 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11610) );
  NAND2_X1 U14792 ( .A1(n14113), .A2(n11610), .ZN(n11611) );
  AOI21_X1 U14793 ( .B1(n11408), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11611), .ZN(
        n11612) );
  OAI21_X1 U14794 ( .B1(n11861), .B2(n11613), .A(n11612), .ZN(n11615) );
  XNOR2_X1 U14795 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n11631), .ZN(
        n15763) );
  NAND2_X1 U14796 ( .A1(n15763), .A2(n11858), .ZN(n11614) );
  NAND2_X1 U14797 ( .A1(n11615), .A2(n11614), .ZN(n14422) );
  AOI22_X1 U14798 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14799 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11847), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14800 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13274), .B1(
        n9971), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14801 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U14802 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11626) );
  AOI22_X1 U14803 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11659), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14804 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11846), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14805 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14806 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11840), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11621) );
  NAND4_X1 U14807 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11625) );
  NOR2_X1 U14808 ( .A1(n11626), .A2(n11625), .ZN(n11630) );
  NAND2_X1 U14809 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U14810 ( .A1(n14113), .A2(n11627), .ZN(n11628) );
  AOI21_X1 U14811 ( .B1(n11408), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11628), .ZN(
        n11629) );
  OAI21_X1 U14812 ( .B1(n11861), .B2(n11630), .A(n11629), .ZN(n11635) );
  OAI21_X1 U14813 ( .B1(n11633), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n11651), .ZN(n14606) );
  OR2_X1 U14814 ( .A1(n14606), .A2(n14113), .ZN(n11634) );
  AOI22_X1 U14815 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14816 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14817 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14818 ( .A1(n9649), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11637) );
  NAND4_X1 U14819 ( .A1(n11640), .A2(n11639), .A3(n11638), .A4(n11637), .ZN(
        n11647) );
  AOI22_X1 U14820 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14821 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14822 ( .A1(n11641), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14823 ( .A1(n9971), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11752), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11642) );
  NAND4_X1 U14824 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11646) );
  NOR2_X1 U14825 ( .A1(n11647), .A2(n11646), .ZN(n11650) );
  AOI21_X1 U14826 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20839), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11648) );
  AOI21_X1 U14827 ( .B1(n11408), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11648), .ZN(
        n11649) );
  OAI21_X1 U14828 ( .B1(n11861), .B2(n11650), .A(n11649), .ZN(n11654) );
  AND2_X1 U14829 ( .A1(n11651), .A2(n20839), .ZN(n11652) );
  NOR2_X1 U14830 ( .A1(n11671), .A2(n11652), .ZN(n15752) );
  NAND2_X1 U14831 ( .A1(n15752), .A2(n11858), .ZN(n11653) );
  INV_X2 U14832 ( .A(n14586), .ZN(n11677) );
  AOI22_X1 U14833 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14834 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14835 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11656) );
  NAND4_X1 U14836 ( .A1(n11658), .A2(n11657), .A3(n11656), .A4(n11655), .ZN(
        n11666) );
  AOI22_X1 U14837 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14838 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14839 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14840 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11661) );
  NAND4_X1 U14841 ( .A1(n11664), .A2(n11663), .A3(n11662), .A4(n11661), .ZN(
        n11665) );
  NOR2_X1 U14842 ( .A1(n11666), .A2(n11665), .ZN(n11670) );
  OAI21_X1 U14843 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20757), .A(
        n20750), .ZN(n11667) );
  INV_X1 U14844 ( .A(n11667), .ZN(n11668) );
  AOI21_X1 U14845 ( .B1(n11865), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11668), .ZN(
        n11669) );
  OAI21_X1 U14846 ( .B1(n11861), .B2(n11670), .A(n11669), .ZN(n11675) );
  INV_X1 U14847 ( .A(n11671), .ZN(n11672) );
  INV_X1 U14848 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U14849 ( .A1(n11672), .A2(n14589), .ZN(n11673) );
  NAND2_X1 U14850 ( .A1(n11721), .A2(n11673), .ZN(n14588) );
  NAND2_X1 U14851 ( .A1(n11675), .A2(n11674), .ZN(n14587) );
  AOI22_X1 U14852 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14853 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14854 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14855 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11678) );
  NAND4_X1 U14856 ( .A1(n11681), .A2(n11680), .A3(n11679), .A4(n11678), .ZN(
        n11687) );
  AOI22_X1 U14857 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14858 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14859 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11683) );
  NAND4_X1 U14860 ( .A1(n11685), .A2(n11684), .A3(n11683), .A4(n11682), .ZN(
        n11686) );
  NOR2_X1 U14861 ( .A1(n11687), .A2(n11686), .ZN(n11705) );
  AOI22_X1 U14862 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14863 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14864 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14865 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(
        n11697) );
  AOI22_X1 U14866 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14867 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14868 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14869 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11692) );
  NAND4_X1 U14870 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11696) );
  NOR2_X1 U14871 ( .A1(n11697), .A2(n11696), .ZN(n11706) );
  XOR2_X1 U14872 ( .A(n11705), .B(n11706), .Z(n11698) );
  NAND2_X1 U14873 ( .A1(n11698), .A2(n11829), .ZN(n11702) );
  NAND2_X1 U14874 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11699) );
  NAND2_X1 U14875 ( .A1(n14113), .A2(n11699), .ZN(n11700) );
  AOI21_X1 U14876 ( .B1(n11408), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11700), .ZN(
        n11701) );
  NAND2_X1 U14877 ( .A1(n11702), .A2(n11701), .ZN(n11704) );
  XNOR2_X1 U14878 ( .A(n11721), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14573) );
  NAND2_X1 U14879 ( .A1(n14573), .A2(n11858), .ZN(n11703) );
  NAND2_X1 U14880 ( .A1(n11704), .A2(n11703), .ZN(n14330) );
  NOR2_X1 U14881 ( .A1(n11706), .A2(n11705), .ZN(n11728) );
  AOI22_X1 U14882 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14883 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14884 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14885 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11708) );
  NAND4_X1 U14886 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11717) );
  AOI22_X1 U14887 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14888 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14889 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11713) );
  INV_X1 U14890 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20910) );
  NAND4_X1 U14891 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11716) );
  OR2_X1 U14892 ( .A1(n11717), .A2(n11716), .ZN(n11727) );
  INV_X1 U14893 ( .A(n11727), .ZN(n11718) );
  XNOR2_X1 U14894 ( .A(n11728), .B(n11718), .ZN(n11719) );
  NAND2_X1 U14895 ( .A1(n11719), .A2(n11829), .ZN(n11726) );
  INV_X1 U14896 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14322) );
  AOI21_X1 U14897 ( .B1(n14322), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11720) );
  AOI21_X1 U14898 ( .B1(n11408), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11720), .ZN(
        n11725) );
  INV_X1 U14899 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14575) );
  NAND2_X1 U14900 ( .A1(n11722), .A2(n14322), .ZN(n11723) );
  NAND2_X1 U14901 ( .A1(n11764), .A2(n11723), .ZN(n14567) );
  NOR2_X1 U14902 ( .A1(n14567), .A2(n14113), .ZN(n11724) );
  AOI21_X1 U14903 ( .B1(n11726), .B2(n11725), .A(n11724), .ZN(n14317) );
  NAND2_X1 U14904 ( .A1(n11728), .A2(n11727), .ZN(n11745) );
  AOI22_X1 U14905 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14906 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14907 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14908 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U14909 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11738) );
  AOI22_X1 U14910 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14911 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14912 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14913 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n11737) );
  NOR2_X1 U14914 ( .A1(n11738), .A2(n11737), .ZN(n11746) );
  XOR2_X1 U14915 ( .A(n11745), .B(n11746), .Z(n11739) );
  NAND2_X1 U14916 ( .A1(n11739), .A2(n11829), .ZN(n11744) );
  NAND2_X1 U14917 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11740) );
  NAND2_X1 U14918 ( .A1(n14113), .A2(n11740), .ZN(n11741) );
  AOI21_X1 U14919 ( .B1(n11408), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11741), .ZN(
        n11743) );
  XNOR2_X1 U14920 ( .A(n11764), .B(n14309), .ZN(n14558) );
  NOR2_X1 U14921 ( .A1(n14558), .A2(n14113), .ZN(n11742) );
  AOI21_X1 U14922 ( .B1(n11744), .B2(n11743), .A(n11742), .ZN(n14304) );
  NOR2_X1 U14923 ( .A1(n11746), .A2(n11745), .ZN(n11773) );
  AOI22_X1 U14924 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11750) );
  AOI22_X1 U14925 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11749) );
  AOI22_X1 U14926 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U14927 ( .A1(n11660), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11747) );
  NAND4_X1 U14928 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11758) );
  AOI22_X1 U14929 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14930 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14931 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11754) );
  NAND4_X1 U14932 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n11757) );
  OR2_X1 U14933 ( .A1(n11758), .A2(n11757), .ZN(n11772) );
  INV_X1 U14934 ( .A(n11772), .ZN(n11759) );
  XNOR2_X1 U14935 ( .A(n11773), .B(n11759), .ZN(n11763) );
  INV_X1 U14936 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n11761) );
  NAND2_X1 U14937 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11760) );
  OAI211_X1 U14938 ( .C1(n11805), .C2(n11761), .A(n14113), .B(n11760), .ZN(
        n11762) );
  AOI21_X1 U14939 ( .B1(n11763), .B2(n11829), .A(n11762), .ZN(n11769) );
  INV_X1 U14940 ( .A(n11765), .ZN(n11766) );
  INV_X1 U14941 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14547) );
  NAND2_X1 U14942 ( .A1(n11766), .A2(n14547), .ZN(n11767) );
  NAND2_X1 U14943 ( .A1(n11808), .A2(n11767), .ZN(n14298) );
  NOR2_X1 U14944 ( .A1(n14298), .A2(n14113), .ZN(n11768) );
  NAND2_X1 U14945 ( .A1(n11773), .A2(n11772), .ZN(n11790) );
  AOI22_X1 U14946 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14947 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9648), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14948 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n13274), .B1(
        n9971), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14949 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11774) );
  NAND4_X1 U14950 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11783) );
  AOI22_X1 U14951 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11659), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14952 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11846), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14953 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14954 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11778) );
  NAND4_X1 U14955 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11782) );
  NOR2_X1 U14956 ( .A1(n11783), .A2(n11782), .ZN(n11791) );
  XOR2_X1 U14957 ( .A(n11790), .B(n11791), .Z(n11784) );
  NAND2_X1 U14958 ( .A1(n11784), .A2(n11829), .ZN(n11787) );
  INV_X1 U14959 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14537) );
  AOI21_X1 U14960 ( .B1(n14537), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11785) );
  AOI21_X1 U14961 ( .B1(n11865), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11785), .ZN(
        n11786) );
  NAND2_X1 U14962 ( .A1(n11787), .A2(n11786), .ZN(n11789) );
  XNOR2_X1 U14963 ( .A(n11808), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14539) );
  NAND2_X1 U14964 ( .A1(n14539), .A2(n11858), .ZN(n11788) );
  NAND2_X1 U14965 ( .A1(n11789), .A2(n11788), .ZN(n14285) );
  NOR2_X1 U14966 ( .A1(n11791), .A2(n11790), .ZN(n11816) );
  AOI22_X1 U14967 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11822), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U14968 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11848), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14969 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14970 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11792) );
  NAND4_X1 U14971 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11801) );
  AOI22_X1 U14972 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14973 ( .A1(n11838), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11849), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14974 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11797) );
  NAND4_X1 U14975 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11800) );
  OR2_X1 U14976 ( .A1(n11801), .A2(n11800), .ZN(n11815) );
  INV_X1 U14977 ( .A(n11815), .ZN(n11802) );
  XNOR2_X1 U14978 ( .A(n11816), .B(n11802), .ZN(n11807) );
  INV_X1 U14979 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U14980 ( .A1(n20750), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11803) );
  OAI211_X1 U14981 ( .C1(n11805), .C2(n11804), .A(n14113), .B(n11803), .ZN(
        n11806) );
  AOI21_X1 U14982 ( .B1(n11807), .B2(n11829), .A(n11806), .ZN(n11814) );
  INV_X1 U14983 ( .A(n11808), .ZN(n11809) );
  INV_X1 U14984 ( .A(n11810), .ZN(n11811) );
  INV_X1 U14985 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14527) );
  NAND2_X1 U14986 ( .A1(n11811), .A2(n14527), .ZN(n11812) );
  NAND2_X1 U14987 ( .A1(n11834), .A2(n11812), .ZN(n14276) );
  NOR2_X1 U14988 ( .A1(n14276), .A2(n14113), .ZN(n11813) );
  NAND2_X1 U14989 ( .A1(n11816), .A2(n11815), .ZN(n11836) );
  AOI22_X1 U14990 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14991 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11660), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14992 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14993 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11818) );
  NAND4_X1 U14994 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11828) );
  AOI22_X1 U14995 ( .A1(n11822), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14996 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14997 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11824) );
  NAND4_X1 U14998 ( .A1(n11826), .A2(n11825), .A3(n11824), .A4(n11823), .ZN(
        n11827) );
  NOR2_X1 U14999 ( .A1(n11828), .A2(n11827), .ZN(n11837) );
  XOR2_X1 U15000 ( .A(n11836), .B(n11837), .Z(n11830) );
  NAND2_X1 U15001 ( .A1(n11830), .A2(n11829), .ZN(n11833) );
  INV_X1 U15002 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14105) );
  NOR2_X1 U15003 ( .A1(n14105), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11831) );
  AOI211_X1 U15004 ( .C1(n11408), .C2(P1_EAX_REG_29__SCAN_IN), .A(n11858), .B(
        n11831), .ZN(n11832) );
  XNOR2_X1 U15005 ( .A(n11834), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14131) );
  AOI22_X1 U15006 ( .A1(n11833), .A2(n11832), .B1(n11858), .B2(n14131), .ZN(
        n14106) );
  INV_X1 U15007 ( .A(n11834), .ZN(n11835) );
  NAND2_X1 U15008 ( .A1(n11835), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11870) );
  XOR2_X1 U15009 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n11870), .Z(
        n14513) );
  NOR2_X1 U15010 ( .A1(n11837), .A2(n11836), .ZN(n11857) );
  AOI22_X1 U15011 ( .A1(n11839), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11838), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U15012 ( .A1(n11840), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13274), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U15013 ( .A1(n11841), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9649), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11843) );
  NAND4_X1 U15014 ( .A1(n11845), .A2(n11844), .A3(n11843), .A4(n11842), .ZN(
        n11855) );
  AOI22_X1 U15015 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11707), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U15016 ( .A1(n11817), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11847), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U15017 ( .A1(n11848), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15018 ( .A1(n11849), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11751), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11850) );
  NAND4_X1 U15019 ( .A1(n11853), .A2(n11852), .A3(n11851), .A4(n11850), .ZN(
        n11854) );
  NOR2_X1 U15020 ( .A1(n11855), .A2(n11854), .ZN(n11856) );
  XOR2_X1 U15021 ( .A(n11857), .B(n11856), .Z(n11862) );
  AOI21_X1 U15022 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20750), .A(
        n11858), .ZN(n11860) );
  NAND2_X1 U15023 ( .A1(n11865), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11859) );
  OAI211_X1 U15024 ( .C1(n11862), .C2(n11861), .A(n11860), .B(n11859), .ZN(
        n11863) );
  OAI21_X1 U15025 ( .B1(n14113), .B2(n14513), .A(n11863), .ZN(n14261) );
  AOI22_X1 U15026 ( .A1(n11865), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11864), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11866) );
  XNOR2_X1 U15027 ( .A(n14259), .B(n11866), .ZN(n14462) );
  NOR2_X1 U15028 ( .A1(n11867), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20725) );
  NOR2_X2 U15029 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20576) );
  NAND2_X1 U15030 ( .A1(n11872), .A2(n20573), .ZN(n20753) );
  AND2_X1 U15031 ( .A1(n20753), .A2(n20759), .ZN(n11868) );
  NAND2_X1 U15032 ( .A1(n20759), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15713) );
  NAND2_X1 U15033 ( .A1(n20757), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U15034 ( .A1(n15713), .A2(n11869), .ZN(n12945) );
  INV_X1 U15035 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14264) );
  INV_X1 U15036 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14247) );
  INV_X1 U15037 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20709) );
  OR2_X1 U15038 ( .A1(n15922), .A2(n20709), .ZN(n14202) );
  OAI21_X1 U15039 ( .B1(n15914), .B2(n14247), .A(n14202), .ZN(n11873) );
  AOI21_X1 U15040 ( .B1(n15909), .B2(n14129), .A(n11873), .ZN(n11874) );
  INV_X1 U15041 ( .A(n11874), .ZN(n11875) );
  OAI21_X1 U15042 ( .B1(n14208), .B2(n15902), .A(n11877), .ZN(P1_U2968) );
  NAND2_X1 U15043 ( .A1(n11889), .A2(n11879), .ZN(n11883) );
  XNOR2_X2 U15044 ( .A(n11883), .B(n11882), .ZN(n11911) );
  BUF_X2 U15045 ( .A(n11911), .Z(n11900) );
  AND2_X1 U15047 ( .A1(n11897), .A2(n18928), .ZN(n11903) );
  NAND2_X1 U15048 ( .A1(n11900), .A2(n11903), .ZN(n11888) );
  OR2_X2 U15049 ( .A1(n9653), .A2(n11888), .ZN(n11969) );
  INV_X2 U15050 ( .A(n11969), .ZN(n12007) );
  INV_X1 U15051 ( .A(n11890), .ZN(n11891) );
  NOR2_X2 U15052 ( .A1(n11892), .A2(n9653), .ZN(n19201) );
  AOI22_X1 U15053 ( .A1(n12007), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n19201), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11893) );
  INV_X1 U15054 ( .A(n11893), .ZN(n11908) );
  NAND2_X1 U15055 ( .A1(n11918), .A2(n11903), .ZN(n11894) );
  NOR2_X1 U15056 ( .A1(n9652), .A2(n11894), .ZN(n11936) );
  NOR2_X1 U15057 ( .A1(n9653), .A2(n11895), .ZN(n11896) );
  INV_X1 U15058 ( .A(n11968), .ZN(n12006) );
  NAND2_X1 U15059 ( .A1(n11898), .A2(n11897), .ZN(n11899) );
  INV_X1 U15060 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11901) );
  AND2_X1 U15061 ( .A1(n9652), .A2(n11902), .ZN(n11916) );
  INV_X2 U15062 ( .A(n11911), .ZN(n11918) );
  AND2_X1 U15063 ( .A1(n9652), .A2(n11903), .ZN(n11917) );
  NAND3_X1 U15064 ( .A1(n11906), .A2(n11905), .A3(n11904), .ZN(n11907) );
  NOR2_X1 U15065 ( .A1(n11908), .A2(n11907), .ZN(n11928) );
  INV_X1 U15066 ( .A(n11913), .ZN(n11910) );
  INV_X1 U15067 ( .A(n11943), .ZN(n12001) );
  INV_X1 U15068 ( .A(n11914), .ZN(n11912) );
  AOI22_X1 U15069 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n12001), .B1(
        n11959), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11924) );
  NOR2_X2 U15070 ( .A1(n11915), .A2(n11914), .ZN(n11958) );
  AOI22_X1 U15071 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n13511), .B1(
        n19464), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11922) );
  AND2_X1 U15072 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11918), .ZN(
        n11920) );
  NAND2_X1 U15073 ( .A1(n11919), .A2(n13427), .ZN(n11925) );
  NAND2_X1 U15074 ( .A1(n11920), .A2(n11950), .ZN(n11921) );
  AOI22_X1 U15075 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11965), .B1(
        n19433), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15076 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19201), .B1(
        n12007), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11935) );
  NAND2_X1 U15077 ( .A1(n13511), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U15078 ( .A1(n13447), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U15079 ( .A1(n11931), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11932) );
  NAND4_X1 U15080 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11941) );
  INV_X1 U15081 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11939) );
  AOI21_X1 U15082 ( .B1(n12006), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n19737), .ZN(n11938) );
  NAND2_X1 U15083 ( .A1(n11936), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11937) );
  OAI211_X1 U15084 ( .C1(n19270), .C2(n11939), .A(n11938), .B(n11937), .ZN(
        n11940) );
  NOR2_X1 U15085 ( .A1(n11941), .A2(n11940), .ZN(n11955) );
  INV_X1 U15086 ( .A(n11942), .ZN(n11948) );
  INV_X1 U15087 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11946) );
  INV_X1 U15088 ( .A(n19464), .ZN(n11945) );
  INV_X1 U15089 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11944) );
  OAI22_X1 U15090 ( .A1(n11946), .A2(n11943), .B1(n11945), .B2(n11944), .ZN(
        n11947) );
  NOR2_X1 U15091 ( .A1(n11948), .A2(n11947), .ZN(n11954) );
  INV_X1 U15092 ( .A(n11949), .ZN(n11973) );
  AOI22_X1 U15093 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11973), .B1(
        n11960), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11952) );
  AND2_X1 U15094 ( .A1(n11952), .A2(n11951), .ZN(n11953) );
  NOR2_X1 U15095 ( .A1(n12676), .A2(n11983), .ZN(n11956) );
  NAND2_X1 U15096 ( .A1(n19737), .A2(n11956), .ZN(n11987) );
  NAND2_X1 U15097 ( .A1(n11987), .A2(n11986), .ZN(n11957) );
  AOI22_X1 U15098 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n12001), .B1(
        n11959), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15099 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n13447), .B1(
        n19464), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11962) );
  NAND2_X1 U15100 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11961) );
  INV_X1 U15101 ( .A(n11965), .ZN(n19081) );
  INV_X1 U15102 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19106) );
  OR2_X1 U15103 ( .A1(n19081), .A2(n19106), .ZN(n11977) );
  AOI22_X1 U15104 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19201), .B1(
        n11936), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15105 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n13511), .B1(
        n11931), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11966) );
  INV_X1 U15106 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11971) );
  INV_X1 U15107 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11970) );
  OAI22_X1 U15108 ( .A1(n11971), .A2(n11968), .B1(n11969), .B2(n11970), .ZN(
        n11972) );
  INV_X1 U15109 ( .A(n11972), .ZN(n11975) );
  AOI22_X1 U15110 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n11973), .B1(
        n19433), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11974) );
  AND3_X1 U15111 ( .A1(n9711), .A2(n11975), .A3(n11974), .ZN(n11976) );
  NAND3_X1 U15112 ( .A1(n9693), .A2(n11977), .A3(n11976), .ZN(n11980) );
  NAND2_X1 U15113 ( .A1(n11978), .A2(n19737), .ZN(n11979) );
  INV_X1 U15114 ( .A(n12064), .ZN(n11981) );
  INV_X1 U15115 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13691) );
  NAND2_X1 U15116 ( .A1(n12676), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12675) );
  NOR2_X1 U15117 ( .A1(n11983), .A2(n12675), .ZN(n11985) );
  INV_X1 U15118 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16202) );
  AND2_X1 U15119 ( .A1(n12676), .A2(n16202), .ZN(n11984) );
  XNOR2_X1 U15120 ( .A(n11984), .B(n11983), .ZN(n12686) );
  NOR2_X1 U15121 ( .A1(n13527), .A2(n12686), .ZN(n12685) );
  NOR2_X1 U15122 ( .A1(n11985), .A2(n12685), .ZN(n11989) );
  XOR2_X1 U15123 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11989), .Z(
        n12754) );
  INV_X1 U15124 ( .A(n12754), .ZN(n11988) );
  XNOR2_X1 U15125 ( .A(n11987), .B(n11986), .ZN(n12752) );
  NAND2_X1 U15126 ( .A1(n11988), .A2(n12752), .ZN(n12756) );
  INV_X1 U15127 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12290) );
  OR2_X1 U15128 ( .A1(n11989), .A2(n12290), .ZN(n11990) );
  NAND2_X1 U15129 ( .A1(n12756), .A2(n11990), .ZN(n11992) );
  INV_X1 U15130 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11991) );
  XNOR2_X1 U15131 ( .A(n11992), .B(n11991), .ZN(n13497) );
  NAND2_X1 U15132 ( .A1(n11992), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11993) );
  NAND2_X1 U15133 ( .A1(n13477), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11998) );
  NAND2_X1 U15134 ( .A1(n11996), .A2(n11995), .ZN(n11997) );
  NAND2_X1 U15135 ( .A1(n11994), .A2(n11997), .ZN(n13475) );
  INV_X1 U15136 ( .A(n13477), .ZN(n11999) );
  INV_X1 U15137 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13690) );
  NAND2_X1 U15138 ( .A1(n12064), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12019) );
  AOI22_X1 U15139 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12001), .B1(
        n11959), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15140 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19464), .B1(
        n13511), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12003) );
  NAND2_X1 U15141 ( .A1(n11960), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12002) );
  AOI22_X1 U15142 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11965), .B1(
        n19433), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15143 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n13447), .B1(
        n11931), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15144 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11936), .B1(
        n12006), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12011) );
  AOI22_X1 U15145 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19201), .B1(
        n12007), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12010) );
  INV_X1 U15146 ( .A(n11973), .ZN(n19235) );
  INV_X1 U15147 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12008) );
  OR2_X1 U15148 ( .A1(n19235), .A2(n12008), .ZN(n12009) );
  NAND3_X1 U15149 ( .A1(n9694), .A2(n12014), .A3(n12013), .ZN(n12017) );
  NAND2_X1 U15150 ( .A1(n12015), .A2(n19737), .ZN(n12016) );
  INV_X1 U15151 ( .A(n12087), .ZN(n12018) );
  NAND2_X1 U15152 ( .A1(n12021), .A2(n12087), .ZN(n12022) );
  XNOR2_X1 U15153 ( .A(n12031), .B(n12025), .ZN(n12026) );
  INV_X1 U15154 ( .A(n12026), .ZN(n12027) );
  NOR2_X1 U15155 ( .A1(n12031), .A2(n12025), .ZN(n12030) );
  INV_X1 U15156 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12103) );
  XNOR2_X1 U15157 ( .A(n12030), .B(n12103), .ZN(n16126) );
  INV_X1 U15158 ( .A(n12031), .ZN(n12032) );
  NAND3_X1 U15159 ( .A1(n12032), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n15043), .ZN(n12033) );
  AND2_X1 U15160 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16170) );
  AND2_X1 U15161 ( .A1(n16170), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15329) );
  NAND3_X1 U15162 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15327) );
  INV_X1 U15163 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U15164 ( .A1(n15327), .A2(n15335), .ZN(n12034) );
  AND2_X1 U15165 ( .A1(n15329), .A2(n12034), .ZN(n12036) );
  AND2_X1 U15166 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15372) );
  NAND2_X1 U15167 ( .A1(n15372), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15357) );
  NAND2_X1 U15168 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12035) );
  NOR2_X1 U15169 ( .A1(n15357), .A2(n12035), .ZN(n15324) );
  AND2_X1 U15170 ( .A1(n12036), .A2(n15324), .ZN(n15310) );
  INV_X1 U15171 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15306) );
  NAND2_X1 U15172 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15238) );
  NOR2_X4 U15173 ( .A1(n15083), .A2(n15238), .ZN(n15068) );
  XNOR2_X1 U15174 ( .A(n12037), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12311) );
  OAI21_X1 U15175 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19714), .A(
        n12038), .ZN(n12231) );
  MUX2_X1 U15176 ( .A(n12231), .B(n12676), .S(n12229), .Z(n12067) );
  INV_X1 U15177 ( .A(n12039), .ZN(n12041) );
  OAI21_X1 U15178 ( .B1(n12067), .B2(n12041), .A(n12040), .ZN(n12045) );
  NAND2_X1 U15179 ( .A1(n12043), .A2(n12042), .ZN(n12227) );
  INV_X1 U15180 ( .A(n12227), .ZN(n12044) );
  NAND2_X1 U15181 ( .A1(n12045), .A2(n12044), .ZN(n12046) );
  NAND2_X1 U15182 ( .A1(n12046), .A2(n12248), .ZN(n19721) );
  INV_X1 U15183 ( .A(n12313), .ZN(n13253) );
  INV_X1 U15184 ( .A(n12047), .ZN(n12217) );
  NAND2_X1 U15185 ( .A1(n13253), .A2(n12217), .ZN(n12260) );
  OAI21_X1 U15186 ( .B1(n12231), .B2(n12048), .A(n13241), .ZN(n12049) );
  INV_X1 U15187 ( .A(n12049), .ZN(n12053) );
  NAND2_X1 U15188 ( .A1(n12050), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12051) );
  NAND2_X1 U15189 ( .A1(n12051), .A2(n12703), .ZN(n12698) );
  INV_X1 U15190 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18758) );
  AND2_X1 U15191 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18758), .ZN(n12052) );
  OAI21_X1 U15192 ( .B1(n10692), .B2(n12698), .A(n12052), .ZN(n19710) );
  OAI21_X1 U15193 ( .B1(n12053), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n19710), 
        .ZN(n19718) );
  NAND2_X1 U15194 ( .A1(n13253), .A2(n10635), .ZN(n12054) );
  AND2_X1 U15195 ( .A1(n13399), .A2(n16213), .ZN(n12055) );
  NAND2_X1 U15196 ( .A1(n13528), .A2(n19731), .ZN(n19680) );
  OR2_X1 U15197 ( .A1(n19682), .A2(n13574), .ZN(n19706) );
  NAND2_X1 U15198 ( .A1(n19706), .A2(n13371), .ZN(n12056) );
  NOR2_X1 U15199 ( .A1(n13528), .A2(n19736), .ZN(n12057) );
  NOR2_X1 U15200 ( .A1(n18885), .A2(n19671), .ZN(n12298) );
  INV_X1 U15201 ( .A(n12337), .ZN(n12059) );
  NAND2_X1 U15202 ( .A1(n19736), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12058) );
  NAND2_X1 U15203 ( .A1(n12059), .A2(n12058), .ZN(n12679) );
  NOR2_X1 U15204 ( .A1(n19052), .A2(n12060), .ZN(n12061) );
  AOI211_X1 U15205 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n19039), .A(
        n12298), .B(n12061), .ZN(n12062) );
  OAI21_X1 U15206 ( .B1(n14889), .B2(n19047), .A(n12062), .ZN(n12063) );
  AOI21_X1 U15207 ( .B1(n12311), .B2(n19042), .A(n12063), .ZN(n12209) );
  NAND2_X1 U15208 ( .A1(n12064), .A2(n12025), .ZN(n12085) );
  XNOR2_X1 U15209 ( .A(n12083), .B(n10100), .ZN(n18902) );
  INV_X1 U15210 ( .A(n18902), .ZN(n12066) );
  NAND2_X1 U15211 ( .A1(n10242), .A2(n12025), .ZN(n13490) );
  MUX2_X1 U15212 ( .A(n12067), .B(n18920), .S(n13389), .Z(n18924) );
  NOR2_X1 U15213 ( .A1(n18924), .A2(n16202), .ZN(n12683) );
  NOR3_X1 U15214 ( .A1(n12270), .A2(n13421), .A3(n18920), .ZN(n12068) );
  NOR2_X1 U15215 ( .A1(n12071), .A2(n12068), .ZN(n13425) );
  NAND2_X1 U15216 ( .A1(n12683), .A2(n13425), .ZN(n12069) );
  NOR2_X1 U15217 ( .A1(n12683), .A2(n13425), .ZN(n12682) );
  AOI21_X1 U15218 ( .B1(n13527), .B2(n12069), .A(n12682), .ZN(n12751) );
  XNOR2_X1 U15219 ( .A(n12071), .B(n12070), .ZN(n13438) );
  XNOR2_X1 U15220 ( .A(n13438), .B(n12290), .ZN(n12749) );
  NAND2_X1 U15221 ( .A1(n12751), .A2(n12749), .ZN(n12073) );
  NAND2_X1 U15222 ( .A1(n13438), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12072) );
  NAND2_X1 U15223 ( .A1(n12073), .A2(n12072), .ZN(n13491) );
  AND2_X1 U15224 ( .A1(n12075), .A2(n12074), .ZN(n12077) );
  OR2_X1 U15225 ( .A1(n12077), .A2(n12076), .ZN(n13489) );
  INV_X1 U15226 ( .A(n13489), .ZN(n12078) );
  AOI21_X1 U15227 ( .B1(n13491), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12078), .ZN(n12080) );
  NOR2_X1 U15228 ( .A1(n13491), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12079) );
  OR2_X1 U15229 ( .A1(n12076), .A2(n12081), .ZN(n12082) );
  NAND2_X1 U15230 ( .A1(n12083), .A2(n12082), .ZN(n13328) );
  NOR2_X1 U15231 ( .A1(n18902), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12084) );
  NAND2_X1 U15232 ( .A1(n12085), .A2(n12084), .ZN(n12086) );
  INV_X1 U15233 ( .A(n13723), .ZN(n12092) );
  AND2_X1 U15234 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  OR2_X1 U15235 ( .A1(n12090), .A2(n12100), .ZN(n18886) );
  NAND2_X1 U15236 ( .A1(n12093), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13823) );
  OR2_X1 U15237 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  NAND2_X1 U15238 ( .A1(n12094), .A2(n12097), .ZN(n13118) );
  NOR2_X1 U15239 ( .A1(n13118), .A2(n12025), .ZN(n12102) );
  NAND2_X1 U15240 ( .A1(n12102), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16119) );
  INV_X1 U15241 ( .A(n12098), .ZN(n12099) );
  XNOR2_X1 U15242 ( .A(n12100), .B(n12099), .ZN(n18875) );
  NAND2_X1 U15243 ( .A1(n18875), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16120) );
  AND2_X1 U15244 ( .A1(n16119), .A2(n16120), .ZN(n15442) );
  AND2_X1 U15245 ( .A1(n13823), .A2(n15442), .ZN(n12101) );
  INV_X1 U15246 ( .A(n12102), .ZN(n12104) );
  NAND2_X1 U15247 ( .A1(n12104), .A2(n12103), .ZN(n16118) );
  OR2_X1 U15248 ( .A1(n18875), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16122) );
  AND2_X1 U15249 ( .A1(n16118), .A2(n16122), .ZN(n15443) );
  NAND2_X1 U15250 ( .A1(n13389), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12105) );
  XNOR2_X1 U15251 ( .A(n12094), .B(n12105), .ZN(n18864) );
  NAND2_X1 U15252 ( .A1(n18864), .A2(n15043), .ZN(n12116) );
  INV_X1 U15253 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15455) );
  NAND2_X1 U15254 ( .A1(n12116), .A2(n15455), .ZN(n15445) );
  AND2_X1 U15255 ( .A1(n15443), .A2(n15445), .ZN(n12106) );
  NAND3_X1 U15256 ( .A1(n12108), .A2(n13389), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n12107) );
  OAI211_X1 U15257 ( .C1(n12108), .C2(P2_EBX_REG_10__SCAN_IN), .A(n12186), .B(
        n12107), .ZN(n18851) );
  OR2_X1 U15258 ( .A1(n18851), .A2(n12025), .ZN(n12110) );
  AND3_X1 U15259 ( .A1(n13389), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n9714), .ZN(
        n12112) );
  NOR2_X1 U15260 ( .A1(n12113), .A2(n12112), .ZN(n18842) );
  NAND2_X1 U15261 ( .A1(n18842), .A2(n15043), .ZN(n12114) );
  INV_X1 U15262 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15434) );
  AND2_X1 U15263 ( .A1(n12114), .A2(n15434), .ZN(n15427) );
  NOR2_X1 U15264 ( .A1(n12114), .A2(n15434), .ZN(n15428) );
  NAND2_X1 U15265 ( .A1(n15043), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12115) );
  OR2_X1 U15266 ( .A1(n18851), .A2(n12115), .ZN(n16102) );
  NAND2_X1 U15267 ( .A1(n16102), .A2(n16101), .ZN(n15424) );
  NOR2_X1 U15268 ( .A1(n15428), .A2(n15424), .ZN(n12117) );
  NAND3_X1 U15269 ( .A1(n13389), .A2(P2_EBX_REG_12__SCAN_IN), .A3(n12118), 
        .ZN(n12119) );
  NAND2_X1 U15270 ( .A1(n12141), .A2(n12119), .ZN(n13465) );
  NOR2_X1 U15271 ( .A1(n12120), .A2(n15418), .ZN(n15409) );
  NAND2_X1 U15272 ( .A1(n12120), .A2(n15418), .ZN(n15408) );
  INV_X1 U15273 ( .A(n12122), .ZN(n12124) );
  NAND3_X1 U15274 ( .A1(n12155), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n13389), 
        .ZN(n12123) );
  OR2_X1 U15275 ( .A1(n18786), .A2(n12025), .ZN(n12125) );
  NAND2_X1 U15276 ( .A1(n12125), .A2(n15306), .ZN(n15106) );
  INV_X1 U15277 ( .A(n12126), .ZN(n12127) );
  XNOR2_X1 U15278 ( .A(n12128), .B(n12127), .ZN(n18821) );
  AOI21_X1 U15279 ( .B1(n18821), .B2(n15043), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15109) );
  OR3_X1 U15280 ( .A1(n12135), .A2(n13663), .A3(n12270), .ZN(n12129) );
  NAND3_X1 U15281 ( .A1(n12130), .A2(n12129), .A3(n12186), .ZN(n18827) );
  INV_X1 U15282 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15393) );
  OAI21_X1 U15283 ( .B1(n18827), .B2(n12025), .A(n15393), .ZN(n12132) );
  NAND2_X1 U15284 ( .A1(n15043), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U15285 ( .A1(n12170), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12133) );
  MUX2_X1 U15286 ( .A(n12170), .B(n12133), .S(n12143), .Z(n12134) );
  OR2_X1 U15287 ( .A1(n12143), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12136) );
  NAND2_X1 U15288 ( .A1(n12134), .A2(n12136), .ZN(n13621) );
  INV_X1 U15289 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16168) );
  NAND2_X1 U15290 ( .A1(n12160), .A2(n16168), .ZN(n15107) );
  INV_X1 U15291 ( .A(n12135), .ZN(n12138) );
  NAND3_X1 U15292 ( .A1(n12136), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n12170), 
        .ZN(n12137) );
  NAND2_X1 U15293 ( .A1(n12138), .A2(n12137), .ZN(n12646) );
  OR2_X1 U15294 ( .A1(n12646), .A2(n12025), .ZN(n12139) );
  INV_X1 U15295 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15370) );
  NAND2_X1 U15296 ( .A1(n12139), .A2(n15370), .ZN(n15176) );
  NAND2_X1 U15297 ( .A1(n12141), .A2(n12140), .ZN(n12142) );
  NAND2_X1 U15298 ( .A1(n12143), .A2(n12142), .ZN(n12658) );
  NAND2_X1 U15299 ( .A1(n12163), .A2(n15395), .ZN(n15191) );
  NAND4_X1 U15300 ( .A1(n15108), .A2(n15107), .A3(n15176), .A4(n15191), .ZN(
        n12144) );
  NOR2_X1 U15301 ( .A1(n15109), .A2(n12144), .ZN(n12157) );
  NAND2_X1 U15302 ( .A1(n13389), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12145) );
  MUX2_X1 U15303 ( .A(n12170), .B(n12145), .S(n12146), .Z(n12147) );
  OR2_X1 U15304 ( .A1(n12146), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12150) );
  NAND2_X1 U15305 ( .A1(n12147), .A2(n12150), .ZN(n13853) );
  OR2_X1 U15306 ( .A1(n13853), .A2(n12025), .ZN(n12148) );
  INV_X1 U15307 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15358) );
  NAND2_X1 U15308 ( .A1(n12148), .A2(n15358), .ZN(n15145) );
  AND2_X1 U15309 ( .A1(n12170), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12149) );
  NAND2_X1 U15310 ( .A1(n12150), .A2(n12149), .ZN(n12151) );
  NAND2_X1 U15311 ( .A1(n12151), .A2(n12153), .ZN(n18803) );
  OR2_X1 U15312 ( .A1(n18803), .A2(n12025), .ZN(n12152) );
  INV_X1 U15313 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15349) );
  NAND2_X1 U15314 ( .A1(n12152), .A2(n15349), .ZN(n15136) );
  AND2_X1 U15315 ( .A1(n15145), .A2(n15136), .ZN(n15111) );
  NAND2_X1 U15316 ( .A1(n13389), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12154) );
  MUX2_X1 U15317 ( .A(n13389), .B(n12154), .S(n12153), .Z(n12156) );
  NAND2_X1 U15318 ( .A1(n12156), .A2(n12155), .ZN(n18798) );
  NAND2_X1 U15319 ( .A1(n12159), .A2(n15335), .ZN(n15120) );
  NAND4_X1 U15320 ( .A1(n15106), .A2(n12157), .A3(n15111), .A4(n15120), .ZN(
        n12169) );
  NAND2_X1 U15321 ( .A1(n15043), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12158) );
  INV_X1 U15322 ( .A(n12160), .ZN(n12161) );
  NAND2_X1 U15323 ( .A1(n12161), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15173) );
  NAND2_X1 U15324 ( .A1(n15043), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12162) );
  OR2_X1 U15325 ( .A1(n12646), .A2(n12162), .ZN(n15175) );
  INV_X1 U15326 ( .A(n12163), .ZN(n12164) );
  NAND2_X1 U15327 ( .A1(n12164), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15189) );
  NAND4_X1 U15328 ( .A1(n15135), .A2(n15173), .A3(n15175), .A4(n15189), .ZN(
        n12166) );
  AND2_X1 U15329 ( .A1(n15043), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12165) );
  NAND2_X1 U15330 ( .A1(n18821), .A2(n12165), .ZN(n15154) );
  NAND2_X1 U15331 ( .A1(n15154), .A2(n15156), .ZN(n15110) );
  NOR2_X1 U15332 ( .A1(n12166), .A2(n15110), .ZN(n12167) );
  AND4_X1 U15333 ( .A1(n15105), .A2(n15121), .A3(n12167), .A4(n15144), .ZN(
        n12168) );
  NAND3_X1 U15334 ( .A1(n12171), .A2(n12170), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n12172) );
  AND2_X1 U15335 ( .A1(n12176), .A2(n12172), .ZN(n15677) );
  NAND2_X1 U15336 ( .A1(n15677), .A2(n15043), .ZN(n12173) );
  INV_X1 U15337 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15296) );
  NAND2_X1 U15338 ( .A1(n12173), .A2(n15296), .ZN(n15291) );
  OR2_X1 U15339 ( .A1(n12173), .A2(n15296), .ZN(n15292) );
  INV_X1 U15340 ( .A(n12174), .ZN(n12175) );
  XNOR2_X1 U15341 ( .A(n12176), .B(n12175), .ZN(n14878) );
  NAND2_X1 U15342 ( .A1(n14878), .A2(n15043), .ZN(n12177) );
  XNOR2_X1 U15343 ( .A(n12177), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15097) );
  INV_X1 U15344 ( .A(n12186), .ZN(n12181) );
  NAND2_X1 U15345 ( .A1(n13389), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12178) );
  NOR2_X1 U15346 ( .A1(n12179), .A2(n12178), .ZN(n12180) );
  OR3_X1 U15347 ( .A1(n12188), .A2(n12181), .A3(n12180), .ZN(n16043) );
  NOR2_X1 U15348 ( .A1(n16043), .A2(n12025), .ZN(n12182) );
  AND2_X1 U15349 ( .A1(n12182), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15086) );
  INV_X1 U15350 ( .A(n12182), .ZN(n12183) );
  NOR2_X1 U15351 ( .A1(n12188), .A2(n14923), .ZN(n12184) );
  NAND2_X1 U15352 ( .A1(n13389), .A2(n12184), .ZN(n12185) );
  NAND2_X1 U15353 ( .A1(n12186), .A2(n12185), .ZN(n12187) );
  AOI21_X1 U15354 ( .B1(n12188), .B2(n14923), .A(n12187), .ZN(n14873) );
  AOI21_X1 U15355 ( .B1(n14873), .B2(n15043), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15075) );
  AND3_X1 U15356 ( .A1(n13389), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n12189), .ZN(
        n12190) );
  NOR2_X1 U15357 ( .A1(n12191), .A2(n12190), .ZN(n16027) );
  NAND2_X1 U15358 ( .A1(n16027), .A2(n15043), .ZN(n12196) );
  XNOR2_X1 U15359 ( .A(n12196), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15067) );
  NAND2_X1 U15360 ( .A1(n16012), .A2(n12192), .ZN(n12193) );
  NAND2_X1 U15361 ( .A1(n12200), .A2(n12193), .ZN(n14852) );
  OAI21_X1 U15362 ( .B1(n15042), .B2(n15227), .A(n15047), .ZN(n12199) );
  INV_X1 U15363 ( .A(n14873), .ZN(n12195) );
  INV_X1 U15364 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15252) );
  INV_X1 U15365 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15241) );
  OR2_X1 U15366 ( .A1(n12196), .A2(n15241), .ZN(n12197) );
  XOR2_X1 U15367 ( .A(n12201), .B(n12200), .Z(n14839) );
  AOI21_X1 U15368 ( .B1(n14839), .B2(n15043), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14209) );
  AND2_X1 U15369 ( .A1(n13389), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12202) );
  XNOR2_X1 U15370 ( .A(n12203), .B(n12202), .ZN(n16003) );
  INV_X1 U15371 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15024) );
  OAI21_X1 U15372 ( .B1(n16003), .B2(n12025), .A(n15024), .ZN(n15020) );
  NAND2_X1 U15373 ( .A1(n15043), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12204) );
  NOR2_X1 U15374 ( .A1(n16003), .A2(n12204), .ZN(n15019) );
  INV_X1 U15375 ( .A(n14839), .ZN(n12205) );
  NOR3_X1 U15376 ( .A1(n12205), .A2(n12025), .A3(n15200), .ZN(n15018) );
  NAND2_X1 U15377 ( .A1(n12206), .A2(n15043), .ZN(n12207) );
  NAND2_X1 U15378 ( .A1(n12315), .A2(n19040), .ZN(n12208) );
  NAND2_X1 U15379 ( .A1(n12209), .A2(n12208), .ZN(P2_U2983) );
  NAND3_X1 U15380 ( .A1(n12222), .A2(n13241), .A3(n13249), .ZN(n12214) );
  NAND2_X1 U15381 ( .A1(n12210), .A2(n13383), .ZN(n12211) );
  NAND2_X1 U15382 ( .A1(n12211), .A2(n9647), .ZN(n12213) );
  NAND3_X1 U15383 ( .A1(n12214), .A2(n12213), .A3(n12212), .ZN(n12221) );
  OAI21_X1 U15384 ( .B1(n10375), .B2(n10635), .A(n12280), .ZN(n12215) );
  NAND2_X1 U15385 ( .A1(n12215), .A2(n12617), .ZN(n12216) );
  AOI21_X1 U15386 ( .B1(n13383), .B2(n12216), .A(n10431), .ZN(n12219) );
  NAND2_X1 U15387 ( .A1(n12218), .A2(n12217), .ZN(n12279) );
  NAND2_X1 U15388 ( .A1(n12219), .A2(n12279), .ZN(n12220) );
  NOR2_X1 U15389 ( .A1(n12221), .A2(n12220), .ZN(n12694) );
  MUX2_X1 U15390 ( .A(n12222), .B(n12252), .S(n19737), .Z(n12223) );
  NAND3_X1 U15391 ( .A1(n12223), .A2(n13241), .A3(n19600), .ZN(n12224) );
  NAND2_X1 U15392 ( .A1(n12694), .A2(n12224), .ZN(n12225) );
  NOR2_X1 U15393 ( .A1(n12226), .A2(n12225), .ZN(n12258) );
  NAND2_X1 U15394 ( .A1(n12227), .A2(n12312), .ZN(n12245) );
  AOI21_X1 U15395 ( .B1(n12249), .B2(n10635), .A(n12228), .ZN(n12239) );
  INV_X1 U15396 ( .A(n12228), .ZN(n12236) );
  OAI21_X1 U15397 ( .B1(n12231), .B2(n12230), .A(n12229), .ZN(n12235) );
  INV_X1 U15398 ( .A(n12231), .ZN(n12233) );
  OAI211_X1 U15399 ( .C1(n10635), .C2(n12233), .A(n12280), .B(n12232), .ZN(
        n12234) );
  OAI211_X1 U15400 ( .C1(n12236), .C2(n12700), .A(n12235), .B(n12234), .ZN(
        n12237) );
  OAI21_X1 U15401 ( .B1(n12239), .B2(n12238), .A(n12237), .ZN(n12241) );
  NAND2_X1 U15402 ( .A1(n12241), .A2(n12240), .ZN(n12244) );
  OAI21_X1 U15403 ( .B1(n12312), .B2(n12242), .A(n12248), .ZN(n12243) );
  AOI21_X1 U15404 ( .B1(n12245), .B2(n12244), .A(n12243), .ZN(n12246) );
  MUX2_X1 U15405 ( .A(n12703), .B(n12246), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12247) );
  INV_X1 U15406 ( .A(n12248), .ZN(n12250) );
  INV_X1 U15407 ( .A(n12249), .ZN(n12793) );
  NAND3_X1 U15408 ( .A1(n12790), .A2(n13249), .A3(n12252), .ZN(n12257) );
  INV_X1 U15409 ( .A(n12790), .ZN(n12255) );
  AOI21_X1 U15410 ( .B1(n12253), .B2(n12280), .A(n10375), .ZN(n12254) );
  NAND2_X1 U15411 ( .A1(n12255), .A2(n12254), .ZN(n12256) );
  NAND3_X1 U15412 ( .A1(n12258), .A2(n12257), .A3(n12256), .ZN(n12259) );
  INV_X1 U15413 ( .A(n12260), .ZN(n19720) );
  INV_X1 U15414 ( .A(n13066), .ZN(n12263) );
  NAND2_X1 U15415 ( .A1(n12261), .A2(n19737), .ZN(n12262) );
  NAND2_X1 U15416 ( .A1(n12263), .A2(n12262), .ZN(n12264) );
  INV_X1 U15417 ( .A(n12265), .ZN(n12267) );
  AND2_X1 U15418 ( .A1(n12267), .A2(n12266), .ZN(n13244) );
  INV_X1 U15419 ( .A(n13244), .ZN(n13074) );
  NAND2_X1 U15420 ( .A1(n13243), .A2(n10635), .ZN(n12268) );
  NAND2_X1 U15421 ( .A1(n13074), .A2(n12268), .ZN(n12269) );
  AND2_X1 U15422 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15273) );
  NAND2_X1 U15423 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15310), .ZN(
        n15281) );
  NAND3_X1 U15424 ( .A1(n12270), .A2(n13383), .A3(n19737), .ZN(n12271) );
  NOR2_X1 U15425 ( .A1(n12265), .A2(n12271), .ZN(n13073) );
  NAND2_X1 U15426 ( .A1(n12314), .A2(n13073), .ZN(n19075) );
  NAND2_X1 U15427 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19063) );
  NAND2_X1 U15428 ( .A1(n12290), .A2(n19063), .ZN(n13480) );
  INV_X1 U15429 ( .A(n13480), .ZN(n12272) );
  OR2_X1 U15430 ( .A1(n19075), .A2(n12272), .ZN(n12292) );
  INV_X1 U15431 ( .A(n12273), .ZN(n12274) );
  MUX2_X1 U15432 ( .A(n12274), .B(n12700), .S(n10420), .Z(n12276) );
  NAND2_X1 U15433 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  NAND2_X1 U15434 ( .A1(n12277), .A2(n10431), .ZN(n12287) );
  NAND2_X1 U15435 ( .A1(n12278), .A2(n10635), .ZN(n13218) );
  NAND2_X1 U15436 ( .A1(n13218), .A2(n12279), .ZN(n12285) );
  OAI22_X1 U15437 ( .A1(n12275), .A2(n10375), .B1(n13383), .B2(n12280), .ZN(
        n12281) );
  INV_X1 U15438 ( .A(n12281), .ZN(n12282) );
  NAND2_X1 U15439 ( .A1(n12283), .A2(n12282), .ZN(n12284) );
  AOI21_X1 U15440 ( .B1(n10414), .B2(n12285), .A(n12284), .ZN(n12286) );
  AND2_X1 U15441 ( .A1(n12287), .A2(n12286), .ZN(n13224) );
  INV_X1 U15442 ( .A(n12288), .ZN(n12763) );
  NAND2_X1 U15443 ( .A1(n13224), .A2(n12763), .ZN(n12289) );
  NAND2_X1 U15444 ( .A1(n12314), .A2(n12289), .ZN(n19059) );
  NOR2_X1 U15445 ( .A1(n12290), .A2(n19063), .ZN(n12300) );
  INV_X1 U15446 ( .A(n12300), .ZN(n19074) );
  OR2_X1 U15447 ( .A1(n19059), .A2(n19074), .ZN(n12291) );
  INV_X1 U15448 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13729) );
  NAND3_X1 U15449 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13724) );
  NOR2_X1 U15450 ( .A1(n13729), .A2(n13724), .ZN(n13727) );
  INV_X1 U15451 ( .A(n13727), .ZN(n12293) );
  NAND3_X1 U15452 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n16194), .ZN(n15433) );
  NOR2_X1 U15453 ( .A1(n15281), .A2(n15433), .ZN(n15276) );
  AND2_X1 U15454 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15276), .ZN(
        n12294) );
  INV_X1 U15455 ( .A(n15238), .ZN(n12295) );
  NAND2_X1 U15456 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12305) );
  INV_X1 U15457 ( .A(n12305), .ZN(n12296) );
  NAND2_X1 U15458 ( .A1(n15214), .A2(n12296), .ZN(n15201) );
  NOR4_X1 U15459 ( .A1(n15201), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15200), .A4(n15024), .ZN(n12297) );
  AOI211_X1 U15460 ( .C1(n18939), .C2(n16200), .A(n12298), .B(n12297), .ZN(
        n12309) );
  NAND2_X1 U15461 ( .A1(n19075), .A2(n19059), .ZN(n15468) );
  INV_X1 U15462 ( .A(n18900), .ZN(n15058) );
  OR2_X1 U15463 ( .A1(n12314), .A2(n15058), .ZN(n19057) );
  NAND2_X1 U15464 ( .A1(n16209), .A2(n19057), .ZN(n15431) );
  NAND4_X1 U15465 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n13727), .A4(n13480), .ZN(
        n12299) );
  NAND2_X1 U15466 ( .A1(n15468), .A2(n12299), .ZN(n12302) );
  OR2_X1 U15467 ( .A1(n19059), .A2(n12300), .ZN(n19062) );
  NAND2_X1 U15468 ( .A1(n19057), .A2(n19062), .ZN(n13481) );
  INV_X1 U15469 ( .A(n13481), .ZN(n12301) );
  INV_X1 U15470 ( .A(n15273), .ZN(n15263) );
  OAI21_X1 U15471 ( .B1(n15263), .B2(n15281), .A(n15468), .ZN(n12303) );
  NAND3_X1 U15472 ( .A1(n15452), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n12303), .ZN(n15265) );
  NAND2_X1 U15473 ( .A1(n15431), .A2(n15265), .ZN(n15253) );
  INV_X1 U15474 ( .A(n15253), .ZN(n12304) );
  AOI21_X1 U15475 ( .B1(n15431), .B2(n15238), .A(n12304), .ZN(n15228) );
  OAI21_X1 U15476 ( .B1(n15200), .B2(n12305), .A(n15431), .ZN(n12306) );
  NAND2_X1 U15477 ( .A1(n15228), .A2(n12306), .ZN(n15205) );
  NOR2_X1 U15478 ( .A1(n16209), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12307) );
  OAI21_X1 U15479 ( .B1(n15205), .B2(n12307), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12308) );
  OAI211_X1 U15480 ( .C1(n14889), .C2(n16188), .A(n12309), .B(n12308), .ZN(
        n12310) );
  AOI21_X1 U15481 ( .B1(n12311), .B2(n19056), .A(n12310), .ZN(n12317) );
  NOR2_X1 U15482 ( .A1(n12313), .A2(n12312), .ZN(n19719) );
  NAND2_X1 U15483 ( .A1(n12315), .A2(n19065), .ZN(n12316) );
  NAND2_X1 U15484 ( .A1(n12317), .A2(n12316), .ZN(P2_U3015) );
  NAND2_X1 U15485 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19196) );
  NAND2_X1 U15486 ( .A1(n19196), .A2(n12319), .ZN(n12321) );
  NAND2_X1 U15487 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19508) );
  INV_X1 U15488 ( .A(n19508), .ZN(n19296) );
  INV_X1 U15489 ( .A(n12338), .ZN(n12320) );
  AND2_X1 U15490 ( .A1(n12321), .A2(n12320), .ZN(n19437) );
  AND2_X1 U15491 ( .A1(n19437), .A2(n19682), .ZN(n19230) );
  AOI21_X1 U15492 ( .B1(n12341), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n19230), .ZN(n12322) );
  INV_X1 U15493 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12324) );
  NOR2_X1 U15494 ( .A1(n13050), .A2(n12324), .ZN(n12325) );
  NAND2_X1 U15495 ( .A1(n12326), .A2(n12325), .ZN(n12335) );
  AOI22_X1 U15496 ( .A1(n12341), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19682), .B2(n19714), .ZN(n12328) );
  NAND2_X1 U15497 ( .A1(n12341), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12330) );
  NAND2_X1 U15498 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19705), .ZN(
        n19356) );
  NAND2_X1 U15499 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19714), .ZN(
        n19387) );
  NAND2_X1 U15500 ( .A1(n19356), .A2(n19387), .ZN(n19229) );
  NAND2_X1 U15501 ( .A1(n19682), .A2(n19229), .ZN(n19389) );
  NAND2_X1 U15502 ( .A1(n12330), .A2(n19389), .ZN(n12331) );
  INV_X1 U15503 ( .A(n12332), .ZN(n12333) );
  NOR2_X1 U15504 ( .A1(n15475), .A2(n12333), .ZN(n12334) );
  NAND2_X1 U15505 ( .A1(n12939), .A2(n12940), .ZN(n12336) );
  NAND2_X1 U15506 ( .A1(n9651), .A2(n12337), .ZN(n12343) );
  NAND2_X1 U15507 ( .A1(n12338), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19080) );
  OAI211_X1 U15508 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n12338), .A(
        n19080), .B(n19682), .ZN(n12339) );
  INV_X1 U15509 ( .A(n12339), .ZN(n12340) );
  AOI21_X1 U15510 ( .B1(n12341), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12340), .ZN(n12342) );
  NAND2_X1 U15511 ( .A1(n12345), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12347) );
  INV_X1 U15512 ( .A(n12347), .ZN(n12350) );
  INV_X1 U15513 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19101) );
  NOR2_X1 U15514 ( .A1(n13050), .A2(n19101), .ZN(n12344) );
  NAND2_X1 U15515 ( .A1(n12345), .A2(n12344), .ZN(n13048) );
  NAND2_X1 U15516 ( .A1(n13062), .A2(n12347), .ZN(n12349) );
  AND3_X1 U15517 ( .A1(n13408), .A2(n10635), .A3(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12348) );
  OAI21_X1 U15518 ( .B1(n13045), .B2(n12350), .A(n10227), .ZN(n12960) );
  INV_X1 U15519 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12352) );
  OR2_X1 U15520 ( .A1(n13506), .A2(n13360), .ZN(n13349) );
  INV_X1 U15521 ( .A(n13352), .ZN(n12353) );
  OR2_X1 U15522 ( .A1(n13349), .A2(n12353), .ZN(n13342) );
  NOR2_X1 U15523 ( .A1(n10237), .A2(n13306), .ZN(n13413) );
  AND2_X1 U15524 ( .A1(n13416), .A2(n13413), .ZN(n12355) );
  AOI22_X1 U15525 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15526 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15527 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15528 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12357) );
  NAND4_X1 U15529 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12357), .ZN(
        n12366) );
  AOI22_X1 U15530 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15531 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15532 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15533 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12361) );
  NAND4_X1 U15534 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n12365) );
  OR2_X1 U15535 ( .A1(n12366), .A2(n12365), .ZN(n13629) );
  AOI22_X1 U15536 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10692), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15537 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12432), .ZN(n12369) );
  AOI22_X1 U15538 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15539 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12367) );
  NAND4_X1 U15540 ( .A1(n12370), .A2(n12369), .A3(n12368), .A4(n12367), .ZN(
        n12376) );
  AOI22_X1 U15541 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n10680), .ZN(n12374) );
  AOI22_X1 U15542 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U15543 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15544 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n13078), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12371) );
  NAND4_X1 U15545 ( .A1(n12374), .A2(n12373), .A3(n12372), .A4(n12371), .ZN(
        n12375) );
  AOI22_X1 U15546 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10692), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15547 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12432), .ZN(n12379) );
  AOI22_X1 U15548 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15549 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12377) );
  NAND4_X1 U15550 ( .A1(n12380), .A2(n12379), .A3(n12378), .A4(n12377), .ZN(
        n12386) );
  AOI22_X1 U15551 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__2__SCAN_IN), .B2(n10680), .ZN(n12384) );
  AOI22_X1 U15552 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15553 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15554 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n13078), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12381) );
  NAND4_X1 U15555 ( .A1(n12384), .A2(n12383), .A3(n12382), .A4(n12381), .ZN(
        n12385) );
  NOR2_X1 U15556 ( .A1(n12386), .A2(n12385), .ZN(n13778) );
  INV_X1 U15557 ( .A(n13778), .ZN(n12387) );
  AOI22_X1 U15558 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10692), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12391) );
  AOI22_X1 U15559 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12432), .ZN(n12390) );
  AOI22_X1 U15560 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U15561 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12388) );
  NAND4_X1 U15562 ( .A1(n12391), .A2(n12390), .A3(n12389), .A4(n12388), .ZN(
        n12397) );
  AOI22_X1 U15563 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n10680), .ZN(n12395) );
  AOI22_X1 U15564 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15565 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15566 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n13078), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12392) );
  NAND4_X1 U15567 ( .A1(n12395), .A2(n12394), .A3(n12393), .A4(n12392), .ZN(
        n12396) );
  NOR2_X1 U15568 ( .A1(n12397), .A2(n12396), .ZN(n13791) );
  AOI22_X1 U15569 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10692), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15570 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12432), .ZN(n12400) );
  AOI22_X1 U15571 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15572 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12398) );
  NAND4_X1 U15573 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n12398), .ZN(
        n12407) );
  AOI22_X1 U15574 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__4__SCAN_IN), .B2(n10680), .ZN(n12405) );
  AOI22_X1 U15575 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15576 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15577 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13078), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12402) );
  NAND4_X1 U15578 ( .A1(n12405), .A2(n12404), .A3(n12403), .A4(n12402), .ZN(
        n12406) );
  OR2_X1 U15579 ( .A1(n12407), .A2(n12406), .ZN(n14954) );
  AOI22_X1 U15580 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15581 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15582 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15583 ( .A1(n10681), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12408) );
  NAND4_X1 U15584 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12419) );
  AOI22_X1 U15585 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10680), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15586 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15587 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15588 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13078), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12414) );
  NAND4_X1 U15589 ( .A1(n12417), .A2(n12416), .A3(n12415), .A4(n12414), .ZN(
        n12418) );
  OR2_X1 U15590 ( .A1(n12419), .A2(n12418), .ZN(n13832) );
  AOI22_X1 U15591 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10692), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U15592 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12432), .ZN(n12422) );
  AOI22_X1 U15593 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15594 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12420) );
  NAND4_X1 U15595 ( .A1(n12423), .A2(n12422), .A3(n12421), .A4(n12420), .ZN(
        n12429) );
  AOI22_X1 U15596 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n10680), .ZN(n12427) );
  AOI22_X1 U15597 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15598 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15599 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n13078), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12424) );
  NAND4_X1 U15600 ( .A1(n12427), .A2(n12426), .A3(n12425), .A4(n12424), .ZN(
        n12428) );
  NOR2_X1 U15601 ( .A1(n12429), .A2(n12428), .ZN(n14944) );
  INV_X1 U15602 ( .A(n14944), .ZN(n12430) );
  AOI22_X1 U15603 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10692), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15604 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12432), .ZN(n12435) );
  AOI22_X1 U15605 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10599), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15606 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10681), .B1(
        n10641), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12433) );
  NAND4_X1 U15607 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n12433), .ZN(
        n12442) );
  AOI22_X1 U15608 ( .A1(n10627), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n10680), .ZN(n12440) );
  AOI22_X1 U15609 ( .A1(n12413), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10626), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15610 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10668), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15611 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n13078), .B1(
        n10621), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12437) );
  NAND4_X1 U15612 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        n12441) );
  NOR2_X1 U15613 ( .A1(n12442), .A2(n12441), .ZN(n12461) );
  AOI22_X1 U15614 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15615 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12445) );
  AND2_X1 U15616 ( .A1(n12446), .A2(n12445), .ZN(n12449) );
  AOI22_X1 U15617 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15618 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12447) );
  XNOR2_X1 U15619 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12570) );
  NAND4_X1 U15620 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12570), .ZN(
        n12456) );
  AOI22_X1 U15621 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15622 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12450) );
  AND2_X1 U15623 ( .A1(n12451), .A2(n12450), .ZN(n12454) );
  AOI22_X1 U15624 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U15625 ( .A1(n12454), .A2(n12578), .A3(n12453), .A4(n12452), .ZN(
        n12455) );
  NAND2_X1 U15626 ( .A1(n12456), .A2(n12455), .ZN(n12478) );
  NOR2_X1 U15627 ( .A1(n19737), .A2(n12478), .ZN(n12457) );
  XOR2_X1 U15628 ( .A(n12461), .B(n12457), .Z(n12479) );
  XNOR2_X2 U15629 ( .A(n12458), .B(n12479), .ZN(n14936) );
  INV_X1 U15630 ( .A(n12478), .ZN(n12462) );
  NAND2_X1 U15631 ( .A1(n19737), .A2(n12462), .ZN(n14935) );
  NOR2_X2 U15632 ( .A1(n14936), .A2(n14935), .ZN(n14934) );
  INV_X1 U15633 ( .A(n12479), .ZN(n12459) );
  INV_X1 U15634 ( .A(n12461), .ZN(n12463) );
  AND2_X1 U15635 ( .A1(n12463), .A2(n12462), .ZN(n12476) );
  AOI22_X1 U15636 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15637 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12464) );
  AND2_X1 U15638 ( .A1(n12465), .A2(n12464), .ZN(n12468) );
  AOI22_X1 U15639 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12466) );
  NAND4_X1 U15640 ( .A1(n12468), .A2(n12467), .A3(n12466), .A4(n12570), .ZN(
        n12475) );
  AOI22_X1 U15641 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15642 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12469) );
  AND2_X1 U15643 ( .A1(n12470), .A2(n12469), .ZN(n12473) );
  AOI22_X1 U15644 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12471) );
  NAND4_X1 U15645 ( .A1(n12473), .A2(n12578), .A3(n12472), .A4(n12471), .ZN(
        n12474) );
  AND2_X1 U15646 ( .A1(n12475), .A2(n12474), .ZN(n12477) );
  NAND2_X1 U15647 ( .A1(n12476), .A2(n12477), .ZN(n12480) );
  OAI211_X1 U15648 ( .C1(n12476), .C2(n12477), .A(n12493), .B(n12480), .ZN(
        n14926) );
  NAND2_X1 U15649 ( .A1(n19737), .A2(n12477), .ZN(n14929) );
  INV_X1 U15650 ( .A(n12480), .ZN(n12494) );
  AOI22_X1 U15651 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15652 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12481) );
  AND2_X1 U15653 ( .A1(n12482), .A2(n12481), .ZN(n12485) );
  AOI22_X1 U15654 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12483) );
  NAND4_X1 U15655 ( .A1(n12485), .A2(n12484), .A3(n12483), .A4(n12570), .ZN(
        n12492) );
  AOI22_X1 U15656 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15657 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12486) );
  AND2_X1 U15658 ( .A1(n12487), .A2(n12486), .ZN(n12490) );
  AOI22_X1 U15659 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12488) );
  NAND4_X1 U15660 ( .A1(n12490), .A2(n12578), .A3(n12489), .A4(n12488), .ZN(
        n12491) );
  AND2_X1 U15661 ( .A1(n12492), .A2(n12491), .ZN(n12495) );
  NAND2_X1 U15662 ( .A1(n12494), .A2(n12495), .ZN(n12514) );
  OAI211_X1 U15663 ( .C1(n12494), .C2(n12495), .A(n12493), .B(n12514), .ZN(
        n12498) );
  INV_X1 U15664 ( .A(n12495), .ZN(n12496) );
  NOR2_X1 U15665 ( .A1(n10635), .A2(n12496), .ZN(n14921) );
  INV_X1 U15666 ( .A(n12497), .ZN(n12500) );
  AOI22_X1 U15667 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12503) );
  AOI22_X1 U15668 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12502) );
  AND2_X1 U15669 ( .A1(n12503), .A2(n12502), .ZN(n12506) );
  AOI22_X1 U15670 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12504) );
  NAND4_X1 U15671 ( .A1(n12506), .A2(n12505), .A3(n12504), .A4(n12570), .ZN(
        n12513) );
  AOI22_X1 U15672 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U15673 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12507) );
  AND2_X1 U15674 ( .A1(n12508), .A2(n12507), .ZN(n12511) );
  AOI22_X1 U15675 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12509) );
  NAND4_X1 U15676 ( .A1(n12511), .A2(n12578), .A3(n12510), .A4(n12509), .ZN(
        n12512) );
  NAND2_X1 U15677 ( .A1(n12513), .A2(n12512), .ZN(n12516) );
  AOI21_X1 U15678 ( .B1(n12514), .B2(n12516), .A(n13050), .ZN(n12515) );
  OR2_X1 U15679 ( .A1(n12514), .A2(n12516), .ZN(n12533) );
  NAND2_X1 U15680 ( .A1(n12515), .A2(n12533), .ZN(n12518) );
  XNOR2_X2 U15681 ( .A(n12517), .B(n12518), .ZN(n14913) );
  NOR2_X1 U15682 ( .A1(n10635), .A2(n12516), .ZN(n14912) );
  AOI22_X1 U15683 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U15684 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12521) );
  AND2_X1 U15685 ( .A1(n12522), .A2(n12521), .ZN(n12525) );
  AOI22_X1 U15686 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12523) );
  NAND4_X1 U15687 ( .A1(n12525), .A2(n12524), .A3(n12523), .A4(n12570), .ZN(
        n12532) );
  AOI22_X1 U15688 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U15689 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12526) );
  AND2_X1 U15690 ( .A1(n12527), .A2(n12526), .ZN(n12530) );
  AOI22_X1 U15691 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12528) );
  NAND4_X1 U15692 ( .A1(n12530), .A2(n12578), .A3(n12529), .A4(n12528), .ZN(
        n12531) );
  NAND2_X1 U15693 ( .A1(n12532), .A2(n12531), .ZN(n12535) );
  NOR2_X1 U15694 ( .A1(n12533), .A2(n12535), .ZN(n14898) );
  NOR2_X1 U15695 ( .A1(n10635), .A2(n12535), .ZN(n14906) );
  AOI22_X1 U15696 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U15697 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12536) );
  AND2_X1 U15698 ( .A1(n12537), .A2(n12536), .ZN(n12540) );
  AOI22_X1 U15699 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12538) );
  NAND4_X1 U15700 ( .A1(n12540), .A2(n12539), .A3(n12538), .A4(n12570), .ZN(
        n12547) );
  AOI22_X1 U15701 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U15702 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12541) );
  AND2_X1 U15703 ( .A1(n12542), .A2(n12541), .ZN(n12545) );
  AOI22_X1 U15704 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9646), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12543) );
  NAND4_X1 U15705 ( .A1(n12545), .A2(n12578), .A3(n12544), .A4(n12543), .ZN(
        n12546) );
  NAND2_X1 U15706 ( .A1(n12547), .A2(n12546), .ZN(n12562) );
  AOI22_X1 U15707 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15708 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12549) );
  AND2_X1 U15709 ( .A1(n12550), .A2(n12549), .ZN(n12553) );
  AOI22_X1 U15710 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12551) );
  NAND4_X1 U15711 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12570), .ZN(
        n12561) );
  INV_X1 U15712 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n19585) );
  AOI22_X1 U15713 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12554), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15714 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12555) );
  AND2_X1 U15715 ( .A1(n12556), .A2(n12555), .ZN(n12559) );
  INV_X1 U15716 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n20940) );
  AOI22_X1 U15717 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12557) );
  NAND4_X1 U15718 ( .A1(n12559), .A2(n12578), .A3(n12558), .A4(n12557), .ZN(
        n12560) );
  NAND2_X1 U15719 ( .A1(n12561), .A2(n12560), .ZN(n12565) );
  INV_X1 U15720 ( .A(n12562), .ZN(n14901) );
  AND2_X1 U15721 ( .A1(n10635), .A2(n14901), .ZN(n12563) );
  NAND2_X1 U15722 ( .A1(n14898), .A2(n12563), .ZN(n12564) );
  NOR2_X1 U15723 ( .A1(n12564), .A2(n12565), .ZN(n12566) );
  AOI21_X1 U15724 ( .B1(n12565), .B2(n12564), .A(n12566), .ZN(n14893) );
  NAND2_X1 U15725 ( .A1(n14894), .A2(n14893), .ZN(n14895) );
  INV_X1 U15726 ( .A(n12566), .ZN(n12567) );
  NAND2_X1 U15727 ( .A1(n14895), .A2(n12567), .ZN(n12590) );
  AOI22_X1 U15728 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9644), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15729 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12571) );
  NAND3_X1 U15730 ( .A1(n12572), .A2(n12571), .A3(n12570), .ZN(n12587) );
  AOI22_X1 U15731 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15732 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12573) );
  NAND2_X1 U15733 ( .A1(n12574), .A2(n12573), .ZN(n12586) );
  AOI22_X1 U15734 ( .A1(n12568), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12575), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15735 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12577), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12579) );
  NAND3_X1 U15736 ( .A1(n12580), .A2(n12579), .A3(n12578), .ZN(n12585) );
  AOI22_X1 U15737 ( .A1(n9634), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12548), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15738 ( .A1(n13067), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12581), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12582) );
  NAND2_X1 U15739 ( .A1(n12583), .A2(n12582), .ZN(n12584) );
  OAI22_X1 U15740 ( .A1(n12587), .A2(n12586), .B1(n12585), .B2(n12584), .ZN(
        n12588) );
  XNOR2_X1 U15741 ( .A(n12590), .B(n12589), .ZN(n14241) );
  AND2_X1 U15742 ( .A1(n12275), .A2(n19600), .ZN(n13250) );
  AND2_X1 U15743 ( .A1(n13252), .A2(n13250), .ZN(n12591) );
  AOI21_X1 U15744 ( .B1(n13248), .B2(n13073), .A(n12591), .ZN(n12695) );
  NAND2_X1 U15745 ( .A1(n12593), .A2(n12592), .ZN(n12594) );
  NAND2_X1 U15746 ( .A1(n12695), .A2(n12594), .ZN(n12595) );
  INV_X1 U15747 ( .A(n12597), .ZN(n12598) );
  NOR4_X1 U15748 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12602) );
  NOR4_X1 U15749 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12601) );
  NOR4_X1 U15750 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12600) );
  NOR4_X1 U15751 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12599) );
  NAND4_X1 U15752 ( .A1(n12602), .A2(n12601), .A3(n12600), .A4(n12599), .ZN(
        n12607) );
  NOR4_X1 U15753 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12605) );
  NOR4_X1 U15754 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12604) );
  NOR4_X1 U15755 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12603) );
  NAND4_X1 U15756 ( .A1(n12605), .A2(n12604), .A3(n12603), .A4(n19624), .ZN(
        n12606) );
  INV_X1 U15757 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12609) );
  OR2_X1 U15758 ( .A1(n13380), .A2(n12609), .ZN(n12611) );
  NAND2_X1 U15759 ( .A1(n13380), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12610) );
  NAND2_X1 U15760 ( .A1(n12611), .A2(n12610), .ZN(n19032) );
  INV_X1 U15761 ( .A(n12612), .ZN(n14215) );
  INV_X1 U15762 ( .A(n12613), .ZN(n12614) );
  NAND2_X1 U15763 ( .A1(n14215), .A2(n12614), .ZN(n12615) );
  NAND2_X1 U15764 ( .A1(n12616), .A2(n12615), .ZN(n16005) );
  INV_X1 U15765 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12618) );
  OAI22_X1 U15766 ( .A1(n16005), .A2(n18967), .B1(n18966), .B2(n12618), .ZN(
        n12619) );
  AOI21_X1 U15767 ( .B1(n16065), .B2(n19032), .A(n12619), .ZN(n12622) );
  NOR2_X2 U15768 ( .A1(n12815), .A2(n13382), .ZN(n18940) );
  NOR2_X2 U15769 ( .A1(n12815), .A2(n13380), .ZN(n18938) );
  AOI22_X1 U15770 ( .A1(n18940), .A2(BUF2_REG_30__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12621) );
  OAI21_X1 U15771 ( .B1(n14241), .B2(n18978), .A(n12623), .ZN(P2_U2889) );
  NOR2_X1 U15772 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12625) );
  NOR4_X1 U15773 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12624) );
  NAND4_X1 U15774 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12625), .A4(n12624), .ZN(n12638) );
  NOR4_X1 U15775 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12629) );
  NOR4_X1 U15776 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12628) );
  NOR4_X1 U15777 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12627) );
  NOR4_X1 U15778 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12626) );
  AND4_X1 U15779 ( .A1(n12629), .A2(n12628), .A3(n12627), .A4(n12626), .ZN(
        n12634) );
  NOR4_X1 U15780 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12632) );
  NOR4_X1 U15781 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n12631) );
  NOR4_X1 U15782 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12630) );
  INV_X1 U15783 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20670) );
  AND4_X1 U15784 ( .A1(n12632), .A2(n12631), .A3(n12630), .A4(n20670), .ZN(
        n12633) );
  NAND2_X1 U15785 ( .A1(n12634), .A2(n12633), .ZN(n12635) );
  INV_X1 U15786 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20748) );
  NOR3_X1 U15787 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20748), .ZN(n12637) );
  NOR4_X1 U15788 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12636) );
  NAND4_X1 U15789 ( .A1(n19996), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12637), .A4(
        n12636), .ZN(U214) );
  NOR2_X1 U15790 ( .A1(n13380), .A2(n12638), .ZN(n16302) );
  NAND2_X1 U15791 ( .A1(n16302), .A2(U214), .ZN(U212) );
  AOI211_X1 U15792 ( .C1(n12645), .C2(n12639), .A(n18830), .B(n18936), .ZN(
        n12654) );
  INV_X1 U15793 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19641) );
  OR3_X1 U15794 ( .A1(n12670), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n12640), .ZN(
        n12641) );
  NAND2_X2 U15795 ( .A1(n12642), .A2(n12641), .ZN(n18917) );
  AOI22_X1 U15796 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n18917), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18906), .ZN(n12643) );
  OAI211_X1 U15797 ( .C1(n19641), .C2(n18918), .A(n12643), .B(n18900), .ZN(
        n12653) );
  INV_X1 U15798 ( .A(n12645), .ZN(n15179) );
  NAND2_X1 U15799 ( .A1(n18912), .A2(n18891), .ZN(n18930) );
  OAI22_X1 U15800 ( .A1(n12646), .A2(n18925), .B1(n15179), .B2(n18930), .ZN(
        n12652) );
  NOR2_X1 U15801 ( .A1(n13566), .A2(n12647), .ZN(n12648) );
  OR2_X1 U15802 ( .A1(n13662), .A2(n12648), .ZN(n13635) );
  OAI21_X1 U15803 ( .B1(n12650), .B2(n13615), .A(n12649), .ZN(n16155) );
  OAI22_X1 U15804 ( .A1(n13635), .A2(n18878), .B1(n18916), .B2(n16155), .ZN(
        n12651) );
  AOI211_X1 U15805 ( .C1(n12657), .C2(n12655), .A(n13612), .B(n18936), .ZN(
        n12664) );
  AOI22_X1 U15806 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18906), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n18917), .ZN(n12656) );
  OAI211_X1 U15807 ( .C1(n20932), .C2(n18918), .A(n12656), .B(n18900), .ZN(
        n12663) );
  INV_X1 U15808 ( .A(n12657), .ZN(n15194) );
  OAI22_X1 U15809 ( .A1(n12658), .A2(n18925), .B1(n15194), .B2(n18930), .ZN(
        n12662) );
  AOI21_X1 U15810 ( .B1(n12659), .B2(n13344), .A(n13565), .ZN(n15398) );
  INV_X1 U15811 ( .A(n15398), .ZN(n15195) );
  OAI21_X1 U15812 ( .B1(n12660), .B2(n13466), .A(n13616), .ZN(n15400) );
  OAI22_X1 U15813 ( .A1(n15195), .A2(n18878), .B1(n18916), .B2(n15400), .ZN(
        n12661) );
  OR4_X1 U15814 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        P2_U2842) );
  OR2_X1 U15815 ( .A1(n9647), .A2(n12665), .ZN(n13444) );
  INV_X1 U15816 ( .A(n13444), .ZN(n18933) );
  INV_X1 U15817 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12666) );
  NAND2_X1 U15818 ( .A1(n19682), .A2(n13528), .ZN(n12668) );
  OAI211_X1 U15819 ( .C1(n18933), .C2(n12666), .A(n12668), .B(n12670), .ZN(
        P2_U2814) );
  NOR2_X1 U15820 ( .A1(n18751), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12669)
         );
  INV_X1 U15821 ( .A(n12275), .ZN(n12667) );
  AOI22_X1 U15822 ( .A1(n12669), .A2(n12668), .B1(n12667), .B2(n18751), .ZN(
        P2_U3612) );
  INV_X1 U15823 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12674) );
  INV_X1 U15824 ( .A(n19600), .ZN(n19734) );
  NOR2_X1 U15825 ( .A1(n12670), .A2(n19734), .ZN(n12671) );
  OR2_X1 U15826 ( .A1(n19035), .A2(n12671), .ZN(n12705) );
  AND2_X1 U15827 ( .A1(n12671), .A2(n10635), .ZN(n19033) );
  INV_X1 U15828 ( .A(n19033), .ZN(n12673) );
  AOI22_X1 U15829 ( .A1(n13382), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13380), .ZN(n13525) );
  INV_X1 U15830 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12672) );
  OAI222_X1 U15831 ( .A1(n12674), .A2(n12705), .B1(n12673), .B2(n13525), .C1(
        n12869), .C2(n12672), .ZN(P2_U2982) );
  OAI21_X1 U15832 ( .B1(n12676), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12675), .ZN(n12677) );
  INV_X1 U15833 ( .A(n12677), .ZN(n16201) );
  NOR2_X1 U15834 ( .A1(n18900), .A2(n18919), .ZN(n16206) );
  XNOR2_X1 U15835 ( .A(n18924), .B(n16202), .ZN(n16203) );
  NOR2_X1 U15836 ( .A1(n16134), .A2(n16203), .ZN(n12678) );
  AOI211_X1 U15837 ( .C1(n19042), .C2(n16201), .A(n16206), .B(n12678), .ZN(
        n12681) );
  OAI21_X1 U15838 ( .B1(n19039), .B2(n12679), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12680) );
  OAI211_X1 U15839 ( .C1(n19047), .C2(n9877), .A(n12681), .B(n12680), .ZN(
        P2_U3014) );
  AOI21_X1 U15840 ( .B1(n12683), .B2(n13425), .A(n12682), .ZN(n12684) );
  XOR2_X1 U15841 ( .A(n12684), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n15465) );
  AOI21_X1 U15842 ( .B1(n13527), .B2(n12686), .A(n12685), .ZN(n15464) );
  NOR2_X1 U15843 ( .A1(n18885), .A2(n19620), .ZN(n15467) );
  AOI21_X1 U15844 ( .B1(n19042), .B2(n15464), .A(n15467), .ZN(n12688) );
  NAND2_X1 U15845 ( .A1(n19039), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12687) );
  OAI211_X1 U15846 ( .C1(n19052), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12688), .B(n12687), .ZN(n12689) );
  AOI21_X1 U15847 ( .B1(n19040), .B2(n15465), .A(n12689), .ZN(n12690) );
  OAI21_X1 U15848 ( .B1(n13427), .B2(n19047), .A(n12690), .ZN(P2_U3013) );
  NOR2_X1 U15849 ( .A1(n9647), .A2(n12691), .ZN(n12692) );
  NAND2_X1 U15850 ( .A1(n12790), .A2(n12692), .ZN(n12696) );
  INV_X1 U15851 ( .A(n13248), .ZN(n12693) );
  NAND2_X1 U15852 ( .A1(n12693), .A2(n13244), .ZN(n12764) );
  AND4_X1 U15853 ( .A1(n12696), .A2(n12695), .A3(n12694), .A4(n12764), .ZN(
        n13240) );
  INV_X1 U15854 ( .A(n16213), .ZN(n18755) );
  NAND2_X1 U15855 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19711), .ZN(n15734) );
  OAI22_X1 U15856 ( .A1(n13240), .A2(n18755), .B1(n18758), .B2(n15734), .ZN(
        n12697) );
  INV_X1 U15857 ( .A(n15477), .ZN(n12704) );
  INV_X1 U15858 ( .A(n12698), .ZN(n12699) );
  NOR2_X1 U15859 ( .A1(n12700), .A2(n12699), .ZN(n12701) );
  OR3_X1 U15860 ( .A1(n15477), .A2(n19680), .A3(n13254), .ZN(n12702) );
  OAI21_X1 U15861 ( .B1(n12704), .B2(n12703), .A(n12702), .ZN(P2_U3595) );
  INV_X2 U15862 ( .A(n12705), .ZN(n19036) );
  AOI22_X1 U15863 ( .A1(n19036), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19035), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15864 ( .A1(n13382), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13380), .ZN(n18975) );
  INV_X1 U15865 ( .A(n18975), .ZN(n12706) );
  NAND2_X1 U15866 ( .A1(n19033), .A2(n12706), .ZN(n12820) );
  NAND2_X1 U15867 ( .A1(n12707), .A2(n12820), .ZN(P2_U2955) );
  AOI22_X1 U15868 ( .A1(n19036), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19035), .ZN(n12708) );
  OAI22_X1 U15869 ( .A1(n13380), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13382), .ZN(n12817) );
  INV_X1 U15870 ( .A(n12817), .ZN(n16051) );
  NAND2_X1 U15871 ( .A1(n19033), .A2(n16051), .ZN(n12838) );
  NAND2_X1 U15872 ( .A1(n12708), .A2(n12838), .ZN(P2_U2958) );
  AOI22_X1 U15873 ( .A1(n19036), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19035), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15874 ( .A1(n13382), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13380), .ZN(n18982) );
  INV_X1 U15875 ( .A(n18982), .ZN(n12709) );
  NAND2_X1 U15876 ( .A1(n19033), .A2(n12709), .ZN(n12824) );
  NAND2_X1 U15877 ( .A1(n12710), .A2(n12824), .ZN(P2_U2953) );
  AOI22_X1 U15878 ( .A1(n19036), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19035), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15879 ( .A1(n13382), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13380), .ZN(n15012) );
  INV_X1 U15880 ( .A(n15012), .ZN(n12711) );
  NAND2_X1 U15881 ( .A1(n19033), .A2(n12711), .ZN(n12840) );
  NAND2_X1 U15882 ( .A1(n12712), .A2(n12840), .ZN(P2_U2959) );
  AOI22_X1 U15883 ( .A1(n19036), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19035), .ZN(n12713) );
  MUX2_X1 U15884 ( .A(BUF1_REG_9__SCAN_IN), .B(BUF2_REG_9__SCAN_IN), .S(n13380), .Z(n14997) );
  NAND2_X1 U15885 ( .A1(n19033), .A2(n14997), .ZN(n12828) );
  NAND2_X1 U15886 ( .A1(n12713), .A2(n12828), .ZN(P2_U2961) );
  AOI22_X1 U15887 ( .A1(n19036), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19035), .ZN(n12714) );
  MUX2_X1 U15888 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n13380), .Z(n14983) );
  NAND2_X1 U15889 ( .A1(n19033), .A2(n14983), .ZN(n12832) );
  NAND2_X1 U15890 ( .A1(n12714), .A2(n12832), .ZN(P2_U2963) );
  AOI22_X1 U15891 ( .A1(n19036), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19035), .ZN(n12716) );
  OAI22_X1 U15892 ( .A1(n13380), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13382), .ZN(n12715) );
  INV_X1 U15893 ( .A(n12715), .ZN(n16064) );
  NAND2_X1 U15894 ( .A1(n19033), .A2(n16064), .ZN(n12830) );
  NAND2_X1 U15895 ( .A1(n12716), .A2(n12830), .ZN(P2_U2954) );
  AOI22_X1 U15896 ( .A1(n19036), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19035), .ZN(n12718) );
  OAI22_X1 U15897 ( .A1(n13380), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13382), .ZN(n12717) );
  INV_X1 U15898 ( .A(n12717), .ZN(n16058) );
  NAND2_X1 U15899 ( .A1(n19033), .A2(n16058), .ZN(n12834) );
  NAND2_X1 U15900 ( .A1(n12718), .A2(n12834), .ZN(P2_U2956) );
  AOI22_X1 U15901 ( .A1(n19036), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19035), .ZN(n12720) );
  AOI22_X1 U15902 ( .A1(n13382), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13380), .ZN(n18993) );
  INV_X1 U15903 ( .A(n18993), .ZN(n12719) );
  NAND2_X1 U15904 ( .A1(n19033), .A2(n12719), .ZN(n12826) );
  NAND2_X1 U15905 ( .A1(n12720), .A2(n12826), .ZN(P2_U2952) );
  AOI22_X1 U15906 ( .A1(n19036), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19035), .ZN(n12724) );
  INV_X1 U15907 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n12721) );
  OR2_X1 U15908 ( .A1(n13380), .A2(n12721), .ZN(n12723) );
  NAND2_X1 U15909 ( .A1(n13380), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12722) );
  NAND2_X1 U15910 ( .A1(n12723), .A2(n12722), .ZN(n14966) );
  NAND2_X1 U15911 ( .A1(n19033), .A2(n14966), .ZN(n12822) );
  NAND2_X1 U15912 ( .A1(n12724), .A2(n12822), .ZN(P2_U2980) );
  AOI22_X1 U15913 ( .A1(n19036), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19035), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15914 ( .A1(n13382), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13380), .ZN(n13837) );
  INV_X1 U15915 ( .A(n13837), .ZN(n18957) );
  NAND2_X1 U15916 ( .A1(n19033), .A2(n18957), .ZN(n12836) );
  NAND2_X1 U15917 ( .A1(n12725), .A2(n12836), .ZN(P2_U2957) );
  NAND2_X1 U15918 ( .A1(n19036), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12728) );
  INV_X1 U15919 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16346) );
  OR2_X1 U15920 ( .A1(n13380), .A2(n16346), .ZN(n12727) );
  NAND2_X1 U15921 ( .A1(n13380), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12726) );
  NAND2_X1 U15922 ( .A1(n12727), .A2(n12726), .ZN(n18954) );
  NAND2_X1 U15923 ( .A1(n19033), .A2(n18954), .ZN(n12865) );
  OAI211_X1 U15924 ( .C1(n15004), .C2(n12869), .A(n12728), .B(n12865), .ZN(
        P2_U2960) );
  NAND2_X1 U15925 ( .A1(n19036), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12731) );
  INV_X1 U15926 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16338) );
  OR2_X1 U15927 ( .A1(n13380), .A2(n16338), .ZN(n12730) );
  NAND2_X1 U15928 ( .A1(n13380), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12729) );
  AND2_X1 U15929 ( .A1(n12730), .A2(n12729), .ZN(n14971) );
  INV_X1 U15930 ( .A(n14971), .ZN(n18947) );
  NAND2_X1 U15931 ( .A1(n19033), .A2(n18947), .ZN(n12863) );
  OAI211_X1 U15932 ( .C1(n14970), .C2(n12869), .A(n12731), .B(n12863), .ZN(
        P2_U2964) );
  INV_X1 U15933 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U15934 ( .A1(n19036), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12734) );
  INV_X1 U15935 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16342) );
  OR2_X1 U15936 ( .A1(n13380), .A2(n16342), .ZN(n12733) );
  NAND2_X1 U15937 ( .A1(n13380), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U15938 ( .A1(n12733), .A2(n12732), .ZN(n18950) );
  NAND2_X1 U15939 ( .A1(n19033), .A2(n18950), .ZN(n12867) );
  OAI211_X1 U15940 ( .C1(n12796), .C2(n12869), .A(n12734), .B(n12867), .ZN(
        P2_U2962) );
  NAND2_X1 U15941 ( .A1(n14128), .A2(n20576), .ZN(n19753) );
  INV_X1 U15942 ( .A(n19753), .ZN(n12735) );
  NOR2_X1 U15943 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(n12735), .ZN(n12748)
         );
  INV_X1 U15944 ( .A(n12738), .ZN(n12742) );
  NOR4_X1 U15945 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12743) );
  NOR2_X1 U15946 ( .A1(n12744), .A2(n12743), .ZN(n12883) );
  NAND2_X1 U15947 ( .A1(n12737), .A2(n12883), .ZN(n12772) );
  INV_X1 U15948 ( .A(n12870), .ZN(n14255) );
  OAI21_X1 U15949 ( .B1(n14381), .B2(n14255), .A(n20752), .ZN(n12747) );
  OAI21_X1 U15950 ( .B1(n12748), .B2(n20752), .A(n12747), .ZN(P1_U3487) );
  INV_X1 U15951 ( .A(n12749), .ZN(n12750) );
  XNOR2_X1 U15952 ( .A(n12751), .B(n12750), .ZN(n19066) );
  INV_X1 U15953 ( .A(n12752), .ZN(n12753) );
  NAND2_X1 U15954 ( .A1(n12754), .A2(n12753), .ZN(n12755) );
  AND2_X1 U15955 ( .A1(n12756), .A2(n12755), .ZN(n19055) );
  NAND2_X1 U15956 ( .A1(n19055), .A2(n19042), .ZN(n12758) );
  NOR2_X1 U15957 ( .A1(n18900), .A2(n19622), .ZN(n19053) );
  AOI21_X1 U15958 ( .B1(n19039), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n19053), .ZN(n12757) );
  OAI211_X1 U15959 ( .C1(n19052), .C2(n13434), .A(n12758), .B(n12757), .ZN(
        n12759) );
  AOI21_X1 U15960 ( .B1(n19066), .B2(n19040), .A(n12759), .ZN(n12760) );
  OAI21_X1 U15961 ( .B1(n11918), .B2(n19047), .A(n12760), .ZN(P2_U3012) );
  NAND2_X1 U15962 ( .A1(n10635), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12761) );
  NAND2_X1 U15963 ( .A1(n12764), .A2(n12763), .ZN(n12765) );
  MUX2_X1 U15964 ( .A(n9877), .B(n18920), .S(n14946), .Z(n12766) );
  OAI21_X1 U15965 ( .B1(n19708), .B2(n14961), .A(n12766), .ZN(P2_U2887) );
  INV_X1 U15966 ( .A(n12767), .ZN(n12768) );
  MUX2_X1 U15967 ( .A(n13427), .B(n13421), .S(n14946), .Z(n12770) );
  OAI21_X1 U15968 ( .B1(n19699), .B2(n14961), .A(n12770), .ZN(P2_U2886) );
  AND2_X1 U15969 ( .A1(n13008), .A2(n12968), .ZN(n12771) );
  AOI21_X1 U15970 ( .B1(n12772), .B2(n12745), .A(n12771), .ZN(n19749) );
  NAND2_X1 U15971 ( .A1(n12773), .A2(n20659), .ZN(n20758) );
  NAND3_X1 U15972 ( .A1(n12968), .A2(n20758), .A3(n12998), .ZN(n12775) );
  NAND2_X1 U15973 ( .A1(n12775), .A2(n20661), .ZN(n12776) );
  AND2_X1 U15974 ( .A1(n19749), .A2(n12776), .ZN(n15701) );
  OR2_X1 U15975 ( .A1(n15701), .A2(n19750), .ZN(n19756) );
  INV_X1 U15976 ( .A(n19756), .ZN(n12788) );
  INV_X1 U15977 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12787) );
  INV_X1 U15978 ( .A(n12737), .ZN(n12777) );
  NOR2_X1 U15979 ( .A1(n12777), .A2(n12883), .ZN(n12785) );
  OR2_X1 U15980 ( .A1(n12780), .A2(n14383), .ZN(n12779) );
  AND2_X1 U15981 ( .A1(n12779), .A2(n12778), .ZN(n12898) );
  NOR2_X1 U15982 ( .A1(n12929), .A2(n13019), .ZN(n13007) );
  OR2_X1 U15983 ( .A1(n12780), .A2(n14381), .ZN(n12781) );
  NAND2_X1 U15984 ( .A1(n12888), .A2(n12781), .ZN(n13015) );
  NAND2_X1 U15985 ( .A1(n13015), .A2(n12782), .ZN(n12783) );
  MUX2_X1 U15986 ( .A(n13032), .B(n12783), .S(n13008), .Z(n12784) );
  OAI21_X1 U15987 ( .B1(n12785), .B2(n12784), .A(n20039), .ZN(n15703) );
  OR2_X1 U15988 ( .A1(n19756), .A2(n15703), .ZN(n12786) );
  OAI21_X1 U15989 ( .B1(n12788), .B2(n12787), .A(n12786), .ZN(P1_U3484) );
  NOR2_X1 U15990 ( .A1(n9647), .A2(n18755), .ZN(n12789) );
  AOI21_X1 U15991 ( .B1(n12790), .B2(n12789), .A(n19035), .ZN(n12792) );
  INV_X1 U15992 ( .A(n12791), .ZN(n19735) );
  INV_X1 U15993 ( .A(n19030), .ZN(n12794) );
  NAND2_X1 U15994 ( .A1(n19711), .A2(n13371), .ZN(n19728) );
  INV_X2 U15995 ( .A(n19728), .ZN(n19025) );
  AOI22_X1 U15996 ( .A1(n19025), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12795) );
  OAI21_X1 U15997 ( .B1(n12796), .B2(n18995), .A(n12795), .ZN(P2_U2925) );
  INV_X1 U15998 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U15999 ( .A1(n19025), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12797) );
  OAI21_X1 U16000 ( .B1(n12798), .B2(n18995), .A(n12797), .ZN(P2_U2931) );
  INV_X1 U16001 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U16002 ( .A1(n19025), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12799) );
  OAI21_X1 U16003 ( .B1(n13630), .B2(n18995), .A(n12799), .ZN(P2_U2935) );
  AOI22_X1 U16004 ( .A1(n19025), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12800) );
  OAI21_X1 U16005 ( .B1(n14963), .B2(n18995), .A(n12800), .ZN(P2_U2922) );
  INV_X1 U16006 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U16007 ( .A1(n19025), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12801) );
  OAI21_X1 U16008 ( .B1(n14995), .B2(n18995), .A(n12801), .ZN(P2_U2926) );
  AOI22_X1 U16009 ( .A1(n19025), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12802) );
  OAI21_X1 U16010 ( .B1(n15004), .B2(n18995), .A(n12802), .ZN(P2_U2927) );
  INV_X1 U16011 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U16012 ( .A1(n19025), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12803) );
  OAI21_X1 U16013 ( .B1(n12804), .B2(n18995), .A(n12803), .ZN(P2_U2933) );
  INV_X1 U16014 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13795) );
  AOI22_X1 U16015 ( .A1(n19025), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12805) );
  OAI21_X1 U16016 ( .B1(n13795), .B2(n18995), .A(n12805), .ZN(P2_U2932) );
  INV_X1 U16017 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13836) );
  AOI22_X1 U16018 ( .A1(n19025), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12806) );
  OAI21_X1 U16019 ( .B1(n13836), .B2(n18995), .A(n12806), .ZN(P2_U2930) );
  AOI22_X1 U16020 ( .A1(n19025), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12807) );
  OAI21_X1 U16021 ( .B1(n15011), .B2(n18995), .A(n12807), .ZN(P2_U2928) );
  AOI22_X1 U16022 ( .A1(n19025), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12808) );
  OAI21_X1 U16023 ( .B1(n14981), .B2(n18995), .A(n12808), .ZN(P2_U2924) );
  AOI22_X1 U16024 ( .A1(n19025), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12809) );
  OAI21_X1 U16025 ( .B1(n14970), .B2(n18995), .A(n12809), .ZN(P2_U2923) );
  INV_X1 U16026 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13648) );
  AOI22_X1 U16027 ( .A1(n19025), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12810) );
  OAI21_X1 U16028 ( .B1(n13648), .B2(n18995), .A(n12810), .ZN(P2_U2934) );
  INV_X1 U16029 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U16030 ( .A1(n19025), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12811) );
  OAI21_X1 U16031 ( .B1(n12812), .B2(n18995), .A(n12811), .ZN(P2_U2929) );
  XNOR2_X1 U16032 ( .A(n12814), .B(n12813), .ZN(n18899) );
  AND2_X1 U16033 ( .A1(n18978), .A2(n18967), .ZN(n18964) );
  INV_X1 U16034 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19017) );
  INV_X1 U16035 ( .A(n12815), .ZN(n12816) );
  OAI222_X1 U16036 ( .A1(n18899), .A2(n18964), .B1(n18966), .B2(n19017), .C1(
        n12817), .C2(n18992), .ZN(P2_U2913) );
  OAI21_X1 U16037 ( .B1(n12819), .B2(n12818), .A(n13111), .ZN(n18879) );
  OAI222_X1 U16038 ( .A1(n18879), .A2(n18964), .B1(n18966), .B2(n19015), .C1(
        n18992), .C2(n15012), .ZN(P2_U2912) );
  AOI22_X1 U16039 ( .A1(n19036), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19035), .ZN(n12821) );
  NAND2_X1 U16040 ( .A1(n12821), .A2(n12820), .ZN(P2_U2970) );
  AOI22_X1 U16041 ( .A1(n19036), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19035), .ZN(n12823) );
  NAND2_X1 U16042 ( .A1(n12823), .A2(n12822), .ZN(P2_U2965) );
  AOI22_X1 U16043 ( .A1(n19036), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19035), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U16044 ( .A1(n12825), .A2(n12824), .ZN(P2_U2968) );
  AOI22_X1 U16045 ( .A1(n19036), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19035), .ZN(n12827) );
  NAND2_X1 U16046 ( .A1(n12827), .A2(n12826), .ZN(P2_U2967) );
  AOI22_X1 U16047 ( .A1(n19036), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n19035), .ZN(n12829) );
  NAND2_X1 U16048 ( .A1(n12829), .A2(n12828), .ZN(P2_U2976) );
  AOI22_X1 U16049 ( .A1(n19036), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19035), .ZN(n12831) );
  NAND2_X1 U16050 ( .A1(n12831), .A2(n12830), .ZN(P2_U2969) );
  AOI22_X1 U16051 ( .A1(n19036), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n19035), .ZN(n12833) );
  NAND2_X1 U16052 ( .A1(n12833), .A2(n12832), .ZN(P2_U2978) );
  AOI22_X1 U16053 ( .A1(n19036), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19035), .ZN(n12835) );
  NAND2_X1 U16054 ( .A1(n12835), .A2(n12834), .ZN(P2_U2971) );
  AOI22_X1 U16055 ( .A1(n19036), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19035), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U16056 ( .A1(n12837), .A2(n12836), .ZN(P2_U2972) );
  AOI22_X1 U16057 ( .A1(n19036), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19035), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12839) );
  NAND2_X1 U16058 ( .A1(n12839), .A2(n12838), .ZN(P2_U2973) );
  AOI22_X1 U16059 ( .A1(n19036), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19035), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12841) );
  NAND2_X1 U16060 ( .A1(n12841), .A2(n12840), .ZN(P2_U2974) );
  INV_X1 U16061 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12845) );
  NAND3_X1 U16062 ( .A1(n13284), .A2(n13012), .A3(n13001), .ZN(n12842) );
  OAI21_X1 U16063 ( .B1(n14243), .B2(n20014), .A(n12842), .ZN(n12843) );
  INV_X1 U16064 ( .A(n20758), .ZN(n14121) );
  INV_X1 U16065 ( .A(n13298), .ZN(n15993) );
  OR2_X1 U16066 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15993), .ZN(n19875) );
  NOR2_X4 U16067 ( .A1(n19877), .A2(n19901), .ZN(n15733) );
  AOI22_X1 U16068 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12844) );
  OAI21_X1 U16069 ( .B1(n12845), .B2(n13139), .A(n12844), .ZN(P1_U2917) );
  INV_X1 U16070 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U16071 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12846) );
  OAI21_X1 U16072 ( .B1(n12847), .B2(n13139), .A(n12846), .ZN(P1_U2912) );
  INV_X1 U16073 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U16074 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12848) );
  OAI21_X1 U16075 ( .B1(n12849), .B2(n13139), .A(n12848), .ZN(P1_U2911) );
  INV_X1 U16076 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U16077 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12850) );
  OAI21_X1 U16078 ( .B1(n12851), .B2(n13139), .A(n12850), .ZN(P1_U2920) );
  INV_X1 U16079 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U16080 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12852) );
  OAI21_X1 U16081 ( .B1(n12853), .B2(n13139), .A(n12852), .ZN(P1_U2919) );
  INV_X1 U16082 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U16083 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U16084 ( .B1(n12855), .B2(n13139), .A(n12854), .ZN(P1_U2918) );
  AOI22_X1 U16085 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12856) );
  OAI21_X1 U16086 ( .B1(n11804), .B2(n13139), .A(n12856), .ZN(P1_U2908) );
  INV_X1 U16087 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U16088 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12857) );
  OAI21_X1 U16089 ( .B1(n12858), .B2(n13139), .A(n12857), .ZN(P1_U2909) );
  INV_X1 U16090 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12860) );
  AOI22_X1 U16091 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12859) );
  OAI21_X1 U16092 ( .B1(n12860), .B2(n13139), .A(n12859), .ZN(P1_U2913) );
  INV_X1 U16093 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U16094 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12861) );
  OAI21_X1 U16095 ( .B1(n12862), .B2(n13139), .A(n12861), .ZN(P1_U2907) );
  INV_X1 U16096 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19006) );
  NAND2_X1 U16097 ( .A1(n19036), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12864) );
  OAI211_X1 U16098 ( .C1(n19006), .C2(n12869), .A(n12864), .B(n12863), .ZN(
        P2_U2979) );
  INV_X1 U16099 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19013) );
  NAND2_X1 U16100 ( .A1(n19036), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12866) );
  OAI211_X1 U16101 ( .C1(n19013), .C2(n12869), .A(n12866), .B(n12865), .ZN(
        P2_U2975) );
  NAND2_X1 U16102 ( .A1(n19036), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12868) );
  OAI211_X1 U16103 ( .C1(n10766), .C2(n12869), .A(n12868), .B(n12867), .ZN(
        P2_U2977) );
  NOR2_X1 U16104 ( .A1(n14180), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12872) );
  INV_X1 U16105 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12871) );
  OR2_X1 U16106 ( .A1(n12872), .A2(n12997), .ZN(n14399) );
  NAND2_X1 U16107 ( .A1(n13032), .A2(n13008), .ZN(n12876) );
  NOR2_X1 U16108 ( .A1(n11033), .A2(n20039), .ZN(n12873) );
  NAND3_X1 U16109 ( .A1(n12874), .A2(n12873), .A3(n13277), .ZN(n12969) );
  NAND2_X1 U16110 ( .A1(n12876), .A2(n12875), .ZN(n12877) );
  INV_X1 U16111 ( .A(n12878), .ZN(n12879) );
  AOI21_X1 U16112 ( .B1(n12881), .B2(n12880), .A(n12879), .ZN(n12948) );
  INV_X1 U16113 ( .A(n12948), .ZN(n14402) );
  NAND2_X2 U16114 ( .A1(n19873), .A2(n20039), .ZN(n14460) );
  OAI222_X1 U16115 ( .A1(n14399), .A2(n14448), .B1(n12871), .B2(n19873), .C1(
        n14402), .C2(n14460), .ZN(P1_U2872) );
  NAND2_X1 U16116 ( .A1(n12883), .A2(n20661), .ZN(n13003) );
  OR2_X1 U16117 ( .A1(n15984), .A2(n13003), .ZN(n12887) );
  NAND2_X1 U16118 ( .A1(n20014), .A2(n20661), .ZN(n12884) );
  NAND2_X1 U16119 ( .A1(n12888), .A2(n14381), .ZN(n12916) );
  OAI21_X1 U16120 ( .B1(n12745), .B2(n12884), .A(n12916), .ZN(n12885) );
  NAND2_X1 U16121 ( .A1(n12885), .A2(n13001), .ZN(n12886) );
  OR2_X1 U16122 ( .A1(n12888), .A2(n12737), .ZN(n12890) );
  OAI211_X1 U16123 ( .C1(n13019), .C2(n12973), .A(n12889), .B(n9956), .ZN(
        n12897) );
  OAI211_X1 U16124 ( .C1(n20018), .C2(n14383), .A(n12971), .B(n13010), .ZN(
        n12891) );
  INV_X1 U16125 ( .A(n12891), .ZN(n12895) );
  INV_X1 U16126 ( .A(n13032), .ZN(n12917) );
  OAI211_X1 U16127 ( .C1(n13284), .C2(n12892), .A(n14121), .B(n20661), .ZN(
        n12893) );
  MUX2_X1 U16128 ( .A(n12917), .B(n12893), .S(n13001), .Z(n12894) );
  NAND2_X1 U16129 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13298), .ZN(n15998) );
  INV_X1 U16130 ( .A(n15998), .ZN(n12896) );
  AOI22_X1 U16131 ( .A1(n13012), .A2(n15688), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n12896), .ZN(n15990) );
  OAI21_X1 U16132 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20301), .A(n15990), 
        .ZN(n15987) );
  AND2_X1 U16133 ( .A1(n12898), .A2(n12897), .ZN(n12905) );
  NAND2_X1 U16134 ( .A1(n12899), .A2(n14381), .ZN(n12904) );
  NAND2_X1 U16135 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  NAND2_X1 U16136 ( .A1(n12902), .A2(n20014), .ZN(n12903) );
  INV_X1 U16137 ( .A(n12892), .ZN(n12908) );
  AND4_X1 U16138 ( .A1(n12908), .A2(n12907), .A3(n12906), .A4(n13030), .ZN(
        n12909) );
  NAND3_X1 U16139 ( .A1(n15984), .A2(n13029), .A3(n12909), .ZN(n13273) );
  INV_X1 U16140 ( .A(n13273), .ZN(n13278) );
  OAI22_X1 U16141 ( .A1(n11380), .A2(n13278), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12929), .ZN(n15687) );
  AOI21_X1 U16142 ( .B1(n15687), .B2(n20301), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n12910) );
  NAND2_X1 U16143 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12933) );
  INV_X1 U16144 ( .A(n12933), .ZN(n12923) );
  OAI22_X1 U16145 ( .A1(n12910), .A2(n12923), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15714), .ZN(n12912) );
  INV_X1 U16146 ( .A(n13284), .ZN(n12911) );
  NOR2_X1 U16147 ( .A1(n12911), .A2(n12914), .ZN(n15686) );
  AOI22_X1 U16148 ( .A1(n15987), .A2(n12912), .B1(n20720), .B2(n15686), .ZN(
        n12913) );
  OAI21_X1 U16149 ( .B1(n15987), .B2(n12914), .A(n12913), .ZN(P1_U3474) );
  INV_X1 U16150 ( .A(n15987), .ZN(n20723) );
  XNOR2_X1 U16151 ( .A(n12918), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12920) );
  NAND2_X1 U16152 ( .A1(n12917), .A2(n12916), .ZN(n13282) );
  INV_X1 U16153 ( .A(n12928), .ZN(n12932) );
  NAND2_X1 U16154 ( .A1(n12932), .A2(n12918), .ZN(n13280) );
  NAND2_X1 U16155 ( .A1(n12928), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13275) );
  AND2_X1 U16156 ( .A1(n13280), .A2(n13275), .ZN(n12924) );
  INV_X1 U16157 ( .A(n12924), .ZN(n12919) );
  AOI22_X1 U16158 ( .A1(n13284), .A2(n12920), .B1(n13282), .B2(n12919), .ZN(
        n12922) );
  NAND3_X1 U16159 ( .A1(n13278), .A2(n13277), .A3(n12924), .ZN(n12921) );
  OAI211_X1 U16160 ( .C1(n12915), .C2(n13278), .A(n12922), .B(n12921), .ZN(
        n13272) );
  INV_X1 U16161 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19984) );
  INV_X1 U16162 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U16163 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19984), .B2(n14192), .ZN(
        n12934) );
  AOI222_X1 U16164 ( .A1(n13272), .A2(n20720), .B1(n20719), .B2(n12924), .C1(
        n12923), .C2(n12934), .ZN(n12926) );
  NAND2_X1 U16165 ( .A1(n20723), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12925) );
  OAI21_X1 U16166 ( .B1(n20723), .B2(n12926), .A(n12925), .ZN(P1_U3472) );
  NOR3_X1 U16167 ( .A1(n12929), .A2(n12928), .A3(n10900), .ZN(n12930) );
  AOI21_X1 U16168 ( .B1(n13284), .B2(n10892), .A(n12930), .ZN(n12931) );
  OAI21_X1 U16169 ( .B1(n20433), .B2(n13278), .A(n12931), .ZN(n15689) );
  NAND2_X1 U16170 ( .A1(n12932), .A2(n20719), .ZN(n12935) );
  OAI22_X1 U16171 ( .A1(n12935), .A2(n10900), .B1(n12934), .B2(n12933), .ZN(
        n12936) );
  AOI21_X1 U16172 ( .B1(n15689), .B2(n20720), .A(n12936), .ZN(n12938) );
  NAND2_X1 U16173 ( .A1(n20723), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12937) );
  OAI21_X1 U16174 ( .B1(n20723), .B2(n12938), .A(n12937), .ZN(P1_U3473) );
  INV_X1 U16175 ( .A(n12940), .ZN(n12941) );
  MUX2_X1 U16176 ( .A(n11918), .B(n10456), .S(n14946), .Z(n12942) );
  OAI21_X1 U16177 ( .B1(n13554), .B2(n14961), .A(n12942), .ZN(P2_U2885) );
  OAI21_X1 U16178 ( .B1(n12944), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12943), .ZN(n13038) );
  NAND2_X1 U16179 ( .A1(n19944), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13026) );
  OAI21_X1 U16180 ( .B1(n19932), .B2(n12945), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12946) );
  OAI211_X1 U16181 ( .C1(n13038), .C2(n15902), .A(n13026), .B(n12946), .ZN(
        n12947) );
  AOI21_X1 U16182 ( .B1(n12948), .B2(n19938), .A(n12947), .ZN(n12949) );
  INV_X1 U16183 ( .A(n12949), .ZN(P1_U2999) );
  OR2_X1 U16184 ( .A1(n12951), .A2(n12950), .ZN(n12952) );
  NAND2_X1 U16185 ( .A1(n12952), .A2(n16175), .ZN(n18866) );
  INV_X1 U16186 ( .A(n14997), .ZN(n12953) );
  INV_X1 U16187 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19011) );
  OAI222_X1 U16188 ( .A1(n18866), .A2(n18964), .B1(n12953), .B2(n18992), .C1(
        n19011), .C2(n18966), .ZN(P2_U2910) );
  AND2_X1 U16189 ( .A1(n12954), .A2(n20751), .ZN(n12955) );
  OR2_X2 U16190 ( .A1(n14243), .A2(n12955), .ZN(n19926) );
  OR2_X1 U16191 ( .A1(n19926), .A2(n20014), .ZN(n13140) );
  INV_X1 U16192 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14499) );
  INV_X1 U16193 ( .A(n19916), .ZN(n12958) );
  INV_X1 U16194 ( .A(n19996), .ZN(n19997) );
  INV_X1 U16195 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12956) );
  NOR2_X1 U16196 ( .A1(n19997), .A2(n12956), .ZN(n12957) );
  AOI21_X1 U16197 ( .B1(DATAI_15_), .B2(n19997), .A(n12957), .ZN(n14498) );
  INV_X1 U16198 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19876) );
  OAI222_X1 U16199 ( .A1(n13140), .A2(n14499), .B1(n12958), .B2(n14498), .C1(
        n13141), .C2(n19876), .ZN(P1_U2967) );
  INV_X1 U16200 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n19889) );
  NAND2_X1 U16201 ( .A1(n19926), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n12959) );
  MUX2_X1 U16202 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n19996), .Z(
        n14479) );
  NAND2_X1 U16203 ( .A1(n19916), .A2(n14479), .ZN(n13165) );
  OAI211_X1 U16204 ( .C1(n13140), .C2(n19889), .A(n12959), .B(n13165), .ZN(
        P1_U2960) );
  OAI211_X1 U16205 ( .C1(n12351), .C2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n14945), .B(n13059), .ZN(n12966) );
  OR2_X1 U16206 ( .A1(n13057), .A2(n12962), .ZN(n12963) );
  AND2_X1 U16207 ( .A1(n12961), .A2(n12963), .ZN(n18911) );
  NAND2_X1 U16208 ( .A1(n18911), .A2(n14890), .ZN(n12965) );
  OAI211_X1 U16209 ( .C1(n14890), .C2(n12967), .A(n12966), .B(n12965), .ZN(
        P2_U2882) );
  AND2_X1 U16210 ( .A1(n12973), .A2(n20039), .ZN(n12974) );
  INV_X1 U16211 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19904) );
  NAND2_X1 U16212 ( .A1(n19997), .A2(DATAI_0_), .ZN(n12976) );
  NAND2_X1 U16213 ( .A1(n19996), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12975) );
  AND2_X1 U16214 ( .A1(n12976), .A2(n12975), .ZN(n20007) );
  OAI222_X1 U16215 ( .A1(n14507), .A2(n14402), .B1(n14505), .B2(n19904), .C1(
        n14504), .C2(n20007), .ZN(P1_U2904) );
  OAI21_X1 U16216 ( .B1(n12978), .B2(n12977), .A(n12981), .ZN(n14395) );
  INV_X1 U16217 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19900) );
  NAND2_X1 U16218 ( .A1(n19997), .A2(DATAI_1_), .ZN(n12980) );
  NAND2_X1 U16219 ( .A1(n19996), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12979) );
  AND2_X1 U16220 ( .A1(n12980), .A2(n12979), .ZN(n20015) );
  OAI222_X1 U16221 ( .A1(n14507), .A2(n14395), .B1(n14505), .B2(n19900), .C1(
        n14504), .C2(n20015), .ZN(P1_U2903) );
  NAND2_X1 U16222 ( .A1(n12982), .A2(n12981), .ZN(n12983) );
  NAND2_X1 U16223 ( .A1(n12984), .A2(n12983), .ZN(n19859) );
  INV_X1 U16224 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n19854) );
  OR2_X1 U16225 ( .A1(n15922), .A2(n19854), .ZN(n19967) );
  OAI21_X1 U16226 ( .B1(n15914), .B2(n12985), .A(n19967), .ZN(n12986) );
  AOI21_X1 U16227 ( .B1(n19851), .B2(n15909), .A(n12986), .ZN(n12990) );
  OR2_X1 U16228 ( .A1(n12988), .A2(n12987), .ZN(n19970) );
  NAND3_X1 U16229 ( .A1(n19970), .A2(n19969), .A3(n19939), .ZN(n12989) );
  OAI211_X1 U16230 ( .C1(n19859), .C2(n19998), .A(n12990), .B(n12989), .ZN(
        P1_U2997) );
  INV_X1 U16231 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20903) );
  NAND2_X1 U16232 ( .A1(n19944), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19979) );
  OAI21_X1 U16233 ( .B1(n15914), .B2(n20903), .A(n19979), .ZN(n12994) );
  OAI21_X1 U16234 ( .B1(n12992), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n12991), .ZN(n19983) );
  NOR2_X1 U16235 ( .A1(n19983), .A2(n15902), .ZN(n12993) );
  AOI211_X1 U16236 ( .C1(n15909), .C2(n20903), .A(n12994), .B(n12993), .ZN(
        n12995) );
  OAI21_X1 U16237 ( .B1(n19998), .B2(n14395), .A(n12995), .ZN(P1_U2998) );
  INV_X1 U16238 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12999) );
  INV_X1 U16239 ( .A(n12998), .ZN(n14165) );
  MUX2_X1 U16240 ( .A(n14166), .B(n14161), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n12996) );
  XNOR2_X1 U16241 ( .A(n13041), .B(n12997), .ZN(n14389) );
  XNOR2_X1 U16242 ( .A(n14389), .B(n14168), .ZN(n19980) );
  OAI222_X1 U16243 ( .A1(n14395), .A2(n14460), .B1(n12999), .B2(n19873), .C1(
        n14448), .C2(n19980), .ZN(P1_U2871) );
  NAND2_X1 U16244 ( .A1(n12892), .A2(n20661), .ZN(n13000) );
  AOI22_X1 U16245 ( .A1(n13000), .A2(n9956), .B1(n20756), .B2(n20758), .ZN(
        n13002) );
  OAI21_X1 U16246 ( .B1(n13002), .B2(n13716), .A(n13001), .ZN(n13006) );
  NAND2_X1 U16247 ( .A1(n20014), .A2(n20758), .ZN(n20755) );
  INV_X1 U16248 ( .A(n13003), .ZN(n13004) );
  NAND2_X1 U16249 ( .A1(n20755), .A2(n13004), .ZN(n13005) );
  MUX2_X1 U16250 ( .A(n13006), .B(n13005), .S(n20018), .Z(n13011) );
  NAND2_X1 U16251 ( .A1(n13008), .A2(n13007), .ZN(n13009) );
  NAND3_X1 U16252 ( .A1(n13011), .A2(n13010), .A3(n13009), .ZN(n13013) );
  NAND2_X1 U16253 ( .A1(n13022), .A2(n11112), .ZN(n13014) );
  NAND2_X1 U16254 ( .A1(n13015), .A2(n13014), .ZN(n13016) );
  OR2_X1 U16255 ( .A1(n13017), .A2(n13016), .ZN(n13018) );
  NAND2_X1 U16256 ( .A1(n13020), .A2(n13019), .ZN(n15711) );
  NAND2_X1 U16257 ( .A1(n13022), .A2(n13021), .ZN(n13023) );
  AND2_X1 U16258 ( .A1(n15711), .A2(n13023), .ZN(n13024) );
  INV_X1 U16259 ( .A(n15943), .ZN(n14749) );
  NOR2_X1 U16260 ( .A1(n19944), .A2(n13033), .ZN(n19991) );
  OAI21_X1 U16261 ( .B1(n14749), .B2(n19991), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13027) );
  OAI211_X1 U16262 ( .C1(n19981), .C2(n14399), .A(n13027), .B(n13026), .ZN(
        n13036) );
  OAI211_X1 U16263 ( .C1(n9956), .C2(n13030), .A(n13029), .B(n13028), .ZN(
        n13031) );
  NAND2_X1 U16264 ( .A1(n13033), .A2(n13031), .ZN(n15938) );
  NAND2_X1 U16265 ( .A1(n15938), .A2(n14767), .ZN(n13035) );
  INV_X1 U16266 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13034) );
  AND2_X1 U16267 ( .A1(n13035), .A2(n13034), .ZN(n19990) );
  NOR2_X1 U16268 ( .A1(n13036), .A2(n19990), .ZN(n13037) );
  OAI21_X1 U16269 ( .B1(n13038), .B2(n14832), .A(n13037), .ZN(P1_U3031) );
  INV_X1 U16270 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19898) );
  NAND2_X1 U16271 ( .A1(n19997), .A2(DATAI_2_), .ZN(n13040) );
  NAND2_X1 U16272 ( .A1(n19996), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13039) );
  AND2_X1 U16273 ( .A1(n13040), .A2(n13039), .ZN(n20019) );
  OAI222_X1 U16274 ( .A1(n14507), .A2(n19859), .B1(n14505), .B2(n19898), .C1(
        n14504), .C2(n20019), .ZN(P1_U2902) );
  MUX2_X1 U16275 ( .A(n14155), .B(n14255), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13043) );
  NOR2_X1 U16276 ( .A1(n14180), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13042) );
  NOR2_X1 U16277 ( .A1(n13043), .A2(n13042), .ZN(n13092) );
  XNOR2_X1 U16278 ( .A(n13093), .B(n13092), .ZN(n19964) );
  INV_X1 U16279 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13044) );
  OAI222_X1 U16280 ( .A1(n19964), .A2(n14448), .B1(n19873), .B2(n13044), .C1(
        n19859), .C2(n14460), .ZN(P1_U2870) );
  INV_X1 U16281 ( .A(n13062), .ZN(n13046) );
  INV_X1 U16282 ( .A(n13064), .ZN(n13053) );
  INV_X1 U16283 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13049) );
  NAND2_X1 U16284 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10373), .ZN(
        n13047) );
  OAI211_X1 U16285 ( .C1(n13050), .C2(n13049), .A(n13048), .B(n13047), .ZN(
        n13052) );
  OAI21_X1 U16286 ( .B1(n13053), .B2(n13052), .A(n13051), .ZN(n18959) );
  NOR2_X1 U16287 ( .A1(n13055), .A2(n13054), .ZN(n13056) );
  OR2_X1 U16288 ( .A1(n13057), .A2(n13056), .ZN(n19046) );
  MUX2_X1 U16289 ( .A(n19046), .B(n10479), .S(n14946), .Z(n13058) );
  OAI21_X1 U16290 ( .B1(n18959), .B2(n14961), .A(n13058), .ZN(P2_U2883) );
  XOR2_X1 U16291 ( .A(n13059), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .Z(n13061)
         );
  OAI21_X1 U16292 ( .B1(n10486), .B2(n10240), .A(n13125), .ZN(n18894) );
  MUX2_X1 U16293 ( .A(n10482), .B(n18894), .S(n14890), .Z(n13060) );
  OAI21_X1 U16294 ( .B1(n13061), .B2(n14961), .A(n13060), .ZN(P2_U2881) );
  INV_X1 U16295 ( .A(n13045), .ZN(n13063) );
  NAND2_X1 U16296 ( .A1(n13063), .A2(n13062), .ZN(n13065) );
  INV_X1 U16297 ( .A(n13224), .ZN(n13228) );
  NAND2_X1 U16298 ( .A1(n9652), .A2(n13228), .ZN(n13082) );
  OR2_X1 U16299 ( .A1(n12288), .A2(n13066), .ZN(n13210) );
  INV_X1 U16300 ( .A(n12050), .ZN(n13068) );
  NAND2_X1 U16301 ( .A1(n12261), .A2(n13068), .ZN(n13213) );
  INV_X1 U16302 ( .A(n13069), .ZN(n13071) );
  NAND2_X1 U16303 ( .A1(n13071), .A2(n13070), .ZN(n13206) );
  NAND2_X1 U16304 ( .A1(n13213), .A2(n13206), .ZN(n13072) );
  AOI21_X1 U16305 ( .B1(n13210), .B2(n12444), .A(n13072), .ZN(n13077) );
  INV_X1 U16306 ( .A(n13073), .ZN(n13247) );
  NAND2_X1 U16307 ( .A1(n13074), .A2(n13247), .ZN(n13207) );
  AOI22_X1 U16308 ( .A1(n13207), .A2(n13206), .B1(n12050), .B2(n12261), .ZN(
        n13076) );
  MUX2_X1 U16309 ( .A(n13077), .B(n13076), .S(n13075), .Z(n13080) );
  INV_X1 U16310 ( .A(n13078), .ZN(n13079) );
  AND2_X1 U16311 ( .A1(n13080), .A2(n13079), .ZN(n13081) );
  NAND2_X1 U16312 ( .A1(n13082), .A2(n13081), .ZN(n13233) );
  AOI22_X1 U16313 ( .A1(n13451), .A2(n16215), .B1(n13574), .B2(n13233), .ZN(
        n13084) );
  NAND2_X1 U16314 ( .A1(n15477), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13083) );
  OAI21_X1 U16315 ( .B1(n13084), .B2(n15477), .A(n13083), .ZN(P2_U3596) );
  OR2_X1 U16316 ( .A1(n13086), .A2(n13085), .ZN(n13087) );
  NAND2_X1 U16317 ( .A1(n13333), .A2(n13087), .ZN(n19842) );
  INV_X1 U16318 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n19848) );
  NAND2_X1 U16319 ( .A1(n14163), .A2(n19848), .ZN(n13091) );
  OAI211_X1 U16320 ( .C1(n14168), .C2(P1_EBX_REG_3__SCAN_IN), .A(n13089), .B(
        n14161), .ZN(n13090) );
  AND2_X1 U16321 ( .A1(n13091), .A2(n13090), .ZN(n13096) );
  NAND2_X1 U16322 ( .A1(n13093), .A2(n13092), .ZN(n13095) );
  INV_X1 U16323 ( .A(n19815), .ZN(n13094) );
  AOI21_X1 U16324 ( .B1(n13096), .B2(n13095), .A(n13094), .ZN(n19955) );
  INV_X1 U16325 ( .A(n19873), .ZN(n14458) );
  AOI22_X1 U16326 ( .A1(n19955), .A2(n19869), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14458), .ZN(n13097) );
  OAI21_X1 U16327 ( .B1(n19842), .B2(n14460), .A(n13097), .ZN(P1_U2869) );
  INV_X1 U16328 ( .A(n9653), .ZN(n16146) );
  NOR2_X1 U16329 ( .A1(n16146), .A2(n12964), .ZN(n13098) );
  AOI21_X1 U16330 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n12964), .A(n13098), .ZN(
        n13099) );
  OAI21_X1 U16331 ( .B1(n19683), .B2(n14961), .A(n13099), .ZN(P2_U2884) );
  OR2_X1 U16332 ( .A1(n13101), .A2(n13100), .ZN(n13102) );
  NAND2_X1 U16333 ( .A1(n13102), .A2(n13467), .ZN(n18845) );
  INV_X1 U16334 ( .A(n14983), .ZN(n13103) );
  INV_X1 U16335 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19008) );
  OAI222_X1 U16336 ( .A1(n18845), .A2(n18964), .B1(n13103), .B2(n18992), .C1(
        n19008), .C2(n18966), .ZN(P2_U2908) );
  INV_X1 U16337 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19896) );
  NAND2_X1 U16338 ( .A1(n19997), .A2(DATAI_3_), .ZN(n13105) );
  NAND2_X1 U16339 ( .A1(n19996), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13104) );
  AND2_X1 U16340 ( .A1(n13105), .A2(n13104), .ZN(n20023) );
  OAI222_X1 U16341 ( .A1(n14507), .A2(n19842), .B1(n14505), .B2(n19896), .C1(
        n14504), .C2(n20023), .ZN(P1_U2901) );
  AND2_X1 U16342 ( .A1(n13127), .A2(n13106), .ZN(n13107) );
  NOR2_X1 U16343 ( .A1(n13365), .A2(n13107), .ZN(n16128) );
  INV_X1 U16344 ( .A(n16128), .ZN(n16187) );
  NOR2_X1 U16345 ( .A1(n12060), .A2(n13108), .ZN(n13109) );
  XNOR2_X1 U16346 ( .A(n13109), .B(n16131), .ZN(n13110) );
  NAND2_X1 U16347 ( .A1(n13110), .A2(n18912), .ZN(n13122) );
  INV_X1 U16348 ( .A(n13111), .ZN(n13112) );
  OR2_X1 U16349 ( .A1(n13113), .A2(n13112), .ZN(n13115) );
  INV_X1 U16350 ( .A(n12950), .ZN(n13114) );
  AND2_X1 U16351 ( .A1(n13115), .A2(n13114), .ZN(n18953) );
  OAI21_X1 U16352 ( .B1(n18918), .B2(n13116), .A(n18900), .ZN(n13120) );
  AOI22_X1 U16353 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18906), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n18917), .ZN(n13117) );
  OAI21_X1 U16354 ( .B1(n13118), .B2(n18925), .A(n13117), .ZN(n13119) );
  AOI211_X1 U16355 ( .C1(n18922), .C2(n18953), .A(n13120), .B(n13119), .ZN(
        n13121) );
  OAI211_X1 U16356 ( .C1(n16187), .C2(n18878), .A(n13122), .B(n13121), .ZN(
        P2_U2847) );
  XNOR2_X1 U16357 ( .A(n13123), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U16358 ( .A1(n13125), .A2(n13124), .ZN(n13126) );
  NAND2_X1 U16359 ( .A1(n13127), .A2(n13126), .ZN(n18877) );
  MUX2_X1 U16360 ( .A(n18877), .B(n10869), .S(n14946), .Z(n13128) );
  OAI21_X1 U16361 ( .B1(n13129), .B2(n14961), .A(n13128), .ZN(P2_U2880) );
  INV_X1 U16362 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16363 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19901), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15733), .ZN(n13130) );
  OAI21_X1 U16364 ( .B1(n13131), .B2(n13139), .A(n13130), .ZN(P1_U2906) );
  INV_X1 U16365 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13133) );
  AOI22_X1 U16366 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13132) );
  OAI21_X1 U16367 ( .B1(n13133), .B2(n13139), .A(n13132), .ZN(P1_U2914) );
  INV_X1 U16368 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U16369 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13134) );
  OAI21_X1 U16370 ( .B1(n13135), .B2(n13139), .A(n13134), .ZN(P1_U2916) );
  INV_X1 U16371 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16372 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13136) );
  OAI21_X1 U16373 ( .B1(n13137), .B2(n13139), .A(n13136), .ZN(P1_U2915) );
  AOI22_X1 U16374 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13138) );
  OAI21_X1 U16375 ( .B1(n11761), .B2(n13139), .A(n13138), .ZN(P1_U2910) );
  AOI22_X1 U16376 ( .A1(n19929), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19926), .ZN(n13144) );
  NAND2_X1 U16377 ( .A1(n19997), .A2(DATAI_4_), .ZN(n13143) );
  NAND2_X1 U16378 ( .A1(n19996), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13142) );
  AND2_X1 U16379 ( .A1(n13143), .A2(n13142), .ZN(n20026) );
  INV_X1 U16380 ( .A(n20026), .ZN(n14490) );
  NAND2_X1 U16381 ( .A1(n19916), .A2(n14490), .ZN(n13174) );
  NAND2_X1 U16382 ( .A1(n13144), .A2(n13174), .ZN(P1_U2941) );
  AOI22_X1 U16383 ( .A1(n19929), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19926), .ZN(n13145) );
  INV_X1 U16384 ( .A(n20007), .ZN(n15864) );
  NAND2_X1 U16385 ( .A1(n19916), .A2(n15864), .ZN(n13167) );
  NAND2_X1 U16386 ( .A1(n13145), .A2(n13167), .ZN(P1_U2952) );
  AOI22_X1 U16387 ( .A1(n19929), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19926), .ZN(n13148) );
  NAND2_X1 U16388 ( .A1(n19997), .A2(DATAI_5_), .ZN(n13147) );
  NAND2_X1 U16389 ( .A1(n19996), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13146) );
  AND2_X1 U16390 ( .A1(n13147), .A2(n13146), .ZN(n20030) );
  INV_X1 U16391 ( .A(n20030), .ZN(n14486) );
  NAND2_X1 U16392 ( .A1(n19916), .A2(n14486), .ZN(n13159) );
  NAND2_X1 U16393 ( .A1(n13148), .A2(n13159), .ZN(P1_U2957) );
  AOI22_X1 U16394 ( .A1(n19929), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19926), .ZN(n13151) );
  NAND2_X1 U16395 ( .A1(n19997), .A2(DATAI_6_), .ZN(n13150) );
  NAND2_X1 U16396 ( .A1(n19996), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13149) );
  AND2_X1 U16397 ( .A1(n13150), .A2(n13149), .ZN(n20034) );
  INV_X1 U16398 ( .A(n20034), .ZN(n15855) );
  NAND2_X1 U16399 ( .A1(n19916), .A2(n15855), .ZN(n13161) );
  NAND2_X1 U16400 ( .A1(n13151), .A2(n13161), .ZN(P1_U2958) );
  AOI22_X1 U16401 ( .A1(n19929), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19926), .ZN(n13154) );
  NAND2_X1 U16402 ( .A1(n19997), .A2(DATAI_7_), .ZN(n13153) );
  NAND2_X1 U16403 ( .A1(n19996), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13152) );
  AND2_X1 U16404 ( .A1(n13153), .A2(n13152), .ZN(n20042) );
  INV_X1 U16405 ( .A(n20042), .ZN(n14482) );
  NAND2_X1 U16406 ( .A1(n19916), .A2(n14482), .ZN(n13163) );
  NAND2_X1 U16407 ( .A1(n13154), .A2(n13163), .ZN(P1_U2959) );
  AOI22_X1 U16408 ( .A1(n19929), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19926), .ZN(n13155) );
  INV_X1 U16409 ( .A(n20019), .ZN(n15859) );
  NAND2_X1 U16410 ( .A1(n19916), .A2(n15859), .ZN(n13172) );
  NAND2_X1 U16411 ( .A1(n13155), .A2(n13172), .ZN(P1_U2939) );
  AOI22_X1 U16412 ( .A1(n19929), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19926), .ZN(n13156) );
  INV_X1 U16413 ( .A(n20023), .ZN(n14494) );
  NAND2_X1 U16414 ( .A1(n19916), .A2(n14494), .ZN(n13157) );
  NAND2_X1 U16415 ( .A1(n13156), .A2(n13157), .ZN(P1_U2940) );
  AOI22_X1 U16416 ( .A1(n19929), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19926), .ZN(n13158) );
  NAND2_X1 U16417 ( .A1(n13158), .A2(n13157), .ZN(P1_U2955) );
  AOI22_X1 U16418 ( .A1(n19929), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19926), .ZN(n13160) );
  NAND2_X1 U16419 ( .A1(n13160), .A2(n13159), .ZN(P1_U2942) );
  AOI22_X1 U16420 ( .A1(n19929), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19926), .ZN(n13162) );
  NAND2_X1 U16421 ( .A1(n13162), .A2(n13161), .ZN(P1_U2943) );
  AOI22_X1 U16422 ( .A1(n19929), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19926), .ZN(n13164) );
  NAND2_X1 U16423 ( .A1(n13164), .A2(n13163), .ZN(P1_U2944) );
  AOI22_X1 U16424 ( .A1(n19929), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19926), .ZN(n13166) );
  NAND2_X1 U16425 ( .A1(n13166), .A2(n13165), .ZN(P1_U2945) );
  AOI22_X1 U16426 ( .A1(n19929), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19926), .ZN(n13168) );
  NAND2_X1 U16427 ( .A1(n13168), .A2(n13167), .ZN(P1_U2937) );
  AOI22_X1 U16428 ( .A1(n19929), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19926), .ZN(n13169) );
  INV_X1 U16429 ( .A(n20015), .ZN(n13718) );
  NAND2_X1 U16430 ( .A1(n19916), .A2(n13718), .ZN(n13170) );
  NAND2_X1 U16431 ( .A1(n13169), .A2(n13170), .ZN(P1_U2938) );
  AOI22_X1 U16432 ( .A1(n19929), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19926), .ZN(n13171) );
  NAND2_X1 U16433 ( .A1(n13171), .A2(n13170), .ZN(P1_U2953) );
  AOI22_X1 U16434 ( .A1(n19929), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19926), .ZN(n13173) );
  NAND2_X1 U16435 ( .A1(n13173), .A2(n13172), .ZN(P1_U2954) );
  AOI22_X1 U16436 ( .A1(n19929), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19926), .ZN(n13175) );
  NAND2_X1 U16437 ( .A1(n13175), .A2(n13174), .ZN(P1_U2956) );
  NAND2_X1 U16438 ( .A1(n13177), .A2(n13176), .ZN(n13180) );
  INV_X1 U16439 ( .A(n13178), .ZN(n13179) );
  XNOR2_X1 U16440 ( .A(n13554), .B(n19692), .ZN(n13188) );
  XNOR2_X1 U16441 ( .A(n13182), .B(n13181), .ZN(n15466) );
  NAND2_X1 U16442 ( .A1(n19699), .A2(n15466), .ZN(n13185) );
  OAI21_X1 U16443 ( .B1(n19699), .B2(n15466), .A(n13185), .ZN(n18977) );
  XNOR2_X1 U16444 ( .A(n13184), .B(n13183), .ZN(n16199) );
  NOR2_X1 U16445 ( .A1(n19708), .A2(n16199), .ZN(n18985) );
  NOR2_X1 U16446 ( .A1(n18977), .A2(n18985), .ZN(n18976) );
  INV_X1 U16447 ( .A(n13185), .ZN(n13186) );
  NOR2_X1 U16448 ( .A1(n18976), .A2(n13186), .ZN(n13187) );
  NOR2_X1 U16449 ( .A1(n13188), .A2(n13187), .ZN(n13553) );
  AOI21_X1 U16450 ( .B1(n13188), .B2(n13187), .A(n13553), .ZN(n13192) );
  AOI22_X1 U16451 ( .A1(n18958), .A2(n16064), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n18983), .ZN(n13191) );
  INV_X1 U16452 ( .A(n19692), .ZN(n13189) );
  NAND2_X1 U16453 ( .A1(n13189), .A2(n18984), .ZN(n13190) );
  OAI211_X1 U16454 ( .C1(n13192), .C2(n18978), .A(n13191), .B(n13190), .ZN(
        P2_U2917) );
  NAND2_X1 U16455 ( .A1(n9642), .A2(n13193), .ZN(n13194) );
  XNOR2_X1 U16456 ( .A(n16141), .B(n13194), .ZN(n13204) );
  OAI22_X1 U16457 ( .A1(n16152), .A2(n18931), .B1(n10675), .B2(n18918), .ZN(
        n13200) );
  OR2_X1 U16458 ( .A1(n13196), .A2(n13195), .ZN(n13198) );
  NAND2_X1 U16459 ( .A1(n13198), .A2(n13197), .ZN(n19686) );
  OAI22_X1 U16460 ( .A1(n13489), .A2(n18925), .B1(n18916), .B2(n19686), .ZN(
        n13199) );
  AOI211_X1 U16461 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n18917), .A(n13200), .B(
        n13199), .ZN(n13202) );
  NAND2_X1 U16462 ( .A1(n9652), .A2(n18927), .ZN(n13201) );
  OAI211_X1 U16463 ( .C1(n19683), .C2(n13444), .A(n13202), .B(n13201), .ZN(
        n13203) );
  AOI21_X1 U16464 ( .B1(n13204), .B2(n18912), .A(n13203), .ZN(n13205) );
  INV_X1 U16465 ( .A(n13205), .ZN(P2_U2852) );
  NAND2_X1 U16466 ( .A1(n11911), .A2(n13228), .ZN(n13217) );
  NOR2_X1 U16467 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13214) );
  NAND2_X1 U16468 ( .A1(n12444), .A2(n13206), .ZN(n13208) );
  NAND2_X1 U16469 ( .A1(n13207), .A2(n13208), .ZN(n13212) );
  INV_X1 U16470 ( .A(n13208), .ZN(n13209) );
  NAND2_X1 U16471 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  OAI211_X1 U16472 ( .C1(n13214), .C2(n13213), .A(n13212), .B(n13211), .ZN(
        n13215) );
  INV_X1 U16473 ( .A(n13215), .ZN(n13216) );
  NAND2_X1 U16474 ( .A1(n13217), .A2(n13216), .ZN(n13575) );
  INV_X1 U16475 ( .A(n13575), .ZN(n13232) );
  NAND2_X1 U16476 ( .A1(n13218), .A2(n12265), .ZN(n13226) );
  OAI21_X1 U16477 ( .B1(n13220), .B2(n13219), .A(n13226), .ZN(n13223) );
  NAND2_X1 U16478 ( .A1(n12261), .A2(n13221), .ZN(n13222) );
  OAI211_X1 U16479 ( .C1(n13427), .C2(n13224), .A(n13223), .B(n13222), .ZN(
        n13530) );
  INV_X1 U16480 ( .A(n13530), .ZN(n13225) );
  INV_X1 U16481 ( .A(n19196), .ZN(n19294) );
  AOI21_X1 U16482 ( .B1(n13225), .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n19294), .ZN(n13230) );
  MUX2_X1 U16483 ( .A(n13226), .B(n12261), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13227) );
  AOI21_X1 U16484 ( .B1(n18928), .B2(n13228), .A(n13227), .ZN(n15474) );
  INV_X1 U16485 ( .A(n15474), .ZN(n13229) );
  OAI22_X1 U16486 ( .A1(n13230), .A2(n13229), .B1(n19705), .B2(n13530), .ZN(
        n13231) );
  AOI211_X1 U16487 ( .C1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n13232), .A(
        n13240), .B(n13231), .ZN(n13237) );
  INV_X1 U16488 ( .A(n13240), .ZN(n13234) );
  MUX2_X1 U16489 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13233), .S(
        n13234), .Z(n13262) );
  INV_X1 U16490 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19690) );
  AOI22_X1 U16491 ( .A1(n13240), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n13575), .B2(n13234), .ZN(n13239) );
  NOR2_X1 U16492 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n13239), .ZN(
        n13235) );
  OR3_X1 U16493 ( .A1(n13237), .A2(n13262), .A3(n13235), .ZN(n13236) );
  AOI22_X1 U16494 ( .A1(n13237), .A2(n13262), .B1(n19690), .B2(n13236), .ZN(
        n13238) );
  OR2_X1 U16495 ( .A1(n13238), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n13264) );
  INV_X1 U16496 ( .A(n13239), .ZN(n13261) );
  NAND2_X1 U16497 ( .A1(n13240), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13259) );
  INV_X1 U16498 ( .A(n13241), .ZN(n13242) );
  NAND2_X1 U16499 ( .A1(n13243), .A2(n13242), .ZN(n13246) );
  NAND2_X1 U16500 ( .A1(n13248), .A2(n13244), .ZN(n13245) );
  OAI211_X1 U16501 ( .C1(n13248), .C2(n13247), .A(n13246), .B(n13245), .ZN(
        n19722) );
  NOR2_X1 U16502 ( .A1(n13250), .A2(n13249), .ZN(n13251) );
  AND2_X1 U16503 ( .A1(n13252), .A2(n13251), .ZN(n18756) );
  OAI21_X1 U16504 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n18756), .ZN(n13256) );
  NAND2_X1 U16505 ( .A1(n13253), .A2(n13399), .ZN(n13255) );
  NAND3_X1 U16506 ( .A1(n13256), .A2(n13255), .A3(n13254), .ZN(n13257) );
  NOR2_X1 U16507 ( .A1(n19722), .A2(n13257), .ZN(n13258) );
  NAND2_X1 U16508 ( .A1(n13259), .A2(n13258), .ZN(n13260) );
  AOI21_X1 U16509 ( .B1(n13262), .B2(n13261), .A(n13260), .ZN(n13263) );
  NAND2_X1 U16510 ( .A1(n13264), .A2(n13263), .ZN(n16212) );
  OAI21_X1 U16511 ( .B1(n16212), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13270) );
  INV_X1 U16512 ( .A(n13265), .ZN(n13267) );
  OR2_X1 U16513 ( .A1(n13266), .A2(n19733), .ZN(n19730) );
  AOI21_X1 U16514 ( .B1(n13268), .B2(n13267), .A(n19730), .ZN(n13269) );
  OAI21_X1 U16515 ( .B1(n16214), .B2(n13371), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13271) );
  NAND2_X1 U16516 ( .A1(n13271), .A2(n15734), .ZN(P2_U3593) );
  NOR2_X1 U16517 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n14128), .ZN(n13295) );
  MUX2_X1 U16518 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13272), .S(
        n15688), .Z(n15694) );
  AOI22_X1 U16519 ( .A1(n13295), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15694), .B2(n14128), .ZN(n13292) );
  NAND2_X1 U16520 ( .A1(n20727), .A2(n13273), .ZN(n13288) );
  NAND2_X1 U16521 ( .A1(n13275), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13276) );
  NAND2_X1 U16522 ( .A1(n11184), .A2(n13276), .ZN(n20718) );
  NAND3_X1 U16523 ( .A1(n13278), .A2(n13277), .A3(n20718), .ZN(n13286) );
  NAND2_X1 U16524 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13279) );
  XNOR2_X1 U16525 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13279), .ZN(
        n13283) );
  XNOR2_X1 U16526 ( .A(n13280), .B(n10891), .ZN(n13281) );
  AOI22_X1 U16527 ( .A1(n13284), .A2(n13283), .B1(n13282), .B2(n13281), .ZN(
        n13285) );
  AND2_X1 U16528 ( .A1(n13286), .A2(n13285), .ZN(n13287) );
  NAND2_X1 U16529 ( .A1(n13288), .A2(n13287), .ZN(n20721) );
  NAND2_X1 U16530 ( .A1(n20721), .A2(n15688), .ZN(n13290) );
  OR2_X1 U16531 ( .A1(n15688), .A2(n10890), .ZN(n13289) );
  NAND2_X1 U16532 ( .A1(n13290), .A2(n13289), .ZN(n15695) );
  AOI22_X1 U16533 ( .A1(n15695), .A2(n14128), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13295), .ZN(n13291) );
  XNOR2_X1 U16534 ( .A(n13293), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19821) );
  OAI21_X1 U16535 ( .B1(n19821), .B2(n15984), .A(n15688), .ZN(n13297) );
  INV_X1 U16536 ( .A(n15688), .ZN(n13294) );
  AOI21_X1 U16537 ( .B1(n13294), .B2(n15988), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13296) );
  AOI22_X1 U16538 ( .A1(n13297), .A2(n13296), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13295), .ZN(n15705) );
  OAI21_X1 U16539 ( .B1(n15699), .B2(n10900), .A(n15705), .ZN(n13300) );
  NOR2_X1 U16540 ( .A1(n13300), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13299) );
  NAND2_X1 U16541 ( .A1(n20750), .A2(n14128), .ZN(n15994) );
  INV_X1 U16542 ( .A(n15994), .ZN(n20765) );
  NOR2_X1 U16543 ( .A1(n13300), .A2(n15993), .ZN(n15717) );
  NAND2_X1 U16544 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20301), .ZN(n20728) );
  INV_X1 U16545 ( .A(n20728), .ZN(n14837) );
  OAI22_X1 U16546 ( .A1(n9650), .A2(n20573), .B1(n11380), .B2(n14837), .ZN(
        n13301) );
  OAI21_X1 U16547 ( .B1(n15717), .B2(n13301), .A(n20738), .ZN(n13302) );
  OAI21_X1 U16548 ( .B1(n20738), .B2(n20464), .A(n13302), .ZN(P1_U3478) );
  NOR2_X1 U16549 ( .A1(n13371), .A2(n19680), .ZN(n18752) );
  AOI21_X1 U16550 ( .B1(n19600), .B2(n18752), .A(n16213), .ZN(n13305) );
  NOR2_X1 U16551 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13371), .ZN(n13303) );
  OAI211_X1 U16552 ( .C1(n16214), .C2(n13303), .A(n19734), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13304) );
  OAI211_X1 U16553 ( .C1(n16214), .C2(n13305), .A(n13304), .B(n18883), .ZN(
        P2_U3177) );
  NAND2_X1 U16554 ( .A1(n13123), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13307) );
  INV_X1 U16555 ( .A(n13307), .ZN(n13414) );
  OAI211_X1 U16556 ( .C1(n13414), .C2(n13308), .A(n14945), .B(n13361), .ZN(
        n13310) );
  NAND2_X1 U16557 ( .A1(n12964), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13309) );
  OAI211_X1 U16558 ( .C1(n16187), .C2(n12964), .A(n13310), .B(n13309), .ZN(
        P2_U2879) );
  OAI21_X1 U16559 ( .B1(n13313), .B2(n13312), .A(n13311), .ZN(n13314) );
  INV_X1 U16560 ( .A(n13314), .ZN(n19957) );
  NAND2_X1 U16561 ( .A1(n19957), .A2(n19939), .ZN(n13318) );
  INV_X1 U16562 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n19839) );
  NOR2_X1 U16563 ( .A1(n15922), .A2(n19839), .ZN(n19954) );
  NOR2_X1 U16564 ( .A1(n15914), .A2(n13315), .ZN(n13316) );
  AOI211_X1 U16565 ( .C1(n15909), .C2(n19835), .A(n19954), .B(n13316), .ZN(
        n13317) );
  OAI211_X1 U16566 ( .C1(n19998), .C2(n19842), .A(n13318), .B(n13317), .ZN(
        P1_U2996) );
  INV_X1 U16567 ( .A(n19051), .ZN(n13322) );
  NOR2_X1 U16568 ( .A1(n18891), .A2(n13319), .ZN(n13321) );
  AOI21_X1 U16569 ( .B1(n13322), .B2(n13321), .A(n18883), .ZN(n13320) );
  OAI21_X1 U16570 ( .B1(n13322), .B2(n13321), .A(n13320), .ZN(n13332) );
  INV_X1 U16571 ( .A(n19046), .ZN(n13330) );
  AOI22_X1 U16572 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18906), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n18917), .ZN(n13327) );
  INV_X1 U16573 ( .A(n13197), .ZN(n13323) );
  XNOR2_X1 U16574 ( .A(n13324), .B(n13323), .ZN(n13556) );
  INV_X1 U16575 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19625) );
  OAI21_X1 U16576 ( .B1(n18918), .B2(n19625), .A(n18885), .ZN(n13325) );
  AOI21_X1 U16577 ( .B1(n18922), .B2(n13556), .A(n13325), .ZN(n13326) );
  OAI211_X1 U16578 ( .C1(n13328), .C2(n18925), .A(n13327), .B(n13326), .ZN(
        n13329) );
  AOI21_X1 U16579 ( .B1(n13330), .B2(n18927), .A(n13329), .ZN(n13331) );
  OAI211_X1 U16580 ( .C1(n18959), .C2(n13444), .A(n13332), .B(n13331), .ZN(
        P2_U2851) );
  XOR2_X1 U16581 ( .A(n13334), .B(n13333), .Z(n19937) );
  INV_X1 U16582 ( .A(n19937), .ZN(n13335) );
  INV_X1 U16583 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19894) );
  OAI222_X1 U16584 ( .A1(n14504), .A2(n20026), .B1(n14489), .B2(n13335), .C1(
        n19894), .C2(n14505), .ZN(P1_U2900) );
  OR2_X1 U16585 ( .A1(n13337), .A2(n13336), .ZN(n13338) );
  AND2_X1 U16586 ( .A1(n13589), .A2(n13338), .ZN(n19867) );
  INV_X1 U16587 ( .A(n19867), .ZN(n13340) );
  INV_X1 U16588 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13339) );
  OAI222_X1 U16589 ( .A1(n13340), .A2(n14507), .B1(n13339), .B2(n14505), .C1(
        n14504), .C2(n20030), .ZN(P1_U2899) );
  INV_X1 U16590 ( .A(n14966), .ZN(n13341) );
  INV_X1 U16591 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19004) );
  OAI222_X1 U16592 ( .A1(n15400), .A2(n18964), .B1(n13341), .B2(n18992), .C1(
        n19004), .C2(n18966), .ZN(P2_U2906) );
  NOR2_X1 U16593 ( .A1(n13361), .A2(n13342), .ZN(n13350) );
  XNOR2_X1 U16594 ( .A(n13350), .B(n13343), .ZN(n13348) );
  OAI21_X1 U16595 ( .B1(n13345), .B2(n13355), .A(n13344), .ZN(n15412) );
  INV_X1 U16596 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13346) );
  MUX2_X1 U16597 ( .A(n15412), .B(n13346), .S(n14946), .Z(n13347) );
  OAI21_X1 U16598 ( .B1(n13348), .B2(n14961), .A(n13347), .ZN(P2_U2875) );
  NOR2_X1 U16599 ( .A1(n13361), .A2(n13349), .ZN(n13504) );
  INV_X1 U16600 ( .A(n13350), .ZN(n13351) );
  OAI211_X1 U16601 ( .C1(n13504), .C2(n13352), .A(n13351), .B(n14945), .ZN(
        n13359) );
  NAND2_X1 U16602 ( .A1(n13354), .A2(n13353), .ZN(n13357) );
  INV_X1 U16603 ( .A(n13355), .ZN(n13356) );
  NAND2_X1 U16604 ( .A1(n14890), .A2(n18844), .ZN(n13358) );
  OAI211_X1 U16605 ( .C1(n14890), .C2(n10500), .A(n13359), .B(n13358), .ZN(
        P2_U2876) );
  INV_X1 U16606 ( .A(n13361), .ZN(n13363) );
  OR2_X1 U16607 ( .A1(n13361), .A2(n13360), .ZN(n13505) );
  OAI211_X1 U16608 ( .C1(n13363), .C2(n13362), .A(n14945), .B(n13505), .ZN(
        n13368) );
  NOR2_X1 U16609 ( .A1(n13365), .A2(n13364), .ZN(n13366) );
  OR2_X1 U16610 ( .A1(n13502), .A2(n13366), .ZN(n18867) );
  INV_X1 U16611 ( .A(n18867), .ZN(n16114) );
  NAND2_X1 U16612 ( .A1(n16114), .A2(n14890), .ZN(n13367) );
  OAI211_X1 U16613 ( .C1(n14890), .C2(n10496), .A(n13368), .B(n13367), .ZN(
        P2_U2878) );
  INV_X1 U16614 ( .A(n19682), .ZN(n19684) );
  NAND2_X1 U16615 ( .A1(n19690), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19268) );
  INV_X1 U16616 ( .A(n19268), .ZN(n19295) );
  NAND2_X1 U16617 ( .A1(n19295), .A2(n19705), .ZN(n19231) );
  NOR2_X1 U16618 ( .A1(n19684), .A2(n19231), .ZN(n13370) );
  NOR2_X1 U16619 ( .A1(n19356), .A2(n19268), .ZN(n13409) );
  INV_X1 U16620 ( .A(n13409), .ZN(n13377) );
  AOI21_X1 U16621 ( .B1(n11969), .B2(n13377), .A(n19733), .ZN(n13369) );
  NOR2_X1 U16622 ( .A1(n13370), .A2(n13369), .ZN(n13412) );
  OAI21_X1 U16623 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n13371), .ZN(n19732) );
  INV_X1 U16624 ( .A(n19732), .ZN(n13373) );
  INV_X1 U16625 ( .A(n19711), .ZN(n13372) );
  NAND2_X1 U16626 ( .A1(n13373), .A2(n13372), .ZN(n13374) );
  NAND2_X1 U16627 ( .A1(n16064), .A2(n19516), .ZN(n19528) );
  NAND2_X1 U16628 ( .A1(n19298), .A2(n19472), .ZN(n13378) );
  OAI21_X1 U16629 ( .B1(n12007), .B2(n19733), .A(n19731), .ZN(n13376) );
  AOI22_X1 U16630 ( .A1(n13378), .A2(n19231), .B1(n13377), .B2(n13376), .ZN(
        n13379) );
  NAND2_X1 U16631 ( .A1(n13379), .A2(n19516), .ZN(n13404) );
  AOI22_X1 U16632 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n13406), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n13405), .ZN(n19484) );
  INV_X1 U16633 ( .A(n19484), .ZN(n19560) );
  AOI22_X1 U16634 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13404), .B1(
        n19290), .B2(n19560), .ZN(n13385) );
  INV_X1 U16635 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16313) );
  INV_X1 U16636 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18091) );
  OAI22_X2 U16637 ( .A1(n16313), .A2(n13403), .B1(n18091), .B2(n13402), .ZN(
        n19561) );
  NOR2_X2 U16638 ( .A1(n13383), .A2(n13407), .ZN(n19558) );
  AOI22_X1 U16639 ( .A1(n19251), .A2(n19561), .B1(n13409), .B2(n19558), .ZN(
        n13384) );
  OAI211_X1 U16640 ( .C1(n13412), .C2(n19528), .A(n13385), .B(n13384), .ZN(
        P2_U3090) );
  INV_X1 U16641 ( .A(n19588), .ZN(n19549) );
  AOI22_X1 U16642 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n13406), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n13405), .ZN(n19505) );
  INV_X1 U16643 ( .A(n19505), .ZN(n19590) );
  AOI22_X1 U16644 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13404), .B1(
        n19290), .B2(n19590), .ZN(n13388) );
  INV_X1 U16645 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16304) );
  INV_X1 U16646 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18116) );
  OAI22_X2 U16647 ( .A1(n16304), .A2(n13403), .B1(n18116), .B2(n13402), .ZN(
        n19592) );
  NOR2_X2 U16648 ( .A1(n13386), .A2(n13407), .ZN(n19586) );
  AOI22_X1 U16649 ( .A1(n19251), .A2(n19592), .B1(n13409), .B2(n19586), .ZN(
        n13387) );
  OAI211_X1 U16650 ( .C1(n13412), .C2(n19549), .A(n13388), .B(n13387), .ZN(
        P2_U3095) );
  INV_X1 U16651 ( .A(n19573), .ZN(n19540) );
  AOI22_X1 U16652 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n13406), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n13405), .ZN(n19495) );
  INV_X1 U16653 ( .A(n19495), .ZN(n19574) );
  AOI22_X1 U16654 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n13404), .B1(
        n19251), .B2(n19574), .ZN(n13391) );
  INV_X1 U16655 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16323) );
  INV_X1 U16656 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18106) );
  OAI22_X2 U16657 ( .A1(n16323), .A2(n13403), .B1(n18106), .B2(n13402), .ZN(
        n19575) );
  NOR2_X2 U16658 ( .A1(n13389), .A2(n13407), .ZN(n19572) );
  AOI22_X1 U16659 ( .A1(n19290), .A2(n19575), .B1(n13409), .B2(n19572), .ZN(
        n13390) );
  OAI211_X1 U16660 ( .C1(n13412), .C2(n19540), .A(n13391), .B(n13390), .ZN(
        P2_U3093) );
  INV_X1 U16661 ( .A(n19552), .ZN(n19525) );
  AOI22_X1 U16662 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n13406), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n13405), .ZN(n19481) );
  INV_X1 U16663 ( .A(n19481), .ZN(n19553) );
  AOI22_X1 U16664 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13404), .B1(
        n19290), .B2(n19553), .ZN(n13393) );
  INV_X1 U16665 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16315) );
  INV_X1 U16666 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18086) );
  OAI22_X2 U16667 ( .A1(n16315), .A2(n13403), .B1(n18086), .B2(n13402), .ZN(
        n19554) );
  AOI22_X1 U16668 ( .A1(n19251), .A2(n19554), .B1(n13409), .B2(n19551), .ZN(
        n13392) );
  OAI211_X1 U16669 ( .C1(n13412), .C2(n19525), .A(n13393), .B(n13392), .ZN(
        P2_U3089) );
  NAND2_X1 U16670 ( .A1(n16058), .A2(n19516), .ZN(n19537) );
  AOI22_X1 U16671 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n13406), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n13405), .ZN(n19491) );
  AOI22_X1 U16672 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13404), .B1(
        n19290), .B2(n19568), .ZN(n13395) );
  AOI22_X1 U16673 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13406), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n13405), .ZN(n19452) );
  NOR2_X2 U16674 ( .A1(n10375), .A2(n13407), .ZN(n19565) );
  AOI22_X1 U16675 ( .A1(n19251), .A2(n19567), .B1(n13409), .B2(n19565), .ZN(
        n13394) );
  OAI211_X1 U16676 ( .C1(n13412), .C2(n19537), .A(n13395), .B(n13394), .ZN(
        P2_U3092) );
  INV_X1 U16677 ( .A(n19485), .ZN(n19534) );
  INV_X1 U16678 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16327) );
  INV_X1 U16679 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18094) );
  OAI22_X2 U16680 ( .A1(n16327), .A2(n13403), .B1(n18094), .B2(n13402), .ZN(
        n19531) );
  AOI22_X1 U16681 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13404), .B1(
        n19290), .B2(n19531), .ZN(n13397) );
  INV_X1 U16682 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16311) );
  INV_X1 U16683 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n20933) );
  AOI22_X1 U16684 ( .A1(n19251), .A2(n19530), .B1(n13409), .B2(n19529), .ZN(
        n13396) );
  OAI211_X1 U16685 ( .C1(n13412), .C2(n19534), .A(n13397), .B(n13396), .ZN(
        P2_U3091) );
  INV_X1 U16686 ( .A(n19467), .ZN(n19522) );
  INV_X1 U16687 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16333) );
  INV_X1 U16688 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18077) );
  OAI22_X2 U16689 ( .A1(n16333), .A2(n13403), .B1(n18077), .B2(n13402), .ZN(
        n19519) );
  AOI22_X1 U16690 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13404), .B1(
        n19290), .B2(n19519), .ZN(n13401) );
  AOI22_X1 U16691 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n13405), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n13406), .ZN(n19478) );
  INV_X1 U16692 ( .A(n19478), .ZN(n19512) );
  AND2_X1 U16693 ( .A1(n13399), .A2(n13398), .ZN(n19511) );
  AOI22_X1 U16694 ( .A1(n19251), .A2(n19512), .B1(n19511), .B2(n13409), .ZN(
        n13400) );
  OAI211_X1 U16695 ( .C1(n13412), .C2(n19522), .A(n13401), .B(n13400), .ZN(
        P2_U3088) );
  NAND2_X1 U16696 ( .A1(n16051), .A2(n19516), .ZN(n19543) );
  INV_X1 U16697 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16305) );
  INV_X1 U16698 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18110) );
  OAI22_X2 U16699 ( .A1(n16305), .A2(n13403), .B1(n18110), .B2(n13402), .ZN(
        n19582) );
  AOI22_X1 U16700 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13404), .B1(
        n19251), .B2(n19582), .ZN(n13411) );
  AOI22_X1 U16701 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n13406), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n13405), .ZN(n19498) );
  INV_X1 U16702 ( .A(n19498), .ZN(n19581) );
  NOR2_X2 U16703 ( .A1(n13408), .A2(n13407), .ZN(n19579) );
  AOI22_X1 U16704 ( .A1(n19290), .A2(n19581), .B1(n13409), .B2(n19579), .ZN(
        n13410) );
  OAI211_X1 U16705 ( .C1(n13412), .C2(n19543), .A(n13411), .B(n13410), .ZN(
        P2_U3094) );
  INV_X1 U16706 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13420) );
  AND2_X1 U16707 ( .A1(n13414), .A2(n13413), .ZN(n13417) );
  NAND2_X1 U16708 ( .A1(n13123), .A2(n13415), .ZN(n13560) );
  OAI211_X1 U16709 ( .C1(n13417), .C2(n13416), .A(n13560), .B(n14945), .ZN(
        n13419) );
  NAND2_X1 U16710 ( .A1(n15398), .A2(n14890), .ZN(n13418) );
  OAI211_X1 U16711 ( .C1(n14890), .C2(n13420), .A(n13419), .B(n13418), .ZN(
        P2_U2874) );
  INV_X1 U16712 ( .A(n18917), .ZN(n18887) );
  OAI22_X1 U16713 ( .A1(n18887), .A2(n13421), .B1(n15466), .B2(n18916), .ZN(
        n13424) );
  OAI22_X1 U16714 ( .A1(n13422), .A2(n18931), .B1(n19620), .B2(n18918), .ZN(
        n13423) );
  AOI211_X1 U16715 ( .C1(n18901), .C2(n13425), .A(n13424), .B(n13423), .ZN(
        n13426) );
  OAI21_X1 U16716 ( .B1(n13427), .B2(n18878), .A(n13426), .ZN(n13431) );
  NOR2_X1 U16717 ( .A1(n18891), .A2(n13428), .ZN(n13435) );
  OAI21_X1 U16718 ( .B1(n18937), .B2(n13429), .A(n13435), .ZN(n13526) );
  OAI22_X1 U16719 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18930), .B1(
        n13526), .B2(n18883), .ZN(n13430) );
  AOI211_X1 U16720 ( .C1(n18933), .C2(n19076), .A(n13431), .B(n13430), .ZN(
        n13432) );
  INV_X1 U16721 ( .A(n13432), .ZN(P2_U2854) );
  INV_X1 U16722 ( .A(n13434), .ZN(n13436) );
  INV_X1 U16723 ( .A(n13435), .ZN(n13433) );
  AOI221_X1 U16724 ( .B1(n13436), .B2(n13435), .C1(n13434), .C2(n13433), .A(
        n18883), .ZN(n13437) );
  INV_X1 U16725 ( .A(n13437), .ZN(n13443) );
  AOI22_X1 U16726 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n18917), .B1(n13438), .B2(
        n18901), .ZN(n13440) );
  AOI22_X1 U16727 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18906), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n18829), .ZN(n13439) );
  OAI211_X1 U16728 ( .C1(n19692), .C2(n18916), .A(n13440), .B(n13439), .ZN(
        n13441) );
  AOI21_X1 U16729 ( .B1(n11900), .B2(n18927), .A(n13441), .ZN(n13442) );
  OAI211_X1 U16730 ( .C1(n13554), .C2(n13444), .A(n13443), .B(n13442), .ZN(
        P2_U2853) );
  INV_X1 U16731 ( .A(n19208), .ZN(n19679) );
  NAND2_X1 U16732 ( .A1(n12319), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19390) );
  INV_X1 U16733 ( .A(n19390), .ZN(n13445) );
  AND2_X1 U16734 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n13445), .ZN(
        n13452) );
  AOI21_X1 U16735 ( .B1(n19471), .B2(n19679), .A(n13452), .ZN(n13450) );
  NAND2_X1 U16736 ( .A1(n19294), .A2(n13445), .ZN(n13448) );
  NAND2_X1 U16737 ( .A1(n13448), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13446) );
  NOR2_X1 U16738 ( .A1(n13447), .A2(n13446), .ZN(n13454) );
  INV_X1 U16739 ( .A(n13448), .ZN(n19427) );
  OAI21_X1 U16740 ( .B1(n19427), .B2(n19731), .A(n19516), .ZN(n13449) );
  INV_X1 U16741 ( .A(n19430), .ZN(n13461) );
  INV_X1 U16742 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U16743 ( .A1(n19460), .A2(n19531), .B1(n19429), .B2(n19530), .ZN(
        n13456) );
  AOI21_X1 U16744 ( .B1(n19731), .B2(n13452), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13453) );
  NOR2_X1 U16745 ( .A1(n13454), .A2(n13453), .ZN(n19428) );
  AOI22_X1 U16746 ( .A1(n19428), .A2(n19485), .B1(n19529), .B2(n19427), .ZN(
        n13455) );
  OAI211_X1 U16747 ( .C1(n13461), .C2(n13457), .A(n13456), .B(n13455), .ZN(
        P2_U3139) );
  INV_X1 U16748 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13460) );
  AOI22_X1 U16749 ( .A1(n19460), .A2(n19519), .B1(n19429), .B2(n19512), .ZN(
        n13459) );
  AOI22_X1 U16750 ( .A1(n19428), .A2(n19467), .B1(n19511), .B2(n19427), .ZN(
        n13458) );
  OAI211_X1 U16751 ( .C1(n13461), .C2(n13460), .A(n13459), .B(n13458), .ZN(
        P2_U3136) );
  NOR2_X1 U16752 ( .A1(n18891), .A2(n13462), .ZN(n13463) );
  XNOR2_X1 U16753 ( .A(n13463), .B(n16093), .ZN(n13473) );
  AOI22_X1 U16754 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18906), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n18917), .ZN(n13464) );
  OAI21_X1 U16755 ( .B1(n13465), .B2(n18925), .A(n13464), .ZN(n13472) );
  AOI21_X1 U16756 ( .B1(n18829), .B2(P2_REIP_REG_12__SCAN_IN), .A(n15058), 
        .ZN(n13470) );
  AOI21_X1 U16757 ( .B1(n13468), .B2(n13467), .A(n13466), .ZN(n18946) );
  NAND2_X1 U16758 ( .A1(n18922), .A2(n18946), .ZN(n13469) );
  OAI211_X1 U16759 ( .C1(n15412), .C2(n18878), .A(n13470), .B(n13469), .ZN(
        n13471) );
  AOI211_X1 U16760 ( .C1(n13473), .C2(n18912), .A(n13472), .B(n13471), .ZN(
        n13474) );
  INV_X1 U16761 ( .A(n13474), .ZN(P2_U2843) );
  XNOR2_X1 U16762 ( .A(n13475), .B(n13690), .ZN(n13476) );
  XNOR2_X1 U16763 ( .A(n13477), .B(n13476), .ZN(n19043) );
  INV_X1 U16764 ( .A(n19043), .ZN(n13488) );
  XNOR2_X1 U16765 ( .A(n13478), .B(n9742), .ZN(n19041) );
  NOR2_X1 U16766 ( .A1(n19046), .A2(n16188), .ZN(n13486) );
  INV_X1 U16767 ( .A(n13725), .ZN(n13479) );
  NAND2_X1 U16768 ( .A1(n13479), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13689) );
  NOR2_X1 U16769 ( .A1(n19075), .A2(n13480), .ZN(n19054) );
  NOR2_X1 U16770 ( .A1(n19054), .A2(n13481), .ZN(n13726) );
  OAI21_X1 U16771 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16209), .A(
        n13726), .ZN(n13694) );
  NOR2_X1 U16772 ( .A1(n19625), .A2(n18900), .ZN(n13482) );
  AOI21_X1 U16773 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13694), .A(
        n13482), .ZN(n13484) );
  NAND2_X1 U16774 ( .A1(n16200), .A2(n13556), .ZN(n13483) );
  OAI211_X1 U16775 ( .C1(n13689), .C2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13484), .B(n13483), .ZN(n13485) );
  AOI211_X1 U16776 ( .C1(n19041), .C2(n19065), .A(n13486), .B(n13485), .ZN(
        n13487) );
  OAI21_X1 U16777 ( .B1(n13488), .B2(n16189), .A(n13487), .ZN(P2_U3042) );
  NAND2_X1 U16778 ( .A1(n13490), .A2(n13489), .ZN(n13493) );
  XNOR2_X1 U16779 ( .A(n13491), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13492) );
  XNOR2_X1 U16780 ( .A(n13493), .B(n13492), .ZN(n16148) );
  MUX2_X1 U16781 ( .A(n13725), .B(n13726), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13496) );
  OAI22_X1 U16782 ( .A1(n19686), .A2(n19070), .B1(n10675), .B2(n18900), .ZN(
        n13494) );
  INV_X1 U16783 ( .A(n13494), .ZN(n13495) );
  OAI211_X1 U16784 ( .C1(n16188), .C2(n16146), .A(n13496), .B(n13495), .ZN(
        n13499) );
  OR2_X1 U16785 ( .A1(n10242), .A2(n13497), .ZN(n16144) );
  AND3_X1 U16786 ( .A1(n16144), .A2(n19056), .A3(n16143), .ZN(n13498) );
  AOI211_X1 U16787 ( .C1(n16148), .C2(n19065), .A(n13499), .B(n13498), .ZN(
        n13500) );
  INV_X1 U16788 ( .A(n13500), .ZN(P2_U3043) );
  OR2_X1 U16789 ( .A1(n13502), .A2(n13501), .ZN(n13503) );
  NAND2_X1 U16790 ( .A1(n13503), .A2(n13353), .ZN(n16107) );
  INV_X1 U16791 ( .A(n16107), .ZN(n18857) );
  NOR2_X1 U16792 ( .A1(n14890), .A2(n10499), .ZN(n13508) );
  AOI211_X1 U16793 ( .C1(n13506), .C2(n13505), .A(n14961), .B(n13504), .ZN(
        n13507) );
  AOI211_X1 U16794 ( .C1(n18857), .C2(n14890), .A(n13508), .B(n13507), .ZN(
        n13509) );
  INV_X1 U16795 ( .A(n13509), .ZN(P2_U2877) );
  AND2_X1 U16796 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19296), .ZN(
        n13514) );
  AOI21_X1 U16797 ( .B1(n19471), .B2(n19303), .A(n13514), .ZN(n13513) );
  NAND2_X1 U16798 ( .A1(n19080), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13510) );
  INV_X1 U16799 ( .A(n19080), .ZN(n19587) );
  OAI21_X1 U16800 ( .B1(n19587), .B2(n19731), .A(n19516), .ZN(n13512) );
  NOR3_X2 U16801 ( .A1(n13513), .A2(n13516), .A3(n13512), .ZN(n19597) );
  INV_X1 U16802 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13520) );
  AOI21_X1 U16803 ( .B1(n19731), .B2(n13514), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13515) );
  NOR2_X1 U16804 ( .A1(n13516), .A2(n13515), .ZN(n19589) );
  INV_X1 U16805 ( .A(n19511), .ZN(n19118) );
  AOI22_X1 U16806 ( .A1(n19591), .A2(n19519), .B1(n19593), .B2(n19512), .ZN(
        n13517) );
  OAI21_X1 U16807 ( .B1(n19118), .B2(n19080), .A(n13517), .ZN(n13518) );
  AOI21_X1 U16808 ( .B1(n19589), .B2(n19467), .A(n13518), .ZN(n13519) );
  OAI21_X1 U16809 ( .B1(n19597), .B2(n13520), .A(n13519), .ZN(P2_U3168) );
  INV_X1 U16810 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13524) );
  INV_X1 U16811 ( .A(n19529), .ZN(n19135) );
  AOI22_X1 U16812 ( .A1(n19591), .A2(n19531), .B1(n19593), .B2(n19530), .ZN(
        n13521) );
  OAI21_X1 U16813 ( .B1(n19135), .B2(n19080), .A(n13521), .ZN(n13522) );
  AOI21_X1 U16814 ( .B1(n19589), .B2(n19485), .A(n13522), .ZN(n13523) );
  OAI21_X1 U16815 ( .B1(n19597), .B2(n13524), .A(n13523), .ZN(P2_U3171) );
  OAI222_X1 U16816 ( .A1(n16155), .A2(n18964), .B1(n18992), .B2(n13525), .C1(
        n12672), .C2(n18966), .ZN(P2_U2904) );
  OAI21_X1 U16817 ( .B1(n9642), .B2(n13527), .A(n13526), .ZN(n13573) );
  INV_X1 U16818 ( .A(n13573), .ZN(n13531) );
  OAI22_X1 U16819 ( .A1(n9642), .A2(n16202), .B1(n18937), .B2(n18891), .ZN(
        n15473) );
  INV_X1 U16820 ( .A(n15473), .ZN(n13529) );
  NOR2_X1 U16821 ( .A1(n13529), .A2(n13528), .ZN(n13572) );
  AOI222_X1 U16822 ( .A1(n13531), .A2(n13572), .B1(n19076), .B2(n16215), .C1(
        n13530), .C2(n13574), .ZN(n13533) );
  NAND2_X1 U16823 ( .A1(n15477), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13532) );
  OAI21_X1 U16824 ( .B1(n13533), .B2(n15477), .A(n13532), .ZN(P2_U3600) );
  OR2_X1 U16825 ( .A1(n13588), .A2(n13534), .ZN(n13579) );
  NAND2_X1 U16826 ( .A1(n13588), .A2(n13534), .ZN(n13535) );
  INV_X1 U16827 ( .A(n19790), .ZN(n13552) );
  OAI222_X1 U16828 ( .A1(n13552), .A2(n14507), .B1(n13536), .B2(n14505), .C1(
        n14504), .C2(n20042), .ZN(P1_U2897) );
  INV_X1 U16829 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13551) );
  INV_X1 U16830 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19872) );
  NAND2_X1 U16831 ( .A1(n14155), .A2(n19872), .ZN(n13539) );
  NAND2_X1 U16832 ( .A1(n14161), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13537) );
  NAND2_X1 U16833 ( .A1(n13539), .A2(n13538), .ZN(n19816) );
  MUX2_X1 U16834 ( .A(n14163), .B(n14158), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n13540) );
  INV_X1 U16835 ( .A(n13540), .ZN(n13543) );
  NAND2_X1 U16836 ( .A1(n14158), .A2(n14168), .ZN(n13758) );
  NAND2_X1 U16837 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14168), .ZN(
        n13541) );
  AND2_X1 U16838 ( .A1(n13758), .A2(n13541), .ZN(n13542) );
  NAND2_X1 U16839 ( .A1(n13543), .A2(n13542), .ZN(n15976) );
  INV_X1 U16840 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20895) );
  NAND2_X1 U16841 ( .A1(n14155), .A2(n20895), .ZN(n13546) );
  NAND2_X1 U16842 ( .A1(n14161), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13544) );
  AND2_X1 U16843 ( .A1(n13546), .A2(n13545), .ZN(n13591) );
  AND2_X1 U16844 ( .A1(n15976), .A2(n13591), .ZN(n13547) );
  MUX2_X1 U16845 ( .A(n14163), .B(n14158), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n13550) );
  NAND2_X1 U16846 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n14168), .ZN(
        n13548) );
  NAND2_X1 U16847 ( .A1(n13758), .A2(n13548), .ZN(n13549) );
  OAI21_X1 U16848 ( .B1(n9740), .B2(n9748), .A(n13585), .ZN(n19785) );
  OAI222_X1 U16849 ( .A1(n13552), .A2(n14460), .B1(n13551), .B2(n19873), .C1(
        n14448), .C2(n19785), .ZN(P1_U2865) );
  AOI21_X1 U16850 ( .B1(n19692), .B2(n13554), .A(n13553), .ZN(n18971) );
  XNOR2_X1 U16851 ( .A(n19683), .B(n19686), .ZN(n18970) );
  NOR2_X1 U16852 ( .A1(n18971), .A2(n18970), .ZN(n18969) );
  AOI21_X1 U16853 ( .B1(n19686), .B2(n19683), .A(n18969), .ZN(n13555) );
  NOR2_X1 U16854 ( .A1(n13555), .A2(n13556), .ZN(n18960) );
  XNOR2_X1 U16855 ( .A(n18960), .B(n18959), .ZN(n13559) );
  AOI22_X1 U16856 ( .A1(n18984), .A2(n13556), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n18983), .ZN(n13558) );
  NAND2_X1 U16857 ( .A1(n18958), .A2(n16058), .ZN(n13557) );
  OAI211_X1 U16858 ( .C1(n13559), .C2(n18978), .A(n13558), .B(n13557), .ZN(
        P2_U2915) );
  INV_X1 U16859 ( .A(n13560), .ZN(n13563) );
  OAI211_X1 U16860 ( .C1(n13563), .C2(n13562), .A(n14945), .B(n13561), .ZN(
        n13570) );
  INV_X1 U16861 ( .A(n13564), .ZN(n13568) );
  INV_X1 U16862 ( .A(n13565), .ZN(n13567) );
  AOI21_X1 U16863 ( .B1(n13568), .B2(n13567), .A(n13566), .ZN(n16165) );
  NAND2_X1 U16864 ( .A1(n16165), .A2(n14890), .ZN(n13569) );
  OAI211_X1 U16865 ( .C1(n14890), .C2(n13571), .A(n13570), .B(n13569), .ZN(
        P2_U2873) );
  AOI222_X1 U16866 ( .A1(n13575), .A2(n13574), .B1(n13573), .B2(n13572), .C1(
        n16215), .C2(n19697), .ZN(n13577) );
  NAND2_X1 U16867 ( .A1(n15477), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13576) );
  OAI21_X1 U16868 ( .B1(n13577), .B2(n15477), .A(n13576), .ZN(P2_U3599) );
  NOR2_X1 U16869 ( .A1(n13588), .A2(n13578), .ZN(n13595) );
  AOI21_X1 U16870 ( .B1(n13580), .B2(n13579), .A(n13595), .ZN(n13788) );
  INV_X1 U16871 ( .A(n13788), .ZN(n14380) );
  AOI22_X1 U16872 ( .A1(n14234), .A2(n14479), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15863), .ZN(n13581) );
  OAI21_X1 U16873 ( .B1(n14380), .B2(n14489), .A(n13581), .ZN(P1_U2896) );
  INV_X1 U16874 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14376) );
  NAND2_X1 U16875 ( .A1(n14155), .A2(n14376), .ZN(n13584) );
  NAND2_X1 U16876 ( .A1(n14161), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13582) );
  NAND2_X1 U16877 ( .A1(n13584), .A2(n13583), .ZN(n13586) );
  AOI21_X1 U16878 ( .B1(n13586), .B2(n13585), .A(n13603), .ZN(n15966) );
  AOI22_X1 U16879 ( .A1(n15966), .A2(n19869), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14458), .ZN(n13587) );
  OAI21_X1 U16880 ( .B1(n14380), .B2(n14460), .A(n13587), .ZN(P1_U2864) );
  AOI21_X1 U16881 ( .B1(n13590), .B2(n13589), .A(n10112), .ZN(n19798) );
  INV_X1 U16882 ( .A(n19798), .ZN(n13597) );
  AOI21_X1 U16883 ( .B1(n19814), .B2(n15976), .A(n13591), .ZN(n13592) );
  NOR2_X1 U16884 ( .A1(n9740), .A2(n13592), .ZN(n19794) );
  AOI22_X1 U16885 ( .A1(n19794), .A2(n19869), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14458), .ZN(n13593) );
  OAI21_X1 U16886 ( .B1(n13597), .B2(n14460), .A(n13593), .ZN(P1_U2866) );
  OAI21_X1 U16887 ( .B1(n13595), .B2(n13594), .A(n11478), .ZN(n19777) );
  MUX2_X1 U16888 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n19996), .Z(
        n19905) );
  AOI22_X1 U16889 ( .A1(n14234), .A2(n19905), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15863), .ZN(n13596) );
  OAI21_X1 U16890 ( .B1(n19777), .B2(n14507), .A(n13596), .ZN(P1_U2895) );
  OAI222_X1 U16891 ( .A1(n13597), .A2(n14507), .B1(n14505), .B2(n11411), .C1(
        n14504), .C2(n20034), .ZN(P1_U2898) );
  INV_X1 U16892 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13605) );
  MUX2_X1 U16893 ( .A(n14163), .B(n14158), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n13598) );
  INV_X1 U16894 ( .A(n13598), .ZN(n13601) );
  NAND2_X1 U16895 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n14168), .ZN(
        n13599) );
  AND2_X1 U16896 ( .A1(n13758), .A2(n13599), .ZN(n13600) );
  NAND2_X1 U16897 ( .A1(n13601), .A2(n13600), .ZN(n13602) );
  NOR2_X1 U16898 ( .A1(n13603), .A2(n13602), .ZN(n13604) );
  OR2_X1 U16899 ( .A1(n13659), .A2(n13604), .ZN(n19773) );
  OAI222_X1 U16900 ( .A1(n19777), .A2(n14460), .B1(n13605), .B2(n19873), .C1(
        n14448), .C2(n19773), .ZN(P1_U2863) );
  XOR2_X1 U16901 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13607), .Z(
        n13608) );
  XNOR2_X1 U16902 ( .A(n13606), .B(n13608), .ZN(n14831) );
  INV_X1 U16903 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20674) );
  NOR2_X1 U16904 ( .A1(n15922), .A2(n20674), .ZN(n14829) );
  AOI21_X1 U16905 ( .B1(n19932), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n14829), .ZN(n13609) );
  OAI21_X1 U16906 ( .B1(n19943), .B2(n19805), .A(n13609), .ZN(n13610) );
  AOI21_X1 U16907 ( .B1(n19798), .B2(n19938), .A(n13610), .ZN(n13611) );
  OAI21_X1 U16908 ( .B1(n14831), .B2(n15902), .A(n13611), .ZN(P1_U2993) );
  NOR2_X1 U16909 ( .A1(n18891), .A2(n13612), .ZN(n13613) );
  XNOR2_X1 U16910 ( .A(n13613), .B(n16087), .ZN(n13614) );
  NAND2_X1 U16911 ( .A1(n13614), .A2(n18912), .ZN(n13625) );
  AOI21_X1 U16912 ( .B1(n13617), .B2(n13616), .A(n13615), .ZN(n18943) );
  NAND2_X1 U16913 ( .A1(n18922), .A2(n18943), .ZN(n13618) );
  OAI211_X1 U16914 ( .C1(n13619), .C2(n18918), .A(n13618), .B(n18900), .ZN(
        n13623) );
  AOI22_X1 U16915 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18906), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n18917), .ZN(n13620) );
  OAI21_X1 U16916 ( .B1(n13621), .B2(n18925), .A(n13620), .ZN(n13622) );
  AOI211_X1 U16917 ( .C1(n16165), .C2(n18927), .A(n13623), .B(n13622), .ZN(
        n13624) );
  NAND2_X1 U16918 ( .A1(n13625), .A2(n13624), .ZN(P2_U2841) );
  INV_X1 U16919 ( .A(n13627), .ZN(n13628) );
  OAI21_X1 U16920 ( .B1(n13626), .B2(n13629), .A(n13628), .ZN(n13665) );
  XNOR2_X1 U16921 ( .A(n13644), .B(n13643), .ZN(n18833) );
  INV_X1 U16922 ( .A(n18833), .ZN(n13632) );
  INV_X1 U16923 ( .A(n16065), .ZN(n15013) );
  OAI22_X1 U16924 ( .A1(n15013), .A2(n18993), .B1(n18966), .B2(n13630), .ZN(
        n13631) );
  AOI21_X1 U16925 ( .B1(n18984), .B2(n13632), .A(n13631), .ZN(n13634) );
  AOI22_X1 U16926 ( .A1(n18940), .A2(BUF2_REG_16__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n13633) );
  OAI211_X1 U16927 ( .C1(n13665), .C2(n18978), .A(n13634), .B(n13633), .ZN(
        P2_U2903) );
  NOR2_X1 U16928 ( .A1(n14890), .A2(n10871), .ZN(n13638) );
  AOI211_X1 U16929 ( .C1(n13636), .C2(n13561), .A(n14961), .B(n13626), .ZN(
        n13637) );
  AOI211_X1 U16930 ( .C1(n16159), .C2(n14890), .A(n13638), .B(n13637), .ZN(
        n13639) );
  INV_X1 U16931 ( .A(n13639), .ZN(P2_U2872) );
  OAI21_X1 U16932 ( .B1(n13627), .B2(n13641), .A(n13640), .ZN(n13709) );
  INV_X1 U16933 ( .A(n13642), .ZN(n13646) );
  NAND2_X1 U16934 ( .A1(n13644), .A2(n13643), .ZN(n13645) );
  NAND2_X1 U16935 ( .A1(n13646), .A2(n13645), .ZN(n13647) );
  NAND2_X1 U16936 ( .A1(n13647), .A2(n13855), .ZN(n15374) );
  INV_X1 U16937 ( .A(n15374), .ZN(n18822) );
  OAI22_X1 U16938 ( .A1(n15013), .A2(n18982), .B1(n18966), .B2(n13648), .ZN(
        n13649) );
  AOI21_X1 U16939 ( .B1(n18984), .B2(n18822), .A(n13649), .ZN(n13651) );
  AOI22_X1 U16940 ( .A1(n18940), .A2(BUF2_REG_17__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13650) );
  OAI211_X1 U16941 ( .C1(n13709), .C2(n18978), .A(n13651), .B(n13650), .ZN(
        P2_U2902) );
  NOR2_X1 U16942 ( .A1(n13654), .A2(n13653), .ZN(n13655) );
  INV_X1 U16943 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13660) );
  MUX2_X1 U16944 ( .A(n14155), .B(n14255), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13657) );
  NOR2_X1 U16945 ( .A1(n14180), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13656) );
  NOR2_X1 U16946 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  NAND2_X1 U16947 ( .A1(n13659), .A2(n13658), .ZN(n13769) );
  OAI21_X1 U16948 ( .B1(n13659), .B2(n13658), .A(n13769), .ZN(n15839) );
  OAI222_X1 U16949 ( .A1(n15843), .A2(n14460), .B1(n13660), .B2(n19873), .C1(
        n14448), .C2(n15839), .ZN(P1_U2862) );
  OAI21_X1 U16950 ( .B1(n13662), .B2(n13661), .A(n13705), .ZN(n18834) );
  MUX2_X1 U16951 ( .A(n13663), .B(n18834), .S(n14890), .Z(n13664) );
  OAI21_X1 U16952 ( .B1(n13665), .B2(n14961), .A(n13664), .ZN(P2_U2871) );
  NAND2_X1 U16953 ( .A1(n13667), .A2(n13666), .ZN(n13668) );
  NAND2_X1 U16954 ( .A1(n13669), .A2(n13668), .ZN(n15911) );
  INV_X1 U16955 ( .A(n15911), .ZN(n13680) );
  INV_X1 U16956 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14827) );
  NAND2_X1 U16957 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19949) );
  NOR2_X1 U16958 ( .A1(n15982), .A2(n19949), .ZN(n13670) );
  AOI21_X1 U16959 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19946) );
  NAND2_X1 U16960 ( .A1(n15943), .A2(n13034), .ZN(n19985) );
  NAND2_X1 U16961 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14185) );
  OAI22_X1 U16962 ( .A1(n14767), .A2(n19946), .B1(n19965), .B2(n14185), .ZN(
        n19953) );
  NAND2_X1 U16963 ( .A1(n13670), .A2(n19953), .ZN(n14826) );
  NOR2_X1 U16964 ( .A1(n14827), .A2(n14826), .ZN(n15972) );
  INV_X1 U16965 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13678) );
  NAND2_X1 U16966 ( .A1(n19944), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n15912) );
  OAI21_X1 U16967 ( .B1(n19785), .B2(n19981), .A(n15912), .ZN(n13677) );
  INV_X1 U16968 ( .A(n19965), .ZN(n13675) );
  NOR2_X1 U16969 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19949), .ZN(
        n15978) );
  INV_X1 U16970 ( .A(n13670), .ZN(n14184) );
  NOR2_X1 U16971 ( .A1(n19946), .A2(n14184), .ZN(n14187) );
  INV_X1 U16972 ( .A(n15938), .ZN(n14725) );
  NAND2_X1 U16973 ( .A1(n14725), .A2(n13034), .ZN(n13672) );
  INV_X1 U16974 ( .A(n19991), .ZN(n13671) );
  OAI21_X1 U16975 ( .B1(n14187), .B2(n14767), .A(n19977), .ZN(n14808) );
  NAND2_X1 U16976 ( .A1(n19961), .A2(n14185), .ZN(n19947) );
  INV_X1 U16977 ( .A(n19947), .ZN(n13673) );
  AOI211_X1 U16978 ( .C1(n19961), .C2(n19949), .A(n14808), .B(n13673), .ZN(
        n15983) );
  INV_X1 U16979 ( .A(n15983), .ZN(n13674) );
  AOI211_X1 U16980 ( .C1(n13675), .C2(n15978), .A(n14827), .B(n13674), .ZN(
        n15968) );
  NAND2_X1 U16981 ( .A1(n14805), .A2(n14767), .ZN(n19986) );
  INV_X1 U16982 ( .A(n19986), .ZN(n14768) );
  NAND2_X1 U16983 ( .A1(n14768), .A2(n19977), .ZN(n14201) );
  INV_X1 U16984 ( .A(n14201), .ZN(n15967) );
  NOR3_X1 U16985 ( .A1(n15968), .A2(n15967), .A3(n13678), .ZN(n13676) );
  AOI211_X1 U16986 ( .C1(n15972), .C2(n13678), .A(n13677), .B(n13676), .ZN(
        n13679) );
  OAI21_X1 U16987 ( .B1(n13680), .B2(n14832), .A(n13679), .ZN(P1_U3024) );
  XNOR2_X1 U16988 ( .A(n13681), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13682) );
  XNOR2_X1 U16989 ( .A(n13683), .B(n13682), .ZN(n16135) );
  OAI21_X1 U16990 ( .B1(n13687), .B2(n13685), .A(n13684), .ZN(n13686) );
  OAI21_X1 U16991 ( .B1(n13688), .B2(n13687), .A(n13686), .ZN(n16132) );
  NOR2_X1 U16992 ( .A1(n10703), .A2(n18885), .ZN(n13693) );
  AOI221_X1 U16993 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13691), .C2(n13690), .A(
        n13689), .ZN(n13692) );
  AOI211_X1 U16994 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n13694), .A(
        n13693), .B(n13692), .ZN(n13701) );
  OAI21_X1 U16995 ( .B1(n13697), .B2(n13696), .A(n13695), .ZN(n18963) );
  INV_X1 U16996 ( .A(n18911), .ZN(n13698) );
  OAI22_X1 U16997 ( .A1(n18963), .A2(n19070), .B1(n16188), .B2(n13698), .ZN(
        n13699) );
  INV_X1 U16998 ( .A(n13699), .ZN(n13700) );
  OAI211_X1 U16999 ( .C1(n16132), .C2(n16189), .A(n13701), .B(n13700), .ZN(
        n13702) );
  INV_X1 U17000 ( .A(n13702), .ZN(n13703) );
  OAI21_X1 U17001 ( .B1(n16135), .B2(n16204), .A(n13703), .ZN(P2_U3041) );
  NAND2_X1 U17002 ( .A1(n12964), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13708) );
  NAND2_X1 U17003 ( .A1(n13705), .A2(n13704), .ZN(n13706) );
  NAND2_X1 U17004 ( .A1(n18823), .A2(n14890), .ZN(n13707) );
  OAI211_X1 U17005 ( .C1(n13709), .C2(n14961), .A(n13708), .B(n13707), .ZN(
        P2_U2870) );
  AND2_X1 U17006 ( .A1(n13710), .A2(n13711), .ZN(n14430) );
  OAI21_X1 U17007 ( .B1(n14430), .B2(n13712), .A(n14622), .ZN(n15783) );
  NOR3_X1 U17008 ( .A1(n15863), .A2(n19996), .A3(n13713), .ZN(n13714) );
  AOI22_X1 U17009 ( .A1(n15866), .A2(DATAI_17_), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n15863), .ZN(n13720) );
  NOR3_X1 U17010 ( .A1(n15863), .A2(n14461), .A3(n20029), .ZN(n13715) );
  NAND2_X1 U17011 ( .A1(n13716), .A2(n19996), .ZN(n13717) );
  AOI22_X1 U17012 ( .A1(n15865), .A2(n13718), .B1(n14493), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13719) );
  OAI211_X1 U17013 ( .C1(n15783), .C2(n14507), .A(n13720), .B(n13719), .ZN(
        P1_U2887) );
  XNOR2_X1 U17014 ( .A(n13721), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13740) );
  XOR2_X1 U17015 ( .A(n13722), .B(n13723), .Z(n13738) );
  NOR2_X1 U17016 ( .A1(n13725), .A2(n13724), .ZN(n13730) );
  OAI21_X1 U17017 ( .B1(n16209), .B2(n13727), .A(n13726), .ZN(n16185) );
  INV_X1 U17018 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19628) );
  NOR2_X1 U17019 ( .A1(n19628), .A2(n18885), .ZN(n13728) );
  AOI221_X1 U17020 ( .B1(n13730), .B2(n13729), .C1(n16185), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n13728), .ZN(n13731) );
  INV_X1 U17021 ( .A(n13731), .ZN(n13733) );
  OAI22_X1 U17022 ( .A1(n18899), .A2(n19070), .B1(n16188), .B2(n18894), .ZN(
        n13732) );
  AOI211_X1 U17023 ( .C1(n13738), .C2(n19065), .A(n13733), .B(n13732), .ZN(
        n13734) );
  OAI21_X1 U17024 ( .B1(n13740), .B2(n16189), .A(n13734), .ZN(P2_U3040) );
  OAI22_X1 U17025 ( .A1(n19628), .A2(n18900), .B1(n19052), .B2(n18892), .ZN(
        n13735) );
  AOI21_X1 U17026 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19039), .A(
        n13735), .ZN(n13736) );
  OAI21_X1 U17027 ( .B1(n18894), .B2(n19047), .A(n13736), .ZN(n13737) );
  AOI21_X1 U17028 ( .B1(n13738), .B2(n19040), .A(n13737), .ZN(n13739) );
  OAI21_X1 U17029 ( .B1(n13740), .B2(n16133), .A(n13739), .ZN(P2_U3008) );
  INV_X1 U17030 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n13763) );
  MUX2_X1 U17031 ( .A(n14163), .B(n14158), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13743) );
  NAND2_X1 U17032 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14168), .ZN(
        n13741) );
  NAND2_X1 U17033 ( .A1(n13758), .A2(n13741), .ZN(n13742) );
  NOR2_X1 U17034 ( .A1(n13743), .A2(n13742), .ZN(n13768) );
  INV_X1 U17035 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15819) );
  NAND2_X1 U17036 ( .A1(n14155), .A2(n15819), .ZN(n13746) );
  NAND2_X1 U17037 ( .A1(n14161), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13744) );
  NAND2_X1 U17038 ( .A1(n13746), .A2(n13745), .ZN(n14457) );
  INV_X1 U17039 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U17040 ( .A1(n14163), .A2(n14447), .ZN(n13750) );
  INV_X1 U17041 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13747) );
  OAI211_X1 U17042 ( .C1(n14168), .C2(P1_EBX_REG_13__SCAN_IN), .A(n13748), .B(
        n14161), .ZN(n13749) );
  NAND2_X1 U17043 ( .A1(n13750), .A2(n13749), .ZN(n14360) );
  MUX2_X1 U17044 ( .A(n14155), .B(n14255), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13752) );
  NOR2_X1 U17045 ( .A1(n14180), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13751) );
  NOR2_X1 U17046 ( .A1(n13752), .A2(n13751), .ZN(n13803) );
  INV_X1 U17047 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15802) );
  NAND2_X1 U17048 ( .A1(n14163), .A2(n15802), .ZN(n13755) );
  OAI211_X1 U17049 ( .C1(n14168), .C2(P1_EBX_REG_15__SCAN_IN), .A(n13753), .B(
        n14161), .ZN(n13754) );
  MUX2_X1 U17050 ( .A(n14166), .B(n14161), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13756) );
  OAI21_X1 U17051 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n14180), .A(
        n13756), .ZN(n14432) );
  MUX2_X1 U17052 ( .A(n14163), .B(n14158), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13760) );
  NAND2_X1 U17053 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n14168), .ZN(
        n13757) );
  NAND2_X1 U17054 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  NOR2_X1 U17055 ( .A1(n13760), .A2(n13759), .ZN(n13761) );
  AND2_X1 U17056 ( .A1(n14434), .A2(n13761), .ZN(n13762) );
  OR2_X1 U17057 ( .A1(n13762), .A2(n14771), .ZN(n15793) );
  OAI222_X1 U17058 ( .A1(n14460), .A2(n15783), .B1(n19873), .B2(n13763), .C1(
        n15793), .C2(n14448), .ZN(P1_U2855) );
  NAND2_X1 U17059 ( .A1(n13764), .A2(n13766), .ZN(n14356) );
  XNOR2_X1 U17060 ( .A(n14356), .B(n14354), .ZN(n15904) );
  INV_X1 U17061 ( .A(n15904), .ZN(n13772) );
  MUX2_X1 U17062 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n19996), .Z(
        n19909) );
  AOI22_X1 U17063 ( .A1(n14234), .A2(n19909), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15863), .ZN(n13767) );
  OAI21_X1 U17064 ( .B1(n13772), .B2(n14489), .A(n13767), .ZN(P1_U2893) );
  INV_X1 U17065 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n13771) );
  NAND2_X1 U17066 ( .A1(n13769), .A2(n13768), .ZN(n13770) );
  NAND2_X1 U17067 ( .A1(n14456), .A2(n13770), .ZN(n15829) );
  OAI222_X1 U17068 ( .A1(n13772), .A2(n14460), .B1(n13771), .B2(n19873), .C1(
        n14448), .C2(n15829), .ZN(P1_U2861) );
  NAND2_X1 U17069 ( .A1(n13774), .A2(n13773), .ZN(n13775) );
  NAND2_X1 U17070 ( .A1(n13863), .A2(n13775), .ZN(n15365) );
  INV_X1 U17071 ( .A(n13776), .ZN(n13777) );
  AOI21_X1 U17072 ( .B1(n13778), .B2(n13640), .A(n13777), .ZN(n16067) );
  NAND2_X1 U17073 ( .A1(n16067), .A2(n14945), .ZN(n13780) );
  NAND2_X1 U17074 ( .A1(n12964), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13779) );
  OAI211_X1 U17075 ( .C1(n15365), .C2(n12964), .A(n13780), .B(n13779), .ZN(
        P2_U2869) );
  INV_X1 U17076 ( .A(n13781), .ZN(n13782) );
  NOR2_X1 U17077 ( .A1(n13783), .A2(n13782), .ZN(n13784) );
  XNOR2_X1 U17078 ( .A(n13785), .B(n13784), .ZN(n15970) );
  INV_X1 U17079 ( .A(n15970), .ZN(n13790) );
  NAND2_X1 U17080 ( .A1(n19944), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15964) );
  NAND2_X1 U17081 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13786) );
  OAI211_X1 U17082 ( .C1(n19943), .C2(n14373), .A(n15964), .B(n13786), .ZN(
        n13787) );
  AOI21_X1 U17083 ( .B1(n13788), .B2(n19938), .A(n13787), .ZN(n13789) );
  OAI21_X1 U17084 ( .B1(n13790), .B2(n15902), .A(n13789), .ZN(P1_U2991) );
  AOI21_X1 U17085 ( .B1(n13791), .B2(n13776), .A(n9655), .ZN(n13792) );
  INV_X1 U17086 ( .A(n13792), .ZN(n13867) );
  AND2_X1 U17087 ( .A1(n13857), .A2(n13793), .ZN(n13794) );
  OR2_X1 U17088 ( .A1(n13794), .A2(n15320), .ZN(n18814) );
  INV_X1 U17089 ( .A(n18814), .ZN(n15347) );
  OAI22_X1 U17090 ( .A1(n15013), .A2(n18975), .B1(n18966), .B2(n13795), .ZN(
        n13796) );
  AOI21_X1 U17091 ( .B1(n18984), .B2(n15347), .A(n13796), .ZN(n13798) );
  AOI22_X1 U17092 ( .A1(n18940), .A2(BUF2_REG_19__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n13797) );
  OAI211_X1 U17093 ( .C1(n13867), .C2(n18978), .A(n13798), .B(n13797), .ZN(
        P2_U2900) );
  NAND2_X1 U17094 ( .A1(n13710), .A2(n13799), .ZN(n14357) );
  INV_X1 U17095 ( .A(n14438), .ZN(n13800) );
  AOI21_X1 U17096 ( .B1(n13801), .B2(n14357), .A(n13800), .ZN(n15893) );
  INV_X1 U17097 ( .A(n15893), .ZN(n13806) );
  MUX2_X1 U17098 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n19996), .Z(
        n19915) );
  AOI22_X1 U17099 ( .A1(n14234), .A2(n19915), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15863), .ZN(n13802) );
  OAI21_X1 U17100 ( .B1(n13806), .B2(n14507), .A(n13802), .ZN(P1_U2890) );
  INV_X1 U17101 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13805) );
  OR2_X1 U17102 ( .A1(n14362), .A2(n13803), .ZN(n13804) );
  NAND2_X1 U17103 ( .A1(n14442), .A2(n13804), .ZN(n15812) );
  OAI222_X1 U17104 ( .A1(n13806), .A2(n14460), .B1(n13805), .B2(n19873), .C1(
        n14448), .C2(n15812), .ZN(P1_U2858) );
  XNOR2_X1 U17105 ( .A(n14628), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13808) );
  XNOR2_X1 U17106 ( .A(n13807), .B(n13808), .ZN(n13820) );
  NAND3_X1 U17107 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n15972), .ZN(n15956) );
  INV_X1 U17108 ( .A(n15956), .ZN(n13814) );
  NAND2_X1 U17109 ( .A1(n19944), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n13816) );
  OAI21_X1 U17110 ( .B1(n19773), .B2(n19981), .A(n13816), .ZN(n13813) );
  INV_X1 U17111 ( .A(n14808), .ZN(n13811) );
  NAND2_X1 U17112 ( .A1(n14187), .A2(n19947), .ZN(n13809) );
  NAND3_X1 U17113 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14186) );
  OAI21_X1 U17114 ( .B1(n13809), .B2(n14186), .A(n19986), .ZN(n13810) );
  AND2_X1 U17115 ( .A1(n13811), .A2(n13810), .ZN(n15963) );
  NOR2_X1 U17116 ( .A1(n15963), .A2(n15957), .ZN(n13812) );
  AOI211_X1 U17117 ( .C1(n13814), .C2(n15957), .A(n13813), .B(n13812), .ZN(
        n13815) );
  OAI21_X1 U17118 ( .B1(n13820), .B2(n14832), .A(n13815), .ZN(P1_U3022) );
  OAI21_X1 U17119 ( .B1(n15914), .B2(n19774), .A(n13816), .ZN(n13818) );
  NOR2_X1 U17120 ( .A1(n19777), .A2(n19998), .ZN(n13817) );
  AOI211_X1 U17121 ( .C1(n15909), .C2(n19778), .A(n13818), .B(n13817), .ZN(
        n13819) );
  OAI21_X1 U17122 ( .B1(n13820), .B2(n15902), .A(n13819), .ZN(P1_U2990) );
  XNOR2_X1 U17123 ( .A(n13821), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13848) );
  NAND2_X1 U17124 ( .A1(n13822), .A2(n13823), .ZN(n16123) );
  NAND2_X1 U17125 ( .A1(n16122), .A2(n16120), .ZN(n13824) );
  XNOR2_X1 U17126 ( .A(n16123), .B(n13824), .ZN(n13845) );
  OAI22_X1 U17127 ( .A1(n16151), .A2(n13825), .B1(n19630), .B2(n18900), .ZN(
        n13826) );
  AOI21_X1 U17128 ( .B1(n16142), .B2(n18873), .A(n13826), .ZN(n13827) );
  OAI21_X1 U17129 ( .B1(n18877), .B2(n19047), .A(n13827), .ZN(n13828) );
  AOI21_X1 U17130 ( .B1(n13845), .B2(n19040), .A(n13828), .ZN(n13829) );
  OAI21_X1 U17131 ( .B1(n13848), .B2(n16133), .A(n13829), .ZN(P2_U3007) );
  OAI21_X1 U17132 ( .B1(n13830), .B2(n13832), .A(n14943), .ZN(n14953) );
  OR2_X1 U17133 ( .A1(n15322), .A2(n13833), .ZN(n13835) );
  AND2_X1 U17134 ( .A1(n13835), .A2(n13834), .ZN(n18778) );
  OAI22_X1 U17135 ( .A1(n15013), .A2(n13837), .B1(n18966), .B2(n13836), .ZN(
        n13838) );
  AOI21_X1 U17136 ( .B1(n18984), .B2(n18778), .A(n13838), .ZN(n13840) );
  AOI22_X1 U17137 ( .A1(n18940), .A2(BUF2_REG_21__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n13839) );
  OAI211_X1 U17138 ( .C1(n14953), .C2(n18978), .A(n13840), .B(n13839), .ZN(
        P2_U2898) );
  INV_X1 U17139 ( .A(n18877), .ZN(n13841) );
  AOI22_X1 U17140 ( .A1(n13841), .A2(n19067), .B1(n15058), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n13843) );
  NAND2_X1 U17141 ( .A1(n16194), .A2(n20776), .ZN(n13842) );
  OAI211_X1 U17142 ( .C1(n18879), .C2(n19070), .A(n13843), .B(n13842), .ZN(
        n13844) );
  AOI21_X1 U17143 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16185), .A(
        n13844), .ZN(n13847) );
  NAND2_X1 U17144 ( .A1(n13845), .A2(n19065), .ZN(n13846) );
  OAI211_X1 U17145 ( .C1(n13848), .C2(n16189), .A(n13847), .B(n13846), .ZN(
        P2_U3039) );
  AOI211_X1 U17146 ( .C1(n15149), .C2(n13850), .A(n13849), .B(n18883), .ZN(
        n13861) );
  AOI21_X1 U17147 ( .B1(P2_REIP_REG_18__SCAN_IN), .B2(n18829), .A(n15058), 
        .ZN(n13852) );
  AOI22_X1 U17148 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18906), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n18917), .ZN(n13851) );
  OAI211_X1 U17149 ( .C1(n13853), .C2(n18925), .A(n13852), .B(n13851), .ZN(
        n13860) );
  NAND2_X1 U17150 ( .A1(n13855), .A2(n13854), .ZN(n13856) );
  AND2_X1 U17151 ( .A1(n13857), .A2(n13856), .ZN(n16066) );
  INV_X1 U17152 ( .A(n16066), .ZN(n13858) );
  OAI22_X1 U17153 ( .A1(n15365), .A2(n18878), .B1(n18916), .B2(n13858), .ZN(
        n13859) );
  OR3_X1 U17154 ( .A1(n13861), .A2(n13860), .A3(n13859), .ZN(P2_U2837) );
  AND2_X1 U17155 ( .A1(n13863), .A2(n13862), .ZN(n13864) );
  OR2_X1 U17156 ( .A1(n13864), .A2(n14958), .ZN(n18806) );
  MUX2_X1 U17157 ( .A(n18806), .B(n13865), .S(n14946), .Z(n13866) );
  OAI21_X1 U17158 ( .B1(n13867), .B2(n14961), .A(n13866), .ZN(P2_U2868) );
  INV_X2 U17159 ( .A(n9678), .ZN(n17040) );
  AOI22_X1 U17160 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17040), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13872) );
  NOR2_X1 U17161 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U17162 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13871) );
  NAND4_X1 U17163 ( .A1(n18695), .A2(n18702), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U17164 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13870) );
  AOI22_X1 U17165 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13869) );
  NAND4_X1 U17166 ( .A1(n13872), .A2(n13871), .A3(n13870), .A4(n13869), .ZN(
        n13883) );
  AOI22_X1 U17167 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13881) );
  CLKBUF_X3 U17168 ( .A(n13884), .Z(n17060) );
  AOI22_X1 U17169 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13880) );
  CLKBUF_X3 U17170 ( .A(n13937), .Z(n17061) );
  AOI22_X1 U17171 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13879) );
  NOR2_X2 U17172 ( .A1(n18695), .A2(n13877), .ZN(n15537) );
  INV_X2 U17173 ( .A(n15487), .ZN(n17046) );
  AOI22_X1 U17174 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13878) );
  NAND4_X1 U17175 ( .A1(n13881), .A2(n13880), .A3(n13879), .A4(n13878), .ZN(
        n13882) );
  NOR2_X1 U17176 ( .A1(n13883), .A2(n13882), .ZN(n17196) );
  INV_X1 U17177 ( .A(n17196), .ZN(n13987) );
  NAND3_X1 U17178 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .ZN(n13983) );
  CLKBUF_X3 U17179 ( .A(n15572), .Z(n17045) );
  AOI22_X1 U17180 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U17181 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17182 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13893) );
  NOR2_X1 U17183 ( .A1(n16903), .A2(n20943), .ZN(n13891) );
  INV_X2 U17184 ( .A(n9678), .ZN(n16999) );
  AOI22_X1 U17185 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13889) );
  AOI22_X1 U17186 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U17187 ( .A1(n15509), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13887) );
  AOI22_X1 U17188 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16976), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13886) );
  NAND4_X1 U17189 ( .A1(n13889), .A2(n13888), .A3(n13887), .A4(n13886), .ZN(
        n13890) );
  AOI211_X2 U17190 ( .C1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .C2(n17044), .A(
        n13891), .B(n13890), .ZN(n13892) );
  AOI22_X1 U17191 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U17192 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U17193 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17194 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13896) );
  NAND4_X1 U17195 ( .A1(n13899), .A2(n13898), .A3(n13897), .A4(n13896), .ZN(
        n13905) );
  AOI22_X1 U17196 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U17197 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U17198 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17199 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13900) );
  NAND4_X1 U17200 ( .A1(n13903), .A2(n13902), .A3(n13901), .A4(n13900), .ZN(
        n13904) );
  AOI22_X1 U17201 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17040), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17202 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U17203 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U17204 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13906) );
  NAND4_X1 U17205 ( .A1(n13909), .A2(n13908), .A3(n13907), .A4(n13906), .ZN(
        n13916) );
  AOI22_X1 U17206 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13914) );
  AOI22_X1 U17207 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17208 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U17209 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13911) );
  NAND4_X1 U17210 ( .A1(n13914), .A2(n13913), .A3(n13912), .A4(n13911), .ZN(
        n13915) );
  AOI22_X1 U17211 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U17212 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13925) );
  INV_X4 U17213 ( .A(n15558), .ZN(n15509) );
  AOI22_X1 U17214 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13917) );
  OAI21_X1 U17215 ( .B1(n15487), .B2(n20929), .A(n13917), .ZN(n13923) );
  AOI22_X1 U17216 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13921) );
  AOI22_X1 U17217 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13920) );
  AOI22_X1 U17218 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13919) );
  AOI22_X1 U17219 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13918) );
  NAND4_X1 U17220 ( .A1(n13921), .A2(n13920), .A3(n13919), .A4(n13918), .ZN(
        n13922) );
  AOI211_X1 U17221 ( .C1(n15537), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n13923), .B(n13922), .ZN(n13924) );
  NAND3_X1 U17222 ( .A1(n13926), .A2(n13925), .A3(n13924), .ZN(n18104) );
  NAND2_X1 U17223 ( .A1(n18109), .A2(n17118), .ZN(n14009) );
  AOI22_X1 U17224 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U17225 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13935) );
  AOI22_X1 U17226 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13927) );
  OAI21_X1 U17227 ( .B1(n13939), .B2(n20848), .A(n13927), .ZN(n13933) );
  AOI22_X1 U17228 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U17229 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13930) );
  AOI22_X1 U17230 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U17231 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13928) );
  NAND4_X1 U17232 ( .A1(n13931), .A2(n13930), .A3(n13929), .A4(n13928), .ZN(
        n13932) );
  AOI211_X1 U17233 ( .C1(n16976), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n13933), .B(n13932), .ZN(n13934) );
  NAND3_X1 U17234 ( .A1(n13936), .A2(n13935), .A3(n13934), .ZN(n18096) );
  AOI22_X1 U17235 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U17236 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U17237 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13938) );
  OAI21_X1 U17238 ( .B1(n13939), .B2(n20899), .A(n13938), .ZN(n13945) );
  AOI22_X1 U17239 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13943) );
  AOI22_X1 U17240 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13942) );
  AOI22_X1 U17241 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13941) );
  AOI22_X1 U17242 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13940) );
  NAND4_X1 U17243 ( .A1(n13943), .A2(n13942), .A3(n13941), .A4(n13940), .ZN(
        n13944) );
  AOI211_X1 U17244 ( .C1(n15537), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n13945), .B(n13944), .ZN(n13946) );
  NAND3_X1 U17245 ( .A1(n13948), .A2(n13947), .A3(n13946), .ZN(n18089) );
  INV_X1 U17246 ( .A(n18089), .ZN(n15626) );
  NAND2_X1 U17247 ( .A1(n13989), .A2(n15626), .ZN(n18520) );
  AOI22_X1 U17248 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13958) );
  AOI22_X1 U17249 ( .A1(n15509), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U17250 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13949) );
  OAI21_X1 U17251 ( .B1(n13971), .B2(n17091), .A(n13949), .ZN(n13955) );
  AOI22_X1 U17252 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U17253 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U17254 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U17255 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13950) );
  NAND4_X1 U17256 ( .A1(n13953), .A2(n13952), .A3(n13951), .A4(n13950), .ZN(
        n13954) );
  AOI211_X1 U17257 ( .C1(n9638), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n13955), .B(n13954), .ZN(n13956) );
  NAND3_X1 U17258 ( .A1(n13958), .A2(n13957), .A3(n13956), .ZN(n18099) );
  NAND2_X1 U17259 ( .A1(n14013), .A2(n17197), .ZN(n13969) );
  AOI22_X1 U17260 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18541), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18702), .ZN(n14002) );
  AND2_X1 U17261 ( .A1(n14002), .A2(n14003), .ZN(n13959) );
  AOI22_X1 U17262 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18561), .B2(n18695), .ZN(
        n13963) );
  NOR2_X1 U17263 ( .A1(n13964), .A2(n13963), .ZN(n13960) );
  AOI22_X1 U17264 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18572), .B1(
        n13961), .B2(n18685), .ZN(n13967) );
  NAND2_X1 U17265 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18572), .ZN(
        n13962) );
  OAI22_X1 U17266 ( .A1(n13967), .A2(n18562), .B1(n13965), .B2(n13962), .ZN(
        n13968) );
  AOI211_X1 U17267 ( .C1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n18708), .A(
        n14003), .B(n13968), .ZN(n15623) );
  XNOR2_X1 U17268 ( .A(n13964), .B(n13963), .ZN(n15625) );
  OAI21_X1 U17269 ( .B1(n13968), .B2(n15625), .A(n14006), .ZN(n14004) );
  AOI21_X1 U17270 ( .B1(n14002), .B2(n15623), .A(n14004), .ZN(n18510) );
  NOR2_X1 U17271 ( .A1(n18109), .A2(n14013), .ZN(n13988) );
  NOR2_X2 U17272 ( .A1(n17197), .A2(n13989), .ZN(n15635) );
  AND3_X1 U17273 ( .A1(n13988), .A2(n15635), .A3(n15629), .ZN(n15641) );
  NAND2_X1 U17274 ( .A1(n18510), .A2(n15641), .ZN(n14020) );
  NAND2_X1 U17275 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18688), .ZN(n16423) );
  INV_X1 U17276 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U17277 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13970) );
  OAI21_X1 U17278 ( .B1(n13971), .B2(n17102), .A(n13970), .ZN(n13977) );
  AOI22_X1 U17279 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U17280 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17281 ( .A1(n13884), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13973) );
  AOI22_X1 U17282 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13972) );
  NAND4_X1 U17283 ( .A1(n13975), .A2(n13974), .A3(n13973), .A4(n13972), .ZN(
        n13976) );
  NAND2_X1 U17284 ( .A1(n18727), .A2(n18085), .ZN(n16223) );
  NOR3_X4 U17285 ( .A1(n16752), .A2(n13981), .A3(n16223), .ZN(n17107) );
  INV_X1 U17286 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17108) );
  INV_X1 U17287 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17103) );
  NOR2_X1 U17288 ( .A1(n17108), .A2(n17103), .ZN(n17097) );
  NAND2_X1 U17289 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17097), .ZN(n17035) );
  INV_X1 U17290 ( .A(n17035), .ZN(n13982) );
  INV_X1 U17291 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16715) );
  INV_X1 U17292 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17079) );
  INV_X1 U17293 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16738) );
  INV_X1 U17294 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17078) );
  NOR4_X1 U17295 ( .A1(n16715), .A2(n17079), .A3(n16738), .A4(n17078), .ZN(
        n17038) );
  NAND4_X1 U17296 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17107), .A3(n13982), .A4(
        n17038), .ZN(n17075) );
  NAND2_X1 U17297 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17034), .ZN(n17020) );
  NAND2_X1 U17298 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17007), .ZN(n14023) );
  INV_X1 U17299 ( .A(n14023), .ZN(n16968) );
  NAND2_X1 U17300 ( .A1(n17197), .A2(n16968), .ZN(n16967) );
  NOR2_X1 U17301 ( .A1(n13983), .A2(n16967), .ZN(n16964) );
  INV_X1 U17302 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20777) );
  INV_X1 U17303 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16637) );
  NOR2_X1 U17304 ( .A1(n20777), .A2(n16637), .ZN(n13984) );
  AOI21_X1 U17305 ( .B1(n16968), .B2(n13984), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n13985) );
  NOR2_X1 U17306 ( .A1(n16964), .A2(n13985), .ZN(n13986) );
  MUX2_X1 U17307 ( .A(n13987), .B(n13986), .S(n17101), .Z(P3_U2688) );
  NAND2_X1 U17308 ( .A1(n18688), .A2(n18679), .ZN(n18683) );
  NAND2_X1 U17309 ( .A1(n18109), .A2(n18104), .ZN(n13991) );
  NOR4_X1 U17310 ( .A1(n18099), .A2(n18096), .A3(n13998), .A4(n13991), .ZN(
        n14000) );
  INV_X1 U17311 ( .A(n13988), .ZN(n18521) );
  NAND2_X1 U17312 ( .A1(n15626), .A2(n18521), .ZN(n13995) );
  NAND2_X1 U17313 ( .A1(n18104), .A2(n17115), .ZN(n18536) );
  NOR2_X1 U17314 ( .A1(n16752), .A2(n18085), .ZN(n15639) );
  OAI21_X1 U17315 ( .B1(n17197), .B2(n15742), .A(n15639), .ZN(n14016) );
  OAI21_X1 U17316 ( .B1(n15629), .B2(n13999), .A(n14016), .ZN(n13996) );
  NAND2_X1 U17317 ( .A1(n16752), .A2(n14009), .ZN(n13994) );
  AOI22_X1 U17318 ( .A1(n14013), .A2(n15742), .B1(n13989), .B2(n13998), .ZN(
        n13993) );
  OR2_X1 U17319 ( .A1(n18089), .A2(n15640), .ZN(n14010) );
  AOI21_X1 U17320 ( .B1(n18114), .B2(n13991), .A(n14013), .ZN(n13990) );
  AOI21_X1 U17321 ( .B1(n13991), .B2(n14010), .A(n13990), .ZN(n13992) );
  OAI211_X1 U17322 ( .C1(n13995), .C2(n13994), .A(n13993), .B(n13992), .ZN(
        n14015) );
  AOI21_X1 U17323 ( .B1(n18096), .B2(n13996), .A(n14015), .ZN(n15636) );
  NAND2_X1 U17324 ( .A1(n14000), .A2(n15636), .ZN(n15634) );
  NOR2_X1 U17325 ( .A1(n13998), .A2(n13997), .ZN(n14001) );
  NAND2_X1 U17326 ( .A1(n14000), .A2(n18089), .ZN(n14014) );
  NAND2_X1 U17327 ( .A1(n17302), .A2(n14014), .ZN(n16405) );
  NAND2_X1 U17328 ( .A1(n15640), .A2(n16405), .ZN(n14008) );
  INV_X1 U17329 ( .A(n18553), .ZN(n18529) );
  OAI21_X1 U17330 ( .B1(n18529), .B2(n18685), .A(n18572), .ZN(n15479) );
  NAND2_X1 U17331 ( .A1(n18530), .A2(n15479), .ZN(n18518) );
  NOR2_X1 U17332 ( .A1(n18683), .A2(n18518), .ZN(n14022) );
  XNOR2_X1 U17333 ( .A(n14003), .B(n14002), .ZN(n14007) );
  INV_X1 U17334 ( .A(n14004), .ZN(n14005) );
  NAND2_X1 U17335 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18733) );
  NOR2_X1 U17336 ( .A1(n16222), .A2(n18599), .ZN(n14018) );
  INV_X1 U17337 ( .A(n17302), .ZN(n17305) );
  NAND2_X1 U17338 ( .A1(n18732), .A2(n17305), .ZN(n18576) );
  NAND2_X2 U17339 ( .A1(n18669), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18672) );
  OAI211_X1 U17340 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18607), .B(n18672), .ZN(n18730) );
  AOI21_X1 U17341 ( .B1(n14008), .B2(n18576), .A(n18730), .ZN(n17265) );
  INV_X1 U17342 ( .A(n14009), .ZN(n14011) );
  NOR2_X1 U17343 ( .A1(n14011), .A2(n14010), .ZN(n14012) );
  OAI211_X1 U17344 ( .C1(n14013), .C2(n15742), .A(n15635), .B(n14012), .ZN(
        n15621) );
  OAI21_X1 U17345 ( .B1(n15621), .B2(n14015), .A(n14014), .ZN(n14017) );
  NAND2_X1 U17346 ( .A1(n14017), .A2(n14016), .ZN(n15622) );
  AOI21_X1 U17347 ( .B1(n14018), .B2(n17265), .A(n15622), .ZN(n14021) );
  NOR2_X1 U17348 ( .A1(n18732), .A2(n17302), .ZN(n14019) );
  NAND3_X1 U17349 ( .A1(n14021), .A2(n15741), .A3(n14020), .ZN(n18558) );
  INV_X1 U17350 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18584) );
  NAND2_X1 U17351 ( .A1(n18584), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18081) );
  NOR3_X1 U17352 ( .A1(n18688), .A2(n18584), .A3(n18742), .ZN(n18588) );
  NAND2_X1 U17353 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18588), .ZN(n15480) );
  OAI211_X1 U17354 ( .C1(n18581), .C2(n18535), .A(n18081), .B(n15480), .ZN(
        n18706) );
  INV_X1 U17355 ( .A(n18706), .ZN(n18709) );
  MUX2_X1 U17356 ( .A(n14022), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18709), .Z(P3_U3284) );
  AND2_X1 U17357 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16848) );
  NAND2_X1 U17358 ( .A1(n17197), .A2(n17107), .ZN(n17109) );
  INV_X1 U17359 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16508) );
  INV_X1 U17360 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16529) );
  INV_X1 U17361 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16583) );
  INV_X1 U17362 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16593) );
  NAND4_X1 U17363 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(P3_EBX_REG_13__SCAN_IN), .ZN(n16929)
         );
  NAND2_X1 U17364 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n9643), .ZN(n16927) );
  INV_X1 U17365 ( .A(n16927), .ZN(n16902) );
  NOR2_X1 U17366 ( .A1(n18114), .A2(n16900), .ZN(n16876) );
  NAND2_X1 U17367 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16876), .ZN(n16870) );
  NAND2_X1 U17368 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16875), .ZN(n16860) );
  NAND2_X1 U17369 ( .A1(n17101), .A2(n16858), .ZN(n14024) );
  OAI21_X1 U17370 ( .B1(n16848), .B2(n17109), .A(n14024), .ZN(n16849) );
  AOI22_X1 U17371 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14028) );
  AOI22_X1 U17372 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14027) );
  AOI22_X1 U17373 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14026) );
  AOI22_X1 U17374 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14025) );
  NAND4_X1 U17375 ( .A1(n14028), .A2(n14027), .A3(n14026), .A4(n14025), .ZN(
        n14034) );
  AOI22_X1 U17376 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14032) );
  AOI22_X1 U17377 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14031) );
  AOI22_X1 U17378 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U17379 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14029) );
  NAND4_X1 U17380 ( .A1(n14032), .A2(n14031), .A3(n14030), .A4(n14029), .ZN(
        n14033) );
  NOR2_X1 U17381 ( .A1(n14034), .A2(n14033), .ZN(n14098) );
  AOI22_X1 U17382 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14038) );
  AOI22_X1 U17383 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14037) );
  AOI22_X1 U17384 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14036) );
  AOI22_X1 U17385 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14035) );
  NAND4_X1 U17386 ( .A1(n14038), .A2(n14037), .A3(n14036), .A4(n14035), .ZN(
        n14044) );
  AOI22_X1 U17387 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14042) );
  AOI22_X1 U17388 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U17389 ( .A1(n13937), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U17390 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14039) );
  NAND4_X1 U17391 ( .A1(n14042), .A2(n14041), .A3(n14040), .A4(n14039), .ZN(
        n14043) );
  NOR2_X1 U17392 ( .A1(n14044), .A2(n14043), .ZN(n16856) );
  AOI22_X1 U17393 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17040), .ZN(n14048) );
  AOI22_X1 U17394 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14047) );
  AOI22_X1 U17395 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n15536), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15537), .ZN(n14046) );
  AOI22_X1 U17396 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16976), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13910), .ZN(n14045) );
  NAND4_X1 U17397 ( .A1(n14048), .A2(n14047), .A3(n14046), .A4(n14045), .ZN(
        n14054) );
  AOI22_X1 U17398 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U17399 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17067), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n13884), .ZN(n14051) );
  AOI22_X1 U17400 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17061), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17045), .ZN(n14050) );
  AOI22_X1 U17401 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17046), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14049) );
  NAND4_X1 U17402 ( .A1(n14052), .A2(n14051), .A3(n14050), .A4(n14049), .ZN(
        n14053) );
  NOR2_X1 U17403 ( .A1(n14054), .A2(n14053), .ZN(n16866) );
  AOI22_X1 U17404 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14065) );
  INV_X1 U17405 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15571) );
  AOI22_X1 U17406 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14057) );
  AOI22_X1 U17407 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14056) );
  OAI211_X1 U17408 ( .C1(n16832), .C2(n15571), .A(n14057), .B(n14056), .ZN(
        n14063) );
  AOI22_X1 U17409 ( .A1(n13937), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U17410 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14060) );
  AOI22_X1 U17411 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U17412 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14058) );
  NAND4_X1 U17413 ( .A1(n14061), .A2(n14060), .A3(n14059), .A4(n14058), .ZN(
        n14062) );
  AOI211_X1 U17414 ( .C1(n15502), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n14063), .B(n14062), .ZN(n14064) );
  NAND2_X1 U17415 ( .A1(n14065), .A2(n14064), .ZN(n16872) );
  AOI22_X1 U17416 ( .A1(n15509), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14075) );
  AOI22_X1 U17417 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14074) );
  AOI22_X1 U17418 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14066) );
  OAI21_X1 U17419 ( .B1(n9678), .B2(n20943), .A(n14066), .ZN(n14072) );
  AOI22_X1 U17420 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14070) );
  AOI22_X1 U17421 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14069) );
  AOI22_X1 U17422 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U17423 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14067) );
  NAND4_X1 U17424 ( .A1(n14070), .A2(n14069), .A3(n14068), .A4(n14067), .ZN(
        n14071) );
  AOI211_X1 U17425 ( .C1(n17066), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n14072), .B(n14071), .ZN(n14073) );
  NAND3_X1 U17426 ( .A1(n14075), .A2(n14074), .A3(n14073), .ZN(n16873) );
  NAND2_X1 U17427 ( .A1(n16872), .A2(n16873), .ZN(n16871) );
  NOR2_X1 U17428 ( .A1(n16866), .A2(n16871), .ZN(n16865) );
  AOI22_X1 U17429 ( .A1(n13937), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U17430 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14085) );
  AOI22_X1 U17431 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14084) );
  AND2_X1 U17432 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n14082) );
  AOI22_X1 U17433 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U17434 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14079) );
  AOI22_X1 U17435 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U17436 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14077) );
  NAND4_X1 U17437 ( .A1(n14080), .A2(n14079), .A3(n14078), .A4(n14077), .ZN(
        n14081) );
  AOI211_X1 U17438 ( .C1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .C2(n9633), .A(
        n14082), .B(n14081), .ZN(n14083) );
  NAND4_X1 U17439 ( .A1(n14086), .A2(n14085), .A3(n14084), .A4(n14083), .ZN(
        n16862) );
  NAND2_X1 U17440 ( .A1(n16865), .A2(n16862), .ZN(n16861) );
  NOR2_X1 U17441 ( .A1(n16856), .A2(n16861), .ZN(n16855) );
  AOI22_X1 U17442 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14097) );
  AOI22_X1 U17443 ( .A1(n13937), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U17444 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14088) );
  OAI211_X1 U17445 ( .C1(n16832), .C2(n17091), .A(n14089), .B(n14088), .ZN(
        n14095) );
  AOI22_X1 U17446 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14093) );
  AOI22_X1 U17447 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U17448 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U17449 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14090) );
  NAND4_X1 U17450 ( .A1(n14093), .A2(n14092), .A3(n14091), .A4(n14090), .ZN(
        n14094) );
  AOI211_X1 U17451 ( .C1(n15536), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n14095), .B(n14094), .ZN(n14096) );
  NAND2_X1 U17452 ( .A1(n14097), .A2(n14096), .ZN(n16852) );
  NAND2_X1 U17453 ( .A1(n16855), .A2(n16852), .ZN(n16851) );
  NOR2_X1 U17454 ( .A1(n14098), .A2(n16851), .ZN(n16846) );
  AOI21_X1 U17455 ( .B1(n14098), .B2(n16851), .A(n16846), .ZN(n17128) );
  AOI22_X1 U17456 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16849), .B1(n17128), 
        .B2(n17105), .ZN(n14102) );
  INV_X1 U17457 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14100) );
  INV_X1 U17458 ( .A(n16858), .ZN(n14099) );
  NAND3_X1 U17459 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14100), .A3(n14099), 
        .ZN(n14101) );
  NAND2_X1 U17460 ( .A1(n14102), .A2(n14101), .ZN(P3_U2675) );
  XNOR2_X1 U17461 ( .A(n14628), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14103) );
  INV_X1 U17462 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20705) );
  OR2_X1 U17463 ( .A1(n15922), .A2(n20705), .ZN(n14660) );
  OAI21_X1 U17464 ( .B1(n15914), .B2(n14105), .A(n14660), .ZN(n14109) );
  NAND2_X2 U17465 ( .A1(n14260), .A2(n14107), .ZN(n14111) );
  NOR2_X1 U17466 ( .A1(n14111), .A2(n19998), .ZN(n14108) );
  OAI21_X1 U17467 ( .B1(n15902), .B2(n14666), .A(n14110), .ZN(P1_U2970) );
  INV_X1 U17468 ( .A(n20754), .ZN(n14114) );
  NOR2_X1 U17469 ( .A1(n20301), .A2(n15994), .ZN(n15716) );
  NAND2_X1 U17470 ( .A1(n15716), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14112) );
  OAI211_X1 U17471 ( .C1(n14114), .C2(n14113), .A(n14112), .B(n15922), .ZN(
        n14115) );
  INV_X1 U17472 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20689) );
  INV_X1 U17473 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20687) );
  INV_X1 U17474 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20684) );
  INV_X1 U17475 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20677) );
  INV_X1 U17476 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20669) );
  NAND4_X1 U17477 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19799)
         );
  NOR3_X1 U17478 ( .A1(n20669), .A2(n20674), .A3(n19799), .ZN(n19789) );
  NAND2_X1 U17479 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19789), .ZN(n14366) );
  NOR2_X1 U17480 ( .A1(n20677), .A2(n14366), .ZN(n14371) );
  NAND3_X1 U17481 ( .A1(n14371), .A2(P1_REIP_REG_10__SCAN_IN), .A3(
        P1_REIP_REG_9__SCAN_IN), .ZN(n15828) );
  NAND2_X1 U17482 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14368) );
  NOR2_X1 U17483 ( .A1(n15828), .A2(n14368), .ZN(n14359) );
  NAND3_X1 U17484 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n14359), .ZN(n15804) );
  NOR2_X1 U17485 ( .A1(n20684), .A2(n15804), .ZN(n15798) );
  NAND2_X1 U17486 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n15798), .ZN(n15771) );
  NOR2_X1 U17487 ( .A1(n20687), .A2(n15771), .ZN(n15770) );
  NAND2_X1 U17488 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15770), .ZN(n15764) );
  NOR2_X1 U17489 ( .A1(n20689), .A2(n15764), .ZN(n14346) );
  AND2_X1 U17490 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14117) );
  AND2_X1 U17491 ( .A1(n14346), .A2(n14117), .ZN(n14334) );
  AND2_X1 U17492 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14118) );
  NAND2_X1 U17493 ( .A1(n14334), .A2(n14118), .ZN(n14323) );
  NAND2_X1 U17494 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14119) );
  OR2_X1 U17495 ( .A1(n14323), .A2(n14119), .ZN(n14126) );
  NAND2_X1 U17496 ( .A1(n19827), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14124) );
  NAND2_X1 U17497 ( .A1(n20661), .A2(n20757), .ZN(n15709) );
  INV_X1 U17498 ( .A(n15709), .ZN(n14120) );
  OAI21_X1 U17499 ( .B1(n20014), .B2(n14121), .A(n14120), .ZN(n14132) );
  NOR2_X1 U17500 ( .A1(n14132), .A2(n14122), .ZN(n14123) );
  NAND2_X1 U17501 ( .A1(n19826), .A2(n19827), .ZN(n19801) );
  OAI21_X1 U17502 ( .B1(n14126), .B2(n14124), .A(n19801), .ZN(n14286) );
  NAND3_X1 U17503 ( .A1(n14286), .A2(P1_REIP_REG_28__SCAN_IN), .A3(
        P1_REIP_REG_27__SCAN_IN), .ZN(n14125) );
  NAND2_X1 U17504 ( .A1(n14125), .A2(n19801), .ZN(n14246) );
  INV_X1 U17505 ( .A(n14246), .ZN(n14274) );
  NOR2_X1 U17506 ( .A1(n14126), .A2(n19826), .ZN(n14297) );
  AND2_X1 U17507 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14127) );
  AND2_X1 U17508 ( .A1(n14297), .A2(n14127), .ZN(n14275) );
  NAND2_X1 U17509 ( .A1(n14275), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14263) );
  NOR2_X1 U17510 ( .A1(n14129), .A2(n14128), .ZN(n14130) );
  AOI22_X1 U17511 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19853), .B1(
        n19850), .B2(n14131), .ZN(n14136) );
  NOR2_X1 U17512 ( .A1(n12998), .A2(n20811), .ZN(n14171) );
  NAND2_X1 U17513 ( .A1(n14132), .A2(n9956), .ZN(n14133) );
  OR2_X1 U17514 ( .A1(n14171), .A2(n14133), .ZN(n14134) );
  NOR2_X2 U17515 ( .A1(n14173), .A2(n14134), .ZN(n19849) );
  NAND2_X1 U17516 ( .A1(n19849), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14135) );
  OAI211_X1 U17517 ( .C1(n14263), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14136), 
        .B(n14135), .ZN(n14175) );
  INV_X1 U17518 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15854) );
  NAND2_X1 U17519 ( .A1(n14155), .A2(n15854), .ZN(n14139) );
  NAND2_X1 U17520 ( .A1(n14161), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14137) );
  INV_X1 U17521 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14426) );
  NAND2_X1 U17522 ( .A1(n14163), .A2(n14426), .ZN(n14142) );
  OAI211_X1 U17523 ( .C1(n14168), .C2(P1_EBX_REG_19__SCAN_IN), .A(n14140), .B(
        n14161), .ZN(n14141) );
  NAND2_X1 U17524 ( .A1(n14142), .A2(n14141), .ZN(n14423) );
  INV_X1 U17525 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14419) );
  NAND2_X1 U17526 ( .A1(n14155), .A2(n14419), .ZN(n14145) );
  NAND2_X1 U17527 ( .A1(n14161), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14143) );
  INV_X1 U17528 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15753) );
  NAND2_X1 U17529 ( .A1(n14163), .A2(n15753), .ZN(n14148) );
  OAI211_X1 U17530 ( .C1(n14168), .C2(P1_EBX_REG_21__SCAN_IN), .A(n14146), .B(
        n14161), .ZN(n14147) );
  INV_X1 U17531 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15851) );
  NAND2_X1 U17532 ( .A1(n14155), .A2(n15851), .ZN(n14151) );
  NAND2_X1 U17533 ( .A1(n14161), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14149) );
  NAND2_X1 U17534 ( .A1(n14151), .A2(n14150), .ZN(n14722) );
  INV_X1 U17535 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14412) );
  NAND2_X1 U17536 ( .A1(n14163), .A2(n14412), .ZN(n14154) );
  OAI211_X1 U17537 ( .C1(n12998), .C2(P1_EBX_REG_23__SCAN_IN), .A(n14152), .B(
        n14161), .ZN(n14153) );
  NAND2_X1 U17538 ( .A1(n14154), .A2(n14153), .ZN(n14333) );
  MUX2_X1 U17539 ( .A(n14155), .B(n14255), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14157) );
  NOR2_X1 U17540 ( .A1(n14180), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14156) );
  NOR2_X1 U17541 ( .A1(n14157), .A2(n14156), .ZN(n14319) );
  MUX2_X1 U17542 ( .A(n14163), .B(n14158), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14160) );
  AND2_X1 U17543 ( .A1(n14168), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14159) );
  NOR2_X1 U17544 ( .A1(n14160), .A2(n14159), .ZN(n14305) );
  MUX2_X1 U17545 ( .A(n14166), .B(n14161), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14162) );
  OAI21_X1 U17546 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14180), .A(
        n14162), .ZN(n14295) );
  INV_X1 U17547 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14520) );
  INV_X1 U17548 ( .A(n14163), .ZN(n14169) );
  OAI21_X1 U17549 ( .B1(n14165), .B2(n14520), .A(n14164), .ZN(n14282) );
  MUX2_X1 U17550 ( .A(n14166), .B(n14161), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14167) );
  OAI21_X1 U17551 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14180), .A(
        n14167), .ZN(n14273) );
  OAI22_X1 U17552 ( .A1(n14180), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n14168), .ZN(n14253) );
  OAI22_X1 U17553 ( .A1(n14253), .A2(n14255), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14169), .ZN(n14170) );
  NAND2_X1 U17554 ( .A1(n14272), .A2(n14170), .ZN(n14256) );
  OAI21_X1 U17555 ( .B1(n14272), .B2(n14170), .A(n14256), .ZN(n14657) );
  NAND2_X1 U17556 ( .A1(n14171), .A2(n15709), .ZN(n14172) );
  NOR2_X1 U17557 ( .A1(n14657), .A2(n19865), .ZN(n14174) );
  AOI211_X1 U17558 ( .C1(n14274), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14175), 
        .B(n14174), .ZN(n14176) );
  OAI21_X1 U17559 ( .B1(n14111), .B2(n15842), .A(n14176), .ZN(P1_U2811) );
  AOI22_X1 U17560 ( .A1(n15866), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15863), .ZN(n14178) );
  MUX2_X1 U17561 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n19996), .Z(
        n19913) );
  AOI22_X1 U17562 ( .A1(n15865), .A2(n19913), .B1(BUF1_REG_29__SCAN_IN), .B2(
        n14493), .ZN(n14177) );
  OAI211_X1 U17563 ( .C1(n14111), .C2(n14489), .A(n14178), .B(n14177), .ZN(
        P1_U2875) );
  INV_X1 U17564 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14179) );
  OAI222_X1 U17565 ( .A1(n14460), .A2(n14111), .B1(n14179), .B2(n19873), .C1(
        n14657), .C2(n14448), .ZN(P1_U2843) );
  AOI22_X1 U17566 ( .A1(n14180), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12998), .ZN(n14181) );
  AOI22_X1 U17567 ( .A1(n14180), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12998), .ZN(n14257) );
  XNOR2_X1 U17568 ( .A(n14181), .B(n14257), .ZN(n14183) );
  OR2_X1 U17569 ( .A1(n14181), .A2(n14255), .ZN(n14182) );
  MUX2_X1 U17570 ( .A(n14183), .B(n14182), .S(n14256), .Z(n14403) );
  INV_X1 U17571 ( .A(n14403), .ZN(n14206) );
  NOR2_X1 U17572 ( .A1(n14185), .A2(n14184), .ZN(n14807) );
  NAND2_X1 U17573 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15958) );
  NOR2_X1 U17574 ( .A1(n14186), .A2(n15958), .ZN(n14806) );
  NAND2_X1 U17575 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14806), .ZN(
        n14810) );
  NOR2_X1 U17576 ( .A1(n14813), .A2(n14810), .ZN(n14194) );
  AND2_X1 U17577 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14194), .ZN(
        n14795) );
  NAND2_X1 U17578 ( .A1(n14807), .A2(n14795), .ZN(n14765) );
  INV_X1 U17579 ( .A(n14765), .ZN(n15944) );
  NAND2_X1 U17580 ( .A1(n15944), .A2(n13675), .ZN(n14703) );
  NAND2_X1 U17581 ( .A1(n14194), .A2(n14187), .ZN(n15941) );
  NOR2_X1 U17582 ( .A1(n14767), .A2(n15941), .ZN(n14724) );
  NAND2_X1 U17583 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14724), .ZN(
        n14188) );
  AND2_X1 U17584 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14730) );
  INV_X1 U17585 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14781) );
  NAND2_X1 U17586 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15925) );
  NOR2_X1 U17587 ( .A1(n14781), .A2(n15925), .ZN(n14774) );
  NAND3_X1 U17588 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n14774), .ZN(n14195) );
  INV_X1 U17589 ( .A(n14195), .ZN(n14189) );
  NAND3_X1 U17590 ( .A1(n14729), .A2(n14730), .A3(n14189), .ZN(n14190) );
  INV_X1 U17591 ( .A(n14518), .ZN(n14684) );
  NAND2_X1 U17592 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14191) );
  NOR2_X1 U17593 ( .A1(n14715), .A2(n14191), .ZN(n14667) );
  NAND2_X1 U17594 ( .A1(n14667), .A2(n14193), .ZN(n14661) );
  NAND3_X1 U17595 ( .A1(n14192), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14204) );
  INV_X1 U17596 ( .A(n14193), .ZN(n14200) );
  INV_X1 U17597 ( .A(n14687), .ZN(n14198) );
  NAND2_X1 U17598 ( .A1(n14807), .A2(n14194), .ZN(n15945) );
  OR2_X1 U17599 ( .A1(n13747), .A2(n14195), .ZN(n14756) );
  NOR2_X1 U17600 ( .A1(n15945), .A2(n14756), .ZN(n14726) );
  INV_X1 U17601 ( .A(n14767), .ZN(n19962) );
  OAI21_X1 U17602 ( .B1(n14756), .B2(n15941), .A(n19962), .ZN(n14196) );
  OAI211_X1 U17603 ( .C1(n14805), .C2(n14726), .A(n19977), .B(n14196), .ZN(
        n14758) );
  INV_X1 U17604 ( .A(n14729), .ZN(n14197) );
  OAI21_X1 U17605 ( .B1(n14758), .B2(n14197), .A(n14201), .ZN(n14738) );
  OAI21_X1 U17606 ( .B1(n14768), .B2(n14730), .A(n14738), .ZN(n14712) );
  AOI21_X1 U17607 ( .B1(n14198), .B2(n19986), .A(n14712), .ZN(n14685) );
  INV_X1 U17608 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14683) );
  OAI21_X1 U17609 ( .B1(n14683), .B2(n14686), .A(n19986), .ZN(n14199) );
  NAND2_X1 U17610 ( .A1(n14685), .A2(n14199), .ZN(n14680) );
  AOI21_X1 U17611 ( .B1(n14200), .B2(n19986), .A(n14680), .ZN(n14659) );
  OAI211_X1 U17612 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14768), .A(
        n14659), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14655) );
  NAND3_X1 U17613 ( .A1(n14655), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14201), .ZN(n14203) );
  OAI211_X1 U17614 ( .C1(n14661), .C2(n14204), .A(n14203), .B(n14202), .ZN(
        n14205) );
  AOI21_X1 U17615 ( .B1(n14206), .B2(n19974), .A(n14205), .ZN(n14207) );
  OAI21_X1 U17616 ( .B1(n14208), .B2(n14832), .A(n14207), .ZN(P1_U3000) );
  NAND2_X1 U17617 ( .A1(n14855), .A2(n14211), .ZN(n14212) );
  NAND2_X1 U17618 ( .A1(n9698), .A2(n14212), .ZN(n15035) );
  NAND2_X1 U17619 ( .A1(n15214), .A2(n15227), .ZN(n15230) );
  NAND2_X1 U17620 ( .A1(n15228), .A2(n15230), .ZN(n15221) );
  AOI21_X1 U17621 ( .B1(n15214), .B2(n15213), .A(n15221), .ZN(n14219) );
  NAND2_X1 U17622 ( .A1(n14858), .A2(n14213), .ZN(n14214) );
  INV_X1 U17623 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19666) );
  NOR2_X1 U17624 ( .A1(n18885), .A2(n19666), .ZN(n15033) );
  INV_X1 U17625 ( .A(n15033), .ZN(n14216) );
  INV_X1 U17626 ( .A(n14217), .ZN(n14218) );
  OAI21_X1 U17627 ( .B1(n14219), .B2(n15200), .A(n14218), .ZN(n14220) );
  INV_X1 U17628 ( .A(n14220), .ZN(n14221) );
  NAND2_X1 U17629 ( .A1(n14222), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14225) );
  XNOR2_X1 U17630 ( .A(n14223), .B(n14226), .ZN(n14224) );
  MUX2_X1 U17631 ( .A(n14225), .B(n14224), .S(n11289), .Z(n14228) );
  INV_X1 U17632 ( .A(n14222), .ZN(n14227) );
  NAND3_X1 U17633 ( .A1(n14227), .A2(n14788), .A3(n14226), .ZN(n14817) );
  NAND2_X1 U17634 ( .A1(n14228), .A2(n14817), .ZN(n15960) );
  NAND2_X1 U17635 ( .A1(n15960), .A2(n19939), .ZN(n14233) );
  INV_X1 U17636 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14229) );
  NOR2_X1 U17637 ( .A1(n15922), .A2(n14229), .ZN(n15954) );
  INV_X1 U17638 ( .A(n15846), .ZN(n14230) );
  NOR2_X1 U17639 ( .A1(n19943), .A2(n14230), .ZN(n14231) );
  AOI211_X1 U17640 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15954), .B(n14231), .ZN(n14232) );
  OAI211_X1 U17641 ( .C1(n19998), .C2(n15843), .A(n14233), .B(n14232), .ZN(
        P1_U2989) );
  MUX2_X1 U17642 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n19996), .Z(
        n19907) );
  AOI22_X1 U17643 ( .A1(n14234), .A2(n19907), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15863), .ZN(n14235) );
  OAI21_X1 U17644 ( .B1(n15843), .B2(n14507), .A(n14235), .ZN(P1_U2894) );
  NAND2_X1 U17645 ( .A1(n9698), .A2(n10052), .ZN(n14237) );
  NAND2_X1 U17646 ( .A1(n14238), .A2(n14237), .ZN(n16006) );
  NOR2_X1 U17647 ( .A1(n16006), .A2(n12964), .ZN(n14239) );
  AOI21_X1 U17648 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n12964), .A(n14239), .ZN(
        n14240) );
  OAI21_X1 U17649 ( .B1(n14241), .B2(n14961), .A(n14240), .ZN(P2_U2857) );
  NAND2_X1 U17650 ( .A1(n14242), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14244)
         );
  NAND3_X1 U17651 ( .A1(n14244), .A2(n19753), .A3(n14243), .ZN(P1_U2801) );
  NAND2_X1 U17652 ( .A1(n14462), .A2(n19797), .ZN(n14252) );
  NAND2_X1 U17653 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14248) );
  NAND2_X1 U17654 ( .A1(n19837), .A2(n14248), .ZN(n14245) );
  NAND2_X1 U17655 ( .A1(n14246), .A2(n14245), .ZN(n14267) );
  OAI22_X1 U17656 ( .A1(n19847), .A2(n20811), .B1(n14247), .B2(n19819), .ZN(
        n14250) );
  NOR3_X1 U17657 ( .A1(n14263), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14248), 
        .ZN(n14249) );
  AOI211_X1 U17658 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14267), .A(n14250), 
        .B(n14249), .ZN(n14251) );
  OAI211_X1 U17659 ( .C1(n14403), .C2(n19865), .A(n14252), .B(n14251), .ZN(
        P1_U2809) );
  INV_X1 U17660 ( .A(n14253), .ZN(n14254) );
  AOI22_X1 U17661 ( .A1(n14256), .A2(n14255), .B1(n14254), .B2(n14272), .ZN(
        n14258) );
  AOI21_X1 U17662 ( .B1(n14261), .B2(n14260), .A(n14259), .ZN(n14515) );
  NAND2_X1 U17663 ( .A1(n14515), .A2(n19797), .ZN(n14270) );
  INV_X1 U17664 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14262) );
  OAI21_X1 U17665 ( .B1(n14263), .B2(n20705), .A(n14262), .ZN(n14268) );
  INV_X1 U17666 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14404) );
  NOR2_X1 U17667 ( .A1(n19847), .A2(n14404), .ZN(n14266) );
  OAI22_X1 U17668 ( .A1(n14264), .A2(n19819), .B1(n19833), .B2(n14513), .ZN(
        n14265) );
  AOI211_X1 U17669 ( .C1(n14268), .C2(n14267), .A(n14266), .B(n14265), .ZN(
        n14269) );
  OAI211_X1 U17670 ( .C1(n19865), .C2(n14652), .A(n14270), .B(n14269), .ZN(
        P1_U2810) );
  AOI21_X1 U17671 ( .B1(n14271), .B2(n14283), .A(n9663), .ZN(n14525) );
  INV_X1 U17672 ( .A(n14525), .ZN(n14470) );
  AOI21_X1 U17673 ( .B1(n14273), .B2(n14281), .A(n14272), .ZN(n14672) );
  INV_X1 U17674 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14406) );
  OAI21_X1 U17675 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14275), .A(n14274), 
        .ZN(n14278) );
  INV_X1 U17676 ( .A(n14276), .ZN(n14529) );
  AOI22_X1 U17677 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19853), .B1(
        n19850), .B2(n14529), .ZN(n14277) );
  OAI211_X1 U17678 ( .C1(n19847), .C2(n14406), .A(n14278), .B(n14277), .ZN(
        n14279) );
  AOI21_X1 U17679 ( .B1(n14672), .B2(n19834), .A(n14279), .ZN(n14280) );
  OAI21_X1 U17680 ( .B1(n14470), .B2(n15842), .A(n14280), .ZN(P1_U2812) );
  OAI21_X1 U17681 ( .B1(n9717), .B2(n14282), .A(n14281), .ZN(n14677) );
  INV_X1 U17682 ( .A(n14283), .ZN(n14284) );
  AOI21_X1 U17683 ( .B1(n14285), .B2(n14293), .A(n14284), .ZN(n14535) );
  NAND2_X1 U17684 ( .A1(n14535), .A2(n19797), .ZN(n14291) );
  INV_X1 U17685 ( .A(n14286), .ZN(n14296) );
  INV_X1 U17686 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14536) );
  NAND3_X1 U17687 ( .A1(n14297), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n14536), 
        .ZN(n14288) );
  AOI22_X1 U17688 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19853), .B1(
        n19850), .B2(n14539), .ZN(n14287) );
  OAI211_X1 U17689 ( .C1(n9970), .C2(n19847), .A(n14288), .B(n14287), .ZN(
        n14289) );
  AOI21_X1 U17690 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14296), .A(n14289), 
        .ZN(n14290) );
  OAI211_X1 U17691 ( .C1(n19865), .C2(n14677), .A(n14291), .B(n14290), .ZN(
        P1_U2813) );
  AOI21_X1 U17692 ( .B1(n14294), .B2(n14303), .A(n10124), .ZN(n14545) );
  INV_X1 U17693 ( .A(n14545), .ZN(n14476) );
  AOI21_X1 U17694 ( .B1(n14295), .B2(n14307), .A(n9717), .ZN(n14693) );
  INV_X1 U17695 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14408) );
  OAI21_X1 U17696 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n14297), .A(n14296), 
        .ZN(n14300) );
  INV_X1 U17697 ( .A(n14298), .ZN(n14549) );
  AOI22_X1 U17698 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19853), .B1(
        n19850), .B2(n14549), .ZN(n14299) );
  OAI211_X1 U17699 ( .C1(n19847), .C2(n14408), .A(n14300), .B(n14299), .ZN(
        n14301) );
  AOI21_X1 U17700 ( .B1(n14693), .B2(n19834), .A(n14301), .ZN(n14302) );
  OAI21_X1 U17701 ( .B1(n14476), .B2(n15842), .A(n14302), .ZN(P1_U2814) );
  OAI21_X1 U17702 ( .B1(n9707), .B2(n14304), .A(n14303), .ZN(n14562) );
  NAND2_X1 U17703 ( .A1(n14321), .A2(n14305), .ZN(n14306) );
  NAND2_X1 U17704 ( .A1(n14307), .A2(n14306), .ZN(n14701) );
  INV_X1 U17705 ( .A(n14701), .ZN(n14315) );
  OR2_X1 U17706 ( .A1(n19836), .A2(n14323), .ZN(n14308) );
  NAND2_X1 U17707 ( .A1(n19801), .A2(n14308), .ZN(n14337) );
  INV_X1 U17708 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14557) );
  OAI22_X1 U17709 ( .A1(n14309), .A2(n19819), .B1(n19833), .B2(n14558), .ZN(
        n14310) );
  AOI21_X1 U17710 ( .B1(n19849), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14310), .ZN(
        n14313) );
  OAI21_X1 U17711 ( .B1(n14323), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14311) );
  OAI211_X1 U17712 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n19837), .B(n14311), .ZN(n14312) );
  OAI211_X1 U17713 ( .C1(n14337), .C2(n14557), .A(n14313), .B(n14312), .ZN(
        n14314) );
  AOI21_X1 U17714 ( .B1(n14315), .B2(n19834), .A(n14314), .ZN(n14316) );
  OAI21_X1 U17715 ( .B1(n14562), .B2(n15842), .A(n14316), .ZN(P1_U2815) );
  NOR2_X1 U17716 ( .A1(n9708), .A2(n14317), .ZN(n14318) );
  OR2_X1 U17717 ( .A1(n14331), .A2(n14319), .ZN(n14320) );
  NAND2_X1 U17718 ( .A1(n14321), .A2(n14320), .ZN(n14711) );
  INV_X1 U17719 ( .A(n14711), .ZN(n14328) );
  INV_X1 U17720 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20696) );
  OAI22_X1 U17721 ( .A1(n14322), .A2(n19819), .B1(n19833), .B2(n14567), .ZN(
        n14325) );
  NOR3_X1 U17722 ( .A1(n19826), .A2(n14323), .A3(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14324) );
  AOI211_X1 U17723 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n19849), .A(n14325), .B(
        n14324), .ZN(n14326) );
  OAI21_X1 U17724 ( .B1(n20696), .B2(n14337), .A(n14326), .ZN(n14327) );
  AOI21_X1 U17725 ( .B1(n14328), .B2(n19834), .A(n14327), .ZN(n14329) );
  OAI21_X1 U17726 ( .B1(n14571), .B2(n15842), .A(n14329), .ZN(P1_U2816) );
  AOI21_X1 U17727 ( .B1(n14330), .B2(n14584), .A(n9708), .ZN(n14577) );
  INV_X1 U17728 ( .A(n14577), .ZN(n14485) );
  INV_X1 U17729 ( .A(n14331), .ZN(n14332) );
  OAI21_X1 U17730 ( .B1(n14720), .B2(n14333), .A(n14332), .ZN(n14411) );
  INV_X1 U17731 ( .A(n14411), .ZN(n14717) );
  AND2_X1 U17732 ( .A1(n19837), .A2(n14334), .ZN(n15745) );
  AOI21_X1 U17733 ( .B1(n15745), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U17734 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19853), .B1(
        n19850), .B2(n14573), .ZN(n14336) );
  NAND2_X1 U17735 ( .A1(n19849), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n14335) );
  OAI211_X1 U17736 ( .C1(n14338), .C2(n14337), .A(n14336), .B(n14335), .ZN(
        n14339) );
  AOI21_X1 U17737 ( .B1(n14717), .B2(n19834), .A(n14339), .ZN(n14340) );
  OAI21_X1 U17738 ( .B1(n14485), .B2(n15842), .A(n14340), .ZN(P1_U2817) );
  NOR2_X1 U17739 ( .A1(n14341), .A2(n14342), .ZN(n14343) );
  OR2_X1 U17740 ( .A1(n14425), .A2(n14344), .ZN(n14345) );
  AND2_X1 U17741 ( .A1(n14345), .A2(n14416), .ZN(n14748) );
  INV_X1 U17742 ( .A(n14346), .ZN(n14351) );
  INV_X1 U17743 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14604) );
  NOR2_X1 U17744 ( .A1(n14351), .A2(n14604), .ZN(n15760) );
  OR2_X1 U17745 ( .A1(n19826), .A2(n15760), .ZN(n14350) );
  NAND2_X1 U17746 ( .A1(n14350), .A2(n19827), .ZN(n15751) );
  NAND2_X1 U17747 ( .A1(n15751), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14349) );
  OAI22_X1 U17748 ( .A1(n14606), .A2(n19833), .B1(n14419), .B2(n19847), .ZN(
        n14347) );
  AOI21_X1 U17749 ( .B1(n19853), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14347), .ZN(n14348) );
  OAI211_X1 U17750 ( .C1(n14351), .C2(n14350), .A(n14349), .B(n14348), .ZN(
        n14352) );
  AOI21_X1 U17751 ( .B1(n14748), .B2(n19834), .A(n14352), .ZN(n14353) );
  OAI21_X1 U17752 ( .B1(n14603), .B2(n15842), .A(n14353), .ZN(P1_U2820) );
  INV_X1 U17753 ( .A(n14354), .ZN(n14355) );
  OAI21_X1 U17754 ( .B1(n14356), .B2(n14355), .A(n13764), .ZN(n14452) );
  AND2_X1 U17755 ( .A1(n14452), .A2(n14451), .ZN(n14454) );
  OAI21_X1 U17756 ( .B1(n14454), .B2(n14358), .A(n14357), .ZN(n14645) );
  OAI21_X1 U17757 ( .B1(n19826), .B2(n14359), .A(n19827), .ZN(n15825) );
  NOR2_X1 U17758 ( .A1(n14455), .A2(n14360), .ZN(n14361) );
  OR2_X1 U17759 ( .A1(n14362), .A2(n14361), .ZN(n15948) );
  OAI22_X1 U17760 ( .A1(n14447), .A2(n19847), .B1(n19865), .B2(n15948), .ZN(
        n14363) );
  AOI21_X1 U17761 ( .B1(n14648), .B2(n19850), .A(n14363), .ZN(n14364) );
  OAI211_X1 U17762 ( .C1(n19819), .C2(n14644), .A(n14364), .B(n19817), .ZN(
        n14365) );
  AOI21_X1 U17763 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15825), .A(n14365), 
        .ZN(n14370) );
  NOR2_X1 U17764 ( .A1(n19826), .A2(n14366), .ZN(n14374) );
  INV_X1 U17765 ( .A(n14374), .ZN(n14367) );
  NOR2_X1 U17766 ( .A1(n14367), .A2(n20677), .ZN(n19781) );
  NAND3_X1 U17767 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n19781), .ZN(n15836) );
  NOR2_X1 U17768 ( .A1(n14368), .A2(n15836), .ZN(n15811) );
  NAND2_X1 U17769 ( .A1(n15811), .A2(n14643), .ZN(n14369) );
  OAI211_X1 U17770 ( .C1(n14645), .C2(n15842), .A(n14370), .B(n14369), .ZN(
        P1_U2827) );
  OAI21_X1 U17771 ( .B1(n19826), .B2(n14371), .A(n19827), .ZN(n15837) );
  NAND2_X1 U17772 ( .A1(n19853), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14372) );
  OAI211_X1 U17773 ( .C1(n19833), .C2(n14373), .A(n19817), .B(n14372), .ZN(
        n14378) );
  AOI22_X1 U17774 ( .A1(n19834), .A2(n15966), .B1(n14374), .B2(n20677), .ZN(
        n14375) );
  OAI21_X1 U17775 ( .B1(n14376), .B2(n19847), .A(n14375), .ZN(n14377) );
  AOI211_X1 U17776 ( .C1(P1_REIP_REG_8__SCAN_IN), .C2(n15837), .A(n14378), .B(
        n14377), .ZN(n14379) );
  OAI21_X1 U17777 ( .B1(n14380), .B2(n15842), .A(n14379), .ZN(P1_U2832) );
  NAND2_X1 U17778 ( .A1(n14385), .A2(n14381), .ZN(n14382) );
  NAND2_X1 U17779 ( .A1(n15842), .A2(n14382), .ZN(n19830) );
  INV_X1 U17780 ( .A(n14383), .ZN(n14384) );
  NAND2_X1 U17781 ( .A1(n14385), .A2(n14384), .ZN(n19820) );
  NAND2_X1 U17782 ( .A1(n19850), .A2(n20903), .ZN(n14388) );
  NAND2_X1 U17783 ( .A1(n19853), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14387) );
  AOI22_X1 U17784 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n19849), .B1(n19836), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14386) );
  AND3_X1 U17785 ( .A1(n14388), .A2(n14387), .A3(n14386), .ZN(n14392) );
  INV_X1 U17786 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14390) );
  AOI22_X1 U17787 ( .A1(n19837), .A2(n14390), .B1(n19834), .B2(n14389), .ZN(
        n14391) );
  OAI211_X1 U17788 ( .C1(n20433), .C2(n19820), .A(n14392), .B(n14391), .ZN(
        n14393) );
  INV_X1 U17789 ( .A(n14393), .ZN(n14394) );
  OAI21_X1 U17790 ( .B1(n14395), .B2(n19858), .A(n14394), .ZN(P1_U2839) );
  INV_X1 U17791 ( .A(n19820), .ZN(n19862) );
  NAND2_X1 U17792 ( .A1(n19819), .A2(n19833), .ZN(n14396) );
  AOI22_X1 U17793 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n14396), .B1(
        n19849), .B2(P1_EBX_REG_0__SCAN_IN), .ZN(n14398) );
  NAND2_X1 U17794 ( .A1(n19801), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14397) );
  OAI211_X1 U17795 ( .C1(n14399), .C2(n19865), .A(n14398), .B(n14397), .ZN(
        n14400) );
  AOI21_X1 U17796 ( .B1(n20111), .B2(n19862), .A(n14400), .ZN(n14401) );
  OAI21_X1 U17797 ( .B1(n14402), .B2(n19858), .A(n14401), .ZN(P1_U2840) );
  INV_X1 U17798 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n20811) );
  OAI22_X1 U17799 ( .A1(n14403), .A2(n14448), .B1(n19873), .B2(n20811), .ZN(
        P1_U2841) );
  INV_X1 U17800 ( .A(n14515), .ZN(n14467) );
  OAI222_X1 U17801 ( .A1(n14460), .A2(n14467), .B1(n14404), .B2(n19873), .C1(
        n14652), .C2(n14448), .ZN(P1_U2842) );
  INV_X1 U17802 ( .A(n14672), .ZN(n14405) );
  OAI222_X1 U17803 ( .A1(n14460), .A2(n14470), .B1(n14406), .B2(n19873), .C1(
        n14405), .C2(n14448), .ZN(P1_U2844) );
  INV_X1 U17804 ( .A(n14535), .ZN(n14473) );
  OAI222_X1 U17805 ( .A1(n14460), .A2(n14473), .B1(n9970), .B2(n19873), .C1(
        n14677), .C2(n14448), .ZN(P1_U2845) );
  INV_X1 U17806 ( .A(n14693), .ZN(n14407) );
  OAI222_X1 U17807 ( .A1(n14460), .A2(n14476), .B1(n14408), .B2(n19873), .C1(
        n14407), .C2(n14448), .ZN(P1_U2846) );
  INV_X1 U17808 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14409) );
  OAI222_X1 U17809 ( .A1(n14460), .A2(n14562), .B1(n14409), .B2(n19873), .C1(
        n14701), .C2(n14448), .ZN(P1_U2847) );
  INV_X1 U17810 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14410) );
  OAI222_X1 U17811 ( .A1(n14460), .A2(n14571), .B1(n14410), .B2(n19873), .C1(
        n14711), .C2(n14448), .ZN(P1_U2848) );
  OAI222_X1 U17812 ( .A1(n14460), .A2(n14485), .B1(n14412), .B2(n19873), .C1(
        n14411), .C2(n14448), .ZN(P1_U2849) );
  OAI21_X1 U17813 ( .B1(n14414), .B2(n14413), .A(n14586), .ZN(n15756) );
  NAND2_X1 U17814 ( .A1(n14416), .A2(n14415), .ZN(n14417) );
  AND2_X1 U17815 ( .A1(n14721), .A2(n14417), .ZN(n15754) );
  AOI22_X1 U17816 ( .A1(n15754), .A2(n19869), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14458), .ZN(n14418) );
  OAI21_X1 U17817 ( .B1(n15756), .B2(n14460), .A(n14418), .ZN(P1_U2851) );
  NOR2_X1 U17818 ( .A1(n19873), .A2(n14419), .ZN(n14420) );
  AOI21_X1 U17819 ( .B1(n14748), .B2(n19869), .A(n14420), .ZN(n14421) );
  OAI21_X1 U17820 ( .B1(n14603), .B2(n14460), .A(n14421), .ZN(P1_U2852) );
  AOI21_X1 U17821 ( .B1(n14422), .B2(n14620), .A(n14341), .ZN(n15769) );
  INV_X1 U17822 ( .A(n14460), .ZN(n19870) );
  NOR2_X1 U17823 ( .A1(n14769), .A2(n14423), .ZN(n14424) );
  OR2_X1 U17824 ( .A1(n14425), .A2(n14424), .ZN(n15775) );
  OAI22_X1 U17825 ( .A1(n15775), .A2(n14448), .B1(n14426), .B2(n19873), .ZN(
        n14427) );
  AOI21_X1 U17826 ( .B1(n15769), .B2(n19870), .A(n14427), .ZN(n14428) );
  INV_X1 U17827 ( .A(n14428), .ZN(P1_U2853) );
  NAND2_X1 U17828 ( .A1(n13710), .A2(n14429), .ZN(n14440) );
  AOI21_X1 U17829 ( .B1(n14431), .B2(n14440), .A(n14430), .ZN(n15880) );
  INV_X1 U17830 ( .A(n15880), .ZN(n14436) );
  INV_X1 U17831 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14435) );
  NAND2_X1 U17832 ( .A1(n14444), .A2(n14432), .ZN(n14433) );
  NAND2_X1 U17833 ( .A1(n14434), .A2(n14433), .ZN(n15923) );
  OAI222_X1 U17834 ( .A1(n14436), .A2(n14460), .B1(n14435), .B2(n19873), .C1(
        n14448), .C2(n15923), .ZN(P1_U2856) );
  NAND2_X1 U17835 ( .A1(n14438), .A2(n14437), .ZN(n14439) );
  NAND2_X1 U17836 ( .A1(n15889), .A2(n19870), .ZN(n14446) );
  NAND2_X1 U17837 ( .A1(n14442), .A2(n14441), .ZN(n14443) );
  AND2_X1 U17838 ( .A1(n14444), .A2(n14443), .ZN(n15932) );
  NAND2_X1 U17839 ( .A1(n15932), .A2(n19869), .ZN(n14445) );
  OAI211_X1 U17840 ( .C1(n15802), .C2(n19873), .A(n14446), .B(n14445), .ZN(
        P1_U2857) );
  OAI22_X1 U17841 ( .A1(n15948), .A2(n14448), .B1(n14447), .B2(n19873), .ZN(
        n14449) );
  INV_X1 U17842 ( .A(n14449), .ZN(n14450) );
  OAI21_X1 U17843 ( .B1(n14645), .B2(n14460), .A(n14450), .ZN(P1_U2859) );
  NOR2_X1 U17844 ( .A1(n14452), .A2(n14451), .ZN(n14453) );
  AOI21_X1 U17845 ( .B1(n14457), .B2(n14456), .A(n14455), .ZN(n15822) );
  AOI22_X1 U17846 ( .A1(n15822), .A2(n19869), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n14458), .ZN(n14459) );
  OAI21_X1 U17847 ( .B1(n15897), .B2(n14460), .A(n14459), .ZN(P1_U2860) );
  NAND3_X1 U17848 ( .A1(n14462), .A2(n14461), .A3(n14505), .ZN(n14464) );
  AOI22_X1 U17849 ( .A1(n15866), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15863), .ZN(n14463) );
  OAI211_X1 U17850 ( .C1(n15870), .C2(n16304), .A(n14464), .B(n14463), .ZN(
        P1_U2873) );
  AOI22_X1 U17851 ( .A1(n15866), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n15863), .ZN(n14466) );
  AOI22_X1 U17852 ( .A1(n15865), .A2(n19915), .B1(BUF1_REG_30__SCAN_IN), .B2(
        n14493), .ZN(n14465) );
  OAI211_X1 U17853 ( .C1(n14467), .C2(n14507), .A(n14466), .B(n14465), .ZN(
        P1_U2874) );
  AOI22_X1 U17854 ( .A1(n15866), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n15863), .ZN(n14469) );
  MUX2_X1 U17855 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n19996), .Z(
        n19911) );
  AOI22_X1 U17856 ( .A1(n15865), .A2(n19911), .B1(BUF1_REG_28__SCAN_IN), .B2(
        n14493), .ZN(n14468) );
  OAI211_X1 U17857 ( .C1(n14470), .C2(n14489), .A(n14469), .B(n14468), .ZN(
        P1_U2876) );
  AOI22_X1 U17858 ( .A1(n15866), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15863), .ZN(n14472) );
  AOI22_X1 U17859 ( .A1(n15865), .A2(n19909), .B1(BUF1_REG_27__SCAN_IN), .B2(
        n14493), .ZN(n14471) );
  OAI211_X1 U17860 ( .C1(n14473), .C2(n14489), .A(n14472), .B(n14471), .ZN(
        P1_U2877) );
  AOI22_X1 U17861 ( .A1(n15866), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n15863), .ZN(n14475) );
  AOI22_X1 U17862 ( .A1(n15865), .A2(n19907), .B1(BUF1_REG_26__SCAN_IN), .B2(
        n14493), .ZN(n14474) );
  OAI211_X1 U17863 ( .C1(n14476), .C2(n14489), .A(n14475), .B(n14474), .ZN(
        P1_U2878) );
  AOI22_X1 U17864 ( .A1(n15866), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n15863), .ZN(n14478) );
  AOI22_X1 U17865 ( .A1(n15865), .A2(n19905), .B1(n14493), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14477) );
  OAI211_X1 U17866 ( .C1(n14562), .C2(n14489), .A(n14478), .B(n14477), .ZN(
        P1_U2879) );
  AOI22_X1 U17867 ( .A1(n15866), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n15863), .ZN(n14481) );
  AOI22_X1 U17868 ( .A1(n15865), .A2(n14479), .B1(n14493), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14480) );
  OAI211_X1 U17869 ( .C1(n14571), .C2(n14489), .A(n14481), .B(n14480), .ZN(
        P1_U2880) );
  AOI22_X1 U17870 ( .A1(n15866), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n15863), .ZN(n14484) );
  AOI22_X1 U17871 ( .A1(n15865), .A2(n14482), .B1(n14493), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14483) );
  OAI211_X1 U17872 ( .C1(n14485), .C2(n14489), .A(n14484), .B(n14483), .ZN(
        P1_U2881) );
  AOI22_X1 U17873 ( .A1(n15866), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n15863), .ZN(n14488) );
  AOI22_X1 U17874 ( .A1(n15865), .A2(n14486), .B1(n14493), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14487) );
  OAI211_X1 U17875 ( .C1(n15756), .C2(n14489), .A(n14488), .B(n14487), .ZN(
        P1_U2883) );
  AOI22_X1 U17876 ( .A1(n15866), .A2(DATAI_20_), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15863), .ZN(n14492) );
  AOI22_X1 U17877 ( .A1(n15865), .A2(n14490), .B1(n14493), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14491) );
  OAI211_X1 U17878 ( .C1(n14603), .C2(n14507), .A(n14492), .B(n14491), .ZN(
        P1_U2884) );
  INV_X1 U17879 ( .A(n15769), .ZN(n14497) );
  AOI22_X1 U17880 ( .A1(n15866), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15863), .ZN(n14496) );
  AOI22_X1 U17881 ( .A1(n15865), .A2(n14494), .B1(n14493), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14495) );
  OAI211_X1 U17882 ( .C1(n14497), .C2(n14507), .A(n14496), .B(n14495), .ZN(
        P1_U2885) );
  INV_X1 U17883 ( .A(n15889), .ZN(n14500) );
  OAI222_X1 U17884 ( .A1(n14507), .A2(n14500), .B1(n14505), .B2(n14499), .C1(
        n14504), .C2(n14498), .ZN(P1_U2889) );
  INV_X1 U17885 ( .A(n19913), .ZN(n14502) );
  OAI222_X1 U17886 ( .A1(n14507), .A2(n14645), .B1(n14504), .B2(n14502), .C1(
        n14501), .C2(n14505), .ZN(P1_U2891) );
  INV_X1 U17887 ( .A(n19911), .ZN(n14503) );
  OAI222_X1 U17888 ( .A1(n15897), .A2(n14507), .B1(n14506), .B2(n14505), .C1(
        n14504), .C2(n14503), .ZN(P1_U2892) );
  NAND2_X1 U17889 ( .A1(n14628), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14509) );
  OAI21_X1 U17890 ( .B1(n14510), .B2(n14509), .A(n14508), .ZN(n14511) );
  XNOR2_X1 U17891 ( .A(n14511), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14656) );
  NAND2_X1 U17892 ( .A1(n19944), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14651) );
  NAND2_X1 U17893 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14512) );
  OAI211_X1 U17894 ( .C1(n19943), .C2(n14513), .A(n14651), .B(n14512), .ZN(
        n14514) );
  AOI21_X1 U17895 ( .B1(n14515), .B2(n19938), .A(n14514), .ZN(n14516) );
  OAI21_X1 U17896 ( .B1(n14656), .B2(n15902), .A(n14516), .ZN(P1_U2969) );
  NAND2_X1 U17897 ( .A1(n11289), .A2(n14518), .ZN(n14542) );
  NAND2_X1 U17898 ( .A1(n14517), .A2(n14542), .ZN(n14523) );
  OAI21_X1 U17899 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14519), .A(
        n14523), .ZN(n14522) );
  MUX2_X1 U17900 ( .A(n14520), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n11289), .Z(n14521) );
  OAI211_X1 U17901 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14523), .A(
        n14522), .B(n14521), .ZN(n14524) );
  XOR2_X1 U17902 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14524), .Z(
        n14674) );
  NAND2_X1 U17903 ( .A1(n14525), .A2(n19938), .ZN(n14531) );
  INV_X1 U17904 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14526) );
  OR2_X1 U17905 ( .A1(n15922), .A2(n14526), .ZN(n14668) );
  OAI21_X1 U17906 ( .B1(n15914), .B2(n14527), .A(n14668), .ZN(n14528) );
  AOI21_X1 U17907 ( .B1(n14529), .B2(n15909), .A(n14528), .ZN(n14530) );
  OAI211_X1 U17908 ( .C1(n14674), .C2(n15902), .A(n14531), .B(n14530), .ZN(
        P1_U2971) );
  INV_X1 U17909 ( .A(n14532), .ZN(n14534) );
  NAND2_X1 U17910 ( .A1(n14535), .A2(n19938), .ZN(n14541) );
  OR2_X1 U17911 ( .A1(n15922), .A2(n14536), .ZN(n14675) );
  OAI21_X1 U17912 ( .B1(n15914), .B2(n14537), .A(n14675), .ZN(n14538) );
  AOI21_X1 U17913 ( .B1(n14539), .B2(n15909), .A(n14538), .ZN(n14540) );
  OAI211_X1 U17914 ( .C1(n14682), .C2(n15902), .A(n14541), .B(n14540), .ZN(
        P1_U2972) );
  NAND3_X1 U17915 ( .A1(n14543), .A2(n14542), .A3(n14553), .ZN(n14544) );
  XNOR2_X1 U17916 ( .A(n14544), .B(n14683), .ZN(n14695) );
  NAND2_X1 U17917 ( .A1(n14545), .A2(n19938), .ZN(n14551) );
  INV_X1 U17918 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14546) );
  OR2_X1 U17919 ( .A1(n15922), .A2(n14546), .ZN(n14689) );
  OAI21_X1 U17920 ( .B1(n15914), .B2(n14547), .A(n14689), .ZN(n14548) );
  AOI21_X1 U17921 ( .B1(n14549), .B2(n15909), .A(n14548), .ZN(n14550) );
  OAI211_X1 U17922 ( .C1(n14695), .C2(n15902), .A(n14551), .B(n14550), .ZN(
        P1_U2973) );
  INV_X1 U17923 ( .A(n14517), .ZN(n14552) );
  NAND3_X1 U17924 ( .A1(n14552), .A2(n14705), .A3(n14565), .ZN(n14555) );
  NAND2_X1 U17925 ( .A1(n14564), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14554) );
  MUX2_X1 U17926 ( .A(n14555), .B(n14554), .S(n11289), .Z(n14556) );
  NOR2_X1 U17927 ( .A1(n15922), .A2(n14557), .ZN(n14697) );
  NOR2_X1 U17928 ( .A1(n19943), .A2(n14558), .ZN(n14559) );
  AOI211_X1 U17929 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14697), .B(n14559), .ZN(n14560) );
  OAI211_X1 U17930 ( .C1(n14562), .C2(n19998), .A(n14561), .B(n14560), .ZN(
        P1_U2974) );
  NOR2_X1 U17931 ( .A1(n14564), .A2(n14517), .ZN(n14563) );
  MUX2_X1 U17932 ( .A(n14564), .B(n14563), .S(n14788), .Z(n14566) );
  XNOR2_X1 U17933 ( .A(n14566), .B(n14565), .ZN(n14702) );
  NAND2_X1 U17934 ( .A1(n14702), .A2(n19939), .ZN(n14570) );
  NOR2_X1 U17935 ( .A1(n15922), .A2(n20696), .ZN(n14707) );
  NOR2_X1 U17936 ( .A1(n19943), .A2(n14567), .ZN(n14568) );
  AOI211_X1 U17937 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14707), .B(n14568), .ZN(n14569) );
  OAI211_X1 U17938 ( .C1(n19998), .C2(n14571), .A(n14570), .B(n14569), .ZN(
        P1_U2975) );
  XNOR2_X1 U17939 ( .A(n14628), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14572) );
  XNOR2_X1 U17940 ( .A(n14517), .B(n14572), .ZN(n14719) );
  NAND2_X1 U17941 ( .A1(n15909), .A2(n14573), .ZN(n14574) );
  NAND2_X1 U17942 ( .A1(n19944), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14713) );
  OAI211_X1 U17943 ( .C1(n15914), .C2(n14575), .A(n14574), .B(n14713), .ZN(
        n14576) );
  AOI21_X1 U17944 ( .B1(n14577), .B2(n19938), .A(n14576), .ZN(n14578) );
  OAI21_X1 U17945 ( .B1(n14719), .B2(n15902), .A(n14578), .ZN(P1_U2976) );
  AND2_X1 U17946 ( .A1(n14580), .A2(n14579), .ZN(n14583) );
  INV_X1 U17947 ( .A(n14580), .ZN(n14582) );
  OAI22_X1 U17948 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n14583), .B1(
        n14582), .B2(n14581), .ZN(n14735) );
  INV_X1 U17949 ( .A(n14584), .ZN(n14585) );
  AOI21_X1 U17950 ( .B1(n14587), .B2(n14586), .A(n14585), .ZN(n15856) );
  NAND2_X1 U17951 ( .A1(n15856), .A2(n19938), .ZN(n14592) );
  INV_X1 U17952 ( .A(n14588), .ZN(n15746) );
  INV_X1 U17953 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20694) );
  OR2_X1 U17954 ( .A1(n15922), .A2(n20694), .ZN(n14723) );
  OAI21_X1 U17955 ( .B1(n15914), .B2(n14589), .A(n14723), .ZN(n14590) );
  AOI21_X1 U17956 ( .B1(n15746), .B2(n15909), .A(n14590), .ZN(n14591) );
  OAI211_X1 U17957 ( .C1(n14735), .C2(n15902), .A(n14592), .B(n14591), .ZN(
        P1_U2977) );
  NAND2_X1 U17958 ( .A1(n14628), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14594) );
  NOR2_X1 U17959 ( .A1(n14617), .A2(n14594), .ZN(n14596) );
  AOI21_X1 U17960 ( .B1(n14595), .B2(n14788), .A(n14596), .ZN(n14602) );
  NOR2_X1 U17961 ( .A1(n14602), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14601) );
  AOI22_X1 U17962 ( .A1(n14601), .A2(n14788), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14596), .ZN(n14597) );
  XNOR2_X1 U17963 ( .A(n14597), .B(n14737), .ZN(n14743) );
  NAND2_X1 U17964 ( .A1(n19944), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14736) );
  OAI21_X1 U17965 ( .B1(n15914), .B2(n20839), .A(n14736), .ZN(n14599) );
  NOR2_X1 U17966 ( .A1(n15756), .A2(n19998), .ZN(n14598) );
  AOI211_X1 U17967 ( .C1(n15909), .C2(n15752), .A(n14599), .B(n14598), .ZN(
        n14600) );
  OAI21_X1 U17968 ( .B1(n14743), .B2(n15902), .A(n14600), .ZN(P1_U2978) );
  AOI21_X1 U17969 ( .B1(n14602), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14601), .ZN(n14755) );
  INV_X1 U17970 ( .A(n14603), .ZN(n14608) );
  NOR2_X1 U17971 ( .A1(n15922), .A2(n14604), .ZN(n14747) );
  AOI21_X1 U17972 ( .B1(n19932), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14747), .ZN(n14605) );
  OAI21_X1 U17973 ( .B1(n19943), .B2(n14606), .A(n14605), .ZN(n14607) );
  AOI21_X1 U17974 ( .B1(n14608), .B2(n19938), .A(n14607), .ZN(n14609) );
  OAI21_X1 U17975 ( .B1(n14755), .B2(n15902), .A(n14609), .ZN(P1_U2979) );
  NAND2_X1 U17976 ( .A1(n14617), .A2(n14610), .ZN(n14611) );
  MUX2_X1 U17977 ( .A(n14611), .B(n14617), .S(n11289), .Z(n14612) );
  XNOR2_X1 U17978 ( .A(n14612), .B(n14751), .ZN(n14764) );
  NOR2_X1 U17979 ( .A1(n15922), .A2(n20689), .ZN(n14757) );
  INV_X1 U17980 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14613) );
  NOR2_X1 U17981 ( .A1(n15914), .A2(n14613), .ZN(n14614) );
  AOI211_X1 U17982 ( .C1(n15909), .C2(n15763), .A(n14757), .B(n14614), .ZN(
        n14616) );
  NAND2_X1 U17983 ( .A1(n15769), .A2(n19938), .ZN(n14615) );
  OAI211_X1 U17984 ( .C1(n14764), .C2(n15902), .A(n14616), .B(n14615), .ZN(
        P1_U2980) );
  OAI21_X1 U17985 ( .B1(n14619), .B2(n14618), .A(n14617), .ZN(n14780) );
  INV_X1 U17986 ( .A(n14620), .ZN(n14621) );
  AOI21_X1 U17987 ( .B1(n14623), .B2(n14622), .A(n14621), .ZN(n15860) );
  INV_X1 U17988 ( .A(n15776), .ZN(n14625) );
  NAND2_X1 U17989 ( .A1(n19944), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U17990 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14624) );
  OAI211_X1 U17991 ( .C1(n19943), .C2(n14625), .A(n14776), .B(n14624), .ZN(
        n14626) );
  AOI21_X1 U17992 ( .B1(n15860), .B2(n19938), .A(n14626), .ZN(n14627) );
  OAI21_X1 U17993 ( .B1(n15902), .B2(n14780), .A(n14627), .ZN(P1_U2981) );
  NOR2_X1 U17994 ( .A1(n14628), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14633) );
  NAND2_X1 U17995 ( .A1(n14223), .A2(n15873), .ZN(n14790) );
  INV_X1 U17996 ( .A(n14629), .ZN(n14631) );
  OAI21_X1 U17997 ( .B1(n14790), .B2(n14631), .A(n14630), .ZN(n14632) );
  MUX2_X1 U17998 ( .A(n11289), .B(n14633), .S(n14632), .Z(n14634) );
  XOR2_X1 U17999 ( .A(n14781), .B(n14634), .Z(n14787) );
  NAND2_X1 U18000 ( .A1(n19944), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n14782) );
  OAI21_X1 U18001 ( .B1(n15914), .B2(n15786), .A(n14782), .ZN(n14636) );
  NOR2_X1 U18002 ( .A1(n15783), .A2(n19998), .ZN(n14635) );
  AOI211_X1 U18003 ( .C1(n15909), .C2(n15784), .A(n14636), .B(n14635), .ZN(
        n14637) );
  OAI21_X1 U18004 ( .B1(n14787), .B2(n15902), .A(n14637), .ZN(P1_U2982) );
  INV_X1 U18005 ( .A(n14223), .ZN(n14816) );
  AOI22_X1 U18006 ( .A1(n14816), .A2(n14639), .B1(n14788), .B2(n14638), .ZN(
        n14803) );
  INV_X1 U18007 ( .A(n14641), .ZN(n14640) );
  AOI21_X1 U18008 ( .B1(n14788), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14640), .ZN(n14802) );
  NAND2_X1 U18009 ( .A1(n14803), .A2(n14802), .ZN(n14801) );
  NAND2_X1 U18010 ( .A1(n14801), .A2(n14641), .ZN(n14642) );
  INV_X1 U18011 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14643) );
  OAI22_X1 U18012 ( .A1(n15914), .A2(n14644), .B1(n15922), .B2(n14643), .ZN(
        n14647) );
  NOR2_X1 U18013 ( .A1(n14645), .A2(n19998), .ZN(n14646) );
  AOI211_X1 U18014 ( .C1(n15909), .C2(n14648), .A(n14647), .B(n14646), .ZN(
        n14649) );
  OAI21_X1 U18015 ( .B1(n15942), .B2(n15902), .A(n14649), .ZN(P1_U2986) );
  INV_X1 U18016 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14650) );
  OAI21_X1 U18017 ( .B1(n14661), .B2(n14658), .A(n14650), .ZN(n14654) );
  INV_X1 U18018 ( .A(n14651), .ZN(n14653) );
  INV_X1 U18019 ( .A(n14657), .ZN(n14664) );
  NOR2_X1 U18020 ( .A1(n14659), .A2(n14658), .ZN(n14663) );
  OAI21_X1 U18021 ( .B1(n14661), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14660), .ZN(n14662) );
  AOI211_X1 U18022 ( .C1(n14664), .C2(n19974), .A(n14663), .B(n14662), .ZN(
        n14665) );
  OAI21_X1 U18023 ( .B1(n14666), .B2(n14832), .A(n14665), .ZN(P1_U3002) );
  INV_X1 U18024 ( .A(n14667), .ZN(n14676) );
  XNOR2_X1 U18025 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U18026 ( .A1(n14680), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14669) );
  OAI211_X1 U18027 ( .C1(n14676), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14671) );
  AOI21_X1 U18028 ( .B1(n14672), .B2(n19974), .A(n14671), .ZN(n14673) );
  OAI21_X1 U18029 ( .B1(n14674), .B2(n14832), .A(n14673), .ZN(P1_U3003) );
  OAI21_X1 U18030 ( .B1(n14676), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14675), .ZN(n14679) );
  NOR2_X1 U18031 ( .A1(n14677), .A2(n19981), .ZN(n14678) );
  AOI211_X1 U18032 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14680), .A(
        n14679), .B(n14678), .ZN(n14681) );
  OAI21_X1 U18033 ( .B1(n14682), .B2(n14832), .A(n14681), .ZN(P1_U3004) );
  NAND2_X1 U18034 ( .A1(n14684), .A2(n14683), .ZN(n14691) );
  INV_X1 U18035 ( .A(n14685), .ZN(n14698) );
  NAND2_X1 U18036 ( .A1(n14687), .A2(n14686), .ZN(n14688) );
  NOR2_X1 U18037 ( .A1(n14715), .A2(n14688), .ZN(n14696) );
  OAI21_X1 U18038 ( .B1(n14698), .B2(n14696), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14690) );
  OAI211_X1 U18039 ( .C1(n14715), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        n14692) );
  AOI21_X1 U18040 ( .B1(n14693), .B2(n19974), .A(n14692), .ZN(n14694) );
  OAI21_X1 U18041 ( .B1(n14695), .B2(n14832), .A(n14694), .ZN(P1_U3005) );
  AOI211_X1 U18042 ( .C1(n14698), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14697), .B(n14696), .ZN(n14699) );
  OAI211_X1 U18043 ( .C1(n19981), .C2(n14701), .A(n14700), .B(n14699), .ZN(
        P1_U3006) );
  NAND2_X1 U18044 ( .A1(n14702), .A2(n19988), .ZN(n14710) );
  AOI21_X1 U18045 ( .B1(n14767), .B2(n14703), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14704) );
  OR2_X1 U18046 ( .A1(n14712), .A2(n14704), .ZN(n14708) );
  NOR3_X1 U18047 ( .A1(n14715), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n14705), .ZN(n14706) );
  AOI211_X1 U18048 ( .C1(n14708), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14707), .B(n14706), .ZN(n14709) );
  OAI211_X1 U18049 ( .C1(n19981), .C2(n14711), .A(n14710), .B(n14709), .ZN(
        P1_U3007) );
  NAND2_X1 U18050 ( .A1(n14712), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14714) );
  OAI211_X1 U18051 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14715), .A(
        n14714), .B(n14713), .ZN(n14716) );
  AOI21_X1 U18052 ( .B1(n14717), .B2(n19974), .A(n14716), .ZN(n14718) );
  OAI21_X1 U18053 ( .B1(n14719), .B2(n14832), .A(n14718), .ZN(P1_U3008) );
  AOI21_X1 U18054 ( .B1(n14722), .B2(n14721), .A(n14720), .ZN(n15849) );
  INV_X1 U18055 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14731) );
  OAI21_X1 U18056 ( .B1(n14738), .B2(n14731), .A(n14723), .ZN(n14733) );
  NOR2_X1 U18057 ( .A1(n13034), .A2(n15945), .ZN(n15939) );
  AOI21_X1 U18058 ( .B1(n14725), .B2(n15939), .A(n14724), .ZN(n15953) );
  NOR2_X1 U18059 ( .A1(n15953), .A2(n14756), .ZN(n14750) );
  INV_X1 U18060 ( .A(n14726), .ZN(n14727) );
  NOR2_X1 U18061 ( .A1(n15943), .A2(n14727), .ZN(n14728) );
  OR2_X1 U18062 ( .A1(n14750), .A2(n14728), .ZN(n14745) );
  NAND2_X1 U18063 ( .A1(n14745), .A2(n14729), .ZN(n14739) );
  AOI211_X1 U18064 ( .C1(n14737), .C2(n14731), .A(n14730), .B(n14739), .ZN(
        n14732) );
  AOI211_X1 U18065 ( .C1(n19974), .C2(n15849), .A(n14733), .B(n14732), .ZN(
        n14734) );
  OAI21_X1 U18066 ( .B1(n14735), .B2(n14832), .A(n14734), .ZN(P1_U3009) );
  OAI21_X1 U18067 ( .B1(n14738), .B2(n14737), .A(n14736), .ZN(n14741) );
  NOR2_X1 U18068 ( .A1(n14739), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14740) );
  AOI211_X1 U18069 ( .C1(n19974), .C2(n15754), .A(n14741), .B(n14740), .ZN(
        n14742) );
  OAI21_X1 U18070 ( .B1(n14743), .B2(n14832), .A(n14742), .ZN(P1_U3010) );
  AND3_X1 U18071 ( .A1(n14745), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14744), .ZN(n14746) );
  AOI211_X1 U18072 ( .C1(n19974), .C2(n14748), .A(n14747), .B(n14746), .ZN(
        n14754) );
  OR2_X1 U18073 ( .A1(n14750), .A2(n14749), .ZN(n14752) );
  AND2_X1 U18074 ( .A1(n14752), .A2(n14751), .ZN(n14762) );
  OAI21_X1 U18075 ( .B1(n14762), .B2(n14758), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14753) );
  OAI211_X1 U18076 ( .C1(n14755), .C2(n14832), .A(n14754), .B(n14753), .ZN(
        P1_U3011) );
  AOI21_X1 U18077 ( .B1(n15953), .B2(n15945), .A(n14756), .ZN(n14761) );
  AOI21_X1 U18078 ( .B1(n14758), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n14757), .ZN(n14759) );
  OAI21_X1 U18079 ( .B1(n15775), .B2(n19981), .A(n14759), .ZN(n14760) );
  AOI21_X1 U18080 ( .B1(n14762), .B2(n14761), .A(n14760), .ZN(n14763) );
  OAI21_X1 U18081 ( .B1(n14764), .B2(n14832), .A(n14763), .ZN(P1_U3012) );
  AOI21_X1 U18082 ( .B1(n19961), .B2(n14765), .A(n14808), .ZN(n14766) );
  OAI21_X1 U18083 ( .B1(n14795), .B2(n14767), .A(n14766), .ZN(n14796) );
  AOI21_X1 U18084 ( .B1(n14791), .B2(n19986), .A(n14796), .ZN(n15935) );
  OAI21_X1 U18085 ( .B1(n14768), .B2(n14774), .A(n15935), .ZN(n14785) );
  INV_X1 U18086 ( .A(n14769), .ZN(n14770) );
  OAI21_X1 U18087 ( .B1(n14772), .B2(n14771), .A(n14770), .ZN(n15779) );
  NOR2_X1 U18088 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15937), .ZN(
        n14775) );
  NAND2_X1 U18089 ( .A1(n14775), .A2(n14774), .ZN(n14777) );
  OAI211_X1 U18090 ( .C1(n19981), .C2(n15779), .A(n14777), .B(n14776), .ZN(
        n14778) );
  AOI21_X1 U18091 ( .B1(n14785), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n14778), .ZN(n14779) );
  OAI21_X1 U18092 ( .B1(n14780), .B2(n14832), .A(n14779), .ZN(P1_U3013) );
  OAI21_X1 U18093 ( .B1(n15925), .B2(n15937), .A(n14781), .ZN(n14784) );
  OAI21_X1 U18094 ( .B1(n15793), .B2(n19981), .A(n14782), .ZN(n14783) );
  AOI21_X1 U18095 ( .B1(n14785), .B2(n14784), .A(n14783), .ZN(n14786) );
  OAI21_X1 U18096 ( .B1(n14787), .B2(n14832), .A(n14786), .ZN(P1_U3014) );
  AOI22_X1 U18097 ( .A1(n14790), .A2(n14789), .B1(n14788), .B2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14793) );
  MUX2_X1 U18098 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n14791), .S(
        n11289), .Z(n14792) );
  XNOR2_X1 U18099 ( .A(n14793), .B(n14792), .ZN(n15896) );
  NOR2_X1 U18100 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14826), .ZN(
        n14794) );
  AOI22_X1 U18101 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14796), .B1(
        n14795), .B2(n14794), .ZN(n14800) );
  INV_X1 U18102 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14797) );
  OAI22_X1 U18103 ( .A1(n15812), .A2(n19981), .B1(n15922), .B2(n14797), .ZN(
        n14798) );
  INV_X1 U18104 ( .A(n14798), .ZN(n14799) );
  OAI211_X1 U18105 ( .C1(n15896), .C2(n14832), .A(n14800), .B(n14799), .ZN(
        P1_U3017) );
  OAI21_X1 U18106 ( .B1(n14803), .B2(n14802), .A(n14801), .ZN(n14804) );
  INV_X1 U18107 ( .A(n14804), .ZN(n15903) );
  AOI21_X1 U18108 ( .B1(n14807), .B2(n14806), .A(n14805), .ZN(n14809) );
  AOI211_X1 U18109 ( .C1(n19962), .C2(n14810), .A(n14809), .B(n14808), .ZN(
        n14820) );
  OAI21_X1 U18110 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n19965), .A(
        n14820), .ZN(n14812) );
  OAI21_X1 U18111 ( .B1(n14810), .B2(n14826), .A(n14813), .ZN(n14811) );
  OAI21_X1 U18112 ( .B1(n14813), .B2(n14812), .A(n14811), .ZN(n14815) );
  AOI22_X1 U18113 ( .A1(n15822), .A2(n19974), .B1(n19944), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14814) );
  OAI211_X1 U18114 ( .C1(n15903), .C2(n14832), .A(n14815), .B(n14814), .ZN(
        P1_U3019) );
  NAND3_X1 U18115 ( .A1(n14816), .A2(n11289), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14818) );
  NAND2_X1 U18116 ( .A1(n14818), .A2(n14817), .ZN(n14819) );
  XNOR2_X1 U18117 ( .A(n14819), .B(n11300), .ZN(n15905) );
  NOR2_X1 U18118 ( .A1(n15958), .A2(n15956), .ZN(n14822) );
  INV_X1 U18119 ( .A(n14820), .ZN(n14821) );
  MUX2_X1 U18120 ( .A(n14822), .B(n14821), .S(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(n14824) );
  OAI22_X1 U18121 ( .A1(n15829), .A2(n19981), .B1(n15922), .B2(n15835), .ZN(
        n14823) );
  AOI211_X1 U18122 ( .C1(n15905), .C2(n19988), .A(n14824), .B(n14823), .ZN(
        n14825) );
  INV_X1 U18123 ( .A(n14825), .ZN(P1_U3020) );
  AOI21_X1 U18124 ( .B1(n14827), .B2(n14826), .A(n15968), .ZN(n14828) );
  AOI211_X1 U18125 ( .C1(n19974), .C2(n19794), .A(n14829), .B(n14828), .ZN(
        n14830) );
  OAI21_X1 U18126 ( .B1(n14832), .B2(n14831), .A(n14830), .ZN(P1_U3025) );
  NAND2_X1 U18127 ( .A1(n9654), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20566) );
  NAND2_X1 U18128 ( .A1(n20566), .A2(n20576), .ZN(n20113) );
  NOR2_X1 U18129 ( .A1(n9654), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14834) );
  OAI22_X1 U18130 ( .A1(n20113), .A2(n14834), .B1(n20433), .B2(n14837), .ZN(
        n14835) );
  MUX2_X1 U18131 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14835), .S(
        n20738), .Z(P1_U3477) );
  NAND2_X1 U18132 ( .A1(n9654), .A2(n20725), .ZN(n20258) );
  MUX2_X1 U18133 ( .A(n20258), .B(n20113), .S(n20292), .Z(n14836) );
  OAI21_X1 U18134 ( .B1(n14837), .B2(n12915), .A(n14836), .ZN(n14838) );
  MUX2_X1 U18135 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14838), .S(
        n20738), .Z(P1_U3476) );
  AOI22_X1 U18136 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n18829), .B1(n14839), 
        .B2(n18901), .ZN(n14841) );
  AOI22_X1 U18137 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18906), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n18917), .ZN(n14840) );
  OAI211_X1 U18138 ( .C1(n14964), .C2(n18916), .A(n14841), .B(n14840), .ZN(
        n14846) );
  AOI211_X1 U18139 ( .C1(n14844), .C2(n14843), .A(n14842), .B(n18883), .ZN(
        n14845) );
  NOR2_X1 U18140 ( .A1(n14846), .A2(n14845), .ZN(n14847) );
  OAI21_X1 U18141 ( .B1(n15035), .B2(n18878), .A(n14847), .ZN(P2_U2826) );
  AOI211_X1 U18142 ( .C1(n15053), .C2(n14849), .A(n14848), .B(n18883), .ZN(
        n14861) );
  AOI22_X1 U18143 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18917), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18829), .ZN(n14851) );
  NAND2_X1 U18144 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18906), .ZN(
        n14850) );
  OAI211_X1 U18145 ( .C1(n18925), .C2(n14852), .A(n14851), .B(n14850), .ZN(
        n14860) );
  OR2_X1 U18146 ( .A1(n14907), .A2(n14853), .ZN(n14854) );
  NAND2_X1 U18147 ( .A1(n14855), .A2(n14854), .ZN(n15218) );
  NAND2_X1 U18148 ( .A1(n14978), .A2(n14856), .ZN(n14857) );
  NAND2_X1 U18149 ( .A1(n14858), .A2(n14857), .ZN(n15217) );
  OAI22_X1 U18150 ( .A1(n15218), .A2(n18878), .B1(n15217), .B2(n18916), .ZN(
        n14859) );
  OR3_X1 U18151 ( .A1(n14861), .A2(n14860), .A3(n14859), .ZN(P2_U2827) );
  AOI21_X1 U18152 ( .B1(n14862), .B2(n9662), .A(n10069), .ZN(n15256) );
  INV_X1 U18153 ( .A(n15256), .ZN(n14868) );
  AOI22_X1 U18154 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n18917), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18906), .ZN(n14867) );
  NOR2_X1 U18155 ( .A1(n15001), .A2(n14863), .ZN(n14864) );
  OR2_X1 U18156 ( .A1(n14988), .A2(n14864), .ZN(n15248) );
  INV_X1 U18157 ( .A(n15248), .ZN(n14865) );
  AOI22_X1 U18158 ( .A1(n14865), .A2(n18922), .B1(P2_REIP_REG_25__SCAN_IN), 
        .B2(n18829), .ZN(n14866) );
  OAI211_X1 U18159 ( .C1(n14868), .C2(n18878), .A(n14867), .B(n14866), .ZN(
        n14872) );
  AOI211_X1 U18160 ( .C1(n14870), .C2(n15079), .A(n14869), .B(n18883), .ZN(
        n14871) );
  AOI211_X1 U18161 ( .C1(n14873), .C2(n18901), .A(n14872), .B(n14871), .ZN(
        n14874) );
  INV_X1 U18162 ( .A(n14874), .ZN(P2_U2830) );
  AOI211_X1 U18163 ( .C1(n15100), .C2(n14876), .A(n14875), .B(n18883), .ZN(
        n14877) );
  INV_X1 U18164 ( .A(n14877), .ZN(n14888) );
  AOI22_X1 U18165 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18906), .B1(
        n14878), .B2(n18901), .ZN(n14887) );
  NOR2_X1 U18166 ( .A1(n14940), .A2(n14879), .ZN(n14880) );
  OR2_X1 U18167 ( .A1(n14931), .A2(n14880), .ZN(n15280) );
  INV_X1 U18168 ( .A(n15280), .ZN(n14885) );
  NAND2_X1 U18169 ( .A1(n15301), .A2(n14881), .ZN(n14882) );
  NAND2_X1 U18170 ( .A1(n15002), .A2(n14882), .ZN(n15010) );
  AOI22_X1 U18171 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n18917), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18829), .ZN(n14883) );
  OAI21_X1 U18172 ( .B1(n18916), .B2(n15010), .A(n14883), .ZN(n14884) );
  AOI21_X1 U18173 ( .B1(n14885), .B2(n18927), .A(n14884), .ZN(n14886) );
  NAND3_X1 U18174 ( .A1(n14888), .A2(n14887), .A3(n14886), .ZN(P2_U2832) );
  INV_X1 U18175 ( .A(n14889), .ZN(n14891) );
  NAND2_X1 U18176 ( .A1(n14891), .A2(n14890), .ZN(n14892) );
  OAI21_X1 U18177 ( .B1(n14890), .B2(n10560), .A(n14892), .ZN(P2_U2856) );
  OR2_X1 U18178 ( .A1(n14894), .A2(n14893), .ZN(n14962) );
  NAND3_X1 U18179 ( .A1(n14962), .A2(n14895), .A3(n14945), .ZN(n14897) );
  NAND2_X1 U18180 ( .A1(n12964), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14896) );
  OAI211_X1 U18181 ( .C1(n14946), .C2(n15035), .A(n14897), .B(n14896), .ZN(
        P2_U2858) );
  INV_X1 U18182 ( .A(n14898), .ZN(n14899) );
  NAND2_X1 U18183 ( .A1(n14900), .A2(n14899), .ZN(n14902) );
  XNOR2_X1 U18184 ( .A(n14902), .B(n14901), .ZN(n14976) );
  NOR2_X1 U18185 ( .A1(n15218), .A2(n12964), .ZN(n14903) );
  AOI21_X1 U18186 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n12964), .A(n14903), .ZN(
        n14904) );
  OAI21_X1 U18187 ( .B1(n14976), .B2(n14961), .A(n14904), .ZN(P2_U2859) );
  OAI21_X1 U18188 ( .B1(n9715), .B2(n14906), .A(n14905), .ZN(n14986) );
  NAND2_X1 U18189 ( .A1(n14946), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14910) );
  AOI21_X1 U18190 ( .B1(n14908), .B2(n14917), .A(n14907), .ZN(n16018) );
  NAND2_X1 U18191 ( .A1(n16018), .A2(n14890), .ZN(n14909) );
  OAI211_X1 U18192 ( .C1(n14986), .C2(n14961), .A(n14910), .B(n14909), .ZN(
        P2_U2860) );
  OAI21_X1 U18193 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(n14994) );
  NAND2_X1 U18194 ( .A1(n14915), .A2(n14914), .ZN(n14916) );
  NAND2_X1 U18195 ( .A1(n14917), .A2(n14916), .ZN(n16028) );
  NOR2_X1 U18196 ( .A1(n16028), .A2(n12964), .ZN(n14918) );
  AOI21_X1 U18197 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n12964), .A(n14918), .ZN(
        n14919) );
  OAI21_X1 U18198 ( .B1(n14994), .B2(n14961), .A(n14919), .ZN(P2_U2861) );
  OAI21_X1 U18199 ( .B1(n14922), .B2(n14921), .A(n14920), .ZN(n15000) );
  NOR2_X1 U18200 ( .A1(n14890), .A2(n14923), .ZN(n14924) );
  AOI21_X1 U18201 ( .B1(n15256), .B2(n14890), .A(n14924), .ZN(n14925) );
  OAI21_X1 U18202 ( .B1(n15000), .B2(n14961), .A(n14925), .ZN(P2_U2862) );
  AOI21_X1 U18203 ( .B1(n14927), .B2(n14926), .A(n9712), .ZN(n14928) );
  XOR2_X1 U18204 ( .A(n14929), .B(n14928), .Z(n15009) );
  OAI21_X1 U18205 ( .B1(n14931), .B2(n14930), .A(n9662), .ZN(n16046) );
  MUX2_X1 U18206 ( .A(n14932), .B(n16046), .S(n14890), .Z(n14933) );
  OAI21_X1 U18207 ( .B1(n15009), .B2(n14961), .A(n14933), .ZN(P2_U2863) );
  AOI21_X1 U18208 ( .B1(n14936), .B2(n14935), .A(n14934), .ZN(n14937) );
  INV_X1 U18209 ( .A(n14937), .ZN(n15017) );
  MUX2_X1 U18210 ( .A(n15280), .B(n10535), .S(n14946), .Z(n14938) );
  OAI21_X1 U18211 ( .B1(n15017), .B2(n14961), .A(n14938), .ZN(P2_U2864) );
  AND2_X1 U18212 ( .A1(n9676), .A2(n14939), .ZN(n14941) );
  OR2_X1 U18213 ( .A1(n14941), .A2(n14940), .ZN(n16072) );
  AOI21_X1 U18214 ( .B1(n14944), .B2(n14943), .A(n14942), .ZN(n16054) );
  NAND2_X1 U18215 ( .A1(n16054), .A2(n14945), .ZN(n14948) );
  NAND2_X1 U18216 ( .A1(n14946), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14947) );
  OAI211_X1 U18217 ( .C1(n16072), .C2(n12964), .A(n14948), .B(n14947), .ZN(
        P2_U2865) );
  NAND2_X1 U18218 ( .A1(n14956), .A2(n14949), .ZN(n14950) );
  NAND2_X1 U18219 ( .A1(n9676), .A2(n14950), .ZN(n18780) );
  NOR2_X1 U18220 ( .A1(n18780), .A2(n12964), .ZN(n14951) );
  AOI21_X1 U18221 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n12964), .A(n14951), .ZN(
        n14952) );
  OAI21_X1 U18222 ( .B1(n14953), .B2(n14961), .A(n14952), .ZN(P2_U2866) );
  NOR2_X1 U18223 ( .A1(n9655), .A2(n14954), .ZN(n14955) );
  OR2_X1 U18224 ( .A1(n13830), .A2(n14955), .ZN(n16059) );
  OAI21_X1 U18225 ( .B1(n14958), .B2(n14957), .A(n14956), .ZN(n15318) );
  NOR2_X1 U18226 ( .A1(n15318), .A2(n12964), .ZN(n14959) );
  AOI21_X1 U18227 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n12964), .A(n14959), .ZN(
        n14960) );
  OAI21_X1 U18228 ( .B1(n16059), .B2(n14961), .A(n14960), .ZN(P2_U2867) );
  INV_X1 U18229 ( .A(n18978), .ZN(n18986) );
  NAND3_X1 U18230 ( .A1(n14962), .A2(n14895), .A3(n18986), .ZN(n14969) );
  OAI22_X1 U18231 ( .A1(n14964), .A2(n18967), .B1(n18966), .B2(n14963), .ZN(
        n14965) );
  AOI21_X1 U18232 ( .B1(n16065), .B2(n14966), .A(n14965), .ZN(n14968) );
  AOI22_X1 U18233 ( .A1(n18940), .A2(BUF2_REG_29__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14967) );
  NAND3_X1 U18234 ( .A1(n14969), .A2(n14968), .A3(n14967), .ZN(P2_U2890) );
  INV_X1 U18235 ( .A(n15217), .ZN(n14973) );
  OAI22_X1 U18236 ( .A1(n15013), .A2(n14971), .B1(n18966), .B2(n14970), .ZN(
        n14972) );
  AOI21_X1 U18237 ( .B1(n18984), .B2(n14973), .A(n14972), .ZN(n14975) );
  AOI22_X1 U18238 ( .A1(n18940), .A2(BUF2_REG_28__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14974) );
  OAI211_X1 U18239 ( .C1(n14976), .C2(n18978), .A(n14975), .B(n14974), .ZN(
        P2_U2891) );
  INV_X1 U18240 ( .A(n14990), .ZN(n14980) );
  INV_X1 U18241 ( .A(n14977), .ZN(n14979) );
  OAI21_X1 U18242 ( .B1(n14980), .B2(n14979), .A(n14978), .ZN(n16026) );
  OAI22_X1 U18243 ( .A1(n16026), .A2(n18967), .B1(n18966), .B2(n14981), .ZN(
        n14982) );
  AOI21_X1 U18244 ( .B1(n16065), .B2(n14983), .A(n14982), .ZN(n14985) );
  AOI22_X1 U18245 ( .A1(n18940), .A2(BUF2_REG_27__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14984) );
  OAI211_X1 U18246 ( .C1(n14986), .C2(n18978), .A(n14985), .B(n14984), .ZN(
        P2_U2892) );
  OR2_X1 U18247 ( .A1(n14988), .A2(n14987), .ZN(n14989) );
  NAND2_X1 U18248 ( .A1(n14990), .A2(n14989), .ZN(n15236) );
  OAI22_X1 U18249 ( .A1(n15236), .A2(n18967), .B1(n18966), .B2(n12796), .ZN(
        n14991) );
  AOI21_X1 U18250 ( .B1(n16065), .B2(n18950), .A(n14991), .ZN(n14993) );
  AOI22_X1 U18251 ( .A1(n18940), .A2(BUF2_REG_26__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14992) );
  OAI211_X1 U18252 ( .C1(n14994), .C2(n18978), .A(n14993), .B(n14992), .ZN(
        P2_U2893) );
  OAI22_X1 U18253 ( .A1(n15248), .A2(n18967), .B1(n18966), .B2(n14995), .ZN(
        n14996) );
  AOI21_X1 U18254 ( .B1(n16065), .B2(n14997), .A(n14996), .ZN(n14999) );
  AOI22_X1 U18255 ( .A1(n18940), .A2(BUF2_REG_25__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14998) );
  OAI211_X1 U18256 ( .C1(n15000), .C2(n18978), .A(n14999), .B(n14998), .ZN(
        P2_U2894) );
  AOI21_X1 U18257 ( .B1(n15003), .B2(n15002), .A(n15001), .ZN(n16047) );
  INV_X1 U18258 ( .A(n16047), .ZN(n15005) );
  OAI22_X1 U18259 ( .A1(n15005), .A2(n18967), .B1(n18966), .B2(n15004), .ZN(
        n15006) );
  AOI21_X1 U18260 ( .B1(n16065), .B2(n18954), .A(n15006), .ZN(n15008) );
  AOI22_X1 U18261 ( .A1(n18940), .A2(BUF2_REG_24__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15007) );
  OAI211_X1 U18262 ( .C1(n15009), .C2(n18978), .A(n15008), .B(n15007), .ZN(
        P2_U2895) );
  INV_X1 U18263 ( .A(n15010), .ZN(n15277) );
  OAI22_X1 U18264 ( .A1(n15013), .A2(n15012), .B1(n18966), .B2(n15011), .ZN(
        n15014) );
  AOI21_X1 U18265 ( .B1(n18984), .B2(n15277), .A(n15014), .ZN(n15016) );
  AOI22_X1 U18266 ( .A1(n18940), .A2(BUF2_REG_23__SCAN_IN), .B1(n18938), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15015) );
  OAI211_X1 U18267 ( .C1(n15017), .C2(n18978), .A(n15016), .B(n15015), .ZN(
        P2_U2896) );
  INV_X1 U18268 ( .A(n15019), .ZN(n15021) );
  NAND2_X1 U18269 ( .A1(n15021), .A2(n15020), .ZN(n15022) );
  XNOR2_X1 U18270 ( .A(n15023), .B(n15022), .ZN(n15211) );
  XNOR2_X1 U18271 ( .A(n15025), .B(n15024), .ZN(n15209) );
  NOR2_X1 U18272 ( .A1(n18885), .A2(n15026), .ZN(n15203) );
  NOR2_X1 U18273 ( .A1(n19052), .A2(n16000), .ZN(n15027) );
  AOI211_X1 U18274 ( .C1(n19039), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15203), .B(n15027), .ZN(n15028) );
  OAI21_X1 U18275 ( .B1(n16006), .B2(n19047), .A(n15028), .ZN(n15029) );
  AOI21_X1 U18276 ( .B1(n15209), .B2(n19042), .A(n15029), .ZN(n15030) );
  OAI21_X1 U18277 ( .B1(n15211), .B2(n16134), .A(n15030), .ZN(P2_U2984) );
  NOR2_X1 U18278 ( .A1(n19052), .A2(n15031), .ZN(n15032) );
  AOI211_X1 U18279 ( .C1(n19039), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15033), .B(n15032), .ZN(n15034) );
  OAI21_X1 U18280 ( .B1(n15035), .B2(n19047), .A(n15034), .ZN(n15036) );
  AOI21_X1 U18281 ( .B1(n15037), .B2(n19042), .A(n15036), .ZN(n15038) );
  OAI21_X1 U18282 ( .B1(n15039), .B2(n16134), .A(n15038), .ZN(P2_U2985) );
  OAI21_X1 U18283 ( .B1(n15040), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15041), .ZN(n15224) );
  NAND2_X1 U18284 ( .A1(n15042), .A2(n9682), .ZN(n15044) );
  NAND2_X1 U18285 ( .A1(n16012), .A2(n15043), .ZN(n15045) );
  XNOR2_X1 U18286 ( .A(n15044), .B(n15045), .ZN(n15057) );
  INV_X1 U18287 ( .A(n15044), .ZN(n15046) );
  XOR2_X1 U18288 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15047), .Z(
        n15048) );
  XNOR2_X1 U18289 ( .A(n15049), .B(n15048), .ZN(n15212) );
  NAND2_X1 U18290 ( .A1(n15212), .A2(n19040), .ZN(n15055) );
  NAND2_X1 U18291 ( .A1(n15058), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15216) );
  OAI21_X1 U18292 ( .B1(n16151), .B2(n15050), .A(n15216), .ZN(n15052) );
  NOR2_X1 U18293 ( .A1(n15218), .A2(n19047), .ZN(n15051) );
  AOI211_X1 U18294 ( .C1(n16142), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15054) );
  OAI211_X1 U18295 ( .C1(n16133), .C2(n15224), .A(n15055), .B(n15054), .ZN(
        P2_U2986) );
  INV_X1 U18296 ( .A(n15040), .ZN(n15056) );
  OAI21_X1 U18297 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15068), .A(
        n15056), .ZN(n15235) );
  NAND3_X1 U18298 ( .A1(n15226), .A2(n15225), .A3(n19040), .ZN(n15063) );
  NAND2_X1 U18299 ( .A1(n16142), .A2(n16022), .ZN(n15059) );
  NAND2_X1 U18300 ( .A1(n15058), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15229) );
  OAI211_X1 U18301 ( .C1(n16151), .C2(n15060), .A(n15059), .B(n15229), .ZN(
        n15061) );
  AOI21_X1 U18302 ( .B1(n16018), .B2(n16137), .A(n15061), .ZN(n15062) );
  OAI211_X1 U18303 ( .C1(n16133), .C2(n15235), .A(n15063), .B(n15062), .ZN(
        P2_U2987) );
  INV_X1 U18304 ( .A(n15065), .ZN(n15077) );
  NOR2_X1 U18305 ( .A1(n15064), .A2(n15077), .ZN(n15066) );
  XOR2_X1 U18306 ( .A(n15067), .B(n15066), .Z(n15247) );
  INV_X1 U18307 ( .A(n15083), .ZN(n15090) );
  NAND2_X1 U18308 ( .A1(n15090), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15258) );
  AOI21_X1 U18309 ( .B1(n15241), .B2(n15258), .A(n15068), .ZN(n15245) );
  NOR2_X1 U18310 ( .A1(n18900), .A2(n19660), .ZN(n15237) );
  NOR2_X1 U18311 ( .A1(n19052), .A2(n15069), .ZN(n15070) );
  AOI211_X1 U18312 ( .C1(n19039), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15237), .B(n15070), .ZN(n15071) );
  OAI21_X1 U18313 ( .B1(n16028), .B2(n19047), .A(n15071), .ZN(n15072) );
  AOI21_X1 U18314 ( .B1(n15245), .B2(n19042), .A(n15072), .ZN(n15073) );
  OAI21_X1 U18315 ( .B1(n15247), .B2(n16134), .A(n15073), .ZN(P2_U2988) );
  INV_X1 U18316 ( .A(n15064), .ZN(n15078) );
  OAI21_X1 U18317 ( .B1(n15075), .B2(n15077), .A(n15074), .ZN(n15076) );
  OAI21_X1 U18318 ( .B1(n15078), .B2(n15077), .A(n15076), .ZN(n15261) );
  NAND2_X1 U18319 ( .A1(n16142), .A2(n15079), .ZN(n15080) );
  OR2_X1 U18320 ( .A1(n18900), .A2(n19658), .ZN(n15251) );
  OAI211_X1 U18321 ( .C1(n16151), .C2(n15081), .A(n15080), .B(n15251), .ZN(
        n15082) );
  AOI21_X1 U18322 ( .B1(n15256), .B2(n16137), .A(n15082), .ZN(n15085) );
  NAND2_X1 U18323 ( .A1(n15083), .A2(n15252), .ZN(n15257) );
  NAND3_X1 U18324 ( .A1(n15258), .A2(n19042), .A3(n15257), .ZN(n15084) );
  OAI211_X1 U18325 ( .C1(n15261), .C2(n16134), .A(n15085), .B(n15084), .ZN(
        P2_U2989) );
  NOR2_X1 U18326 ( .A1(n9722), .A2(n15086), .ZN(n15087) );
  XNOR2_X1 U18327 ( .A(n15088), .B(n15087), .ZN(n15272) );
  AOI21_X1 U18328 ( .B1(n15262), .B2(n15089), .A(n15090), .ZN(n15270) );
  INV_X1 U18329 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19656) );
  NOR2_X1 U18330 ( .A1(n18885), .A2(n19656), .ZN(n15266) );
  NOR2_X1 U18331 ( .A1(n19052), .A2(n15091), .ZN(n15092) );
  AOI211_X1 U18332 ( .C1(n19039), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15266), .B(n15092), .ZN(n15093) );
  OAI21_X1 U18333 ( .B1(n16046), .B2(n19047), .A(n15093), .ZN(n15094) );
  AOI21_X1 U18334 ( .B1(n15270), .B2(n19042), .A(n15094), .ZN(n15095) );
  OAI21_X1 U18335 ( .B1(n15272), .B2(n16134), .A(n15095), .ZN(P2_U2990) );
  OAI21_X1 U18336 ( .B1(n9656), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15089), .ZN(n15290) );
  NOR2_X1 U18337 ( .A1(n15096), .A2(n15097), .ZN(n15287) );
  NOR2_X1 U18338 ( .A1(n15287), .A2(n16134), .ZN(n15103) );
  INV_X1 U18339 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19654) );
  OAI22_X1 U18340 ( .A1(n16151), .A2(n10246), .B1(n19654), .B2(n18900), .ZN(
        n15099) );
  AOI21_X1 U18341 ( .B1(n16142), .B2(n15100), .A(n15099), .ZN(n15101) );
  OAI21_X1 U18342 ( .B1(n15280), .B2(n19047), .A(n15101), .ZN(n15102) );
  AOI21_X1 U18343 ( .B1(n15103), .B2(n15098), .A(n15102), .ZN(n15104) );
  OAI21_X1 U18344 ( .B1(n15290), .B2(n16133), .A(n15104), .ZN(P2_U2991) );
  NAND2_X1 U18345 ( .A1(n15188), .A2(n15189), .ZN(n15187) );
  INV_X1 U18346 ( .A(n15107), .ZN(n16081) );
  INV_X1 U18347 ( .A(n15109), .ZN(n15155) );
  OAI21_X1 U18348 ( .B1(n15385), .B2(n15110), .A(n15155), .ZN(n15147) );
  INV_X1 U18349 ( .A(n15135), .ZN(n15112) );
  INV_X1 U18350 ( .A(n15120), .ZN(n15113) );
  AOI21_X1 U18351 ( .B1(n15306), .B2(n15126), .A(n15114), .ZN(n15315) );
  NOR2_X1 U18352 ( .A1(n18885), .A2(n19651), .ZN(n15308) );
  NOR2_X1 U18353 ( .A1(n16151), .A2(n15115), .ZN(n15116) );
  AOI211_X1 U18354 ( .C1(n18784), .C2(n16142), .A(n15308), .B(n15116), .ZN(
        n15117) );
  OAI21_X1 U18355 ( .B1(n18780), .B2(n19047), .A(n15117), .ZN(n15118) );
  AOI21_X1 U18356 ( .B1(n15315), .B2(n19042), .A(n15118), .ZN(n15119) );
  OAI21_X1 U18357 ( .B1(n15317), .B2(n16134), .A(n15119), .ZN(P2_U2993) );
  NAND2_X1 U18358 ( .A1(n15121), .A2(n15120), .ZN(n15122) );
  XNOR2_X1 U18359 ( .A(n15123), .B(n15122), .ZN(n15341) );
  INV_X1 U18360 ( .A(n15327), .ZN(n15125) );
  INV_X1 U18361 ( .A(n15126), .ZN(n15127) );
  NOR2_X1 U18362 ( .A1(n18885), .A2(n15128), .ZN(n15323) );
  NOR2_X1 U18363 ( .A1(n19052), .A2(n15129), .ZN(n15130) );
  AOI211_X1 U18364 ( .C1(n19039), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15323), .B(n15130), .ZN(n15131) );
  OAI21_X1 U18365 ( .B1(n15318), .B2(n19047), .A(n15131), .ZN(n15132) );
  AOI21_X1 U18366 ( .B1(n15338), .B2(n19042), .A(n15132), .ZN(n15133) );
  OAI21_X1 U18367 ( .B1(n15341), .B2(n16134), .A(n15133), .ZN(P2_U2994) );
  NAND2_X1 U18368 ( .A1(n15134), .A2(n15145), .ZN(n15138) );
  NAND2_X1 U18369 ( .A1(n15136), .A2(n15135), .ZN(n15137) );
  XNOR2_X1 U18370 ( .A(n15138), .B(n15137), .ZN(n15354) );
  AOI21_X1 U18371 ( .B1(n15349), .B2(n15139), .A(n9695), .ZN(n15352) );
  NOR2_X1 U18372 ( .A1(n18885), .A2(n19648), .ZN(n15342) );
  AOI21_X1 U18373 ( .B1(n19039), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15342), .ZN(n15141) );
  NAND2_X1 U18374 ( .A1(n18808), .A2(n16142), .ZN(n15140) );
  OAI211_X1 U18375 ( .C1(n18806), .C2(n19047), .A(n15141), .B(n15140), .ZN(
        n15142) );
  AOI21_X1 U18376 ( .B1(n15352), .B2(n19042), .A(n15142), .ZN(n15143) );
  OAI21_X1 U18377 ( .B1(n16134), .B2(n15354), .A(n15143), .ZN(P2_U2995) );
  NAND2_X1 U18378 ( .A1(n15145), .A2(n15144), .ZN(n15146) );
  XNOR2_X1 U18379 ( .A(n15147), .B(n15146), .ZN(n15369) );
  AOI21_X1 U18380 ( .B1(n15358), .B2(n15162), .A(n15148), .ZN(n15367) );
  NOR2_X1 U18381 ( .A1(n18885), .A2(n19646), .ZN(n15356) );
  AOI21_X1 U18382 ( .B1(n19039), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15356), .ZN(n15151) );
  NAND2_X1 U18383 ( .A1(n15149), .A2(n16142), .ZN(n15150) );
  OAI211_X1 U18384 ( .C1(n15365), .C2(n19047), .A(n15151), .B(n15150), .ZN(
        n15152) );
  AOI21_X1 U18385 ( .B1(n15367), .B2(n19042), .A(n15152), .ZN(n15153) );
  OAI21_X1 U18386 ( .B1(n16134), .B2(n15369), .A(n15153), .ZN(P2_U2996) );
  NAND2_X1 U18387 ( .A1(n15155), .A2(n15154), .ZN(n15159) );
  INV_X1 U18388 ( .A(n15385), .ZN(n15157) );
  NAND2_X1 U18389 ( .A1(n15157), .A2(n15156), .ZN(n15158) );
  XOR2_X1 U18390 ( .A(n15159), .B(n15158), .Z(n15382) );
  NOR2_X1 U18391 ( .A1(n18885), .A2(n19644), .ZN(n15376) );
  AOI21_X1 U18392 ( .B1(n19039), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15376), .ZN(n15160) );
  OAI21_X1 U18393 ( .B1(n19052), .B2(n18826), .A(n15160), .ZN(n15161) );
  AOI21_X1 U18394 ( .B1(n16137), .B2(n18823), .A(n15161), .ZN(n15164) );
  OAI211_X1 U18395 ( .C1(n15373), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15162), .B(n19042), .ZN(n15163) );
  OAI211_X1 U18396 ( .C1(n15382), .C2(n16134), .A(n15164), .B(n15163), .ZN(
        P2_U2997) );
  INV_X1 U18397 ( .A(n15389), .ZN(n16079) );
  AOI21_X1 U18398 ( .B1(n16079), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15172) );
  NAND2_X1 U18399 ( .A1(n10012), .A2(n19042), .ZN(n15171) );
  INV_X1 U18400 ( .A(n18834), .ZN(n15388) );
  NAND2_X1 U18401 ( .A1(n15058), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15383) );
  NAND2_X1 U18402 ( .A1(n19039), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15165) );
  OAI211_X1 U18403 ( .C1(n19052), .C2(n18832), .A(n15383), .B(n15165), .ZN(
        n15169) );
  AND2_X1 U18404 ( .A1(n15167), .A2(n15166), .ZN(n15384) );
  NOR3_X1 U18405 ( .A1(n15385), .A2(n15384), .A3(n16134), .ZN(n15168) );
  AOI211_X1 U18406 ( .C1(n15388), .C2(n16137), .A(n15169), .B(n15168), .ZN(
        n15170) );
  OAI21_X1 U18407 ( .B1(n15172), .B2(n15171), .A(n15170), .ZN(P2_U2998) );
  XNOR2_X1 U18408 ( .A(n15389), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16160) );
  INV_X1 U18409 ( .A(n15173), .ZN(n16082) );
  OR2_X1 U18410 ( .A1(n15174), .A2(n16082), .ZN(n15178) );
  AND2_X1 U18411 ( .A1(n15176), .A2(n15175), .ZN(n15177) );
  XNOR2_X1 U18412 ( .A(n15178), .B(n15177), .ZN(n16163) );
  AOI22_X1 U18413 ( .A1(n16159), .A2(n16137), .B1(P2_REIP_REG_15__SCAN_IN), 
        .B2(n15058), .ZN(n15183) );
  OAI22_X1 U18414 ( .A1(n16151), .A2(n15180), .B1(n19052), .B2(n15179), .ZN(
        n15181) );
  INV_X1 U18415 ( .A(n15181), .ZN(n15182) );
  OAI211_X1 U18416 ( .C1(n16163), .C2(n16134), .A(n15183), .B(n15182), .ZN(
        n15184) );
  AOI21_X1 U18417 ( .B1(n19042), .B2(n16160), .A(n15184), .ZN(n15185) );
  INV_X1 U18418 ( .A(n15185), .ZN(P2_U2999) );
  NOR2_X1 U18419 ( .A1(n15423), .A2(n15418), .ZN(n15407) );
  INV_X1 U18420 ( .A(n15186), .ZN(n16080) );
  OAI21_X1 U18421 ( .B1(n15407), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16080), .ZN(n15406) );
  INV_X1 U18422 ( .A(n15187), .ZN(n15192) );
  AOI21_X1 U18423 ( .B1(n15191), .B2(n15189), .A(n15188), .ZN(n15190) );
  AOI21_X1 U18424 ( .B1(n15192), .B2(n15191), .A(n15190), .ZN(n15401) );
  INV_X1 U18425 ( .A(n15401), .ZN(n15198) );
  OAI22_X1 U18426 ( .A1(n16151), .A2(n15193), .B1(n20932), .B2(n18885), .ZN(
        n15197) );
  OAI22_X1 U18427 ( .A1(n15195), .A2(n19047), .B1(n19052), .B2(n15194), .ZN(
        n15196) );
  AOI211_X1 U18428 ( .C1(n15198), .C2(n19040), .A(n15197), .B(n15196), .ZN(
        n15199) );
  OAI21_X1 U18429 ( .B1(n16133), .B2(n15406), .A(n15199), .ZN(P2_U3001) );
  INV_X1 U18430 ( .A(n16005), .ZN(n15204) );
  NOR3_X1 U18431 ( .A1(n15201), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15200), .ZN(n15202) );
  NAND2_X1 U18432 ( .A1(n15205), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15206) );
  OAI211_X1 U18433 ( .C1(n16006), .C2(n16188), .A(n15207), .B(n15206), .ZN(
        n15208) );
  AOI21_X1 U18434 ( .B1(n15209), .B2(n19056), .A(n15208), .ZN(n15210) );
  OAI21_X1 U18435 ( .B1(n15211), .B2(n16204), .A(n15210), .ZN(P2_U3016) );
  NAND2_X1 U18436 ( .A1(n15212), .A2(n19065), .ZN(n15223) );
  NAND3_X1 U18437 ( .A1(n15214), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15213), .ZN(n15215) );
  OAI211_X1 U18438 ( .C1(n19070), .C2(n15217), .A(n15216), .B(n15215), .ZN(
        n15220) );
  NOR2_X1 U18439 ( .A1(n15218), .A2(n16188), .ZN(n15219) );
  AOI211_X1 U18440 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15221), .A(
        n15220), .B(n15219), .ZN(n15222) );
  OAI211_X1 U18441 ( .C1(n15224), .C2(n16189), .A(n15223), .B(n15222), .ZN(
        P2_U3018) );
  NAND3_X1 U18442 ( .A1(n15226), .A2(n15225), .A3(n19065), .ZN(n15234) );
  NOR2_X1 U18443 ( .A1(n15228), .A2(n15227), .ZN(n15232) );
  OAI211_X1 U18444 ( .C1(n19070), .C2(n16026), .A(n15230), .B(n15229), .ZN(
        n15231) );
  AOI211_X1 U18445 ( .C1(n16018), .C2(n19067), .A(n15232), .B(n15231), .ZN(
        n15233) );
  OAI211_X1 U18446 ( .C1(n15235), .C2(n16189), .A(n15234), .B(n15233), .ZN(
        P2_U3019) );
  INV_X1 U18447 ( .A(n15236), .ZN(n16029) );
  INV_X1 U18448 ( .A(n15237), .ZN(n15240) );
  OAI211_X1 U18449 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15249), .B(n15238), .ZN(
        n15239) );
  OAI211_X1 U18450 ( .C1(n15253), .C2(n15241), .A(n15240), .B(n15239), .ZN(
        n15242) );
  AOI21_X1 U18451 ( .B1(n16200), .B2(n16029), .A(n15242), .ZN(n15243) );
  OAI21_X1 U18452 ( .B1(n16028), .B2(n16188), .A(n15243), .ZN(n15244) );
  AOI21_X1 U18453 ( .B1(n15245), .B2(n19056), .A(n15244), .ZN(n15246) );
  OAI21_X1 U18454 ( .B1(n15247), .B2(n16204), .A(n15246), .ZN(P2_U3020) );
  NOR2_X1 U18455 ( .A1(n19070), .A2(n15248), .ZN(n15255) );
  NAND2_X1 U18456 ( .A1(n15249), .A2(n15252), .ZN(n15250) );
  OAI211_X1 U18457 ( .C1(n15253), .C2(n15252), .A(n15251), .B(n15250), .ZN(
        n15254) );
  AOI211_X1 U18458 ( .C1(n15256), .C2(n19067), .A(n15255), .B(n15254), .ZN(
        n15260) );
  NAND3_X1 U18459 ( .A1(n15258), .A2(n19056), .A3(n15257), .ZN(n15259) );
  OAI211_X1 U18460 ( .C1(n15261), .C2(n16204), .A(n15260), .B(n15259), .ZN(
        P2_U3021) );
  INV_X1 U18461 ( .A(n15276), .ZN(n15297) );
  OAI21_X1 U18462 ( .B1(n15263), .B2(n15297), .A(n15262), .ZN(n15264) );
  NAND2_X1 U18463 ( .A1(n15265), .A2(n15264), .ZN(n15268) );
  AOI21_X1 U18464 ( .B1(n16200), .B2(n16047), .A(n15266), .ZN(n15267) );
  OAI211_X1 U18465 ( .C1(n16046), .C2(n16188), .A(n15268), .B(n15267), .ZN(
        n15269) );
  AOI21_X1 U18466 ( .B1(n15270), .B2(n19056), .A(n15269), .ZN(n15271) );
  OAI21_X1 U18467 ( .B1(n15272), .B2(n16204), .A(n15271), .ZN(P2_U3022) );
  AOI21_X1 U18468 ( .B1(n15283), .B2(n15296), .A(n15273), .ZN(n15275) );
  NOR2_X1 U18469 ( .A1(n19654), .A2(n18900), .ZN(n15274) );
  AOI21_X1 U18470 ( .B1(n15276), .B2(n15275), .A(n15274), .ZN(n15279) );
  NAND2_X1 U18471 ( .A1(n16200), .A2(n15277), .ZN(n15278) );
  OAI211_X1 U18472 ( .C1(n15280), .C2(n16188), .A(n15279), .B(n15278), .ZN(
        n15285) );
  NAND2_X1 U18473 ( .A1(n15468), .A2(n15281), .ZN(n15282) );
  AND2_X1 U18474 ( .A1(n15452), .A2(n15282), .ZN(n15307) );
  NOR2_X1 U18475 ( .A1(n15307), .A2(n15283), .ZN(n15284) );
  NOR2_X1 U18476 ( .A1(n15285), .A2(n15284), .ZN(n15289) );
  INV_X1 U18477 ( .A(n15098), .ZN(n15286) );
  OR3_X1 U18478 ( .A1(n15287), .A2(n15286), .A3(n16204), .ZN(n15288) );
  OAI211_X1 U18479 ( .C1(n15290), .C2(n16189), .A(n15289), .B(n15288), .ZN(
        P2_U3023) );
  NAND2_X1 U18480 ( .A1(n15292), .A2(n15291), .ZN(n15294) );
  XOR2_X1 U18481 ( .A(n15294), .B(n15293), .Z(n16073) );
  NOR2_X1 U18482 ( .A1(n15114), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16071) );
  OR3_X1 U18483 ( .A1(n16071), .A2(n9656), .A3(n16189), .ZN(n15305) );
  NAND2_X1 U18484 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n15058), .ZN(n15295) );
  OAI221_X1 U18485 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15297), 
        .C1(n15296), .C2(n15307), .A(n15295), .ZN(n15303) );
  OR2_X1 U18486 ( .A1(n15299), .A2(n15298), .ZN(n15300) );
  NAND2_X1 U18487 ( .A1(n15301), .A2(n15300), .ZN(n16052) );
  OAI22_X1 U18488 ( .A1(n16072), .A2(n16188), .B1(n19070), .B2(n16052), .ZN(
        n15302) );
  NOR2_X1 U18489 ( .A1(n15303), .A2(n15302), .ZN(n15304) );
  OAI211_X1 U18490 ( .C1(n16073), .C2(n16204), .A(n15305), .B(n15304), .ZN(
        P2_U3024) );
  NOR2_X1 U18491 ( .A1(n15307), .A2(n15306), .ZN(n15314) );
  NOR2_X1 U18492 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15433), .ZN(
        n15309) );
  AOI21_X1 U18493 ( .B1(n15310), .B2(n15309), .A(n15308), .ZN(n15312) );
  NAND2_X1 U18494 ( .A1(n16200), .A2(n18778), .ZN(n15311) );
  OAI211_X1 U18495 ( .C1(n18780), .C2(n16188), .A(n15312), .B(n15311), .ZN(
        n15313) );
  AOI211_X1 U18496 ( .C1(n15315), .C2(n19056), .A(n15314), .B(n15313), .ZN(
        n15316) );
  OAI21_X1 U18497 ( .B1(n15317), .B2(n16204), .A(n15316), .ZN(P2_U3025) );
  INV_X1 U18498 ( .A(n15318), .ZN(n18793) );
  NOR2_X1 U18499 ( .A1(n15320), .A2(n15319), .ZN(n15321) );
  OR2_X1 U18500 ( .A1(n15322), .A2(n15321), .ZN(n18791) );
  INV_X1 U18501 ( .A(n15323), .ZN(n15326) );
  NOR2_X1 U18502 ( .A1(n15327), .A2(n15433), .ZN(n16169) );
  NAND3_X1 U18503 ( .A1(n16153), .A2(n15324), .A3(n15335), .ZN(n15325) );
  OAI211_X1 U18504 ( .C1(n19070), .C2(n18791), .A(n15326), .B(n15325), .ZN(
        n15337) );
  NAND2_X1 U18505 ( .A1(n15468), .A2(n15327), .ZN(n15328) );
  NAND2_X1 U18506 ( .A1(n15452), .A2(n15328), .ZN(n15396) );
  INV_X1 U18507 ( .A(n15329), .ZN(n15330) );
  AND2_X1 U18508 ( .A1(n15468), .A2(n15330), .ZN(n15331) );
  OR2_X1 U18509 ( .A1(n15396), .A2(n15331), .ZN(n16158) );
  AND2_X1 U18510 ( .A1(n15468), .A2(n15357), .ZN(n15332) );
  OR2_X1 U18511 ( .A1(n16158), .A2(n15332), .ZN(n15355) );
  AOI21_X1 U18512 ( .B1(n15358), .B2(n15468), .A(n15355), .ZN(n15350) );
  NAND2_X1 U18513 ( .A1(n15349), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15333) );
  NOR2_X1 U18514 ( .A1(n15357), .A2(n15333), .ZN(n15334) );
  NAND2_X1 U18515 ( .A1(n16153), .A2(n15334), .ZN(n15343) );
  AOI21_X1 U18516 ( .B1(n15350), .B2(n15343), .A(n15335), .ZN(n15336) );
  AOI211_X1 U18517 ( .C1(n18793), .C2(n19067), .A(n15337), .B(n15336), .ZN(
        n15340) );
  NAND2_X1 U18518 ( .A1(n15338), .A2(n19056), .ZN(n15339) );
  OAI211_X1 U18519 ( .C1(n15341), .C2(n16204), .A(n15340), .B(n15339), .ZN(
        P2_U3026) );
  INV_X1 U18520 ( .A(n15342), .ZN(n15344) );
  NAND2_X1 U18521 ( .A1(n15344), .A2(n15343), .ZN(n15346) );
  NOR2_X1 U18522 ( .A1(n18806), .A2(n16188), .ZN(n15345) );
  AOI211_X1 U18523 ( .C1(n16200), .C2(n15347), .A(n15346), .B(n15345), .ZN(
        n15348) );
  OAI21_X1 U18524 ( .B1(n15350), .B2(n15349), .A(n15348), .ZN(n15351) );
  AOI21_X1 U18525 ( .B1(n15352), .B2(n19056), .A(n15351), .ZN(n15353) );
  OAI21_X1 U18526 ( .B1(n16204), .B2(n15354), .A(n15353), .ZN(P2_U3027) );
  NAND2_X1 U18527 ( .A1(n15355), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15364) );
  INV_X1 U18528 ( .A(n15356), .ZN(n15361) );
  INV_X1 U18529 ( .A(n15357), .ZN(n15359) );
  NAND3_X1 U18530 ( .A1(n16153), .A2(n15359), .A3(n15358), .ZN(n15360) );
  NAND2_X1 U18531 ( .A1(n15361), .A2(n15360), .ZN(n15362) );
  AOI21_X1 U18532 ( .B1(n16200), .B2(n16066), .A(n15362), .ZN(n15363) );
  OAI211_X1 U18533 ( .C1(n15365), .C2(n16188), .A(n15364), .B(n15363), .ZN(
        n15366) );
  AOI21_X1 U18534 ( .B1(n15367), .B2(n19056), .A(n15366), .ZN(n15368) );
  OAI21_X1 U18535 ( .B1(n16204), .B2(n15369), .A(n15368), .ZN(P2_U3028) );
  INV_X1 U18536 ( .A(n19059), .ZN(n15371) );
  OAI21_X1 U18537 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16209), .A(
        n15394), .ZN(n15380) );
  AOI22_X1 U18538 ( .A1(n15373), .A2(n19056), .B1(n15372), .B2(n16153), .ZN(
        n15378) );
  NOR2_X1 U18539 ( .A1(n19070), .A2(n15374), .ZN(n15375) );
  AOI211_X1 U18540 ( .C1(n18823), .C2(n19067), .A(n15376), .B(n15375), .ZN(
        n15377) );
  OAI21_X1 U18541 ( .B1(n15378), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15377), .ZN(n15379) );
  AOI21_X1 U18542 ( .B1(n15380), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15379), .ZN(n15381) );
  OAI21_X1 U18543 ( .B1(n15382), .B2(n16204), .A(n15381), .ZN(P2_U3029) );
  OAI21_X1 U18544 ( .B1(n19070), .B2(n18833), .A(n15383), .ZN(n15387) );
  NOR3_X1 U18545 ( .A1(n15385), .A2(n15384), .A3(n16204), .ZN(n15386) );
  AOI211_X1 U18546 ( .C1(n19067), .C2(n15388), .A(n15387), .B(n15386), .ZN(
        n15392) );
  NOR2_X1 U18547 ( .A1(n15389), .A2(n16189), .ZN(n15390) );
  OAI211_X1 U18548 ( .C1(n15390), .C2(n16153), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n15393), .ZN(n15391) );
  OAI211_X1 U18549 ( .C1(n15394), .C2(n15393), .A(n15392), .B(n15391), .ZN(
        P2_U3030) );
  INV_X1 U18550 ( .A(n16169), .ZN(n15415) );
  OAI21_X1 U18551 ( .B1(n15418), .B2(n15415), .A(n15395), .ZN(n15404) );
  INV_X1 U18552 ( .A(n15396), .ZN(n15419) );
  OAI21_X1 U18553 ( .B1(n16170), .B2(n15415), .A(n15419), .ZN(n16164) );
  AOI22_X1 U18554 ( .A1(n15398), .A2(n19067), .B1(n15397), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n15399) );
  OAI21_X1 U18555 ( .B1(n19070), .B2(n15400), .A(n15399), .ZN(n15403) );
  NOR2_X1 U18556 ( .A1(n15401), .A2(n16204), .ZN(n15402) );
  AOI211_X1 U18557 ( .C1(n15404), .C2(n16164), .A(n15403), .B(n15402), .ZN(
        n15405) );
  OAI21_X1 U18558 ( .B1(n16189), .B2(n15406), .A(n15405), .ZN(P2_U3033) );
  AOI21_X1 U18559 ( .B1(n15418), .B2(n15423), .A(n15407), .ZN(n16088) );
  INV_X1 U18560 ( .A(n16088), .ZN(n15422) );
  OR2_X1 U18561 ( .A1(n15409), .A2(n9827), .ZN(n15410) );
  XNOR2_X1 U18562 ( .A(n15411), .B(n15410), .ZN(n16090) );
  INV_X1 U18563 ( .A(n15412), .ZN(n16089) );
  NAND2_X1 U18564 ( .A1(n16200), .A2(n18946), .ZN(n15414) );
  NAND2_X1 U18565 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n15058), .ZN(n15413) );
  OAI211_X1 U18566 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15415), .A(
        n15414), .B(n15413), .ZN(n15416) );
  AOI21_X1 U18567 ( .B1(n19067), .B2(n16089), .A(n15416), .ZN(n15417) );
  OAI21_X1 U18568 ( .B1(n15419), .B2(n15418), .A(n15417), .ZN(n15420) );
  AOI21_X1 U18569 ( .B1(n16090), .B2(n19065), .A(n15420), .ZN(n15421) );
  OAI21_X1 U18570 ( .B1(n15422), .B2(n16189), .A(n15421), .ZN(P2_U3034) );
  NAND2_X1 U18571 ( .A1(n15124), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16100) );
  NOR2_X1 U18572 ( .A1(n16100), .A2(n12109), .ZN(n16099) );
  OAI21_X1 U18573 ( .B1(n16099), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15423), .ZN(n16095) );
  INV_X1 U18574 ( .A(n15424), .ZN(n15425) );
  NAND2_X1 U18575 ( .A1(n15426), .A2(n15425), .ZN(n15430) );
  NOR2_X1 U18576 ( .A1(n15428), .A2(n15427), .ZN(n15429) );
  XNOR2_X1 U18577 ( .A(n15430), .B(n15429), .ZN(n16094) );
  INV_X1 U18578 ( .A(n15431), .ZN(n15432) );
  AOI21_X1 U18579 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15452), .A(
        n15432), .ZN(n16180) );
  INV_X1 U18580 ( .A(n15433), .ZN(n15456) );
  NAND2_X1 U18581 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15456), .ZN(
        n16177) );
  AOI221_X1 U18582 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n12109), .C2(n15434), .A(
        n16177), .ZN(n15436) );
  NOR2_X1 U18583 ( .A1(n10781), .A2(n18900), .ZN(n15435) );
  AOI211_X1 U18584 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16180), .A(
        n15436), .B(n15435), .ZN(n15439) );
  INV_X1 U18585 ( .A(n18845), .ZN(n15437) );
  AOI22_X1 U18586 ( .A1(n19067), .A2(n18844), .B1(n16200), .B2(n15437), .ZN(
        n15438) );
  OAI211_X1 U18587 ( .C1(n16094), .C2(n16204), .A(n15439), .B(n15438), .ZN(
        n15440) );
  INV_X1 U18588 ( .A(n15440), .ZN(n15441) );
  OAI21_X1 U18589 ( .B1(n16095), .B2(n16189), .A(n15441), .ZN(P2_U3035) );
  OAI21_X1 U18590 ( .B1(n15124), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16100), .ZN(n16112) );
  INV_X1 U18591 ( .A(n15442), .ZN(n15444) );
  OAI21_X1 U18592 ( .B1(n16123), .B2(n15444), .A(n15443), .ZN(n15447) );
  NAND2_X1 U18593 ( .A1(n16101), .A2(n15445), .ZN(n15446) );
  NAND2_X1 U18594 ( .A1(n15447), .A2(n15446), .ZN(n15451) );
  INV_X1 U18595 ( .A(n16101), .ZN(n15449) );
  OR2_X1 U18596 ( .A1(n15448), .A2(n15449), .ZN(n15450) );
  NAND2_X1 U18597 ( .A1(n15451), .A2(n15450), .ZN(n16111) );
  INV_X1 U18598 ( .A(n15452), .ZN(n15454) );
  NOR2_X1 U18599 ( .A1(n10755), .A2(n18885), .ZN(n15453) );
  AOI221_X1 U18600 ( .B1(n15456), .B2(n15455), .C1(n15454), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15453), .ZN(n15459) );
  OAI22_X1 U18601 ( .A1(n18867), .A2(n16188), .B1(n19070), .B2(n18866), .ZN(
        n15457) );
  INV_X1 U18602 ( .A(n15457), .ZN(n15458) );
  OAI211_X1 U18603 ( .C1(n16111), .C2(n16204), .A(n15459), .B(n15458), .ZN(
        n15460) );
  INV_X1 U18604 ( .A(n15460), .ZN(n15461) );
  OAI21_X1 U18605 ( .B1(n16112), .B2(n16189), .A(n15461), .ZN(P2_U3037) );
  INV_X1 U18606 ( .A(n19057), .ZN(n15463) );
  AOI22_X1 U18607 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15463), .B1(
        n15462), .B2(n19067), .ZN(n15472) );
  AOI22_X1 U18608 ( .A1(n15465), .A2(n19065), .B1(n19056), .B2(n15464), .ZN(
        n15471) );
  INV_X1 U18609 ( .A(n15466), .ZN(n19703) );
  AOI21_X1 U18610 ( .B1(n16200), .B2(n19703), .A(n15467), .ZN(n15470) );
  OAI211_X1 U18611 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15468), .B(n19063), .ZN(n15469) );
  NAND4_X1 U18612 ( .A1(n15472), .A2(n15471), .A3(n15470), .A4(n15469), .ZN(
        P2_U3045) );
  INV_X1 U18613 ( .A(n16215), .ZN(n15476) );
  OAI222_X1 U18614 ( .A1(n15476), .A2(n15475), .B1(n19680), .B2(n15474), .C1(
        n13528), .C2(n15473), .ZN(n15478) );
  MUX2_X1 U18615 ( .A(n15478), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15477), .Z(P2_U3601) );
  NOR2_X1 U18616 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18679), .ZN(
        n18122) );
  INV_X1 U18617 ( .A(n18122), .ZN(n15481) );
  INV_X1 U18618 ( .A(n18588), .ZN(n18677) );
  NOR2_X1 U18619 ( .A1(n15479), .A2(n9633), .ZN(n18070) );
  OAI211_X1 U18620 ( .C1(n18677), .C2(n18070), .A(n18426), .B(n15480), .ZN(
        n18076) );
  NAND2_X1 U18621 ( .A1(n15481), .A2(n18076), .ZN(n15484) );
  INV_X1 U18622 ( .A(n15484), .ZN(n15483) );
  NAND3_X1 U18623 ( .A1(n18742), .A2(n18679), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18324) );
  NAND2_X1 U18624 ( .A1(n18742), .A2(n18679), .ZN(n16402) );
  AND2_X1 U18625 ( .A1(n18683), .A2(n16402), .ZN(n18726) );
  INV_X1 U18626 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18731) );
  NOR2_X1 U18627 ( .A1(n18688), .A2(n18731), .ZN(n17532) );
  INV_X1 U18628 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18540) );
  OAI22_X1 U18629 ( .A1(n18726), .A2(n17532), .B1(n18540), .B2(n18679), .ZN(
        n15486) );
  NAND3_X1 U18630 ( .A1(n18541), .A2(n18076), .A3(n15486), .ZN(n15482) );
  OAI221_X1 U18631 ( .B1(n18541), .B2(n15483), .C1(n18541), .C2(n18324), .A(
        n15482), .ZN(P3_U2864) );
  NAND2_X1 U18632 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18253) );
  NOR2_X1 U18633 ( .A1(n18726), .A2(n17532), .ZN(n15485) );
  AOI221_X1 U18634 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18253), .C1(n15485), 
        .C2(n18253), .A(n15484), .ZN(n18075) );
  INV_X1 U18635 ( .A(n18324), .ZN(n18370) );
  OAI221_X1 U18636 ( .B1(n18370), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18370), .C2(n15486), .A(n18076), .ZN(n18073) );
  AOI22_X1 U18637 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18075), .B1(
        n18073), .B2(n18561), .ZN(P3_U2865) );
  AOI22_X1 U18638 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U18639 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15496) );
  AOI22_X1 U18640 ( .A1(n15509), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15488) );
  OAI21_X1 U18641 ( .B1(n16832), .B2(n20943), .A(n15488), .ZN(n15494) );
  AOI22_X1 U18642 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15492) );
  AOI22_X1 U18643 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15491) );
  AOI22_X1 U18644 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U18645 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15489) );
  NAND4_X1 U18646 ( .A1(n15492), .A2(n15491), .A3(n15490), .A4(n15489), .ZN(
        n15493) );
  AOI22_X1 U18647 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15501) );
  AOI22_X1 U18648 ( .A1(n13937), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18649 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15499) );
  AOI22_X1 U18650 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15498) );
  NAND4_X1 U18651 ( .A1(n15501), .A2(n15500), .A3(n15499), .A4(n15498), .ZN(
        n15508) );
  AOI22_X1 U18652 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U18653 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15505) );
  AOI22_X1 U18654 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U18655 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15502), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15503) );
  NAND4_X1 U18656 ( .A1(n15506), .A2(n15505), .A3(n15504), .A4(n15503), .ZN(
        n15507) );
  AOI22_X1 U18657 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U18658 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15512) );
  AOI22_X1 U18659 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U18660 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15510) );
  NAND4_X1 U18661 ( .A1(n15513), .A2(n15512), .A3(n15511), .A4(n15510), .ZN(
        n15519) );
  AOI22_X1 U18662 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15517) );
  AOI22_X1 U18663 ( .A1(n17040), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U18664 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15515) );
  AOI22_X1 U18665 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15514) );
  NAND4_X1 U18666 ( .A1(n15517), .A2(n15516), .A3(n15515), .A4(n15514), .ZN(
        n15518) );
  AOI22_X1 U18667 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15530) );
  AOI22_X1 U18668 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n15572), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15529) );
  AOI22_X1 U18669 ( .A1(n13885), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15520) );
  OAI21_X1 U18670 ( .B1(n15487), .B2(n20899), .A(n15520), .ZN(n15527) );
  AOI22_X1 U18671 ( .A1(n14087), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15525) );
  AOI22_X1 U18672 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15524) );
  AOI22_X1 U18673 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15523) );
  AOI22_X1 U18674 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15522) );
  NAND4_X1 U18675 ( .A1(n15525), .A2(n15524), .A3(n15523), .A4(n15522), .ZN(
        n15526) );
  AOI211_X1 U18676 ( .C1(n16976), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n15527), .B(n15526), .ZN(n15528) );
  NAND3_X1 U18677 ( .A1(n15530), .A2(n15529), .A3(n15528), .ZN(n17252) );
  AOI22_X1 U18678 ( .A1(n14087), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U18679 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13884), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15533) );
  AOI22_X1 U18680 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17040), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n15531), .ZN(n15532) );
  OAI211_X1 U18681 ( .C1(n17102), .C2(n15558), .A(n15533), .B(n15532), .ZN(
        n15543) );
  AOI22_X1 U18682 ( .A1(n14076), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13937), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15541) );
  AOI22_X1 U18683 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n15572), .B1(
        n14055), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15540) );
  AOI22_X1 U18684 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n15535), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n15534), .ZN(n15539) );
  AOI22_X1 U18685 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n15537), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15538) );
  NAND4_X1 U18686 ( .A1(n15541), .A2(n15540), .A3(n15539), .A4(n15538), .ZN(
        n15542) );
  AOI211_X1 U18687 ( .C1(n13910), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n15543), .B(n15542), .ZN(n15544) );
  NAND2_X1 U18688 ( .A1(n15545), .A2(n15544), .ZN(n15569) );
  NAND2_X1 U18689 ( .A1(n17252), .A2(n15569), .ZN(n15586) );
  AOI22_X1 U18690 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15555) );
  AOI22_X1 U18691 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15547) );
  AOI22_X1 U18692 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15546) );
  OAI211_X1 U18693 ( .C1(n15558), .C2(n17091), .A(n15547), .B(n15546), .ZN(
        n15553) );
  AOI22_X1 U18694 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15551) );
  AOI22_X1 U18695 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15550) );
  AOI22_X1 U18696 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15549) );
  AOI22_X1 U18697 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15548) );
  NAND4_X1 U18698 ( .A1(n15551), .A2(n15550), .A3(n15549), .A4(n15548), .ZN(
        n15552) );
  AOI211_X1 U18699 ( .C1(n15537), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n15553), .B(n15552), .ZN(n15554) );
  NAND2_X1 U18700 ( .A1(n15555), .A2(n15554), .ZN(n17244) );
  NAND2_X1 U18701 ( .A1(n15568), .A2(n17244), .ZN(n15589) );
  AOI22_X1 U18702 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15566) );
  AOI22_X1 U18703 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15557) );
  AOI22_X1 U18704 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15556) );
  OAI211_X1 U18705 ( .C1(n15558), .C2(n17084), .A(n15557), .B(n15556), .ZN(
        n15564) );
  AOI22_X1 U18706 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U18707 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15561) );
  AOI22_X1 U18708 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n15560) );
  AOI22_X1 U18709 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16976), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n15559) );
  NAND4_X1 U18710 ( .A1(n15562), .A2(n15561), .A3(n15560), .A4(n15559), .ZN(
        n15563) );
  AOI211_X1 U18711 ( .C1(n15536), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n15564), .B(n15563), .ZN(n15565) );
  NAND2_X1 U18712 ( .A1(n15566), .A2(n15565), .ZN(n17235) );
  INV_X1 U18713 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17776) );
  OAI21_X1 U18714 ( .B1(n15567), .B2(n16292), .A(n17648), .ZN(n15594) );
  XOR2_X1 U18715 ( .A(n17244), .B(n15568), .Z(n15587) );
  XOR2_X1 U18716 ( .A(n20898), .B(n15587), .Z(n17697) );
  NOR2_X1 U18717 ( .A1(n15583), .A2(n15584), .ZN(n15585) );
  INV_X1 U18718 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18689) );
  AOI22_X1 U18719 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15570) );
  OAI21_X1 U18720 ( .B1(n15558), .B2(n15571), .A(n15570), .ZN(n15578) );
  AOI22_X1 U18721 ( .A1(n14087), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15576) );
  AOI22_X1 U18722 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15575) );
  AOI22_X1 U18723 ( .A1(n14076), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15572), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U18724 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15534), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15573) );
  NAND4_X1 U18725 ( .A1(n15576), .A2(n15575), .A3(n15574), .A4(n15573), .ZN(
        n15577) );
  AOI211_X1 U18726 ( .C1(n17068), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n15578), .B(n15577), .ZN(n15581) );
  AOI22_X1 U18727 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U18728 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15579) );
  NAND3_X1 U18729 ( .A1(n15581), .A2(n15580), .A3(n15579), .ZN(n17744) );
  NOR2_X1 U18730 ( .A1(n17735), .A2(n17743), .ZN(n17733) );
  NOR2_X1 U18731 ( .A1(n15582), .A2(n17733), .ZN(n17724) );
  NOR2_X1 U18732 ( .A1(n17724), .A2(n17723), .ZN(n17722) );
  XNOR2_X1 U18733 ( .A(n17248), .B(n15586), .ZN(n17713) );
  XNOR2_X1 U18734 ( .A(n17240), .B(n15589), .ZN(n17684) );
  NOR2_X1 U18735 ( .A1(n17683), .A2(n17684), .ZN(n15590) );
  NAND2_X1 U18736 ( .A1(n17683), .A2(n17684), .ZN(n17682) );
  INV_X1 U18737 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18001) );
  XOR2_X1 U18738 ( .A(n17235), .B(n15591), .Z(n15592) );
  XOR2_X1 U18739 ( .A(n18001), .B(n15592), .Z(n17672) );
  NOR2_X1 U18740 ( .A1(n15595), .A2(n15594), .ZN(n15596) );
  NOR2_X2 U18741 ( .A1(n17662), .A2(n15596), .ZN(n15599) );
  NOR2_X2 U18742 ( .A1(n15601), .A2(n9876), .ZN(n17627) );
  INV_X1 U18743 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17614) );
  NAND2_X1 U18744 ( .A1(n17547), .A2(n17933), .ZN(n17568) );
  INV_X1 U18745 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15598) );
  INV_X1 U18746 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15597) );
  INV_X1 U18747 ( .A(n15601), .ZN(n15602) );
  NAND2_X1 U18748 ( .A1(n17937), .A2(n15601), .ZN(n17981) );
  NAND2_X1 U18749 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17943) );
  INV_X1 U18750 ( .A(n17943), .ZN(n17610) );
  NAND2_X1 U18751 ( .A1(n17610), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17595) );
  NOR2_X1 U18752 ( .A1(n17595), .A2(n17933), .ZN(n17915) );
  NAND2_X1 U18753 ( .A1(n17915), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17903) );
  NOR2_X1 U18754 ( .A1(n15598), .A2(n17903), .ZN(n17875) );
  NAND2_X1 U18755 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17875), .ZN(
        n17858) );
  INV_X1 U18756 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17877) );
  NAND2_X1 U18757 ( .A1(n9876), .A2(n17877), .ZN(n15603) );
  NAND2_X1 U18758 ( .A1(n15604), .A2(n15603), .ZN(n15605) );
  NOR2_X2 U18759 ( .A1(n15606), .A2(n15605), .ZN(n17526) );
  INV_X1 U18760 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17855) );
  NAND2_X1 U18761 ( .A1(n17526), .A2(n17855), .ZN(n17525) );
  NAND2_X2 U18762 ( .A1(n17525), .A2(n17648), .ZN(n17443) );
  NAND2_X1 U18763 ( .A1(n15608), .A2(n15607), .ZN(n17541) );
  NAND2_X1 U18764 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17851) );
  INV_X1 U18765 ( .A(n17851), .ZN(n15613) );
  NAND2_X1 U18766 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17813) );
  INV_X1 U18767 ( .A(n17813), .ZN(n17823) );
  NAND3_X1 U18768 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17823), .ZN(n17457) );
  NOR2_X1 U18769 ( .A1(n17457), .A2(n17820), .ZN(n15614) );
  NAND2_X1 U18770 ( .A1(n15613), .A2(n15614), .ZN(n17798) );
  NOR2_X1 U18771 ( .A1(n17446), .A2(n17798), .ZN(n17436) );
  NAND2_X1 U18772 ( .A1(n17513), .A2(n17845), .ZN(n15609) );
  NOR2_X1 U18773 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15609), .ZN(
        n17476) );
  INV_X1 U18774 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17480) );
  NAND2_X1 U18775 ( .A1(n17476), .A2(n17480), .ZN(n17456) );
  NOR3_X1 U18776 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17456), .ZN(n15610) );
  INV_X1 U18777 ( .A(n15611), .ZN(n15612) );
  NAND2_X1 U18778 ( .A1(n15613), .A2(n17541), .ZN(n17474) );
  NAND2_X1 U18779 ( .A1(n17648), .A2(n9870), .ZN(n15615) );
  OAI221_X1 U18780 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17648), 
        .C1(n17776), .C2(n15616), .A(n15615), .ZN(n17402) );
  INV_X1 U18781 ( .A(n17427), .ZN(n15618) );
  INV_X1 U18782 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17751) );
  NOR2_X1 U18783 ( .A1(n17776), .A2(n17751), .ZN(n15667) );
  INV_X1 U18784 ( .A(n15667), .ZN(n17752) );
  NAND2_X1 U18785 ( .A1(n9876), .A2(n17752), .ZN(n15617) );
  INV_X1 U18786 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15670) );
  NOR2_X1 U18787 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17648), .ZN(
        n16285) );
  NAND2_X1 U18788 ( .A1(n15620), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16224) );
  OAI21_X1 U18789 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15620), .A(
        n16224), .ZN(n16253) );
  NOR2_X1 U18790 ( .A1(n18732), .A2(n18089), .ZN(n15628) );
  NAND2_X1 U18791 ( .A1(n15628), .A2(n18109), .ZN(n15630) );
  AOI21_X1 U18792 ( .B1(n18510), .B2(n15629), .A(n15622), .ZN(n15633) );
  INV_X1 U18793 ( .A(n15623), .ZN(n15624) );
  NOR2_X1 U18794 ( .A1(n15625), .A2(n15624), .ZN(n16221) );
  OAI21_X1 U18795 ( .B1(n15626), .B2(n18085), .A(n18730), .ZN(n15627) );
  OAI21_X1 U18796 ( .B1(n15628), .B2(n15627), .A(n18733), .ZN(n16404) );
  OAI22_X1 U18797 ( .A1(n16221), .A2(n15630), .B1(n15629), .B2(n16404), .ZN(
        n15631) );
  NAND2_X1 U18798 ( .A1(n15631), .A2(n18513), .ZN(n15632) );
  NOR3_X4 U18799 ( .A1(n18515), .A2(n17231), .A3(n18065), .ZN(n17967) );
  NOR2_X1 U18800 ( .A1(n18515), .A2(n16292), .ZN(n17938) );
  NAND2_X1 U18801 ( .A1(n18019), .A2(n17938), .ZN(n17980) );
  INV_X1 U18802 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17760) );
  NOR2_X1 U18803 ( .A1(n17760), .A2(n15670), .ZN(n16256) );
  NAND2_X1 U18804 ( .A1(n16256), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16272) );
  NAND2_X1 U18805 ( .A1(n17436), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17757) );
  NOR2_X1 U18806 ( .A1(n17776), .A2(n17757), .ZN(n17426) );
  NAND2_X1 U18807 ( .A1(n17426), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16283) );
  INV_X1 U18808 ( .A(n17875), .ZN(n17885) );
  INV_X1 U18809 ( .A(n17759), .ZN(n17383) );
  NOR2_X1 U18810 ( .A1(n16272), .A2(n17383), .ZN(n16257) );
  NAND2_X1 U18811 ( .A1(n18526), .A2(n15634), .ZN(n18539) );
  OR2_X1 U18812 ( .A1(n18732), .A2(n15635), .ZN(n15637) );
  OAI21_X1 U18813 ( .B1(n15637), .B2(n16421), .A(n15636), .ZN(n15638) );
  INV_X1 U18814 ( .A(n15638), .ZN(n18519) );
  NOR2_X1 U18815 ( .A1(n15640), .A2(n15639), .ZN(n18744) );
  INV_X1 U18816 ( .A(n17915), .ZN(n17923) );
  NOR2_X1 U18817 ( .A1(n15649), .A2(n17252), .ZN(n15647) );
  NOR2_X1 U18818 ( .A1(n15647), .A2(n17248), .ZN(n15646) );
  NAND2_X1 U18819 ( .A1(n15646), .A2(n17244), .ZN(n15644) );
  NOR2_X1 U18820 ( .A1(n17240), .A2(n15644), .ZN(n15643) );
  NAND2_X1 U18821 ( .A1(n15643), .A2(n17235), .ZN(n15642) );
  NOR2_X1 U18822 ( .A1(n17231), .A2(n15642), .ZN(n15663) );
  XOR2_X1 U18823 ( .A(n15642), .B(n17231), .Z(n17655) );
  XOR2_X1 U18824 ( .A(n15643), .B(n17235), .Z(n15657) );
  XOR2_X1 U18825 ( .A(n15644), .B(n17240), .Z(n15645) );
  NAND2_X1 U18826 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15645), .ZN(
        n15656) );
  XOR2_X1 U18827 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n15645), .Z(
        n17688) );
  XOR2_X1 U18828 ( .A(n15646), .B(n17244), .Z(n17700) );
  XOR2_X1 U18829 ( .A(n17248), .B(n15647), .Z(n15648) );
  NAND2_X1 U18830 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15648), .ZN(
        n15654) );
  XOR2_X1 U18831 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n15648), .Z(
        n17710) );
  OR2_X1 U18832 ( .A1(n15583), .A2(n15650), .ZN(n15653) );
  AOI21_X1 U18833 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n15569), .A(
        n17744), .ZN(n15652) );
  INV_X1 U18834 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18705) );
  AOI221_X1 U18835 ( .B1(n17744), .B2(n15569), .C1(n15652), .C2(n18705), .A(
        n15651), .ZN(n17726) );
  NAND2_X1 U18836 ( .A1(n15653), .A2(n17725), .ZN(n17709) );
  NAND2_X1 U18837 ( .A1(n17710), .A2(n17709), .ZN(n17708) );
  NAND2_X1 U18838 ( .A1(n15654), .A2(n17708), .ZN(n17701) );
  NAND2_X1 U18839 ( .A1(n17700), .A2(n17701), .ZN(n17699) );
  NOR2_X1 U18840 ( .A1(n17700), .A2(n17701), .ZN(n15655) );
  AOI21_X1 U18841 ( .B1(n20898), .B2(n17699), .A(n15655), .ZN(n17687) );
  NAND2_X1 U18842 ( .A1(n17688), .A2(n17687), .ZN(n17686) );
  NAND2_X1 U18843 ( .A1(n15656), .A2(n17686), .ZN(n15658) );
  NAND2_X1 U18844 ( .A1(n15657), .A2(n15658), .ZN(n15659) );
  XOR2_X1 U18845 ( .A(n15658), .B(n15657), .Z(n17669) );
  NAND2_X1 U18846 ( .A1(n17669), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17668) );
  NAND2_X1 U18847 ( .A1(n15663), .A2(n15660), .ZN(n15664) );
  NAND2_X1 U18848 ( .A1(n17655), .A2(n17656), .ZN(n17654) );
  NAND2_X1 U18849 ( .A1(n15663), .A2(n15662), .ZN(n15661) );
  OAI211_X1 U18850 ( .C1(n15663), .C2(n15662), .A(n17654), .B(n15661), .ZN(
        n17641) );
  NAND2_X1 U18851 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17641), .ZN(
        n17640) );
  OAI22_X1 U18852 ( .A1(n17980), .A2(n16257), .B1(n18068), .B2(n16255), .ZN(
        n15665) );
  INV_X1 U18853 ( .A(n15665), .ZN(n15728) );
  NOR2_X1 U18854 ( .A1(n18020), .A2(n18065), .ZN(n16269) );
  NOR2_X1 U18855 ( .A1(n18548), .A2(n18539), .ZN(n17954) );
  INV_X1 U18856 ( .A(n16283), .ZN(n15673) );
  NAND4_X1 U18857 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17974) );
  NOR2_X1 U18858 ( .A1(n17976), .A2(n17974), .ZN(n17856) );
  NAND2_X1 U18859 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17856), .ZN(
        n15666) );
  NAND2_X1 U18860 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17971) );
  NOR2_X1 U18861 ( .A1(n15666), .A2(n17971), .ZN(n17870) );
  NAND2_X1 U18862 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17870), .ZN(
        n17961) );
  NOR2_X1 U18863 ( .A1(n17858), .A2(n17961), .ZN(n17871) );
  NAND3_X1 U18864 ( .A1(n15673), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17871), .ZN(n15669) );
  NAND2_X1 U18865 ( .A1(n16282), .A2(n17870), .ZN(n17807) );
  INV_X1 U18866 ( .A(n17807), .ZN(n17756) );
  AOI21_X1 U18867 ( .B1(n15673), .B2(n17756), .A(n18552), .ZN(n15668) );
  AOI21_X1 U18868 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17973) );
  NOR2_X1 U18869 ( .A1(n17973), .A2(n15666), .ZN(n17873) );
  NAND2_X1 U18870 ( .A1(n16282), .A2(n17873), .ZN(n17850) );
  OAI21_X1 U18871 ( .B1(n17757), .B2(n17850), .A(n18548), .ZN(n17772) );
  OAI21_X1 U18872 ( .B1(n15667), .B2(n18039), .A(n17772), .ZN(n17753) );
  AOI211_X1 U18873 ( .C1(n18524), .C2(n15669), .A(n15668), .B(n17753), .ZN(
        n15726) );
  OAI21_X1 U18874 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17954), .A(
        n15726), .ZN(n16288) );
  AOI22_X1 U18875 ( .A1(n16269), .A2(n15670), .B1(n18019), .B2(n16288), .ZN(
        n15671) );
  NAND3_X1 U18876 ( .A1(n15728), .A2(n15671), .A3(n18035), .ZN(n15672) );
  AOI22_X1 U18877 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15672), .B1(
        n18032), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n15676) );
  INV_X1 U18878 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16258) );
  AOI21_X1 U18879 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18524), .A(
        n18539), .ZN(n18036) );
  OAI22_X1 U18880 ( .A1(n18039), .A2(n17850), .B1(n17807), .B2(n18036), .ZN(
        n17774) );
  NAND3_X1 U18881 ( .A1(n15673), .A2(n18019), .A3(n17774), .ZN(n16271) );
  INV_X1 U18882 ( .A(n17980), .ZN(n17908) );
  NAND2_X1 U18883 ( .A1(n17759), .A2(n17908), .ZN(n15674) );
  OAI211_X1 U18884 ( .C1(n18068), .C2(n17755), .A(n16271), .B(n15674), .ZN(
        n15730) );
  NAND3_X1 U18885 ( .A1(n16256), .A2(n16258), .A3(n15730), .ZN(n15675) );
  OAI211_X1 U18886 ( .C1(n16253), .C2(n17982), .A(n15676), .B(n15675), .ZN(
        P3_U2833) );
  AOI22_X1 U18887 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n18917), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18829), .ZN(n15685) );
  AOI22_X1 U18888 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18906), .B1(
        n15677), .B2(n18901), .ZN(n15684) );
  OAI22_X1 U18889 ( .A1(n16072), .A2(n18878), .B1(n18916), .B2(n16052), .ZN(
        n15678) );
  INV_X1 U18890 ( .A(n15678), .ZN(n15683) );
  AOI21_X1 U18891 ( .B1(n15680), .B2(n15679), .A(n9670), .ZN(n15681) );
  NAND2_X1 U18892 ( .A1(n18912), .A2(n15681), .ZN(n15682) );
  NAND4_X1 U18893 ( .A1(n15685), .A2(n15684), .A3(n15683), .A4(n15682), .ZN(
        P2_U2833) );
  NOR3_X1 U18894 ( .A1(n15687), .A2(n15686), .A3(n20464), .ZN(n15692) );
  INV_X1 U18895 ( .A(n15692), .ZN(n15690) );
  OAI211_X1 U18896 ( .C1(n15690), .C2(n20351), .A(n15689), .B(n15688), .ZN(
        n15691) );
  OAI21_X1 U18897 ( .B1(n15692), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15691), .ZN(n15693) );
  AOI222_X1 U18898 ( .A1(n15694), .A2(n20428), .B1(n15694), .B2(n15693), .C1(
        n20428), .C2(n15693), .ZN(n15698) );
  INV_X1 U18899 ( .A(n15698), .ZN(n15696) );
  OAI21_X1 U18900 ( .B1(n15696), .B2(n20737), .A(n15695), .ZN(n15697) );
  OAI21_X1 U18901 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15698), .A(
        n15697), .ZN(n15708) );
  INV_X1 U18902 ( .A(n15699), .ZN(n15707) );
  INV_X1 U18903 ( .A(n15700), .ZN(n15704) );
  OAI21_X1 U18904 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15701), .ZN(n15702) );
  NAND4_X1 U18905 ( .A1(n15705), .A2(n15704), .A3(n15703), .A4(n15702), .ZN(
        n15706) );
  AOI211_X1 U18906 ( .C1(n15708), .C2(n19995), .A(n15707), .B(n15706), .ZN(
        n15722) );
  OR2_X1 U18907 ( .A1(n20758), .A2(n15709), .ZN(n15710) );
  NOR2_X1 U18908 ( .A1(n15711), .A2(n15710), .ZN(n15712) );
  AOI221_X1 U18909 ( .B1(n15713), .B2(n20649), .C1(n20661), .C2(n20649), .A(
        n15712), .ZN(n15992) );
  OAI221_X1 U18910 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15722), 
        .A(n15992), .ZN(n15999) );
  NOR2_X1 U18911 ( .A1(n15994), .A2(n15714), .ZN(n15715) );
  NOR2_X1 U18912 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15715), .ZN(n15720) );
  AOI211_X1 U18913 ( .C1(n20751), .C2(n20750), .A(n15717), .B(n15716), .ZN(
        n15718) );
  NAND2_X1 U18914 ( .A1(n15999), .A2(n15718), .ZN(n15719) );
  AOI22_X1 U18915 ( .A1(n15999), .A2(n15720), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15719), .ZN(n15721) );
  OAI21_X1 U18916 ( .B1(n15722), .B2(n19750), .A(n15721), .ZN(P1_U3161) );
  NAND2_X1 U18917 ( .A1(n16224), .A2(n9876), .ZN(n16226) );
  OAI21_X1 U18918 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15723), .A(
        n17648), .ZN(n16227) );
  NAND2_X1 U18919 ( .A1(n16226), .A2(n16227), .ZN(n15725) );
  NOR2_X1 U18920 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16272), .ZN(
        n16248) );
  OAI21_X1 U18921 ( .B1(n18065), .B2(n15726), .A(n18035), .ZN(n15727) );
  AOI21_X1 U18922 ( .B1(n16269), .B2(n16272), .A(n15727), .ZN(n16270) );
  AOI21_X1 U18923 ( .B1(n16270), .B2(n15728), .A(n15724), .ZN(n15729) );
  AOI21_X1 U18924 ( .B1(n16248), .B2(n15730), .A(n15729), .ZN(n15731) );
  NAND2_X1 U18925 ( .A1(n18032), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16244) );
  OAI211_X1 U18926 ( .C1(n17982), .C2(n16252), .A(n15731), .B(n16244), .ZN(
        P3_U2832) );
  INV_X1 U18927 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19747) );
  INV_X1 U18928 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20769) );
  NOR2_X1 U18929 ( .A1(n20659), .A2(n20769), .ZN(n20657) );
  INV_X1 U18930 ( .A(HOLD), .ZN(n20660) );
  NOR2_X1 U18931 ( .A1(n19747), .A2(n20660), .ZN(n20652) );
  OAI22_X1 U18932 ( .A1(n20657), .A2(n20652), .B1(n11003), .B2(n20660), .ZN(
        n15732) );
  OAI211_X1 U18933 ( .C1(n19747), .C2(n20661), .A(n20758), .B(n15732), .ZN(
        P1_U3195) );
  AND2_X1 U18934 ( .A1(n15733), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U18935 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15735) );
  NOR3_X1 U18936 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13371), .A3(n19600), 
        .ZN(n16210) );
  INV_X1 U18937 ( .A(n15734), .ZN(n15737) );
  NOR4_X1 U18938 ( .A1(n15736), .A2(n15735), .A3(n16210), .A4(n15737), .ZN(
        P2_U3178) );
  AOI221_X1 U18939 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15737), .C1(n19718), .C2(
        n15737), .A(n19516), .ZN(n19715) );
  INV_X1 U18940 ( .A(n19715), .ZN(n19712) );
  NOR2_X1 U18941 ( .A1(n15738), .A2(n19712), .ZN(P2_U3047) );
  NAND3_X1 U18942 ( .A1(n16752), .A2(n18732), .A3(n15739), .ZN(n15740) );
  INV_X1 U18943 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17338) );
  INV_X2 U18944 ( .A(n17212), .ZN(n17239) );
  AOI22_X1 U18945 ( .A1(n17258), .A2(BUF2_REG_0__SCAN_IN), .B1(n17257), .B2(
        n17744), .ZN(n15744) );
  NOR3_X1 U18946 ( .A1(n17259), .A2(n18114), .A3(P3_EAX_REG_0__SCAN_IN), .ZN(
        n17261) );
  INV_X1 U18947 ( .A(n17261), .ZN(n15743) );
  OAI211_X1 U18948 ( .C1(n17110), .C2(n17338), .A(n15744), .B(n15743), .ZN(
        P3_U2735) );
  AOI22_X1 U18949 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19853), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(n19849), .ZN(n15750) );
  AOI22_X1 U18950 ( .A1(n15746), .A2(n19850), .B1(n15745), .B2(n20694), .ZN(
        n15749) );
  AOI22_X1 U18951 ( .A1(n15856), .A2(n19797), .B1(n19834), .B2(n15849), .ZN(
        n15748) );
  NOR2_X1 U18952 ( .A1(n19826), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15759) );
  OAI21_X1 U18953 ( .B1(n15759), .B2(n15751), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15747) );
  NAND4_X1 U18954 ( .A1(n15750), .A2(n15749), .A3(n15748), .A4(n15747), .ZN(
        P1_U2818) );
  AOI22_X1 U18955 ( .A1(n15752), .A2(n19850), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n15751), .ZN(n15762) );
  OAI22_X1 U18956 ( .A1(n20839), .A2(n19819), .B1(n15753), .B2(n19847), .ZN(
        n15758) );
  INV_X1 U18957 ( .A(n15754), .ZN(n15755) );
  OAI22_X1 U18958 ( .A1(n15756), .A2(n15842), .B1(n15755), .B2(n19865), .ZN(
        n15757) );
  AOI211_X1 U18959 ( .C1(n15760), .C2(n15759), .A(n15758), .B(n15757), .ZN(
        n15761) );
  NAND2_X1 U18960 ( .A1(n15762), .A2(n15761), .ZN(P1_U2819) );
  AOI22_X1 U18961 ( .A1(n15763), .A2(n19850), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n19849), .ZN(n15767) );
  NOR3_X1 U18962 ( .A1(n19826), .A2(P1_REIP_REG_19__SCAN_IN), .A3(n15764), 
        .ZN(n15765) );
  AOI211_X1 U18963 ( .C1(n19853), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19776), .B(n15765), .ZN(n15766) );
  NAND2_X1 U18964 ( .A1(n15767), .A2(n15766), .ZN(n15768) );
  AOI21_X1 U18965 ( .B1(n15769), .B2(n19797), .A(n15768), .ZN(n15774) );
  OAI21_X1 U18966 ( .B1(n19826), .B2(n15770), .A(n19827), .ZN(n15789) );
  NOR2_X1 U18967 ( .A1(n19826), .A2(n15771), .ZN(n15790) );
  INV_X1 U18968 ( .A(n15790), .ZN(n15772) );
  NOR3_X1 U18969 ( .A1(n15772), .A2(P1_REIP_REG_18__SCAN_IN), .A3(n20687), 
        .ZN(n15778) );
  OAI21_X1 U18970 ( .B1(n15789), .B2(n15778), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15773) );
  OAI211_X1 U18971 ( .C1(n15775), .C2(n19865), .A(n15774), .B(n15773), .ZN(
        P1_U2821) );
  AOI22_X1 U18972 ( .A1(n15776), .A2(n19850), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n15789), .ZN(n15782) );
  OAI21_X1 U18973 ( .B1(n19847), .B2(n15854), .A(n19817), .ZN(n15777) );
  AOI211_X1 U18974 ( .C1(n19853), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15778), .B(n15777), .ZN(n15781) );
  INV_X1 U18975 ( .A(n15779), .ZN(n15852) );
  AOI22_X1 U18976 ( .A1(n15860), .A2(n19797), .B1(n19834), .B2(n15852), .ZN(
        n15780) );
  NAND3_X1 U18977 ( .A1(n15782), .A2(n15781), .A3(n15780), .ZN(P1_U2822) );
  INV_X1 U18978 ( .A(n15783), .ZN(n15788) );
  AOI22_X1 U18979 ( .A1(n15784), .A2(n19850), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n19849), .ZN(n15785) );
  OAI211_X1 U18980 ( .C1(n19819), .C2(n15786), .A(n15785), .B(n19817), .ZN(
        n15787) );
  AOI21_X1 U18981 ( .B1(n15788), .B2(n19797), .A(n15787), .ZN(n15792) );
  OAI21_X1 U18982 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15790), .A(n15789), 
        .ZN(n15791) );
  OAI211_X1 U18983 ( .C1(n15793), .C2(n19865), .A(n15792), .B(n15791), .ZN(
        P1_U2823) );
  AOI22_X1 U18984 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19853), .B1(
        P1_EBX_REG_16__SCAN_IN), .B2(n19849), .ZN(n15801) );
  NOR2_X1 U18985 ( .A1(n15923), .A2(n19865), .ZN(n15797) );
  OAI21_X1 U18986 ( .B1(n19836), .B2(n15804), .A(n19801), .ZN(n15818) );
  INV_X1 U18987 ( .A(n15818), .ZN(n15794) );
  AOI21_X1 U18988 ( .B1(n19837), .B2(n20684), .A(n15794), .ZN(n15795) );
  OAI22_X1 U18989 ( .A1(n15795), .A2(n15921), .B1(n15883), .B2(n19833), .ZN(
        n15796) );
  AOI211_X1 U18990 ( .C1(n15880), .C2(n19797), .A(n15797), .B(n15796), .ZN(
        n15800) );
  NAND3_X1 U18991 ( .A1(n19837), .A2(n15921), .A3(n15798), .ZN(n15799) );
  NAND4_X1 U18992 ( .A1(n15801), .A2(n15800), .A3(n19817), .A4(n15799), .ZN(
        P1_U2824) );
  INV_X1 U18993 ( .A(n15932), .ZN(n15808) );
  OAI22_X1 U18994 ( .A1(n20939), .A2(n19819), .B1(n15802), .B2(n19847), .ZN(
        n15803) );
  AOI211_X1 U18995 ( .C1(n19850), .C2(n15888), .A(n19776), .B(n15803), .ZN(
        n15807) );
  INV_X1 U18996 ( .A(n15804), .ZN(n15805) );
  NAND3_X1 U18997 ( .A1(n19837), .A2(n15805), .A3(n20684), .ZN(n15806) );
  OAI211_X1 U18998 ( .C1(n15808), .C2(n19865), .A(n15807), .B(n15806), .ZN(
        n15809) );
  AOI21_X1 U18999 ( .B1(n15889), .B2(n19797), .A(n15809), .ZN(n15810) );
  OAI21_X1 U19000 ( .B1(n15818), .B2(n20684), .A(n15810), .ZN(P1_U2825) );
  AOI21_X1 U19001 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15811), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15817) );
  OAI22_X1 U19002 ( .A1(n15813), .A2(n19819), .B1(n19865), .B2(n15812), .ZN(
        n15814) );
  AOI211_X1 U19003 ( .C1(n19849), .C2(P1_EBX_REG_14__SCAN_IN), .A(n19776), .B(
        n15814), .ZN(n15816) );
  AOI22_X1 U19004 ( .A1(n15893), .A2(n19797), .B1(n19850), .B2(n15892), .ZN(
        n15815) );
  OAI211_X1 U19005 ( .C1(n15818), .C2(n15817), .A(n15816), .B(n15815), .ZN(
        P1_U2826) );
  OAI22_X1 U19006 ( .A1(n15820), .A2(n19819), .B1(n15819), .B2(n19847), .ZN(
        n15821) );
  AOI211_X1 U19007 ( .C1(n15822), .C2(n19834), .A(n19776), .B(n15821), .ZN(
        n15827) );
  INV_X1 U19008 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15835) );
  INV_X1 U19009 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15823) );
  OAI21_X1 U19010 ( .B1(n15835), .B2(n15836), .A(n15823), .ZN(n15824) );
  AOI22_X1 U19011 ( .A1(n15899), .A2(n19850), .B1(n15825), .B2(n15824), .ZN(
        n15826) );
  OAI211_X1 U19012 ( .C1(n15842), .C2(n15897), .A(n15827), .B(n15826), .ZN(
        P1_U2828) );
  NAND2_X1 U19013 ( .A1(n19837), .A2(n15828), .ZN(n15848) );
  AND2_X1 U19014 ( .A1(n15848), .A2(n19827), .ZN(n15841) );
  INV_X1 U19015 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15832) );
  OAI22_X1 U19016 ( .A1(n15908), .A2(n19833), .B1(n19865), .B2(n15829), .ZN(
        n15830) );
  AOI21_X1 U19017 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(n19849), .A(n15830), .ZN(
        n15831) );
  OAI211_X1 U19018 ( .C1(n19819), .C2(n15832), .A(n15831), .B(n19817), .ZN(
        n15833) );
  AOI21_X1 U19019 ( .B1(n19797), .B2(n15904), .A(n15833), .ZN(n15834) );
  OAI221_X1 U19020 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15836), .C1(n15835), 
        .C2(n15841), .A(n15834), .ZN(P1_U2829) );
  INV_X1 U19021 ( .A(n15837), .ZN(n15838) );
  NAND2_X1 U19022 ( .A1(n15838), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n19780) );
  INV_X1 U19023 ( .A(n15839), .ZN(n15955) );
  AOI22_X1 U19024 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(n19849), .B1(n19834), 
        .B2(n15955), .ZN(n15840) );
  OAI211_X1 U19025 ( .C1(n19819), .C2(n11450), .A(n15840), .B(n19817), .ZN(
        n15845) );
  OAI22_X1 U19026 ( .A1(n15843), .A2(n15842), .B1(n14229), .B2(n15841), .ZN(
        n15844) );
  AOI211_X1 U19027 ( .C1(n15846), .C2(n19850), .A(n15845), .B(n15844), .ZN(
        n15847) );
  OAI21_X1 U19028 ( .B1(n15848), .B2(n19780), .A(n15847), .ZN(P1_U2830) );
  AOI22_X1 U19029 ( .A1(n15856), .A2(n19870), .B1(n15849), .B2(n19869), .ZN(
        n15850) );
  OAI21_X1 U19030 ( .B1(n19873), .B2(n15851), .A(n15850), .ZN(P1_U2850) );
  AOI22_X1 U19031 ( .A1(n15860), .A2(n19870), .B1(n19869), .B2(n15852), .ZN(
        n15853) );
  OAI21_X1 U19032 ( .B1(n19873), .B2(n15854), .A(n15853), .ZN(P1_U2854) );
  INV_X1 U19033 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16321) );
  AOI22_X1 U19034 ( .A1(n15865), .A2(n15855), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n15863), .ZN(n15858) );
  AOI22_X1 U19035 ( .A1(n15856), .A2(n15867), .B1(n15866), .B2(DATAI_22_), 
        .ZN(n15857) );
  OAI211_X1 U19036 ( .C1(n15870), .C2(n16321), .A(n15858), .B(n15857), .ZN(
        P1_U2882) );
  INV_X1 U19037 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16329) );
  AOI22_X1 U19038 ( .A1(n15865), .A2(n15859), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15863), .ZN(n15862) );
  AOI22_X1 U19039 ( .A1(n15860), .A2(n15867), .B1(n15866), .B2(DATAI_18_), 
        .ZN(n15861) );
  OAI211_X1 U19040 ( .C1(n15870), .C2(n16329), .A(n15862), .B(n15861), .ZN(
        P1_U2886) );
  AOI22_X1 U19041 ( .A1(n15865), .A2(n15864), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15863), .ZN(n15869) );
  AOI22_X1 U19042 ( .A1(n15880), .A2(n15867), .B1(n15866), .B2(DATAI_16_), 
        .ZN(n15868) );
  OAI211_X1 U19043 ( .C1(n15870), .C2(n16333), .A(n15869), .B(n15868), .ZN(
        P1_U2888) );
  AOI22_X1 U19044 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n19944), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15882) );
  OR2_X1 U19045 ( .A1(n14223), .A2(n15871), .ZN(n15875) );
  AND2_X1 U19046 ( .A1(n15873), .A2(n15872), .ZN(n15874) );
  NAND2_X1 U19047 ( .A1(n15875), .A2(n15874), .ZN(n15885) );
  NAND2_X1 U19048 ( .A1(n15876), .A2(n15877), .ZN(n15884) );
  NAND2_X1 U19049 ( .A1(n15887), .A2(n15877), .ZN(n15879) );
  XNOR2_X1 U19050 ( .A(n15879), .B(n15878), .ZN(n15927) );
  AOI22_X1 U19051 ( .A1(n15927), .A2(n19939), .B1(n19938), .B2(n15880), .ZN(
        n15881) );
  OAI211_X1 U19052 ( .C1(n19943), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        P1_U2983) );
  NAND2_X1 U19053 ( .A1(n15885), .A2(n15884), .ZN(n15886) );
  AOI22_X1 U19054 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19944), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15891) );
  AOI22_X1 U19055 ( .A1(n15889), .A2(n19938), .B1(n15888), .B2(n15909), .ZN(
        n15890) );
  OAI211_X1 U19056 ( .C1(n15931), .C2(n15902), .A(n15891), .B(n15890), .ZN(
        P1_U2984) );
  AOI22_X1 U19057 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19944), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15895) );
  AOI22_X1 U19058 ( .A1(n15893), .A2(n19938), .B1(n15909), .B2(n15892), .ZN(
        n15894) );
  OAI211_X1 U19059 ( .C1(n15896), .C2(n15902), .A(n15895), .B(n15894), .ZN(
        P1_U2985) );
  AOI22_X1 U19060 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19944), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15901) );
  INV_X1 U19061 ( .A(n15897), .ZN(n15898) );
  AOI22_X1 U19062 ( .A1(n15909), .A2(n15899), .B1(n19938), .B2(n15898), .ZN(
        n15900) );
  OAI211_X1 U19063 ( .C1(n15903), .C2(n15902), .A(n15901), .B(n15900), .ZN(
        P1_U2987) );
  AOI22_X1 U19064 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19944), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15907) );
  AOI22_X1 U19065 ( .A1(n19939), .A2(n15905), .B1(n19938), .B2(n15904), .ZN(
        n15906) );
  OAI211_X1 U19066 ( .C1(n19943), .C2(n15908), .A(n15907), .B(n15906), .ZN(
        P1_U2988) );
  INV_X1 U19067 ( .A(n19793), .ZN(n15910) );
  AOI222_X1 U19068 ( .A1(n15911), .A2(n19939), .B1(n15910), .B2(n15909), .C1(
        n19938), .C2(n19790), .ZN(n15913) );
  OAI211_X1 U19069 ( .C1(n20945), .C2(n15914), .A(n15913), .B(n15912), .ZN(
        P1_U2992) );
  AOI22_X1 U19070 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19944), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15920) );
  OAI21_X1 U19071 ( .B1(n15917), .B2(n15916), .A(n15915), .ZN(n15918) );
  INV_X1 U19072 ( .A(n15918), .ZN(n15979) );
  AOI22_X1 U19073 ( .A1(n15979), .A2(n19939), .B1(n19938), .B2(n19867), .ZN(
        n15919) );
  OAI211_X1 U19074 ( .C1(n19943), .C2(n19813), .A(n15920), .B(n15919), .ZN(
        P1_U2994) );
  INV_X1 U19075 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15930) );
  INV_X1 U19076 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15921) );
  OAI22_X1 U19077 ( .A1(n15923), .A2(n19981), .B1(n15922), .B2(n15921), .ZN(
        n15924) );
  INV_X1 U19078 ( .A(n15924), .ZN(n15929) );
  AOI21_X1 U19079 ( .B1(n15936), .B2(n15930), .A(n15937), .ZN(n15926) );
  AOI22_X1 U19080 ( .A1(n15927), .A2(n19988), .B1(n15926), .B2(n15925), .ZN(
        n15928) );
  OAI211_X1 U19081 ( .C1(n15935), .C2(n15930), .A(n15929), .B(n15928), .ZN(
        P1_U3015) );
  INV_X1 U19082 ( .A(n15931), .ZN(n15933) );
  AOI222_X1 U19083 ( .A1(n15933), .A2(n19988), .B1(n19974), .B2(n15932), .C1(
        P1_REIP_REG_15__SCAN_IN), .C2(n19944), .ZN(n15934) );
  OAI221_X1 U19084 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15937), 
        .C1(n15936), .C2(n15935), .A(n15934), .ZN(P1_U3016) );
  NOR2_X1 U19085 ( .A1(n15939), .A2(n15938), .ZN(n15940) );
  AOI211_X1 U19086 ( .C1(n19962), .C2(n15941), .A(n19991), .B(n15940), .ZN(
        n15952) );
  INV_X1 U19087 ( .A(n15942), .ZN(n15950) );
  AOI211_X1 U19088 ( .C1(n13747), .C2(n15945), .A(n15944), .B(n15943), .ZN(
        n15946) );
  AOI21_X1 U19089 ( .B1(n19944), .B2(P1_REIP_REG_13__SCAN_IN), .A(n15946), 
        .ZN(n15947) );
  OAI21_X1 U19090 ( .B1(n15948), .B2(n19981), .A(n15947), .ZN(n15949) );
  AOI21_X1 U19091 ( .B1(n15950), .B2(n19988), .A(n15949), .ZN(n15951) );
  OAI221_X1 U19092 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15953), 
        .C1(n13747), .C2(n15952), .A(n15951), .ZN(P1_U3018) );
  AOI21_X1 U19093 ( .B1(n15955), .B2(n19974), .A(n15954), .ZN(n15962) );
  AOI21_X1 U19094 ( .B1(n14226), .B2(n15957), .A(n15956), .ZN(n15959) );
  AOI22_X1 U19095 ( .A1(n15960), .A2(n19988), .B1(n15959), .B2(n15958), .ZN(
        n15961) );
  OAI211_X1 U19096 ( .C1(n15963), .C2(n14226), .A(n15962), .B(n15961), .ZN(
        P1_U3021) );
  INV_X1 U19097 ( .A(n15964), .ZN(n15965) );
  AOI21_X1 U19098 ( .B1(n15966), .B2(n19974), .A(n15965), .ZN(n15975) );
  NOR3_X1 U19099 ( .A1(n15968), .A2(n15967), .A3(n10002), .ZN(n15969) );
  AOI21_X1 U19100 ( .B1(n15970), .B2(n19988), .A(n15969), .ZN(n15974) );
  NAND2_X1 U19101 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15971) );
  OAI211_X1 U19102 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15972), .B(n15971), .ZN(n15973) );
  NAND3_X1 U19103 ( .A1(n15975), .A2(n15974), .A3(n15973), .ZN(P1_U3023) );
  INV_X1 U19104 ( .A(n15976), .ZN(n15977) );
  XNOR2_X1 U19105 ( .A(n19814), .B(n15977), .ZN(n19866) );
  AOI22_X1 U19106 ( .A1(n19866), .A2(n19974), .B1(n19944), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n15981) );
  AOI22_X1 U19107 ( .A1(n15979), .A2(n19988), .B1(n15978), .B2(n19953), .ZN(
        n15980) );
  OAI211_X1 U19108 ( .C1(n15983), .C2(n15982), .A(n15981), .B(n15980), .ZN(
        P1_U3026) );
  INV_X1 U19109 ( .A(n19821), .ZN(n15986) );
  INV_X1 U19110 ( .A(n15984), .ZN(n15985) );
  NAND3_X1 U19111 ( .A1(n15986), .A2(n15985), .A3(n20720), .ZN(n15989) );
  OAI22_X1 U19112 ( .A1(n15990), .A2(n15989), .B1(n15988), .B2(n15987), .ZN(
        P1_U3468) );
  AOI21_X1 U19113 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n15999), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15997) );
  NOR2_X1 U19114 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20751), .ZN(n15991) );
  OAI221_X1 U19115 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20759), .C2(n15991), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20650) );
  AOI21_X1 U19116 ( .B1(n20650), .B2(n15993), .A(n15992), .ZN(n15996) );
  AOI21_X1 U19117 ( .B1(n20301), .B2(n20661), .A(n15994), .ZN(n15995) );
  NOR3_X1 U19118 ( .A1(n15997), .A2(n15996), .A3(n15995), .ZN(P1_U3162) );
  OAI221_X1 U19119 ( .B1(n20301), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20301), 
        .C2(n15999), .A(n15998), .ZN(P1_U3466) );
  XNOR2_X1 U19120 ( .A(n16001), .B(n16000), .ZN(n16010) );
  AOI22_X1 U19121 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18917), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18829), .ZN(n16002) );
  OAI21_X1 U19122 ( .B1(n16003), .B2(n18925), .A(n16002), .ZN(n16004) );
  AOI21_X1 U19123 ( .B1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18906), .A(
        n16004), .ZN(n16009) );
  OAI22_X1 U19124 ( .A1(n16006), .A2(n18878), .B1(n16005), .B2(n18916), .ZN(
        n16007) );
  INV_X1 U19125 ( .A(n16007), .ZN(n16008) );
  OAI211_X1 U19126 ( .C1(n18883), .C2(n16010), .A(n16009), .B(n16008), .ZN(
        P2_U2825) );
  INV_X1 U19127 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19663) );
  INV_X1 U19128 ( .A(n16011), .ZN(n16013) );
  OAI211_X1 U19129 ( .C1(n16014), .C2(n16013), .A(n16012), .B(n18901), .ZN(
        n16016) );
  AOI22_X1 U19130 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n18917), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18906), .ZN(n16015) );
  OAI211_X1 U19131 ( .C1(n18918), .C2(n19663), .A(n16016), .B(n16015), .ZN(
        n16017) );
  AOI21_X1 U19132 ( .B1(n16018), .B2(n18927), .A(n16017), .ZN(n16019) );
  INV_X1 U19133 ( .A(n16019), .ZN(n16024) );
  AOI211_X1 U19134 ( .C1(n16022), .C2(n16021), .A(n16020), .B(n18883), .ZN(
        n16023) );
  NOR2_X1 U19135 ( .A1(n16024), .A2(n16023), .ZN(n16025) );
  OAI21_X1 U19136 ( .B1(n16026), .B2(n18916), .A(n16025), .ZN(P2_U2828) );
  AOI22_X1 U19137 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n18829), .B1(n16027), 
        .B2(n18901), .ZN(n16038) );
  AOI22_X1 U19138 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18917), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18906), .ZN(n16037) );
  INV_X1 U19139 ( .A(n16028), .ZN(n16030) );
  AOI22_X1 U19140 ( .A1(n16030), .A2(n18927), .B1(n16029), .B2(n18922), .ZN(
        n16036) );
  AOI21_X1 U19141 ( .B1(n16033), .B2(n16032), .A(n16031), .ZN(n16034) );
  NAND2_X1 U19142 ( .A1(n18912), .A2(n16034), .ZN(n16035) );
  NAND4_X1 U19143 ( .A1(n16038), .A2(n16037), .A3(n16036), .A4(n16035), .ZN(
        P2_U2829) );
  AOI211_X1 U19144 ( .C1(n16041), .C2(n16040), .A(n16039), .B(n18883), .ZN(
        n16045) );
  AOI22_X1 U19145 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18917), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18829), .ZN(n16042) );
  OAI21_X1 U19146 ( .B1(n16043), .B2(n18925), .A(n16042), .ZN(n16044) );
  AOI211_X1 U19147 ( .C1(n18906), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16045), .B(n16044), .ZN(n16050) );
  INV_X1 U19148 ( .A(n16046), .ZN(n16048) );
  AOI22_X1 U19149 ( .A1(n16048), .A2(n18927), .B1(n18922), .B2(n16047), .ZN(
        n16049) );
  NAND2_X1 U19150 ( .A1(n16050), .A2(n16049), .ZN(P2_U2831) );
  AOI22_X1 U19151 ( .A1(n16065), .A2(n16051), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n18983), .ZN(n16057) );
  AOI22_X1 U19152 ( .A1(n18938), .A2(BUF1_REG_22__SCAN_IN), .B1(n18940), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16056) );
  INV_X1 U19153 ( .A(n16052), .ZN(n16053) );
  AOI22_X1 U19154 ( .A1(n16054), .A2(n18986), .B1(n18984), .B2(n16053), .ZN(
        n16055) );
  NAND3_X1 U19155 ( .A1(n16057), .A2(n16056), .A3(n16055), .ZN(P2_U2897) );
  AOI22_X1 U19156 ( .A1(n16065), .A2(n16058), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n18983), .ZN(n16063) );
  AOI22_X1 U19157 ( .A1(n18938), .A2(BUF1_REG_20__SCAN_IN), .B1(n18940), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16062) );
  OAI22_X1 U19158 ( .A1(n16059), .A2(n18978), .B1(n18967), .B2(n18791), .ZN(
        n16060) );
  INV_X1 U19159 ( .A(n16060), .ZN(n16061) );
  NAND3_X1 U19160 ( .A1(n16063), .A2(n16062), .A3(n16061), .ZN(P2_U2899) );
  AOI22_X1 U19161 ( .A1(n16065), .A2(n16064), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n18983), .ZN(n16070) );
  AOI22_X1 U19162 ( .A1(n18938), .A2(BUF1_REG_18__SCAN_IN), .B1(n18940), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16069) );
  AOI22_X1 U19163 ( .A1(n16067), .A2(n18986), .B1(n18984), .B2(n16066), .ZN(
        n16068) );
  NAND3_X1 U19164 ( .A1(n16070), .A2(n16069), .A3(n16068), .ZN(P2_U2901) );
  AOI22_X1 U19165 ( .A1(n19039), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n15058), .ZN(n16077) );
  NOR3_X1 U19166 ( .A1(n16071), .A2(n9656), .A3(n16133), .ZN(n16075) );
  OAI22_X1 U19167 ( .A1(n16073), .A2(n16134), .B1(n19047), .B2(n16072), .ZN(
        n16074) );
  NOR2_X1 U19168 ( .A1(n16075), .A2(n16074), .ZN(n16076) );
  OAI211_X1 U19169 ( .C1(n19052), .C2(n16078), .A(n16077), .B(n16076), .ZN(
        P2_U2992) );
  AOI22_X1 U19170 ( .A1(n19039), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n15058), .ZN(n16086) );
  AOI21_X1 U19171 ( .B1(n16168), .B2(n16080), .A(n16079), .ZN(n16167) );
  NOR2_X1 U19172 ( .A1(n16082), .A2(n16081), .ZN(n16083) );
  XNOR2_X1 U19173 ( .A(n16084), .B(n16083), .ZN(n16166) );
  AOI222_X1 U19174 ( .A1(n16167), .A2(n19042), .B1(n19040), .B2(n16166), .C1(
        n16137), .C2(n16165), .ZN(n16085) );
  OAI211_X1 U19175 ( .C1(n19052), .C2(n16087), .A(n16086), .B(n16085), .ZN(
        P2_U3000) );
  AOI22_X1 U19176 ( .A1(n19039), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n15058), .ZN(n16092) );
  AOI222_X1 U19177 ( .A1(n16090), .A2(n19040), .B1(n16137), .B2(n16089), .C1(
        n19042), .C2(n16088), .ZN(n16091) );
  OAI211_X1 U19178 ( .C1(n19052), .C2(n16093), .A(n16092), .B(n16091), .ZN(
        P2_U3002) );
  AOI22_X1 U19179 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n15397), .B1(n16142), 
        .B2(n18840), .ZN(n16098) );
  OAI22_X1 U19180 ( .A1(n16095), .A2(n16133), .B1(n16094), .B2(n16134), .ZN(
        n16096) );
  AOI21_X1 U19181 ( .B1(n16137), .B2(n18844), .A(n16096), .ZN(n16097) );
  OAI211_X1 U19182 ( .C1(n16151), .C2(n20946), .A(n16098), .B(n16097), .ZN(
        P2_U3003) );
  AOI22_X1 U19183 ( .A1(n19039), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n15058), .ZN(n16110) );
  AOI21_X1 U19184 ( .B1(n12109), .B2(n16100), .A(n16099), .ZN(n16181) );
  NAND2_X1 U19185 ( .A1(n15448), .A2(n16101), .ZN(n16106) );
  INV_X1 U19186 ( .A(n16102), .ZN(n16103) );
  NOR2_X1 U19187 ( .A1(n16104), .A2(n16103), .ZN(n16105) );
  XNOR2_X1 U19188 ( .A(n16106), .B(n16105), .ZN(n16184) );
  OAI22_X1 U19189 ( .A1(n16184), .A2(n16134), .B1(n19047), .B2(n16107), .ZN(
        n16108) );
  AOI21_X1 U19190 ( .B1(n16181), .B2(n19042), .A(n16108), .ZN(n16109) );
  OAI211_X1 U19191 ( .C1(n19052), .C2(n18855), .A(n16110), .B(n16109), .ZN(
        P2_U3004) );
  AOI22_X1 U19192 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n15058), .B1(n16142), 
        .B2(n18862), .ZN(n16116) );
  OAI22_X1 U19193 ( .A1(n16112), .A2(n16133), .B1(n16134), .B2(n16111), .ZN(
        n16113) );
  AOI21_X1 U19194 ( .B1(n16137), .B2(n16114), .A(n16113), .ZN(n16115) );
  OAI211_X1 U19195 ( .C1(n16151), .C2(n16117), .A(n16116), .B(n16115), .ZN(
        P2_U3005) );
  AOI22_X1 U19196 ( .A1(n19039), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n15058), .ZN(n16130) );
  NAND2_X1 U19197 ( .A1(n16119), .A2(n16118), .ZN(n16125) );
  INV_X1 U19198 ( .A(n16120), .ZN(n16121) );
  AOI21_X1 U19199 ( .B1(n16123), .B2(n16122), .A(n16121), .ZN(n16124) );
  XOR2_X1 U19200 ( .A(n16125), .B(n16124), .Z(n16192) );
  XOR2_X1 U19201 ( .A(n16127), .B(n16126), .Z(n16186) );
  AOI222_X1 U19202 ( .A1(n16192), .A2(n19040), .B1(n16137), .B2(n16128), .C1(
        n16186), .C2(n19042), .ZN(n16129) );
  OAI211_X1 U19203 ( .C1(n19052), .C2(n16131), .A(n16130), .B(n16129), .ZN(
        P2_U3006) );
  AOI22_X1 U19204 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n15397), .B1(n16142), 
        .B2(n18910), .ZN(n16139) );
  OAI22_X1 U19205 ( .A1(n16135), .A2(n16134), .B1(n16133), .B2(n16132), .ZN(
        n16136) );
  AOI21_X1 U19206 ( .B1(n16137), .B2(n18911), .A(n16136), .ZN(n16138) );
  OAI211_X1 U19207 ( .C1(n16151), .C2(n16140), .A(n16139), .B(n16138), .ZN(
        P2_U3009) );
  AOI22_X1 U19208 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n15058), .B1(n16142), 
        .B2(n16141), .ZN(n16150) );
  NAND3_X1 U19209 ( .A1(n16144), .A2(n16143), .A3(n19042), .ZN(n16145) );
  OAI21_X1 U19210 ( .B1(n19047), .B2(n16146), .A(n16145), .ZN(n16147) );
  AOI21_X1 U19211 ( .B1(n16148), .B2(n19040), .A(n16147), .ZN(n16149) );
  OAI211_X1 U19212 ( .C1(n16152), .C2(n16151), .A(n16150), .B(n16149), .ZN(
        P2_U3011) );
  NOR2_X1 U19213 ( .A1(n19641), .A2(n18885), .ZN(n16157) );
  INV_X1 U19214 ( .A(n16153), .ZN(n16154) );
  OAI22_X1 U19215 ( .A1(n19070), .A2(n16155), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16154), .ZN(n16156) );
  AOI211_X1 U19216 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16158), .A(
        n16157), .B(n16156), .ZN(n16162) );
  AOI22_X1 U19217 ( .A1(n16160), .A2(n19056), .B1(n19067), .B2(n16159), .ZN(
        n16161) );
  OAI211_X1 U19218 ( .C1(n16163), .C2(n16204), .A(n16162), .B(n16161), .ZN(
        P2_U3031) );
  AOI22_X1 U19219 ( .A1(n16164), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16200), .B2(n18943), .ZN(n16174) );
  AOI222_X1 U19220 ( .A1(n16167), .A2(n19056), .B1(n19065), .B2(n16166), .C1(
        n19067), .C2(n16165), .ZN(n16173) );
  NAND2_X1 U19221 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n15058), .ZN(n16172) );
  NAND3_X1 U19222 ( .A1(n16170), .A2(n16169), .A3(n16168), .ZN(n16171) );
  NAND4_X1 U19223 ( .A1(n16174), .A2(n16173), .A3(n16172), .A4(n16171), .ZN(
        P2_U3032) );
  INV_X1 U19224 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19634) );
  NOR2_X1 U19225 ( .A1(n19634), .A2(n18885), .ZN(n16179) );
  XNOR2_X1 U19226 ( .A(n16176), .B(n16175), .ZN(n18952) );
  OAI22_X1 U19227 ( .A1(n16177), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n18952), .B2(n19070), .ZN(n16178) );
  AOI211_X1 U19228 ( .C1(n16180), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16179), .B(n16178), .ZN(n16183) );
  AOI22_X1 U19229 ( .A1(n16181), .A2(n19056), .B1(n19067), .B2(n18857), .ZN(
        n16182) );
  OAI211_X1 U19230 ( .C1(n16184), .C2(n16204), .A(n16183), .B(n16182), .ZN(
        P2_U3036) );
  AOI22_X1 U19231 ( .A1(n16185), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16200), .B2(n18953), .ZN(n16198) );
  INV_X1 U19232 ( .A(n16186), .ZN(n16190) );
  OAI22_X1 U19233 ( .A1(n16190), .A2(n16189), .B1(n16188), .B2(n16187), .ZN(
        n16191) );
  AOI21_X1 U19234 ( .B1(n19065), .B2(n16192), .A(n16191), .ZN(n16197) );
  NAND2_X1 U19235 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n15397), .ZN(n16196) );
  NAND2_X1 U19236 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16193) );
  OAI211_X1 U19237 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16194), .B(n16193), .ZN(n16195) );
  NAND4_X1 U19238 ( .A1(n16198), .A2(n16197), .A3(n16196), .A4(n16195), .ZN(
        P2_U3038) );
  INV_X1 U19239 ( .A(n16199), .ZN(n18988) );
  AOI22_X1 U19240 ( .A1(n19056), .A2(n16201), .B1(n16200), .B2(n18988), .ZN(
        n16208) );
  OAI22_X1 U19241 ( .A1(n16204), .A2(n16203), .B1(n16202), .B2(n19057), .ZN(
        n16205) );
  AOI211_X1 U19242 ( .C1(n19067), .C2(n18928), .A(n16206), .B(n16205), .ZN(
        n16207) );
  OAI211_X1 U19243 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16209), .A(
        n16208), .B(n16207), .ZN(P2_U3046) );
  AOI21_X1 U19244 ( .B1(n19711), .B2(n19710), .A(n16214), .ZN(n16220) );
  AOI211_X1 U19245 ( .C1(n16213), .C2(n16212), .A(n16211), .B(n16210), .ZN(
        n16219) );
  INV_X1 U19246 ( .A(n16214), .ZN(n16217) );
  OAI21_X1 U19247 ( .B1(n16215), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n19732), 
        .ZN(n16216) );
  OAI21_X1 U19248 ( .B1(n16217), .B2(n19600), .A(n16216), .ZN(n16218) );
  OAI211_X1 U19249 ( .C1(n16220), .C2(n13371), .A(n16219), .B(n16218), .ZN(
        P2_U3176) );
  NOR2_X1 U19250 ( .A1(n16222), .A2(n16221), .ZN(n18514) );
  NOR2_X2 U19251 ( .A1(n16232), .A2(n16223), .ZN(n17734) );
  INV_X1 U19252 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18690) );
  AOI22_X1 U19253 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n9876), .B1(
        n17648), .B2(n18690), .ZN(n16231) );
  OAI211_X1 U19254 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n15724), .A(
        n16224), .B(n16227), .ZN(n16225) );
  OAI21_X1 U19255 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18690), .A(
        n16225), .ZN(n16230) );
  NAND2_X1 U19256 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16226), .ZN(
        n16228) );
  NAND3_X1 U19257 ( .A1(n16231), .A2(n16228), .A3(n16227), .ZN(n16229) );
  OAI21_X1 U19258 ( .B1(n16231), .B2(n16230), .A(n16229), .ZN(n16280) );
  INV_X1 U19259 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16447) );
  NAND2_X1 U19260 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16745) );
  NAND2_X1 U19261 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17643) );
  NAND3_X1 U19262 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16233) );
  NOR2_X1 U19263 ( .A1(n17472), .A2(n17462), .ZN(n17461) );
  NOR2_X1 U19264 ( .A1(n17432), .A2(n17422), .ZN(n17417) );
  NAND2_X1 U19265 ( .A1(n17417), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16429) );
  NAND2_X1 U19266 ( .A1(n17374), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17372) );
  INV_X1 U19267 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16234) );
  INV_X1 U19268 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18668) );
  NOR2_X1 U19269 ( .A1(n18668), .A2(n9637), .ZN(n16274) );
  NAND2_X1 U19270 ( .A1(n18584), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17533) );
  INV_X1 U19271 ( .A(n17533), .ZN(n17574) );
  INV_X1 U19272 ( .A(n17588), .ZN(n17507) );
  OR2_X1 U19273 ( .A1(n16236), .A2(n17507), .ZN(n16246) );
  XNOR2_X1 U19274 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16238) );
  NOR2_X1 U19275 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17483), .ZN(
        n16262) );
  NAND2_X1 U19276 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16264), .ZN(
        n16428) );
  AOI22_X1 U19277 ( .A1(n18457), .A2(n16236), .B1(n17574), .B2(n16428), .ZN(
        n16237) );
  NAND2_X1 U19278 ( .A1(n16237), .A2(n17745), .ZN(n16263) );
  NOR2_X1 U19279 ( .A1(n16262), .A2(n16263), .ZN(n16245) );
  OAI22_X1 U19280 ( .A1(n16246), .A2(n16238), .B1(n16245), .B2(n16447), .ZN(
        n16239) );
  AOI211_X1 U19281 ( .C1(n17597), .C2(n16764), .A(n16274), .B(n16239), .ZN(
        n16243) );
  NAND2_X1 U19282 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16255), .ZN(
        n16240) );
  XOR2_X1 U19283 ( .A(n16240), .B(n18690), .Z(n16277) );
  NAND2_X1 U19284 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16257), .ZN(
        n16241) );
  XOR2_X1 U19285 ( .A(n18690), .B(n16241), .Z(n16276) );
  AOI22_X1 U19286 ( .A1(n17738), .A2(n16277), .B1(n17570), .B2(n16276), .ZN(
        n16242) );
  OAI211_X1 U19287 ( .C1(n17650), .C2(n16280), .A(n16243), .B(n16242), .ZN(
        P3_U2799) );
  XNOR2_X1 U19288 ( .A(n9946), .B(n9746), .ZN(n16450) );
  OAI221_X1 U19289 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16246), .C1(
        n9946), .C2(n16245), .A(n16244), .ZN(n16247) );
  AOI21_X1 U19290 ( .B1(n17597), .B2(n16450), .A(n16247), .ZN(n16251) );
  OAI22_X1 U19291 ( .A1(n16255), .A2(n17750), .B1(n16257), .B2(n17649), .ZN(
        n16249) );
  AOI22_X1 U19292 ( .A1(n17602), .A2(n17738), .B1(n17570), .B2(n17914), .ZN(
        n17639) );
  NOR2_X1 U19293 ( .A1(n16283), .A2(n17546), .ZN(n17398) );
  AOI22_X1 U19294 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16249), .B1(
        n16248), .B2(n17398), .ZN(n16250) );
  OAI211_X1 U19295 ( .C1(n17650), .C2(n16252), .A(n16251), .B(n16250), .ZN(
        P3_U2800) );
  INV_X1 U19296 ( .A(n16253), .ZN(n16261) );
  NAND2_X1 U19297 ( .A1(n16254), .A2(n16256), .ZN(n16289) );
  AOI211_X1 U19298 ( .C1(n16258), .C2(n16289), .A(n16255), .B(n17750), .ZN(
        n16260) );
  NAND2_X1 U19299 ( .A1(n16256), .A2(n17759), .ZN(n16287) );
  AOI211_X1 U19300 ( .C1(n16258), .C2(n16287), .A(n16257), .B(n17649), .ZN(
        n16259) );
  AOI211_X1 U19301 ( .C1(n16261), .C2(n17636), .A(n16260), .B(n16259), .ZN(
        n16268) );
  NAND2_X1 U19302 ( .A1(n16286), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16267) );
  AOI21_X1 U19303 ( .B1(n9945), .B2(n16428), .A(n9746), .ZN(n16459) );
  OAI21_X1 U19304 ( .B1(n16262), .B2(n17597), .A(n16459), .ZN(n16266) );
  OAI221_X1 U19305 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16264), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18457), .A(n16263), .ZN(
        n16265) );
  NAND4_X1 U19306 ( .A1(n16268), .A2(n16267), .A3(n16266), .A4(n16265), .ZN(
        P3_U2801) );
  INV_X1 U19307 ( .A(n16269), .ZN(n18053) );
  OAI21_X1 U19308 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18053), .A(
        n16270), .ZN(n16275) );
  NOR4_X1 U19309 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16272), .A3(
        n15724), .A4(n16271), .ZN(n16273) );
  AOI211_X1 U19310 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16275), .A(
        n16274), .B(n16273), .ZN(n16279) );
  INV_X1 U19311 ( .A(n18068), .ZN(n18010) );
  AOI22_X1 U19312 ( .A1(n16277), .A2(n18010), .B1(n16276), .B2(n17908), .ZN(
        n16278) );
  OAI211_X1 U19313 ( .C1(n16280), .C2(n17982), .A(n16279), .B(n16278), .ZN(
        P3_U2831) );
  AOI22_X1 U19314 ( .A1(n17602), .A2(n18509), .B1(n17914), .B2(n17938), .ZN(
        n17857) );
  INV_X1 U19315 ( .A(n17857), .ZN(n16281) );
  AOI21_X1 U19316 ( .B1(n16282), .B2(n16281), .A(n17774), .ZN(n17799) );
  NOR2_X1 U19317 ( .A1(n18065), .A2(n17799), .ZN(n17784) );
  NOR3_X1 U19318 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17760), .A3(
        n16283), .ZN(n17382) );
  AOI22_X1 U19319 ( .A1(n18017), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17784), 
        .B2(n17382), .ZN(n16299) );
  NOR2_X1 U19320 ( .A1(n18065), .A2(n18515), .ZN(n18064) );
  NAND3_X1 U19321 ( .A1(n16285), .A2(n18064), .A3(n16290), .ZN(n16298) );
  AOI21_X1 U19322 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17648), .A(
        n16285), .ZN(n16291) );
  NAND3_X1 U19323 ( .A1(n17391), .A2(n17967), .A3(n16291), .ZN(n16297) );
  INV_X1 U19324 ( .A(n16287), .ZN(n16295) );
  INV_X1 U19325 ( .A(n17938), .ZN(n17913) );
  AOI211_X1 U19326 ( .C1(n18509), .C2(n16289), .A(n18058), .B(n16288), .ZN(
        n16294) );
  INV_X1 U19327 ( .A(n16290), .ZN(n17386) );
  INV_X1 U19328 ( .A(n16291), .ZN(n17385) );
  NAND4_X1 U19329 ( .A1(n16299), .A2(n16298), .A3(n16297), .A4(n16296), .ZN(
        P3_U2834) );
  NOR3_X1 U19330 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16301) );
  NOR4_X1 U19331 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16300) );
  NAND4_X1 U19332 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16301), .A3(n16300), .A4(
        U215), .ZN(U213) );
  INV_X1 U19333 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18994) );
  INV_X2 U19334 ( .A(U214), .ZN(n16361) );
  INV_X1 U19335 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16303) );
  OAI222_X1 U19336 ( .A1(U212), .A2(n18994), .B1(n16363), .B2(n16304), .C1(
        U214), .C2(n16303), .ZN(U216) );
  INV_X1 U19337 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16397) );
  OAI222_X1 U19338 ( .A1(U212), .A2(n18999), .B1(n16363), .B2(n16305), .C1(
        U214), .C2(n16397), .ZN(U217) );
  INV_X1 U19339 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16307) );
  AOI22_X1 U19340 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16360), .ZN(n16306) );
  OAI21_X1 U19341 ( .B1(n16307), .B2(n16363), .A(n16306), .ZN(U218) );
  INV_X1 U19342 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16309) );
  AOI22_X1 U19343 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16360), .ZN(n16308) );
  OAI21_X1 U19344 ( .B1(n16309), .B2(n16363), .A(n16308), .ZN(U219) );
  AOI22_X1 U19345 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16360), .ZN(n16310) );
  OAI21_X1 U19346 ( .B1(n16311), .B2(n16363), .A(n16310), .ZN(U220) );
  AOI22_X1 U19347 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16360), .ZN(n16312) );
  OAI21_X1 U19348 ( .B1(n16313), .B2(n16363), .A(n16312), .ZN(U221) );
  AOI22_X1 U19349 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16360), .ZN(n16314) );
  OAI21_X1 U19350 ( .B1(n16315), .B2(n16363), .A(n16314), .ZN(U222) );
  INV_X1 U19351 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16317) );
  AOI22_X1 U19352 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16360), .ZN(n16316) );
  OAI21_X1 U19353 ( .B1(n16317), .B2(n16363), .A(n16316), .ZN(U223) );
  INV_X1 U19354 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16319) );
  AOI22_X1 U19355 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16360), .ZN(n16318) );
  OAI21_X1 U19356 ( .B1(n16319), .B2(n16363), .A(n16318), .ZN(U224) );
  AOI22_X1 U19357 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16360), .ZN(n16320) );
  OAI21_X1 U19358 ( .B1(n16321), .B2(n16363), .A(n16320), .ZN(U225) );
  AOI22_X1 U19359 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16360), .ZN(n16322) );
  OAI21_X1 U19360 ( .B1(n16323), .B2(n16363), .A(n16322), .ZN(U226) );
  INV_X1 U19361 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16325) );
  AOI22_X1 U19362 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16360), .ZN(n16324) );
  OAI21_X1 U19363 ( .B1(n16325), .B2(n16363), .A(n16324), .ZN(U227) );
  AOI22_X1 U19364 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16360), .ZN(n16326) );
  OAI21_X1 U19365 ( .B1(n16327), .B2(n16363), .A(n16326), .ZN(U228) );
  AOI22_X1 U19366 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16360), .ZN(n16328) );
  OAI21_X1 U19367 ( .B1(n16329), .B2(n16363), .A(n16328), .ZN(U229) );
  INV_X1 U19368 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16331) );
  AOI22_X1 U19369 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16360), .ZN(n16330) );
  OAI21_X1 U19370 ( .B1(n16331), .B2(n16363), .A(n16330), .ZN(U230) );
  AOI22_X1 U19371 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16360), .ZN(n16332) );
  OAI21_X1 U19372 ( .B1(n16333), .B2(n16363), .A(n16332), .ZN(U231) );
  AOI22_X1 U19373 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16360), .ZN(n16334) );
  OAI21_X1 U19374 ( .B1(n12956), .B2(n16363), .A(n16334), .ZN(U232) );
  AOI22_X1 U19375 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16360), .ZN(n16335) );
  OAI21_X1 U19376 ( .B1(n12609), .B2(n16363), .A(n16335), .ZN(U233) );
  AOI22_X1 U19377 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16360), .ZN(n16336) );
  OAI21_X1 U19378 ( .B1(n12721), .B2(n16363), .A(n16336), .ZN(U234) );
  AOI22_X1 U19379 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16360), .ZN(n16337) );
  OAI21_X1 U19380 ( .B1(n16338), .B2(n16363), .A(n16337), .ZN(U235) );
  INV_X1 U19381 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16340) );
  AOI22_X1 U19382 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16360), .ZN(n16339) );
  OAI21_X1 U19383 ( .B1(n16340), .B2(n16363), .A(n16339), .ZN(U236) );
  AOI22_X1 U19384 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16360), .ZN(n16341) );
  OAI21_X1 U19385 ( .B1(n16342), .B2(n16363), .A(n16341), .ZN(U237) );
  INV_X1 U19386 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16344) );
  AOI22_X1 U19387 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16360), .ZN(n16343) );
  OAI21_X1 U19388 ( .B1(n16344), .B2(n16363), .A(n16343), .ZN(U238) );
  AOI22_X1 U19389 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16360), .ZN(n16345) );
  OAI21_X1 U19390 ( .B1(n16346), .B2(n16363), .A(n16345), .ZN(U239) );
  INV_X1 U19391 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16348) );
  AOI22_X1 U19392 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16360), .ZN(n16347) );
  OAI21_X1 U19393 ( .B1(n16348), .B2(n16363), .A(n16347), .ZN(U240) );
  INV_X1 U19394 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16350) );
  AOI22_X1 U19395 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16360), .ZN(n16349) );
  OAI21_X1 U19396 ( .B1(n16350), .B2(n16363), .A(n16349), .ZN(U241) );
  INV_X1 U19397 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16352) );
  AOI22_X1 U19398 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16360), .ZN(n16351) );
  OAI21_X1 U19399 ( .B1(n16352), .B2(n16363), .A(n16351), .ZN(U242) );
  INV_X1 U19400 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16354) );
  AOI22_X1 U19401 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16360), .ZN(n16353) );
  OAI21_X1 U19402 ( .B1(n16354), .B2(n16363), .A(n16353), .ZN(U243) );
  INV_X1 U19403 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16356) );
  AOI22_X1 U19404 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16360), .ZN(n16355) );
  OAI21_X1 U19405 ( .B1(n16356), .B2(n16363), .A(n16355), .ZN(U244) );
  INV_X1 U19406 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20916) );
  AOI22_X1 U19407 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16360), .ZN(n16357) );
  OAI21_X1 U19408 ( .B1(n20916), .B2(n16363), .A(n16357), .ZN(U245) );
  INV_X1 U19409 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16359) );
  AOI22_X1 U19410 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16360), .ZN(n16358) );
  OAI21_X1 U19411 ( .B1(n16359), .B2(n16363), .A(n16358), .ZN(U246) );
  INV_X1 U19412 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16364) );
  AOI22_X1 U19413 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16361), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16360), .ZN(n16362) );
  OAI21_X1 U19414 ( .B1(n16364), .B2(n16363), .A(n16362), .ZN(U247) );
  OAI22_X1 U19415 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16395), .ZN(n16365) );
  INV_X1 U19416 ( .A(n16365), .ZN(U251) );
  OAI22_X1 U19417 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16395), .ZN(n16366) );
  INV_X1 U19418 ( .A(n16366), .ZN(U252) );
  OAI22_X1 U19419 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16395), .ZN(n16367) );
  INV_X1 U19420 ( .A(n16367), .ZN(U253) );
  OAI22_X1 U19421 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16395), .ZN(n16368) );
  INV_X1 U19422 ( .A(n16368), .ZN(U254) );
  INV_X1 U19423 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n20786) );
  INV_X1 U19424 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18101) );
  AOI22_X1 U19425 ( .A1(n16395), .A2(n20786), .B1(n18101), .B2(U215), .ZN(U255) );
  OAI22_X1 U19426 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16395), .ZN(n16369) );
  INV_X1 U19427 ( .A(n16369), .ZN(U256) );
  OAI22_X1 U19428 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16395), .ZN(n16370) );
  INV_X1 U19429 ( .A(n16370), .ZN(U257) );
  OAI22_X1 U19430 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16395), .ZN(n16371) );
  INV_X1 U19431 ( .A(n16371), .ZN(U258) );
  OAI22_X1 U19432 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16395), .ZN(n16372) );
  INV_X1 U19433 ( .A(n16372), .ZN(U259) );
  OAI22_X1 U19434 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16395), .ZN(n16373) );
  INV_X1 U19435 ( .A(n16373), .ZN(U260) );
  OAI22_X1 U19436 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16387), .ZN(n16374) );
  INV_X1 U19437 ( .A(n16374), .ZN(U261) );
  OAI22_X1 U19438 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16387), .ZN(n16375) );
  INV_X1 U19439 ( .A(n16375), .ZN(U262) );
  OAI22_X1 U19440 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16395), .ZN(n16376) );
  INV_X1 U19441 ( .A(n16376), .ZN(U263) );
  OAI22_X1 U19442 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16387), .ZN(n16377) );
  INV_X1 U19443 ( .A(n16377), .ZN(U264) );
  OAI22_X1 U19444 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16395), .ZN(n16378) );
  INV_X1 U19445 ( .A(n16378), .ZN(U265) );
  OAI22_X1 U19446 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16395), .ZN(n16379) );
  INV_X1 U19447 ( .A(n16379), .ZN(U266) );
  OAI22_X1 U19448 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16387), .ZN(n16380) );
  INV_X1 U19449 ( .A(n16380), .ZN(U267) );
  OAI22_X1 U19450 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16387), .ZN(n16381) );
  INV_X1 U19451 ( .A(n16381), .ZN(U268) );
  OAI22_X1 U19452 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16387), .ZN(n16382) );
  INV_X1 U19453 ( .A(n16382), .ZN(U269) );
  OAI22_X1 U19454 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16387), .ZN(n16383) );
  INV_X1 U19455 ( .A(n16383), .ZN(U270) );
  OAI22_X1 U19456 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16387), .ZN(n16384) );
  INV_X1 U19457 ( .A(n16384), .ZN(U271) );
  OAI22_X1 U19458 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16387), .ZN(n16385) );
  INV_X1 U19459 ( .A(n16385), .ZN(U272) );
  OAI22_X1 U19460 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16395), .ZN(n16386) );
  INV_X1 U19461 ( .A(n16386), .ZN(U273) );
  OAI22_X1 U19462 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16387), .ZN(n16388) );
  INV_X1 U19463 ( .A(n16388), .ZN(U274) );
  OAI22_X1 U19464 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16395), .ZN(n16389) );
  INV_X1 U19465 ( .A(n16389), .ZN(U275) );
  OAI22_X1 U19466 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16395), .ZN(n16390) );
  INV_X1 U19467 ( .A(n16390), .ZN(U276) );
  OAI22_X1 U19468 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16395), .ZN(n16391) );
  INV_X1 U19469 ( .A(n16391), .ZN(U277) );
  OAI22_X1 U19470 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16395), .ZN(n16392) );
  INV_X1 U19471 ( .A(n16392), .ZN(U278) );
  OAI22_X1 U19472 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16395), .ZN(n16393) );
  INV_X1 U19473 ( .A(n16393), .ZN(U279) );
  OAI22_X1 U19474 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16395), .ZN(n16394) );
  INV_X1 U19475 ( .A(n16394), .ZN(U280) );
  AOI22_X1 U19476 ( .A1(n16395), .A2(n18999), .B1(n18110), .B2(U215), .ZN(U281) );
  AOI22_X1 U19477 ( .A1(n16395), .A2(n18994), .B1(n18116), .B2(U215), .ZN(U282) );
  INV_X1 U19478 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16396) );
  OAI222_X1 U19479 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n16397), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n18999), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n16396), .ZN(n16398) );
  INV_X2 U19480 ( .A(n20962), .ZN(n20963) );
  INV_X1 U19481 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18628) );
  INV_X1 U19482 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19635) );
  AOI22_X1 U19483 ( .A1(n20963), .A2(n18628), .B1(n19635), .B2(n20962), .ZN(
        U347) );
  INV_X1 U19484 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18626) );
  INV_X1 U19485 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19633) );
  AOI22_X1 U19486 ( .A1(n20963), .A2(n18626), .B1(n19633), .B2(n20962), .ZN(
        U348) );
  INV_X1 U19487 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18623) );
  INV_X1 U19488 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19632) );
  AOI22_X1 U19489 ( .A1(n20963), .A2(n18623), .B1(n19632), .B2(n20962), .ZN(
        U349) );
  INV_X1 U19490 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18622) );
  INV_X1 U19491 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19631) );
  AOI22_X1 U19492 ( .A1(n20963), .A2(n18622), .B1(n19631), .B2(n20962), .ZN(
        U350) );
  INV_X1 U19493 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18620) );
  INV_X1 U19494 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19629) );
  AOI22_X1 U19495 ( .A1(n20963), .A2(n18620), .B1(n19629), .B2(n20962), .ZN(
        U351) );
  INV_X1 U19496 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18617) );
  INV_X1 U19497 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19627) );
  AOI22_X1 U19498 ( .A1(n20963), .A2(n18617), .B1(n19627), .B2(n20962), .ZN(
        U352) );
  INV_X1 U19499 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18616) );
  INV_X1 U19500 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19626) );
  AOI22_X1 U19501 ( .A1(n20963), .A2(n18616), .B1(n19626), .B2(n20962), .ZN(
        U353) );
  INV_X1 U19502 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18614) );
  AOI22_X1 U19503 ( .A1(n20963), .A2(n18614), .B1(n19624), .B2(n20962), .ZN(
        U354) );
  INV_X1 U19504 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18670) );
  INV_X1 U19505 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19670) );
  AOI22_X1 U19506 ( .A1(n20963), .A2(n18670), .B1(n19670), .B2(n16398), .ZN(
        U355) );
  INV_X1 U19507 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18667) );
  INV_X1 U19508 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19667) );
  AOI22_X1 U19509 ( .A1(n20963), .A2(n18667), .B1(n19667), .B2(n16398), .ZN(
        U356) );
  INV_X1 U19510 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18665) );
  INV_X1 U19511 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19665) );
  AOI22_X1 U19512 ( .A1(n20963), .A2(n18665), .B1(n19665), .B2(n20962), .ZN(
        U357) );
  INV_X1 U19513 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18663) );
  INV_X1 U19514 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19662) );
  AOI22_X1 U19515 ( .A1(n20963), .A2(n18663), .B1(n19662), .B2(n20962), .ZN(
        U358) );
  INV_X1 U19516 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18661) );
  INV_X1 U19517 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19661) );
  AOI22_X1 U19518 ( .A1(n20963), .A2(n18661), .B1(n19661), .B2(n20962), .ZN(
        U359) );
  INV_X1 U19519 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18659) );
  INV_X1 U19520 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19659) );
  AOI22_X1 U19521 ( .A1(n20963), .A2(n18659), .B1(n19659), .B2(n20962), .ZN(
        U360) );
  INV_X1 U19522 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18656) );
  INV_X1 U19523 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19657) );
  AOI22_X1 U19524 ( .A1(n20963), .A2(n18656), .B1(n19657), .B2(n20962), .ZN(
        U361) );
  INV_X1 U19525 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18653) );
  INV_X1 U19526 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19655) );
  AOI22_X1 U19527 ( .A1(n20963), .A2(n18653), .B1(n19655), .B2(n20962), .ZN(
        U362) );
  INV_X1 U19528 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18652) );
  INV_X1 U19529 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19653) );
  AOI22_X1 U19530 ( .A1(n20963), .A2(n18652), .B1(n19653), .B2(n20962), .ZN(
        U363) );
  INV_X1 U19531 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18649) );
  INV_X1 U19532 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19652) );
  AOI22_X1 U19533 ( .A1(n20963), .A2(n18649), .B1(n19652), .B2(n20962), .ZN(
        U364) );
  INV_X1 U19534 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18612) );
  INV_X1 U19535 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19623) );
  AOI22_X1 U19536 ( .A1(n20963), .A2(n18612), .B1(n19623), .B2(n16398), .ZN(
        U365) );
  INV_X1 U19537 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18648) );
  INV_X1 U19538 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U19539 ( .A1(n20963), .A2(n18648), .B1(n19650), .B2(n16398), .ZN(
        U366) );
  INV_X1 U19540 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18646) );
  INV_X1 U19541 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19649) );
  AOI22_X1 U19542 ( .A1(n20963), .A2(n18646), .B1(n19649), .B2(n16398), .ZN(
        U367) );
  INV_X1 U19543 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18644) );
  INV_X1 U19544 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19647) );
  AOI22_X1 U19545 ( .A1(n20963), .A2(n18644), .B1(n19647), .B2(n16398), .ZN(
        U368) );
  INV_X1 U19546 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18642) );
  INV_X1 U19547 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19645) );
  AOI22_X1 U19548 ( .A1(n20963), .A2(n18642), .B1(n19645), .B2(n16398), .ZN(
        U369) );
  INV_X1 U19549 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18640) );
  INV_X1 U19550 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19643) );
  AOI22_X1 U19551 ( .A1(n20963), .A2(n18640), .B1(n19643), .B2(n16398), .ZN(
        U370) );
  INV_X1 U19552 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18638) );
  INV_X1 U19553 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19642) );
  AOI22_X1 U19554 ( .A1(n20963), .A2(n18638), .B1(n19642), .B2(n20962), .ZN(
        U371) );
  INV_X1 U19555 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18636) );
  INV_X1 U19556 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U19557 ( .A1(n20963), .A2(n18636), .B1(n19640), .B2(n20962), .ZN(
        U372) );
  INV_X1 U19558 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18634) );
  INV_X1 U19559 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19639) );
  AOI22_X1 U19560 ( .A1(n20963), .A2(n18634), .B1(n19639), .B2(n20962), .ZN(
        U373) );
  INV_X1 U19561 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18632) );
  INV_X1 U19562 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19638) );
  AOI22_X1 U19563 ( .A1(n20963), .A2(n18632), .B1(n19638), .B2(n20962), .ZN(
        U374) );
  INV_X1 U19564 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18610) );
  INV_X1 U19565 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19621) );
  AOI22_X1 U19566 ( .A1(n20963), .A2(n18610), .B1(n19621), .B2(n20962), .ZN(
        U376) );
  INV_X1 U19567 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18609) );
  NAND2_X1 U19568 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18609), .ZN(n18596) );
  AOI22_X1 U19569 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18596), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18607), .ZN(n18676) );
  AOI21_X1 U19570 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18676), .ZN(n16399) );
  INV_X1 U19571 ( .A(n16399), .ZN(P3_U2633) );
  INV_X1 U19572 ( .A(n16405), .ZN(n16400) );
  OAI21_X1 U19573 ( .B1(n16400), .B2(n17303), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16401) );
  OAI21_X1 U19574 ( .B1(n16402), .B2(n16423), .A(n16401), .ZN(P3_U2634) );
  AOI21_X1 U19575 ( .B1(n18607), .B2(n18609), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16403) );
  AOI22_X1 U19576 ( .A1(n18669), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16403), 
        .B2(n18740), .ZN(P3_U2635) );
  NOR2_X1 U19577 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18592) );
  OAI21_X1 U19578 ( .B1(n18592), .B2(BS16), .A(n18676), .ZN(n18674) );
  OAI21_X1 U19579 ( .B1(n18676), .B2(n18731), .A(n18674), .ZN(P3_U2636) );
  AND3_X1 U19580 ( .A1(n16405), .A2(n18513), .A3(n16404), .ZN(n18516) );
  NOR2_X1 U19581 ( .A1(n18516), .A2(n18581), .ZN(n18723) );
  INV_X1 U19582 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16407) );
  OAI21_X1 U19583 ( .B1(n18723), .B2(n16407), .A(n16406), .ZN(P3_U2637) );
  INV_X1 U19584 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18721) );
  NOR4_X1 U19585 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16411) );
  NOR4_X1 U19586 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16410) );
  NOR4_X1 U19587 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16409) );
  NOR4_X1 U19588 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16408) );
  NAND4_X1 U19589 ( .A1(n16411), .A2(n16410), .A3(n16409), .A4(n16408), .ZN(
        n16417) );
  NOR4_X1 U19590 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16415) );
  AOI211_X1 U19591 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_5__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16414) );
  NOR4_X1 U19592 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16413) );
  NOR4_X1 U19593 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16412) );
  NAND4_X1 U19594 ( .A1(n16415), .A2(n16414), .A3(n16413), .A4(n16412), .ZN(
        n16416) );
  NOR2_X1 U19595 ( .A1(n16417), .A2(n16416), .ZN(n18718) );
  INV_X1 U19596 ( .A(n18718), .ZN(n18720) );
  INV_X1 U19597 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18712) );
  NAND2_X1 U19598 ( .A1(n18718), .A2(n18712), .ZN(n18717) );
  NOR3_X1 U19599 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(n18717), .ZN(n16419) );
  AOI21_X1 U19600 ( .B1(P3_BYTEENABLE_REG_1__SCAN_IN), .B2(n18720), .A(n16419), 
        .ZN(n16418) );
  OAI21_X1 U19601 ( .B1(n18721), .B2(n18720), .A(n16418), .ZN(P3_U2638) );
  NAND2_X1 U19602 ( .A1(n18718), .A2(n18721), .ZN(n18710) );
  AOI21_X1 U19603 ( .B1(P3_BYTEENABLE_REG_3__SCAN_IN), .B2(n18720), .A(n16419), 
        .ZN(n16420) );
  OAI21_X1 U19604 ( .B1(P3_DATAWIDTH_REG_1__SCAN_IN), .B2(n18710), .A(n16420), 
        .ZN(P3_U2639) );
  NOR2_X1 U19605 ( .A1(n18679), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18571) );
  INV_X1 U19606 ( .A(n18571), .ZN(n18451) );
  NOR3_X1 U19607 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18590) );
  NOR2_X1 U19608 ( .A1(n16286), .A2(n18585), .ZN(n16422) );
  INV_X1 U19609 ( .A(n18746), .ZN(n18725) );
  AOI211_X1 U19610 ( .C1(n18732), .C2(n18730), .A(n18599), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16424) );
  AOI211_X1 U19611 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18085), .A(n16424), .B(
        n16427), .ZN(n16569) );
  INV_X1 U19612 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18671) );
  INV_X1 U19613 ( .A(n16424), .ZN(n18575) );
  INV_X1 U19614 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18658) );
  INV_X1 U19615 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18654) );
  INV_X1 U19616 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18650) );
  INV_X1 U19617 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18641) );
  INV_X1 U19618 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18639) );
  INV_X1 U19619 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18637) );
  INV_X1 U19620 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18631) );
  INV_X1 U19621 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18618) );
  INV_X1 U19622 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18613) );
  INV_X1 U19623 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18611) );
  NOR2_X1 U19624 ( .A1(n18721), .A2(n18611), .ZN(n16762) );
  INV_X1 U19625 ( .A(n16762), .ZN(n16777) );
  NOR2_X1 U19626 ( .A1(n18613), .A2(n16777), .ZN(n16759) );
  NAND2_X1 U19627 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16759), .ZN(n16658) );
  NOR2_X1 U19628 ( .A1(n18618), .A2(n16658), .ZN(n16675) );
  INV_X1 U19629 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18629) );
  INV_X1 U19630 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18624) );
  NAND2_X1 U19631 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16718) );
  NOR2_X1 U19632 ( .A1(n18624), .A2(n16718), .ZN(n16680) );
  NAND3_X1 U19633 ( .A1(n16680), .A2(P3_REIP_REG_10__SCAN_IN), .A3(
        P3_REIP_REG_9__SCAN_IN), .ZN(n16659) );
  NOR2_X1 U19634 ( .A1(n18629), .A2(n16659), .ZN(n16642) );
  NAND2_X1 U19635 ( .A1(n16675), .A2(n16642), .ZN(n16646) );
  NOR2_X1 U19636 ( .A1(n18631), .A2(n16646), .ZN(n16624) );
  NAND3_X1 U19637 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16624), .ZN(n16602) );
  NOR4_X1 U19638 ( .A1(n18641), .A2(n18639), .A3(n18637), .A4(n16602), .ZN(
        n16570) );
  NAND4_X1 U19639 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n16570), .ZN(n16535) );
  NOR2_X1 U19640 ( .A1(n18650), .A2(n16535), .ZN(n16534) );
  NAND2_X1 U19641 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16534), .ZN(n16525) );
  NOR2_X1 U19642 ( .A1(n18654), .A2(n16525), .ZN(n16523) );
  NAND2_X1 U19643 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16523), .ZN(n16504) );
  NOR2_X1 U19644 ( .A1(n18658), .A2(n16504), .ZN(n16491) );
  NAND2_X1 U19645 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16491), .ZN(n16440) );
  NAND4_X1 U19646 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_28__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16469), .ZN(n16443) );
  NOR3_X1 U19647 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18671), .A3(n16443), 
        .ZN(n16425) );
  AOI21_X1 U19648 ( .B1(n16569), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16425), .ZN(
        n16446) );
  NAND2_X1 U19649 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18085), .ZN(n16426) );
  AOI211_X4 U19650 ( .C1(n18731), .C2(n18733), .A(n16427), .B(n16426), .ZN(
        n16806) );
  NOR3_X1 U19651 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16775) );
  INV_X1 U19652 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16769) );
  NAND2_X1 U19653 ( .A1(n16775), .A2(n16769), .ZN(n16768) );
  NOR2_X1 U19654 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16768), .ZN(n16751) );
  NAND2_X1 U19655 ( .A1(n16751), .A2(n16738), .ZN(n16737) );
  NOR2_X1 U19656 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16737), .ZN(n16722) );
  NAND2_X1 U19657 ( .A1(n16722), .A2(n16715), .ZN(n16708) );
  NOR2_X1 U19658 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16708), .ZN(n16690) );
  NAND2_X1 U19659 ( .A1(n16690), .A2(n17036), .ZN(n16673) );
  NAND2_X1 U19660 ( .A1(n16672), .A2(n16671), .ZN(n16663) );
  NAND2_X1 U19661 ( .A1(n16647), .A2(n16637), .ZN(n16636) );
  INV_X1 U19662 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16620) );
  NAND2_X1 U19663 ( .A1(n16626), .A2(n16620), .ZN(n16619) );
  NAND2_X1 U19664 ( .A1(n16600), .A2(n16593), .ZN(n16592) );
  INV_X1 U19665 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16566) );
  NAND2_X1 U19666 ( .A1(n16577), .A2(n16566), .ZN(n16565) );
  INV_X1 U19667 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20809) );
  NAND2_X1 U19668 ( .A1(n16555), .A2(n20809), .ZN(n16550) );
  NAND2_X1 U19669 ( .A1(n16536), .A2(n16529), .ZN(n16528) );
  NAND2_X1 U19670 ( .A1(n16513), .A2(n16508), .ZN(n16507) );
  NOR2_X1 U19671 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16507), .ZN(n16492) );
  INV_X1 U19672 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16486) );
  NAND2_X1 U19673 ( .A1(n16492), .A2(n16486), .ZN(n16485) );
  NOR2_X1 U19674 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16485), .ZN(n16470) );
  INV_X1 U19675 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16465) );
  NAND2_X1 U19676 ( .A1(n16470), .A2(n16465), .ZN(n16448) );
  NOR2_X1 U19677 ( .A1(n16805), .A2(n16448), .ZN(n16454) );
  INV_X1 U19678 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16818) );
  NOR2_X1 U19679 ( .A1(n17741), .A2(n17372), .ZN(n16430) );
  OAI21_X1 U19680 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16430), .A(
        n16428), .ZN(n17379) );
  INV_X1 U19681 ( .A(n17379), .ZN(n16473) );
  INV_X1 U19682 ( .A(n17419), .ZN(n17416) );
  NAND2_X1 U19683 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17416), .ZN(
        n16434) );
  NOR2_X1 U19684 ( .A1(n16429), .A2(n16434), .ZN(n16432) );
  INV_X1 U19685 ( .A(n16430), .ZN(n16431) );
  OAI21_X1 U19686 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16432), .A(
        n16431), .ZN(n17393) );
  INV_X1 U19687 ( .A(n17393), .ZN(n16482) );
  INV_X1 U19688 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17407) );
  INV_X1 U19689 ( .A(n16434), .ZN(n16435) );
  NAND2_X1 U19690 ( .A1(n17417), .A2(n16435), .ZN(n17376) );
  AOI21_X1 U19691 ( .B1(n17407), .B2(n17376), .A(n16432), .ZN(n17403) );
  NOR2_X1 U19692 ( .A1(n17432), .A2(n16434), .ZN(n16433) );
  OAI21_X1 U19693 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16433), .A(
        n17376), .ZN(n17421) );
  INV_X1 U19694 ( .A(n17421), .ZN(n16502) );
  AOI21_X1 U19695 ( .B1(n17432), .B2(n16434), .A(n16433), .ZN(n17439) );
  NAND2_X1 U19696 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9716), .ZN(
        n16437) );
  INV_X1 U19697 ( .A(n16437), .ZN(n16438) );
  NAND2_X1 U19698 ( .A1(n17461), .A2(n16438), .ZN(n17418) );
  AOI21_X1 U19699 ( .B1(n9952), .B2(n17418), .A(n16435), .ZN(n17441) );
  NOR2_X1 U19700 ( .A1(n17472), .A2(n16437), .ZN(n16436) );
  OAI21_X1 U19701 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16436), .A(
        n17418), .ZN(n17465) );
  INV_X1 U19702 ( .A(n17465), .ZN(n16539) );
  AOI22_X1 U19703 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16437), .B1(
        n16438), .B2(n17472), .ZN(n17469) );
  INV_X1 U19704 ( .A(n17469), .ZN(n16547) );
  NAND3_X1 U19705 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16604), .A3(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16578) );
  INV_X1 U19706 ( .A(n16578), .ZN(n17493) );
  NAND3_X1 U19707 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n17493), .ZN(n17460) );
  AOI21_X1 U19708 ( .B1(n17486), .B2(n17460), .A(n16438), .ZN(n17489) );
  INV_X1 U19709 ( .A(n17460), .ZN(n16439) );
  INV_X1 U19710 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16795) );
  AOI21_X1 U19711 ( .B1(n16439), .B2(n16795), .A(n16734), .ZN(n16558) );
  NOR2_X1 U19712 ( .A1(n17489), .A2(n16558), .ZN(n16557) );
  NOR2_X1 U19713 ( .A1(n16557), .A2(n16734), .ZN(n16546) );
  NOR2_X1 U19714 ( .A1(n17441), .A2(n16522), .ZN(n16521) );
  NOR2_X1 U19715 ( .A1(n16501), .A2(n16734), .ZN(n16494) );
  NOR2_X1 U19716 ( .A1(n17403), .A2(n16494), .ZN(n16493) );
  NOR2_X1 U19717 ( .A1(n16493), .A2(n16734), .ZN(n16481) );
  NOR2_X1 U19718 ( .A1(n16482), .A2(n16481), .ZN(n16480) );
  NOR2_X1 U19719 ( .A1(n16480), .A2(n16734), .ZN(n16472) );
  NOR2_X1 U19720 ( .A1(n16473), .A2(n16472), .ZN(n16471) );
  NOR2_X1 U19721 ( .A1(n16471), .A2(n16734), .ZN(n16458) );
  NOR2_X1 U19722 ( .A1(n16459), .A2(n16458), .ZN(n16457) );
  NAND2_X1 U19723 ( .A1(n16764), .A2(n18585), .ZN(n16794) );
  NAND3_X1 U19724 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(P3_REIP_REG_28__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16442) );
  NAND2_X1 U19725 ( .A1(n16778), .A2(n16440), .ZN(n16441) );
  NAND2_X1 U19726 ( .A1(n16809), .A2(n16441), .ZN(n16484) );
  AOI21_X1 U19727 ( .B1(n16778), .B2(n16442), .A(n16484), .ZN(n16468) );
  NOR2_X1 U19728 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16443), .ZN(n16452) );
  INV_X1 U19729 ( .A(n16452), .ZN(n16444) );
  AOI21_X1 U19730 ( .B1(n16468), .B2(n16444), .A(n18668), .ZN(n16445) );
  NAND2_X1 U19731 ( .A1(n16806), .A2(n16448), .ZN(n16463) );
  XOR2_X1 U19732 ( .A(n16450), .B(n16449), .Z(n16453) );
  OAI22_X1 U19733 ( .A1(n16468), .A2(n18671), .B1(n9946), .B2(n16793), .ZN(
        n16451) );
  AOI211_X1 U19734 ( .C1(n16453), .C2(n18585), .A(n16452), .B(n16451), .ZN(
        n16456) );
  OAI21_X1 U19735 ( .B1(n16807), .B2(n16454), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16455) );
  OAI211_X1 U19736 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16463), .A(n16456), .B(
        n16455), .ZN(P3_U2641) );
  INV_X1 U19737 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18666) );
  AOI211_X1 U19738 ( .C1(n16459), .C2(n16458), .A(n16457), .B(n16757), .ZN(
        n16462) );
  NAND3_X1 U19739 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16469), .ZN(n16460) );
  OAI22_X1 U19740 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16460), .B1(n9945), 
        .B2(n16793), .ZN(n16461) );
  AOI211_X1 U19741 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16807), .A(n16462), .B(
        n16461), .ZN(n16467) );
  INV_X1 U19742 ( .A(n16463), .ZN(n16464) );
  OAI21_X1 U19743 ( .B1(n16470), .B2(n16465), .A(n16464), .ZN(n16466) );
  OAI211_X1 U19744 ( .C1(n16468), .C2(n18666), .A(n16467), .B(n16466), .ZN(
        P3_U2642) );
  NAND2_X1 U19745 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16469), .ZN(n16479) );
  AOI22_X1 U19746 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16784), .B1(
        n16807), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16478) );
  INV_X1 U19747 ( .A(n16484), .ZN(n16500) );
  INV_X1 U19748 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18662) );
  NAND2_X1 U19749 ( .A1(n16469), .A2(n18662), .ZN(n16488) );
  NAND2_X1 U19750 ( .A1(n16500), .A2(n16488), .ZN(n16476) );
  AOI211_X1 U19751 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16485), .A(n16470), .B(
        n16805), .ZN(n16475) );
  AOI211_X1 U19752 ( .C1(n16473), .C2(n16472), .A(n16471), .B(n16757), .ZN(
        n16474) );
  AOI211_X1 U19753 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16476), .A(n16475), 
        .B(n16474), .ZN(n16477) );
  OAI211_X1 U19754 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16479), .A(n16478), 
        .B(n16477), .ZN(P3_U2643) );
  AOI22_X1 U19755 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16784), .B1(
        n16807), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16490) );
  AOI211_X1 U19756 ( .C1(n16482), .C2(n16481), .A(n16480), .B(n16757), .ZN(
        n16483) );
  AOI21_X1 U19757 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16484), .A(n16483), 
        .ZN(n16489) );
  OAI211_X1 U19758 ( .C1(n16492), .C2(n16486), .A(n16806), .B(n16485), .ZN(
        n16487) );
  NAND4_X1 U19759 ( .A1(n16490), .A2(n16489), .A3(n16488), .A4(n16487), .ZN(
        P3_U2644) );
  AOI21_X1 U19760 ( .B1(n16778), .B2(n16491), .A(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n16499) );
  AOI22_X1 U19761 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16784), .B1(
        n16807), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16498) );
  AOI211_X1 U19762 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16507), .A(n16492), .B(
        n16805), .ZN(n16496) );
  AOI211_X1 U19763 ( .C1(n17403), .C2(n16494), .A(n16493), .B(n16757), .ZN(
        n16495) );
  NOR2_X1 U19764 ( .A1(n16496), .A2(n16495), .ZN(n16497) );
  OAI211_X1 U19765 ( .C1(n16500), .C2(n16499), .A(n16498), .B(n16497), .ZN(
        P3_U2645) );
  INV_X1 U19766 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18655) );
  OAI21_X1 U19767 ( .B1(n16523), .B2(n16799), .A(n16809), .ZN(n16520) );
  AOI21_X1 U19768 ( .B1(n16778), .B2(n18655), .A(n16520), .ZN(n16511) );
  AOI211_X1 U19769 ( .C1(n16502), .C2(n9925), .A(n16501), .B(n16757), .ZN(
        n16506) );
  NAND2_X1 U19770 ( .A1(n16778), .A2(n18658), .ZN(n16503) );
  OAI22_X1 U19771 ( .A1(n17422), .A2(n16793), .B1(n16504), .B2(n16503), .ZN(
        n16505) );
  AOI211_X1 U19772 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n16807), .A(n16506), .B(
        n16505), .ZN(n16510) );
  OAI211_X1 U19773 ( .C1(n16513), .C2(n16508), .A(n16806), .B(n16507), .ZN(
        n16509) );
  OAI211_X1 U19774 ( .C1(n16511), .C2(n18658), .A(n16510), .B(n16509), .ZN(
        P3_U2646) );
  NOR2_X1 U19775 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16799), .ZN(n16512) );
  AOI22_X1 U19776 ( .A1(n16807), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16523), 
        .B2(n16512), .ZN(n16519) );
  AOI211_X1 U19777 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16528), .A(n16513), .B(
        n16805), .ZN(n16517) );
  AOI211_X1 U19778 ( .C1(n17439), .C2(n16515), .A(n16514), .B(n16757), .ZN(
        n16516) );
  AOI211_X1 U19779 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16520), .A(n16517), 
        .B(n16516), .ZN(n16518) );
  OAI211_X1 U19780 ( .C1(n17432), .C2(n16793), .A(n16519), .B(n16518), .ZN(
        P3_U2647) );
  INV_X1 U19781 ( .A(n16520), .ZN(n16532) );
  AOI211_X1 U19782 ( .C1(n17441), .C2(n16522), .A(n16521), .B(n16757), .ZN(
        n16527) );
  OR2_X1 U19783 ( .A1(n16799), .A2(n16523), .ZN(n16524) );
  OAI22_X1 U19784 ( .A1(n9952), .A2(n16793), .B1(n16525), .B2(n16524), .ZN(
        n16526) );
  AOI211_X1 U19785 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16807), .A(n16527), .B(
        n16526), .ZN(n16531) );
  OAI211_X1 U19786 ( .C1(n16536), .C2(n16529), .A(n16806), .B(n16528), .ZN(
        n16530) );
  OAI211_X1 U19787 ( .C1(n16532), .C2(n18654), .A(n16531), .B(n16530), .ZN(
        P3_U2648) );
  NOR2_X1 U19788 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16799), .ZN(n16533) );
  AOI22_X1 U19789 ( .A1(n16807), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n16534), 
        .B2(n16533), .ZN(n16544) );
  INV_X1 U19790 ( .A(n16535), .ZN(n16549) );
  OAI221_X1 U19791 ( .B1(n16799), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16799), 
        .C2(n16549), .A(n16809), .ZN(n16542) );
  AOI211_X1 U19792 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16550), .A(n16536), .B(
        n16805), .ZN(n16541) );
  AOI211_X1 U19793 ( .C1(n16539), .C2(n16538), .A(n16537), .B(n16757), .ZN(
        n16540) );
  AOI211_X1 U19794 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16542), .A(n16541), 
        .B(n16540), .ZN(n16543) );
  OAI211_X1 U19795 ( .C1(n17462), .C2(n16793), .A(n16544), .B(n16543), .ZN(
        P3_U2649) );
  AOI22_X1 U19796 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16784), .B1(
        n16807), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16554) );
  OAI21_X1 U19797 ( .B1(n16549), .B2(n16799), .A(n16809), .ZN(n16561) );
  AOI211_X1 U19798 ( .C1(n16547), .C2(n16546), .A(n16545), .B(n16757), .ZN(
        n16548) );
  AOI21_X1 U19799 ( .B1(n16561), .B2(P3_REIP_REG_21__SCAN_IN), .A(n16548), 
        .ZN(n16553) );
  NAND3_X1 U19800 ( .A1(n16778), .A2(n16549), .A3(n18650), .ZN(n16552) );
  OAI211_X1 U19801 ( .C1(n16555), .C2(n20809), .A(n16806), .B(n16550), .ZN(
        n16551) );
  NAND4_X1 U19802 ( .A1(n16554), .A2(n16553), .A3(n16552), .A4(n16551), .ZN(
        P3_U2650) );
  AOI211_X1 U19803 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16565), .A(n16555), .B(
        n16805), .ZN(n16556) );
  AOI21_X1 U19804 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16807), .A(n16556), .ZN(
        n16563) );
  INV_X1 U19805 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18645) );
  INV_X1 U19806 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18643) );
  NOR3_X1 U19807 ( .A1(n16799), .A2(n18637), .A3(n16602), .ZN(n16609) );
  NAND2_X1 U19808 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n16609), .ZN(n16598) );
  NOR2_X1 U19809 ( .A1(n18641), .A2(n16598), .ZN(n16572) );
  INV_X1 U19810 ( .A(n16572), .ZN(n16588) );
  NOR3_X1 U19811 ( .A1(n18645), .A2(n18643), .A3(n16588), .ZN(n16560) );
  INV_X1 U19812 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18647) );
  AOI211_X1 U19813 ( .C1(n17489), .C2(n16558), .A(n16557), .B(n16757), .ZN(
        n16559) );
  AOI221_X1 U19814 ( .B1(n16561), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n16560), 
        .C2(n18647), .A(n16559), .ZN(n16562) );
  OAI211_X1 U19815 ( .C1(n17486), .C2(n16793), .A(n16563), .B(n16562), .ZN(
        P3_U2651) );
  INV_X1 U19816 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17511) );
  NOR2_X1 U19817 ( .A1(n17511), .A2(n16578), .ZN(n16564) );
  OAI21_X1 U19818 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16564), .A(
        n17460), .ZN(n17496) );
  NOR2_X1 U19819 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17741), .ZN(
        n16786) );
  NAND2_X1 U19820 ( .A1(n17495), .A2(n16786), .ZN(n16579) );
  OAI21_X1 U19821 ( .B1(n17511), .B2(n16579), .A(n16764), .ZN(n16582) );
  XNOR2_X1 U19822 ( .A(n17496), .B(n16582), .ZN(n16575) );
  INV_X1 U19823 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17494) );
  OAI211_X1 U19824 ( .C1(n16577), .C2(n16566), .A(n16806), .B(n16565), .ZN(
        n16567) );
  OAI211_X1 U19825 ( .C1(n17494), .C2(n16793), .A(n9637), .B(n16567), .ZN(
        n16568) );
  AOI21_X1 U19826 ( .B1(n16569), .B2(P3_EBX_REG_19__SCAN_IN), .A(n16568), .ZN(
        n16574) );
  OAI21_X1 U19827 ( .B1(n16570), .B2(n16799), .A(n16809), .ZN(n16576) );
  XOR2_X1 U19828 ( .A(n18645), .B(n18643), .Z(n16571) );
  AOI22_X1 U19829 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16576), .B1(n16572), 
        .B2(n16571), .ZN(n16573) );
  OAI211_X1 U19830 ( .C1(n16757), .C2(n16575), .A(n16574), .B(n16573), .ZN(
        P3_U2652) );
  INV_X1 U19831 ( .A(n16576), .ZN(n16599) );
  AOI211_X1 U19832 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16592), .A(n16577), .B(
        n16805), .ZN(n16586) );
  AOI22_X1 U19833 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16578), .B1(
        n17493), .B2(n17511), .ZN(n17508) );
  NOR2_X1 U19834 ( .A1(n16757), .A2(n16764), .ZN(n16797) );
  INV_X1 U19835 ( .A(n16797), .ZN(n16789) );
  INV_X1 U19836 ( .A(n16579), .ZN(n16580) );
  OAI21_X1 U19837 ( .B1(n16580), .B2(n17508), .A(n18585), .ZN(n16581) );
  AOI22_X1 U19838 ( .A1(n17508), .A2(n16582), .B1(n16789), .B2(n16581), .ZN(
        n16585) );
  OAI22_X1 U19839 ( .A1(n17511), .A2(n16793), .B1(n16798), .B2(n16583), .ZN(
        n16584) );
  NOR4_X1 U19840 ( .A1(n18032), .A2(n16586), .A3(n16585), .A4(n16584), .ZN(
        n16587) );
  OAI221_X1 U19841 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16588), .C1(n18643), 
        .C2(n16599), .A(n16587), .ZN(P3_U2653) );
  INV_X1 U19842 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17521) );
  NAND2_X1 U19843 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16604), .ZN(
        n16589) );
  AOI21_X1 U19844 ( .B1(n17521), .B2(n16589), .A(n17493), .ZN(n17524) );
  INV_X1 U19845 ( .A(n17535), .ZN(n17531) );
  NOR2_X1 U19846 ( .A1(n17741), .A2(n17531), .ZN(n17534) );
  NAND2_X1 U19847 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17534), .ZN(
        n16612) );
  OAI21_X1 U19848 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16612), .A(
        n16764), .ZN(n16605) );
  OAI21_X1 U19849 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16734), .A(
        n16605), .ZN(n16591) );
  AOI21_X1 U19850 ( .B1(n17524), .B2(n16591), .A(n16757), .ZN(n16590) );
  OAI21_X1 U19851 ( .B1(n17524), .B2(n16591), .A(n16590), .ZN(n16595) );
  OAI211_X1 U19852 ( .C1(n16600), .C2(n16593), .A(n16806), .B(n16592), .ZN(
        n16594) );
  OAI211_X1 U19853 ( .C1(n16793), .C2(n17521), .A(n16595), .B(n16594), .ZN(
        n16596) );
  AOI211_X1 U19854 ( .C1(n16807), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18017), .B(
        n16596), .ZN(n16597) );
  OAI221_X1 U19855 ( .B1(n16599), .B2(n18641), .C1(n16599), .C2(n16598), .A(
        n16597), .ZN(P3_U2654) );
  INV_X1 U19856 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17536) );
  AOI211_X1 U19857 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16619), .A(n16600), .B(
        n16805), .ZN(n16601) );
  AOI211_X1 U19858 ( .C1(n16807), .C2(P3_EBX_REG_16__SCAN_IN), .A(n18017), .B(
        n16601), .ZN(n16611) );
  AOI21_X1 U19859 ( .B1(n16778), .B2(n16602), .A(n16792), .ZN(n16625) );
  NOR2_X1 U19860 ( .A1(n16799), .A2(n16602), .ZN(n16603) );
  NAND2_X1 U19861 ( .A1(n16603), .A2(n18637), .ZN(n16615) );
  NAND2_X1 U19862 ( .A1(n16625), .A2(n16615), .ZN(n16608) );
  AOI22_X1 U19863 ( .A1(n17536), .A2(n16612), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16604), .ZN(n16606) );
  INV_X1 U19864 ( .A(n16605), .ZN(n16613) );
  INV_X1 U19865 ( .A(n16606), .ZN(n17538) );
  AOI221_X1 U19866 ( .B1(n16606), .B2(n16613), .C1(n17538), .C2(n16605), .A(
        n16757), .ZN(n16607) );
  AOI221_X1 U19867 ( .B1(n16609), .B2(n18639), .C1(n16608), .C2(
        P3_REIP_REG_16__SCAN_IN), .A(n16607), .ZN(n16610) );
  OAI211_X1 U19868 ( .C1(n17536), .C2(n16793), .A(n16611), .B(n16610), .ZN(
        P3_U2655) );
  NOR2_X1 U19869 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16757), .ZN(
        n16796) );
  INV_X1 U19870 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17537) );
  AOI21_X1 U19871 ( .B1(n16796), .B2(n17537), .A(n16797), .ZN(n16623) );
  OAI21_X1 U19872 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17534), .A(
        n16612), .ZN(n17551) );
  INV_X1 U19873 ( .A(n16625), .ZN(n16618) );
  AOI22_X1 U19874 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16784), .B1(
        n16807), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n16616) );
  NAND3_X1 U19875 ( .A1(n18585), .A2(n16613), .A3(n17551), .ZN(n16614) );
  NAND4_X1 U19876 ( .A1(n16616), .A2(n9637), .A3(n16615), .A4(n16614), .ZN(
        n16617) );
  AOI21_X1 U19877 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16618), .A(n16617), 
        .ZN(n16622) );
  OAI211_X1 U19878 ( .C1(n16626), .C2(n16620), .A(n16806), .B(n16619), .ZN(
        n16621) );
  OAI211_X1 U19879 ( .C1(n16623), .C2(n17551), .A(n16622), .B(n16621), .ZN(
        P3_U2656) );
  OR2_X1 U19880 ( .A1(n17741), .A2(n17564), .ZN(n16632) );
  AOI21_X1 U19881 ( .B1(n17563), .B2(n16632), .A(n17534), .ZN(n17566) );
  INV_X1 U19882 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17590) );
  INV_X1 U19883 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16635) );
  NOR2_X1 U19884 ( .A1(n17590), .A2(n16635), .ZN(n17579) );
  INV_X1 U19885 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17617) );
  INV_X1 U19886 ( .A(n17643), .ZN(n17603) );
  INV_X1 U19887 ( .A(n16698), .ZN(n17642) );
  NAND2_X1 U19888 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17642), .ZN(
        n16711) );
  INV_X1 U19889 ( .A(n16711), .ZN(n16721) );
  NAND2_X1 U19890 ( .A1(n17603), .A2(n16721), .ZN(n16697) );
  INV_X1 U19891 ( .A(n16697), .ZN(n16686) );
  NAND2_X1 U19892 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16686), .ZN(
        n16685) );
  NOR2_X1 U19893 ( .A1(n17617), .A2(n16685), .ZN(n16678) );
  AND3_X1 U19894 ( .A1(n16795), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16678), .ZN(n16652) );
  AOI21_X1 U19895 ( .B1(n17579), .B2(n16652), .A(n16734), .ZN(n16633) );
  XNOR2_X1 U19896 ( .A(n17566), .B(n16633), .ZN(n16631) );
  AOI21_X1 U19897 ( .B1(n16807), .B2(P3_EBX_REG_14__SCAN_IN), .A(n18032), .ZN(
        n16630) );
  INV_X1 U19898 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18633) );
  INV_X1 U19899 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18635) );
  NAND2_X1 U19900 ( .A1(n16778), .A2(n16624), .ZN(n16639) );
  AOI221_X1 U19901 ( .B1(n18633), .B2(n18635), .C1(n16639), .C2(n18635), .A(
        n16625), .ZN(n16628) );
  AOI211_X1 U19902 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16636), .A(n16626), .B(
        n16805), .ZN(n16627) );
  AOI211_X1 U19903 ( .C1(n16784), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16628), .B(n16627), .ZN(n16629) );
  OAI211_X1 U19904 ( .C1(n16757), .C2(n16631), .A(n16630), .B(n16629), .ZN(
        P3_U2657) );
  NAND2_X1 U19905 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16678), .ZN(
        n17573) );
  NOR2_X1 U19906 ( .A1(n17590), .A2(n17573), .ZN(n16651) );
  AOI21_X1 U19907 ( .B1(n16651), .B2(n16796), .A(n16797), .ZN(n16645) );
  OAI21_X1 U19908 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16651), .A(
        n16632), .ZN(n17577) );
  NAND3_X1 U19909 ( .A1(n18585), .A2(n16633), .A3(n17577), .ZN(n16634) );
  OAI211_X1 U19910 ( .C1(n16635), .C2(n16793), .A(n9637), .B(n16634), .ZN(
        n16641) );
  OAI211_X1 U19911 ( .C1(n16647), .C2(n16637), .A(n16806), .B(n16636), .ZN(
        n16638) );
  OAI21_X1 U19912 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n16639), .A(n16638), 
        .ZN(n16640) );
  AOI211_X1 U19913 ( .C1(n16807), .C2(P3_EBX_REG_13__SCAN_IN), .A(n16641), .B(
        n16640), .ZN(n16644) );
  OAI221_X1 U19914 ( .B1(n16799), .B2(n16675), .C1(n16799), .C2(n16642), .A(
        n16809), .ZN(n16669) );
  NOR2_X1 U19915 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16799), .ZN(n16649) );
  OAI21_X1 U19916 ( .B1(n16669), .B2(n16649), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n16643) );
  OAI211_X1 U19917 ( .C1(n16645), .C2(n17577), .A(n16644), .B(n16643), .ZN(
        P3_U2658) );
  AOI22_X1 U19918 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16784), .B1(
        n16807), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16657) );
  INV_X1 U19919 ( .A(n16646), .ZN(n16650) );
  AOI211_X1 U19920 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16663), .A(n16647), .B(
        n16805), .ZN(n16648) );
  AOI211_X1 U19921 ( .C1(n16650), .C2(n16649), .A(n18017), .B(n16648), .ZN(
        n16656) );
  AOI21_X1 U19922 ( .B1(n17590), .B2(n17573), .A(n16651), .ZN(n17596) );
  NOR2_X1 U19923 ( .A1(n16652), .A2(n16734), .ZN(n16653) );
  XOR2_X1 U19924 ( .A(n17596), .B(n16653), .Z(n16654) );
  AOI22_X1 U19925 ( .A1(n18585), .A2(n16654), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16669), .ZN(n16655) );
  NAND3_X1 U19926 ( .A1(n16657), .A2(n16656), .A3(n16655), .ZN(P3_U2659) );
  NOR2_X1 U19927 ( .A1(n16799), .A2(n16658), .ZN(n16736) );
  NAND2_X1 U19928 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16736), .ZN(n16701) );
  OAI21_X1 U19929 ( .B1(n16659), .B2(n16701), .A(n18629), .ZN(n16668) );
  INV_X1 U19930 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16666) );
  OAI21_X1 U19931 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16678), .A(
        n17573), .ZN(n16660) );
  INV_X1 U19932 ( .A(n16660), .ZN(n17608) );
  AOI21_X1 U19933 ( .B1(n16678), .B2(n16795), .A(n16734), .ZN(n16662) );
  AOI21_X1 U19934 ( .B1(n17608), .B2(n16662), .A(n16757), .ZN(n16661) );
  OAI21_X1 U19935 ( .B1(n17608), .B2(n16662), .A(n16661), .ZN(n16665) );
  OAI211_X1 U19936 ( .C1(n16672), .C2(n16671), .A(n16806), .B(n16663), .ZN(
        n16664) );
  OAI211_X1 U19937 ( .C1(n16793), .C2(n16666), .A(n16665), .B(n16664), .ZN(
        n16667) );
  AOI21_X1 U19938 ( .B1(n16669), .B2(n16668), .A(n16667), .ZN(n16670) );
  OAI211_X1 U19939 ( .C1(n16798), .C2(n16671), .A(n16670), .B(n9637), .ZN(
        P3_U2660) );
  AOI211_X1 U19940 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16673), .A(n16672), .B(
        n16805), .ZN(n16674) );
  AOI211_X1 U19941 ( .C1(n16807), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18017), .B(
        n16674), .ZN(n16684) );
  NOR2_X1 U19942 ( .A1(n16792), .A2(n16778), .ZN(n16677) );
  INV_X1 U19943 ( .A(n16677), .ZN(n16808) );
  NAND2_X1 U19944 ( .A1(n16675), .A2(n16809), .ZN(n16676) );
  NAND2_X1 U19945 ( .A1(n16808), .A2(n16676), .ZN(n16726) );
  OAI21_X1 U19946 ( .B1(n16680), .B2(n16677), .A(n16726), .ZN(n16702) );
  AOI21_X1 U19947 ( .B1(n17617), .B2(n16685), .A(n16678), .ZN(n17621) );
  NAND2_X1 U19948 ( .A1(n16721), .A2(n16795), .ZN(n16724) );
  NOR2_X1 U19949 ( .A1(n17643), .A2(n16724), .ZN(n16688) );
  AOI21_X1 U19950 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16688), .A(
        n16734), .ZN(n16687) );
  OAI21_X1 U19951 ( .B1(n17621), .B2(n16687), .A(n18585), .ZN(n16679) );
  AOI21_X1 U19952 ( .B1(n17621), .B2(n16687), .A(n16679), .ZN(n16682) );
  INV_X1 U19953 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18627) );
  INV_X1 U19954 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18625) );
  NAND2_X1 U19955 ( .A1(n16680), .A2(n16730), .ZN(n16696) );
  AOI221_X1 U19956 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n18627), .C2(n18625), .A(n16696), .ZN(n16681) );
  AOI211_X1 U19957 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16702), .A(n16682), 
        .B(n16681), .ZN(n16683) );
  OAI211_X1 U19958 ( .C1(n17617), .C2(n16793), .A(n16684), .B(n16683), .ZN(
        P3_U2661) );
  INV_X1 U19959 ( .A(n16702), .ZN(n16695) );
  OR2_X1 U19960 ( .A1(n16805), .A2(n16690), .ZN(n16700) );
  OAI21_X1 U19961 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16686), .A(
        n16685), .ZN(n17633) );
  OAI211_X1 U19962 ( .C1(n16688), .C2(n17633), .A(n18585), .B(n16687), .ZN(
        n16689) );
  OAI211_X1 U19963 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16700), .A(n9637), .B(
        n16689), .ZN(n16693) );
  AOI21_X1 U19964 ( .B1(n16806), .B2(n16690), .A(n16807), .ZN(n16691) );
  OAI22_X1 U19965 ( .A1(n17036), .A2(n16691), .B1(n17633), .B2(n16789), .ZN(
        n16692) );
  AOI211_X1 U19966 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n16784), .A(
        n16693), .B(n16692), .ZN(n16694) );
  OAI221_X1 U19967 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16696), .C1(n18625), 
        .C2(n16695), .A(n16694), .ZN(P3_U2662) );
  INV_X1 U19968 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17660) );
  NOR2_X1 U19969 ( .A1(n17660), .A2(n16711), .ZN(n16710) );
  OAI21_X1 U19970 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16710), .A(
        n16697), .ZN(n17646) );
  NOR2_X1 U19971 ( .A1(n16698), .A2(n17660), .ZN(n17644) );
  AOI21_X1 U19972 ( .B1(n17644), .B2(n16786), .A(n16734), .ZN(n16713) );
  XNOR2_X1 U19973 ( .A(n17646), .B(n16713), .ZN(n16699) );
  AOI21_X1 U19974 ( .B1(n16699), .B2(n18585), .A(n18032), .ZN(n16707) );
  AOI21_X1 U19975 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16708), .A(n16700), .ZN(
        n16705) );
  NOR2_X1 U19976 ( .A1(n16718), .A2(n16701), .ZN(n16703) );
  MUX2_X1 U19977 ( .A(n16703), .B(n16702), .S(P3_REIP_REG_8__SCAN_IN), .Z(
        n16704) );
  AOI211_X1 U19978 ( .C1(n16784), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16705), .B(n16704), .ZN(n16706) );
  OAI211_X1 U19979 ( .C1(n16798), .C2(n17056), .A(n16707), .B(n16706), .ZN(
        P3_U2663) );
  INV_X1 U19980 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18621) );
  OAI211_X1 U19981 ( .C1(n16715), .C2(n16722), .A(n16708), .B(n16806), .ZN(
        n16709) );
  INV_X1 U19982 ( .A(n16709), .ZN(n16717) );
  AOI21_X1 U19983 ( .B1(n17660), .B2(n16711), .A(n16710), .ZN(n17665) );
  AOI21_X1 U19984 ( .B1(n17665), .B2(n16724), .A(n16757), .ZN(n16712) );
  OAI22_X1 U19985 ( .A1(n17665), .A2(n16713), .B1(n16797), .B2(n16712), .ZN(
        n16714) );
  OAI211_X1 U19986 ( .C1(n16798), .C2(n16715), .A(n9637), .B(n16714), .ZN(
        n16716) );
  AOI211_X1 U19987 ( .C1(n16784), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16717), .B(n16716), .ZN(n16720) );
  OAI211_X1 U19988 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16730), .B(n16718), .ZN(n16719) );
  OAI211_X1 U19989 ( .C1(n16726), .C2(n18621), .A(n16720), .B(n16719), .ZN(
        P3_U2664) );
  INV_X1 U19990 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17675) );
  NOR2_X1 U19991 ( .A1(n17741), .A2(n17680), .ZN(n16746) );
  NAND2_X1 U19992 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16746), .ZN(
        n16733) );
  AOI21_X1 U19993 ( .B1(n17675), .B2(n16733), .A(n16721), .ZN(n17678) );
  NOR2_X1 U19994 ( .A1(n17678), .A2(n16794), .ZN(n16725) );
  AOI211_X1 U19995 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16737), .A(n16722), .B(
        n16805), .ZN(n16723) );
  AOI211_X1 U19996 ( .C1(n16725), .C2(n16724), .A(n18032), .B(n16723), .ZN(
        n16732) );
  INV_X1 U19997 ( .A(n16726), .ZN(n16735) );
  INV_X1 U19998 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18619) );
  AOI21_X1 U19999 ( .B1(n16796), .B2(n17675), .A(n16797), .ZN(n16728) );
  INV_X1 U20000 ( .A(n17678), .ZN(n16727) );
  OAI22_X1 U20001 ( .A1(n16728), .A2(n16727), .B1(n17675), .B2(n16793), .ZN(
        n16729) );
  AOI221_X1 U20002 ( .B1(n16735), .B2(P3_REIP_REG_6__SCAN_IN), .C1(n16730), 
        .C2(n18619), .A(n16729), .ZN(n16731) );
  OAI211_X1 U20003 ( .C1(n16798), .C2(n17079), .A(n16732), .B(n16731), .ZN(
        P3_U2665) );
  OAI21_X1 U20004 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16746), .A(
        n16733), .ZN(n17689) );
  AOI21_X1 U20005 ( .B1(n16746), .B2(n16795), .A(n16734), .ZN(n16748) );
  XOR2_X1 U20006 ( .A(n17689), .B(n16748), .Z(n16744) );
  OAI21_X1 U20007 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n16736), .A(n16735), .ZN(
        n16740) );
  OAI211_X1 U20008 ( .C1(n16751), .C2(n16738), .A(n16806), .B(n16737), .ZN(
        n16739) );
  OAI211_X1 U20009 ( .C1(n16793), .C2(n16741), .A(n16740), .B(n16739), .ZN(
        n16742) );
  AOI211_X1 U20010 ( .C1(n16807), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18032), .B(
        n16742), .ZN(n16743) );
  OAI21_X1 U20011 ( .B1(n16757), .B2(n16744), .A(n16743), .ZN(P3_U2666) );
  NOR2_X1 U20012 ( .A1(n16745), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17694) );
  NOR2_X1 U20013 ( .A1(n17741), .A2(n16745), .ZN(n16763) );
  INV_X1 U20014 ( .A(n16746), .ZN(n16747) );
  OAI21_X1 U20015 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16763), .A(
        n16747), .ZN(n17703) );
  AOI22_X1 U20016 ( .A1(n16786), .A2(n17694), .B1(n16748), .B2(n17703), .ZN(
        n16758) );
  INV_X1 U20017 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18615) );
  AND3_X1 U20018 ( .A1(n18615), .A2(n16778), .A3(n16759), .ZN(n16750) );
  OAI22_X1 U20019 ( .A1(n16798), .A2(n17078), .B1(n17703), .B2(n16789), .ZN(
        n16749) );
  AOI211_X1 U20020 ( .C1(n16784), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16750), .B(n16749), .ZN(n16756) );
  OAI21_X1 U20021 ( .B1(n16759), .B2(n16799), .A(n16809), .ZN(n16766) );
  AOI211_X1 U20022 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16768), .A(n16751), .B(
        n16805), .ZN(n16754) );
  NAND2_X1 U20023 ( .A1(n16752), .A2(n18746), .ZN(n16760) );
  OAI221_X1 U20024 ( .B1(n16760), .B2(n15558), .C1(n16760), .C2(n18572), .A(
        n9637), .ZN(n16753) );
  AOI211_X1 U20025 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16766), .A(n16754), .B(
        n16753), .ZN(n16755) );
  OAI211_X1 U20026 ( .C1(n16758), .C2(n16757), .A(n16756), .B(n16755), .ZN(
        P3_U2667) );
  AOI22_X1 U20027 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16784), .B1(
        n16807), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16773) );
  NOR2_X1 U20028 ( .A1(n16759), .A2(n16799), .ZN(n16761) );
  AOI21_X1 U20029 ( .B1(n18685), .B2(n18556), .A(n15509), .ZN(n18680) );
  AOI22_X1 U20030 ( .A1(n16762), .A2(n16761), .B1(n18747), .B2(n18680), .ZN(
        n16772) );
  INV_X1 U20031 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17715) );
  NAND2_X1 U20032 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16774) );
  AOI21_X1 U20033 ( .B1(n17715), .B2(n16774), .A(n16763), .ZN(n17717) );
  OAI21_X1 U20034 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16774), .A(
        n16764), .ZN(n16765) );
  INV_X1 U20035 ( .A(n16765), .ZN(n16785) );
  XOR2_X1 U20036 ( .A(n17717), .B(n16785), .Z(n16767) );
  AOI22_X1 U20037 ( .A1(n18585), .A2(n16767), .B1(P3_REIP_REG_3__SCAN_IN), 
        .B2(n16766), .ZN(n16771) );
  OAI211_X1 U20038 ( .C1(n16775), .C2(n16769), .A(n16806), .B(n16768), .ZN(
        n16770) );
  NAND4_X1 U20039 ( .A1(n16773), .A2(n16772), .A3(n16771), .A4(n16770), .ZN(
        P3_U2668) );
  OAI21_X1 U20040 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16774), .ZN(n17728) );
  NAND2_X1 U20041 ( .A1(n17108), .A2(n17103), .ZN(n16776) );
  AOI211_X1 U20042 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16776), .A(n16775), .B(
        n16805), .ZN(n16783) );
  INV_X1 U20043 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16781) );
  NAND2_X1 U20044 ( .A1(n18695), .A2(n18523), .ZN(n18551) );
  NAND2_X1 U20045 ( .A1(n18556), .A2(n18551), .ZN(n18528) );
  INV_X1 U20046 ( .A(n18528), .ZN(n18691) );
  AOI22_X1 U20047 ( .A1(n16792), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18691), 
        .B2(n18747), .ZN(n16780) );
  OAI211_X1 U20048 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16778), .B(n16777), .ZN(n16779) );
  OAI211_X1 U20049 ( .C1(n16781), .C2(n16798), .A(n16780), .B(n16779), .ZN(
        n16782) );
  AOI211_X1 U20050 ( .C1(n16784), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16783), .B(n16782), .ZN(n16788) );
  OAI211_X1 U20051 ( .C1(n16786), .C2(n17728), .A(n18585), .B(n16785), .ZN(
        n16787) );
  OAI211_X1 U20052 ( .C1(n16789), .C2(n17728), .A(n16788), .B(n16787), .ZN(
        P3_U2669) );
  INV_X1 U20053 ( .A(n17097), .ZN(n16790) );
  OAI21_X1 U20054 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n16790), .ZN(n17104) );
  AND2_X1 U20055 ( .A1(n18523), .A2(n16791), .ZN(n18699) );
  AOI22_X1 U20056 ( .A1(n16792), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18699), 
        .B2(n18747), .ZN(n16804) );
  OAI21_X1 U20057 ( .B1(n16795), .B2(n16794), .A(n16793), .ZN(n16802) );
  OR2_X1 U20058 ( .A1(n16797), .A2(n16796), .ZN(n16801) );
  OAI22_X1 U20059 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16799), .B1(n16798), 
        .B2(n17103), .ZN(n16800) );
  AOI221_X1 U20060 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16802), .C1(
        n17741), .C2(n16801), .A(n16800), .ZN(n16803) );
  OAI211_X1 U20061 ( .C1(n16805), .C2(n17104), .A(n16804), .B(n16803), .ZN(
        P3_U2670) );
  NOR2_X1 U20062 ( .A1(n16807), .A2(n16806), .ZN(n16812) );
  AOI22_X1 U20063 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16808), .B1(n18747), 
        .B2(n18708), .ZN(n16811) );
  NAND3_X1 U20064 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18683), .A3(
        n16809), .ZN(n16810) );
  OAI211_X1 U20065 ( .C1(n16812), .C2(n17108), .A(n16811), .B(n16810), .ZN(
        P3_U2671) );
  NAND4_X1 U20066 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(P3_EBX_REG_25__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n16813)
         );
  NOR2_X1 U20067 ( .A1(n16900), .A2(n16813), .ZN(n16814) );
  NAND4_X1 U20068 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n16848), .A4(n16814), .ZN(n16817) );
  NOR2_X1 U20069 ( .A1(n16818), .A2(n16817), .ZN(n16843) );
  NAND2_X1 U20070 ( .A1(n17101), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16816) );
  NAND2_X1 U20071 ( .A1(n16843), .A2(n17197), .ZN(n16815) );
  OAI22_X1 U20072 ( .A1(n16843), .A2(n16816), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16815), .ZN(P3_U2672) );
  NAND2_X1 U20073 ( .A1(n16818), .A2(n16817), .ZN(n16819) );
  NAND2_X1 U20074 ( .A1(n16819), .A2(n17101), .ZN(n16842) );
  AOI22_X1 U20075 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16823) );
  AOI22_X1 U20076 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16822) );
  AOI22_X1 U20077 ( .A1(n13937), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16821) );
  AOI22_X1 U20078 ( .A1(n15509), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16820) );
  NAND4_X1 U20079 ( .A1(n16823), .A2(n16822), .A3(n16821), .A4(n16820), .ZN(
        n16829) );
  AOI22_X1 U20080 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16827) );
  AOI22_X1 U20081 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16826) );
  AOI22_X1 U20082 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16976), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16825) );
  AOI22_X1 U20083 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16824) );
  NAND4_X1 U20084 ( .A1(n16827), .A2(n16826), .A3(n16825), .A4(n16824), .ZN(
        n16828) );
  NOR2_X1 U20085 ( .A1(n16829), .A2(n16828), .ZN(n16841) );
  AOI22_X1 U20086 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16840) );
  AOI22_X1 U20087 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16831) );
  AOI22_X1 U20088 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16830) );
  OAI211_X1 U20089 ( .C1(n16832), .C2(n17084), .A(n16831), .B(n16830), .ZN(
        n16838) );
  AOI22_X1 U20090 ( .A1(n13937), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16836) );
  AOI22_X1 U20091 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16835) );
  AOI22_X1 U20092 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U20093 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16833) );
  NAND4_X1 U20094 ( .A1(n16836), .A2(n16835), .A3(n16834), .A4(n16833), .ZN(
        n16837) );
  AOI211_X1 U20095 ( .C1(n17046), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n16838), .B(n16837), .ZN(n16839) );
  NAND2_X1 U20096 ( .A1(n16840), .A2(n16839), .ZN(n16845) );
  NAND2_X1 U20097 ( .A1(n16846), .A2(n16845), .ZN(n16844) );
  XNOR2_X1 U20098 ( .A(n16841), .B(n16844), .ZN(n17123) );
  OAI22_X1 U20099 ( .A1(n16843), .A2(n16842), .B1(n17123), .B2(n17101), .ZN(
        P3_U2673) );
  OAI21_X1 U20100 ( .B1(n16846), .B2(n16845), .A(n16844), .ZN(n17127) );
  NOR2_X1 U20101 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16858), .ZN(n16847) );
  AOI22_X1 U20102 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16849), .B1(n16848), 
        .B2(n16847), .ZN(n16850) );
  OAI21_X1 U20103 ( .B1(n17127), .B2(n17101), .A(n16850), .ZN(P3_U2674) );
  OAI21_X1 U20104 ( .B1(n16855), .B2(n16852), .A(n16851), .ZN(n17136) );
  NAND3_X1 U20105 ( .A1(n16858), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17101), 
        .ZN(n16853) );
  OAI221_X1 U20106 ( .B1(n16858), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17101), 
        .C2(n17136), .A(n16853), .ZN(P3_U2676) );
  AOI21_X1 U20107 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17101), .A(n16864), .ZN(
        n16854) );
  INV_X1 U20108 ( .A(n16854), .ZN(n16857) );
  AOI21_X1 U20109 ( .B1(n16856), .B2(n16861), .A(n16855), .ZN(n17137) );
  AOI22_X1 U20110 ( .A1(n16858), .A2(n16857), .B1(n17105), .B2(n17137), .ZN(
        n16859) );
  INV_X1 U20111 ( .A(n16859), .ZN(P3_U2677) );
  INV_X1 U20112 ( .A(n16860), .ZN(n16869) );
  AOI21_X1 U20113 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17101), .A(n16869), .ZN(
        n16863) );
  OAI21_X1 U20114 ( .B1(n16865), .B2(n16862), .A(n16861), .ZN(n17147) );
  OAI22_X1 U20115 ( .A1(n16864), .A2(n16863), .B1(n17101), .B2(n17147), .ZN(
        P3_U2678) );
  AOI21_X1 U20116 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17101), .A(n16875), .ZN(
        n16868) );
  AOI21_X1 U20117 ( .B1(n16866), .B2(n16871), .A(n16865), .ZN(n17148) );
  INV_X1 U20118 ( .A(n17148), .ZN(n16867) );
  OAI22_X1 U20119 ( .A1(n16869), .A2(n16868), .B1(n17101), .B2(n16867), .ZN(
        P3_U2679) );
  INV_X1 U20120 ( .A(n16870), .ZN(n16889) );
  AOI21_X1 U20121 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17101), .A(n16889), .ZN(
        n16874) );
  OAI21_X1 U20122 ( .B1(n16873), .B2(n16872), .A(n16871), .ZN(n17157) );
  OAI22_X1 U20123 ( .A1(n16875), .A2(n16874), .B1(n17101), .B2(n17157), .ZN(
        P3_U2680) );
  AOI21_X1 U20124 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17101), .A(n16876), .ZN(
        n16888) );
  AOI22_X1 U20125 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16886) );
  AOI22_X1 U20126 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16885) );
  AOI22_X1 U20127 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16884) );
  NOR2_X1 U20128 ( .A1(n16903), .A2(n17084), .ZN(n16882) );
  AOI22_X1 U20129 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20130 ( .A1(n13884), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20131 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16878) );
  AOI22_X1 U20132 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16877) );
  NAND4_X1 U20133 ( .A1(n16880), .A2(n16879), .A3(n16878), .A4(n16877), .ZN(
        n16881) );
  AOI211_X1 U20134 ( .C1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .C2(n17044), .A(
        n16882), .B(n16881), .ZN(n16883) );
  NAND4_X1 U20135 ( .A1(n16886), .A2(n16885), .A3(n16884), .A4(n16883), .ZN(
        n17158) );
  INV_X1 U20136 ( .A(n17158), .ZN(n16887) );
  OAI22_X1 U20137 ( .A1(n16889), .A2(n16888), .B1(n16887), .B2(n17101), .ZN(
        P3_U2681) );
  AOI22_X1 U20138 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20139 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16892) );
  AOI22_X1 U20140 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20141 ( .A1(n15535), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16890) );
  NAND4_X1 U20142 ( .A1(n16893), .A2(n16892), .A3(n16891), .A4(n16890), .ZN(
        n16899) );
  AOI22_X1 U20143 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16897) );
  AOI22_X1 U20144 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16896) );
  AOI22_X1 U20145 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16895) );
  AOI22_X1 U20146 ( .A1(n15509), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16894) );
  NAND4_X1 U20147 ( .A1(n16897), .A2(n16896), .A3(n16895), .A4(n16894), .ZN(
        n16898) );
  NOR2_X1 U20148 ( .A1(n16899), .A2(n16898), .ZN(n17166) );
  OAI21_X1 U20149 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16916), .A(n16900), .ZN(
        n16901) );
  AOI22_X1 U20150 ( .A1(n17105), .A2(n17166), .B1(n16901), .B2(n17101), .ZN(
        P3_U2682) );
  OAI21_X1 U20151 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16902), .A(n17101), .ZN(
        n16915) );
  AOI22_X1 U20152 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20153 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20154 ( .A1(n15509), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16911) );
  NOR2_X1 U20155 ( .A1(n16903), .A2(n17091), .ZN(n16909) );
  AOI22_X1 U20156 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U20157 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16906) );
  AOI22_X1 U20158 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20159 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16976), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16904) );
  NAND4_X1 U20160 ( .A1(n16907), .A2(n16906), .A3(n16905), .A4(n16904), .ZN(
        n16908) );
  AOI211_X1 U20161 ( .C1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .C2(n17044), .A(
        n16909), .B(n16908), .ZN(n16910) );
  NAND4_X1 U20162 ( .A1(n16913), .A2(n16912), .A3(n16911), .A4(n16910), .ZN(
        n17167) );
  INV_X1 U20163 ( .A(n17167), .ZN(n16914) );
  OAI22_X1 U20164 ( .A1(n16916), .A2(n16915), .B1(n16914), .B2(n17101), .ZN(
        P3_U2683) );
  AOI22_X1 U20165 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20166 ( .A1(n17060), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U20167 ( .A1(n15535), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20168 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16917) );
  NAND4_X1 U20169 ( .A1(n16920), .A2(n16919), .A3(n16918), .A4(n16917), .ZN(
        n16926) );
  AOI22_X1 U20170 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16924) );
  AOI22_X1 U20171 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20172 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20173 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16921) );
  NAND4_X1 U20174 ( .A1(n16924), .A2(n16923), .A3(n16922), .A4(n16921), .ZN(
        n16925) );
  NOR2_X1 U20175 ( .A1(n16926), .A2(n16925), .ZN(n17176) );
  OAI21_X1 U20176 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n9643), .A(n16927), .ZN(
        n16928) );
  AOI22_X1 U20177 ( .A1(n17105), .A2(n17176), .B1(n16928), .B2(n17101), .ZN(
        P3_U2684) );
  NOR2_X1 U20178 ( .A1(n16929), .A2(n16967), .ZN(n16966) );
  AND2_X1 U20179 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16966), .ZN(n16953) );
  AOI21_X1 U20180 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17101), .A(n16953), .ZN(
        n16940) );
  AOI22_X1 U20181 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20182 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17040), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20183 ( .A1(n15509), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U20184 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16930) );
  NAND4_X1 U20185 ( .A1(n16933), .A2(n16932), .A3(n16931), .A4(n16930), .ZN(
        n16939) );
  AOI22_X1 U20186 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20187 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16936) );
  AOI22_X1 U20188 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U20189 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16934) );
  NAND4_X1 U20190 ( .A1(n16937), .A2(n16936), .A3(n16935), .A4(n16934), .ZN(
        n16938) );
  NOR2_X1 U20191 ( .A1(n16939), .A2(n16938), .ZN(n17181) );
  OAI22_X1 U20192 ( .A1(n9643), .A2(n16940), .B1(n17181), .B2(n17101), .ZN(
        P3_U2685) );
  AOI22_X1 U20193 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n13884), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17067), .ZN(n16945) );
  AOI22_X1 U20194 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17041), .B1(
        n9638), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U20195 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n15509), .B1(
        n15537), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20196 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n15536), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13910), .ZN(n16942) );
  NAND4_X1 U20197 ( .A1(n16945), .A2(n16944), .A3(n16943), .A4(n16942), .ZN(
        n16951) );
  AOI22_X1 U20198 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20199 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17040), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20200 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17045), .ZN(n16947) );
  AOI22_X1 U20201 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17046), .B1(
        n16976), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16946) );
  NAND4_X1 U20202 ( .A1(n16949), .A2(n16948), .A3(n16947), .A4(n16946), .ZN(
        n16950) );
  NOR2_X1 U20203 ( .A1(n16951), .A2(n16950), .ZN(n17186) );
  AOI21_X1 U20204 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17101), .A(n16966), .ZN(
        n16952) );
  OAI22_X1 U20205 ( .A1(n17186), .A2(n17101), .B1(n16953), .B2(n16952), .ZN(
        P3_U2686) );
  AOI22_X1 U20206 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17040), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20207 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16956) );
  AOI22_X1 U20208 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16955) );
  AOI22_X1 U20209 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16954) );
  NAND4_X1 U20210 ( .A1(n16957), .A2(n16956), .A3(n16955), .A4(n16954), .ZN(
        n16963) );
  AOI22_X1 U20211 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U20212 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20213 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16959) );
  AOI22_X1 U20214 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16958) );
  NAND4_X1 U20215 ( .A1(n16961), .A2(n16960), .A3(n16959), .A4(n16958), .ZN(
        n16962) );
  NOR2_X1 U20216 ( .A1(n16963), .A2(n16962), .ZN(n17192) );
  AOI21_X1 U20217 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17101), .A(n16964), .ZN(
        n16965) );
  OAI22_X1 U20218 ( .A1(n17192), .A2(n17101), .B1(n16966), .B2(n16965), .ZN(
        P3_U2687) );
  INV_X1 U20219 ( .A(n16967), .ZN(n16993) );
  NAND2_X1 U20220 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16993), .ZN(n16981) );
  AOI21_X1 U20221 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n16968), .A(n17105), .ZN(
        n16992) );
  AOI22_X1 U20222 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17040), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20223 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16978) );
  AOI22_X1 U20224 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16969) );
  OAI21_X1 U20225 ( .B1(n17043), .B2(n17084), .A(n16969), .ZN(n16975) );
  AOI22_X1 U20226 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20227 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20228 ( .A1(n13884), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20229 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16970) );
  NAND4_X1 U20230 ( .A1(n16973), .A2(n16972), .A3(n16971), .A4(n16970), .ZN(
        n16974) );
  AOI211_X1 U20231 ( .C1(n16976), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16975), .B(n16974), .ZN(n16977) );
  NAND3_X1 U20232 ( .A1(n16979), .A2(n16978), .A3(n16977), .ZN(n17199) );
  AOI22_X1 U20233 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16992), .B1(n17105), 
        .B2(n17199), .ZN(n16980) );
  OAI21_X1 U20234 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16981), .A(n16980), .ZN(
        P3_U2689) );
  AOI22_X1 U20235 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20236 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17040), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U20237 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20238 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16982) );
  NAND4_X1 U20239 ( .A1(n16985), .A2(n16984), .A3(n16983), .A4(n16982), .ZN(
        n16991) );
  AOI22_X1 U20240 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20241 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13884), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20242 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20243 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16986) );
  NAND4_X1 U20244 ( .A1(n16989), .A2(n16988), .A3(n16987), .A4(n16986), .ZN(
        n16990) );
  NOR2_X1 U20245 ( .A1(n16991), .A2(n16990), .ZN(n17204) );
  OAI21_X1 U20246 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n16993), .A(n16992), .ZN(
        n16994) );
  OAI21_X1 U20247 ( .B1(n17204), .B2(n17101), .A(n16994), .ZN(P3_U2690) );
  AOI22_X1 U20248 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20249 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20250 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20251 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16995) );
  NAND4_X1 U20252 ( .A1(n16998), .A2(n16997), .A3(n16996), .A4(n16995), .ZN(
        n17005) );
  AOI22_X1 U20253 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20254 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20255 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13884), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20256 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16976), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17000) );
  NAND4_X1 U20257 ( .A1(n17003), .A2(n17002), .A3(n17001), .A4(n17000), .ZN(
        n17004) );
  NOR2_X1 U20258 ( .A1(n17005), .A2(n17004), .ZN(n17208) );
  NOR2_X1 U20259 ( .A1(n17105), .A2(n17007), .ZN(n17021) );
  NOR2_X1 U20260 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18114), .ZN(n17006) );
  AOI22_X1 U20261 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17021), .B1(n17007), 
        .B2(n17006), .ZN(n17008) );
  OAI21_X1 U20262 ( .B1(n17208), .B2(n17101), .A(n17008), .ZN(P3_U2691) );
  AOI22_X1 U20263 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13884), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20264 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20265 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15536), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20266 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17009) );
  NAND4_X1 U20267 ( .A1(n17012), .A2(n17011), .A3(n17010), .A4(n17009), .ZN(
        n17019) );
  AOI22_X1 U20268 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20269 ( .A1(n17066), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20270 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17061), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20271 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17014) );
  NAND4_X1 U20272 ( .A1(n17017), .A2(n17016), .A3(n17015), .A4(n17014), .ZN(
        n17018) );
  NOR2_X1 U20273 ( .A1(n17019), .A2(n17018), .ZN(n17214) );
  INV_X1 U20274 ( .A(n17020), .ZN(n17022) );
  OAI21_X1 U20275 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17022), .A(n17021), .ZN(
        n17023) );
  OAI21_X1 U20276 ( .B1(n17214), .B2(n17101), .A(n17023), .ZN(P3_U2692) );
  AOI22_X1 U20277 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20278 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20279 ( .A1(n15537), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16976), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20280 ( .A1(n13910), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17024) );
  NAND4_X1 U20281 ( .A1(n17027), .A2(n17026), .A3(n17025), .A4(n17024), .ZN(
        n17033) );
  AOI22_X1 U20282 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20283 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17040), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20284 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20285 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17028) );
  NAND4_X1 U20286 ( .A1(n17031), .A2(n17030), .A3(n17029), .A4(n17028), .ZN(
        n17032) );
  NOR2_X1 U20287 ( .A1(n17033), .A2(n17032), .ZN(n17222) );
  NOR2_X1 U20288 ( .A1(n17105), .A2(n17034), .ZN(n17057) );
  NOR2_X1 U20289 ( .A1(n17035), .A2(n17109), .ZN(n17098) );
  NAND2_X1 U20290 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17098), .ZN(n17090) );
  NOR4_X1 U20291 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17036), .A3(n17056), .A4(
        n17090), .ZN(n17037) );
  AOI22_X1 U20292 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17057), .B1(n17038), 
        .B2(n17037), .ZN(n17039) );
  OAI21_X1 U20293 ( .B1(n17222), .B2(n17101), .A(n17039), .ZN(P3_U2693) );
  AOI22_X1 U20294 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n9638), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17040), .ZN(n17055) );
  AOI22_X1 U20295 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17066), .ZN(n17054) );
  AOI22_X1 U20296 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n15509), .ZN(n17042) );
  OAI21_X1 U20297 ( .B1(n17102), .B2(n17043), .A(n17042), .ZN(n17052) );
  AOI22_X1 U20298 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20299 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17045), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20300 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17067), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n13884), .ZN(n17048) );
  AOI22_X1 U20301 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n15536), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17047) );
  NAND4_X1 U20302 ( .A1(n17050), .A2(n17049), .A3(n17048), .A4(n17047), .ZN(
        n17051) );
  AOI211_X1 U20303 ( .C1(n15537), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n17052), .B(n17051), .ZN(n17053) );
  NAND3_X1 U20304 ( .A1(n17055), .A2(n17054), .A3(n17053), .ZN(n17223) );
  INV_X1 U20305 ( .A(n17223), .ZN(n17059) );
  NOR2_X1 U20306 ( .A1(n17056), .A2(n17075), .ZN(n17077) );
  OAI21_X1 U20307 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17077), .A(n17057), .ZN(
        n17058) );
  OAI21_X1 U20308 ( .B1(n17059), .B2(n17101), .A(n17058), .ZN(P3_U2694) );
  AOI22_X1 U20309 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17060), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20310 ( .A1(n17061), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16999), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17064) );
  AOI22_X1 U20311 ( .A1(n16976), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13910), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17063) );
  AOI22_X1 U20312 ( .A1(n15536), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17046), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17062) );
  NAND4_X1 U20313 ( .A1(n17065), .A2(n17064), .A3(n17063), .A4(n17062), .ZN(
        n17074) );
  AOI22_X1 U20314 ( .A1(n17044), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9633), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20315 ( .A1(n9638), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17066), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20316 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17067), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20317 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15509), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17069) );
  NAND4_X1 U20318 ( .A1(n17072), .A2(n17071), .A3(n17070), .A4(n17069), .ZN(
        n17073) );
  NOR2_X1 U20319 ( .A1(n17074), .A2(n17073), .ZN(n17227) );
  INV_X1 U20320 ( .A(n17075), .ZN(n17082) );
  OAI21_X1 U20321 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17082), .A(n17101), .ZN(
        n17076) );
  OAI22_X1 U20322 ( .A1(n17227), .A2(n17101), .B1(n17077), .B2(n17076), .ZN(
        P3_U2695) );
  NOR2_X1 U20323 ( .A1(n17078), .A2(n17090), .ZN(n17093) );
  NAND2_X1 U20324 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17093), .ZN(n17083) );
  NOR2_X1 U20325 ( .A1(n17079), .A2(n17083), .ZN(n17086) );
  AOI21_X1 U20326 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17101), .A(n17086), .ZN(
        n17081) );
  INV_X1 U20327 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17080) );
  OAI22_X1 U20328 ( .A1(n17082), .A2(n17081), .B1(n17080), .B2(n17101), .ZN(
        P3_U2696) );
  INV_X1 U20329 ( .A(n17083), .ZN(n17089) );
  AOI21_X1 U20330 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17101), .A(n17089), .ZN(
        n17085) );
  OAI22_X1 U20331 ( .A1(n17086), .A2(n17085), .B1(n17084), .B2(n17101), .ZN(
        P3_U2697) );
  AOI21_X1 U20332 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17101), .A(n17093), .ZN(
        n17088) );
  INV_X1 U20333 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17087) );
  OAI22_X1 U20334 ( .A1(n17089), .A2(n17088), .B1(n17087), .B2(n17101), .ZN(
        P3_U2698) );
  INV_X1 U20335 ( .A(n17090), .ZN(n17096) );
  AOI21_X1 U20336 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17101), .A(n17096), .ZN(
        n17092) );
  OAI22_X1 U20337 ( .A1(n17093), .A2(n17092), .B1(n17091), .B2(n17101), .ZN(
        P3_U2699) );
  AOI21_X1 U20338 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17101), .A(n17098), .ZN(
        n17095) );
  INV_X1 U20339 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17094) );
  OAI22_X1 U20340 ( .A1(n17096), .A2(n17095), .B1(n17094), .B2(n17101), .ZN(
        P3_U2700) );
  INV_X1 U20341 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17100) );
  AOI221_X1 U20342 ( .B1(n17097), .B2(n17107), .C1(n18114), .C2(n17107), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17099) );
  AOI211_X1 U20343 ( .C1(n17105), .C2(n17100), .A(n17099), .B(n17098), .ZN(
        P3_U2701) );
  OAI222_X1 U20344 ( .A1(n17104), .A2(n17109), .B1(n17103), .B2(n17107), .C1(
        n17102), .C2(n17101), .ZN(P3_U2702) );
  NAND2_X1 U20345 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17105), .ZN(
        n17106) );
  OAI221_X1 U20346 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17109), .C1(n17108), 
        .C2(n17107), .A(n17106), .ZN(P3_U2703) );
  INV_X1 U20347 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17332) );
  INV_X1 U20348 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17327) );
  INV_X1 U20349 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17371) );
  NAND2_X1 U20350 ( .A1(n17110), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17260) );
  NAND3_X1 U20351 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17112) );
  NAND4_X1 U20352 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17111) );
  NOR3_X2 U20353 ( .A1(n17260), .A2(n17112), .A3(n17111), .ZN(n17226) );
  INV_X1 U20354 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17357) );
  NAND4_X1 U20355 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(P3_EAX_REG_11__SCAN_IN), .ZN(n17113)
         );
  NOR2_X1 U20356 ( .A1(n17357), .A2(n17113), .ZN(n17198) );
  NAND4_X1 U20357 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(n17226), .A4(n17198), .ZN(n17200) );
  NOR2_X2 U20358 ( .A1(n17371), .A2(n17200), .ZN(n17193) );
  INV_X1 U20359 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17319) );
  INV_X1 U20360 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17317) );
  NAND4_X1 U20361 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17114)
         );
  NAND2_X1 U20362 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17154), .ZN(n17153) );
  NAND2_X1 U20363 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17150), .ZN(n17149) );
  NOR2_X2 U20364 ( .A1(n17332), .A2(n17133), .ZN(n17129) );
  NAND2_X1 U20365 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17129), .ZN(n17124) );
  NAND2_X1 U20366 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17120), .ZN(n17119) );
  NAND3_X1 U20367 ( .A1(n17239), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17119), 
        .ZN(n17117) );
  NOR2_X2 U20368 ( .A1(n17115), .A2(n17239), .ZN(n17187) );
  NAND2_X1 U20369 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17187), .ZN(n17116) );
  OAI211_X1 U20370 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17119), .A(n17117), .B(
        n17116), .ZN(P3_U2704) );
  NAND2_X1 U20371 ( .A1(n17118), .A2(n17212), .ZN(n17171) );
  AOI22_X1 U20372 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17187), .ZN(n17122) );
  OAI211_X1 U20373 ( .C1(n17120), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17239), .B(
        n17119), .ZN(n17121) );
  OAI211_X1 U20374 ( .C1(n17123), .C2(n17253), .A(n17122), .B(n17121), .ZN(
        P3_U2705) );
  AOI22_X1 U20375 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17187), .ZN(n17126) );
  OAI211_X1 U20376 ( .C1(n17129), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17239), .B(
        n17124), .ZN(n17125) );
  OAI211_X1 U20377 ( .C1(n17127), .C2(n17253), .A(n17126), .B(n17125), .ZN(
        P3_U2706) );
  INV_X1 U20378 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20379 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17187), .B1(n17257), .B2(
        n17128), .ZN(n17132) );
  AOI211_X1 U20380 ( .C1(n17332), .C2(n17133), .A(n17129), .B(n17212), .ZN(
        n17130) );
  INV_X1 U20381 ( .A(n17130), .ZN(n17131) );
  OAI211_X1 U20382 ( .C1(n17171), .C2(n17211), .A(n17132), .B(n17131), .ZN(
        P3_U2707) );
  AOI22_X1 U20383 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17187), .ZN(n17135) );
  OAI211_X1 U20384 ( .C1(n17138), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17239), .B(
        n17133), .ZN(n17134) );
  OAI211_X1 U20385 ( .C1(n17136), .C2(n17253), .A(n17135), .B(n17134), .ZN(
        P3_U2708) );
  INV_X1 U20386 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20387 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17187), .B1(n17257), .B2(
        n17137), .ZN(n17141) );
  AOI211_X1 U20388 ( .C1(n17327), .C2(n17143), .A(n17138), .B(n17212), .ZN(
        n17139) );
  INV_X1 U20389 ( .A(n17139), .ZN(n17140) );
  OAI211_X1 U20390 ( .C1(n17171), .C2(n17142), .A(n17141), .B(n17140), .ZN(
        P3_U2709) );
  AOI22_X1 U20391 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17187), .ZN(n17146) );
  OAI211_X1 U20392 ( .C1(n17144), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17239), .B(
        n17143), .ZN(n17145) );
  OAI211_X1 U20393 ( .C1(n17147), .C2(n17253), .A(n17146), .B(n17145), .ZN(
        P3_U2710) );
  INV_X1 U20394 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20395 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17187), .B1(n17257), .B2(
        n17148), .ZN(n17152) );
  OAI211_X1 U20396 ( .C1(n17150), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17239), .B(
        n17149), .ZN(n17151) );
  OAI211_X1 U20397 ( .C1(n17171), .C2(n17230), .A(n17152), .B(n17151), .ZN(
        P3_U2711) );
  AOI22_X1 U20398 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17187), .ZN(n17156) );
  OAI211_X1 U20399 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17154), .A(n17239), .B(
        n17153), .ZN(n17155) );
  OAI211_X1 U20400 ( .C1(n17157), .C2(n17253), .A(n17156), .B(n17155), .ZN(
        P3_U2712) );
  INV_X1 U20401 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18111) );
  AOI22_X1 U20402 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17187), .B1(n17257), .B2(
        n17158), .ZN(n17161) );
  INV_X1 U20403 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17313) );
  NOR2_X1 U20404 ( .A1(n18114), .A2(n17189), .ZN(n17183) );
  NAND2_X1 U20405 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17183), .ZN(n17182) );
  NAND2_X1 U20406 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17178), .ZN(n17177) );
  NAND2_X1 U20407 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17172), .ZN(n17168) );
  NAND2_X1 U20408 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17163), .ZN(n17162) );
  OAI21_X1 U20409 ( .B1(n17319), .B2(n17212), .A(n17162), .ZN(n17159) );
  OAI21_X1 U20410 ( .B1(n17319), .B2(n17162), .A(n17159), .ZN(n17160) );
  OAI211_X1 U20411 ( .C1(n18111), .C2(n17171), .A(n17161), .B(n17160), .ZN(
        P3_U2713) );
  AOI22_X1 U20412 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17187), .ZN(n17165) );
  OAI211_X1 U20413 ( .C1(n17163), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17239), .B(
        n17162), .ZN(n17164) );
  OAI211_X1 U20414 ( .C1(n17166), .C2(n17253), .A(n17165), .B(n17164), .ZN(
        P3_U2714) );
  AOI22_X1 U20415 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17187), .B1(n17257), .B2(
        n17167), .ZN(n17170) );
  OAI211_X1 U20416 ( .C1(n17172), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17239), .B(
        n17168), .ZN(n17169) );
  OAI211_X1 U20417 ( .C1(n17171), .C2(n18101), .A(n17170), .B(n17169), .ZN(
        P3_U2715) );
  AOI22_X1 U20418 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17187), .ZN(n17175) );
  AOI211_X1 U20419 ( .C1(n17313), .C2(n17177), .A(n17172), .B(n17212), .ZN(
        n17173) );
  INV_X1 U20420 ( .A(n17173), .ZN(n17174) );
  OAI211_X1 U20421 ( .C1(n17176), .C2(n17253), .A(n17175), .B(n17174), .ZN(
        P3_U2716) );
  AOI22_X1 U20422 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17187), .ZN(n17180) );
  OAI211_X1 U20423 ( .C1(n17178), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17239), .B(
        n17177), .ZN(n17179) );
  OAI211_X1 U20424 ( .C1(n17181), .C2(n17253), .A(n17180), .B(n17179), .ZN(
        P3_U2717) );
  AOI22_X1 U20425 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17187), .ZN(n17185) );
  OAI211_X1 U20426 ( .C1(n17183), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17239), .B(
        n17182), .ZN(n17184) );
  OAI211_X1 U20427 ( .C1(n17186), .C2(n17253), .A(n17185), .B(n17184), .ZN(
        P3_U2718) );
  AOI22_X1 U20428 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17188), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17187), .ZN(n17191) );
  OAI211_X1 U20429 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17193), .A(n17239), .B(
        n17189), .ZN(n17190) );
  OAI211_X1 U20430 ( .C1(n17192), .C2(n17253), .A(n17191), .B(n17190), .ZN(
        P3_U2719) );
  AOI211_X1 U20431 ( .C1(n17371), .C2(n17200), .A(n17212), .B(n17193), .ZN(
        n17194) );
  AOI21_X1 U20432 ( .B1(n17258), .B2(BUF2_REG_15__SCAN_IN), .A(n17194), .ZN(
        n17195) );
  OAI21_X1 U20433 ( .B1(n17196), .B2(n17253), .A(n17195), .ZN(P3_U2720) );
  AND2_X1 U20434 ( .A1(n17197), .A2(n17226), .ZN(n17232) );
  AND2_X1 U20435 ( .A1(n17198), .A2(n17232), .ZN(n17210) );
  NAND2_X1 U20436 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17210), .ZN(n17203) );
  AOI22_X1 U20437 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17258), .B1(n17257), .B2(
        n17199), .ZN(n17202) );
  NAND3_X1 U20438 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17239), .A3(n17200), 
        .ZN(n17201) );
  OAI211_X1 U20439 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17203), .A(n17202), .B(
        n17201), .ZN(P3_U2721) );
  INV_X1 U20440 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17207) );
  INV_X1 U20441 ( .A(n17203), .ZN(n17206) );
  AOI21_X1 U20442 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17239), .A(n17210), .ZN(
        n17205) );
  OAI222_X1 U20443 ( .A1(n17256), .A2(n17207), .B1(n17206), .B2(n17205), .C1(
        n17253), .C2(n17204), .ZN(P3_U2722) );
  INV_X1 U20444 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17361) );
  NAND2_X1 U20445 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17232), .ZN(n17225) );
  NOR2_X1 U20446 ( .A1(n17357), .A2(n17225), .ZN(n17219) );
  NAND2_X1 U20447 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17219), .ZN(n17218) );
  NOR2_X1 U20448 ( .A1(n17361), .A2(n17218), .ZN(n17216) );
  AOI21_X1 U20449 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17239), .A(n17216), .ZN(
        n17209) );
  OAI222_X1 U20450 ( .A1(n17256), .A2(n17211), .B1(n17210), .B2(n17209), .C1(
        n17253), .C2(n17208), .ZN(P3_U2723) );
  INV_X1 U20451 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17217) );
  OAI21_X1 U20452 ( .B1(n17361), .B2(n17212), .A(n17218), .ZN(n17213) );
  INV_X1 U20453 ( .A(n17213), .ZN(n17215) );
  OAI222_X1 U20454 ( .A1(n17256), .A2(n17217), .B1(n17216), .B2(n17215), .C1(
        n17253), .C2(n17214), .ZN(P3_U2724) );
  OAI211_X1 U20455 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17219), .A(n17239), .B(
        n17218), .ZN(n17221) );
  NAND2_X1 U20456 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17258), .ZN(n17220) );
  OAI211_X1 U20457 ( .C1(n17222), .C2(n17253), .A(n17221), .B(n17220), .ZN(
        P3_U2725) );
  NAND2_X1 U20458 ( .A1(n17239), .A2(n17225), .ZN(n17229) );
  AOI22_X1 U20459 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17258), .B1(n17257), .B2(
        n17223), .ZN(n17224) );
  OAI221_X1 U20460 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17225), .C1(n17357), 
        .C2(n17229), .A(n17224), .ZN(P3_U2726) );
  NOR2_X1 U20461 ( .A1(n17226), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n17228) );
  OAI222_X1 U20462 ( .A1(n17256), .A2(n17230), .B1(n17229), .B2(n17228), .C1(
        n17253), .C2(n17227), .ZN(P3_U2727) );
  INV_X1 U20463 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18117) );
  INV_X1 U20464 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17350) );
  INV_X1 U20465 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17346) );
  INV_X1 U20466 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17340) );
  NOR4_X1 U20467 ( .A1(n18114), .A2(n17259), .A3(n17340), .A4(n17338), .ZN(
        n17251) );
  AND2_X1 U20468 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17251), .ZN(n17255) );
  NAND2_X1 U20469 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17255), .ZN(n17243) );
  NOR2_X1 U20470 ( .A1(n17346), .A2(n17243), .ZN(n17247) );
  NAND2_X1 U20471 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17247), .ZN(n17234) );
  NOR2_X1 U20472 ( .A1(n17350), .A2(n17234), .ZN(n17238) );
  AOI21_X1 U20473 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17239), .A(n17238), .ZN(
        n17233) );
  OAI222_X1 U20474 ( .A1(n17256), .A2(n18117), .B1(n17233), .B2(n17232), .C1(
        n17253), .C2(n17231), .ZN(P3_U2728) );
  INV_X1 U20475 ( .A(n17234), .ZN(n17242) );
  AOI21_X1 U20476 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17239), .A(n17242), .ZN(
        n17237) );
  INV_X1 U20477 ( .A(n17235), .ZN(n17236) );
  OAI222_X1 U20478 ( .A1(n18111), .A2(n17256), .B1(n17238), .B2(n17237), .C1(
        n17253), .C2(n17236), .ZN(P3_U2729) );
  INV_X1 U20479 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18105) );
  AOI21_X1 U20480 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17239), .A(n17247), .ZN(
        n17241) );
  OAI222_X1 U20481 ( .A1(n18105), .A2(n17256), .B1(n17242), .B2(n17241), .C1(
        n17253), .C2(n17240), .ZN(P3_U2730) );
  INV_X1 U20482 ( .A(n17243), .ZN(n17250) );
  AOI21_X1 U20483 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17239), .A(n17250), .ZN(
        n17246) );
  INV_X1 U20484 ( .A(n17244), .ZN(n17245) );
  OAI222_X1 U20485 ( .A1(n18101), .A2(n17256), .B1(n17247), .B2(n17246), .C1(
        n17253), .C2(n17245), .ZN(P3_U2731) );
  INV_X1 U20486 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18095) );
  AOI21_X1 U20487 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17239), .A(n17255), .ZN(
        n17249) );
  OAI222_X1 U20488 ( .A1(n18095), .A2(n17256), .B1(n17250), .B2(n17249), .C1(
        n17253), .C2(n17248), .ZN(P3_U2732) );
  INV_X1 U20489 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18090) );
  AOI21_X1 U20490 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17239), .A(n17251), .ZN(
        n17254) );
  OAI222_X1 U20491 ( .A1(n18090), .A2(n17256), .B1(n17255), .B2(n17254), .C1(
        n17253), .C2(n9815), .ZN(P3_U2733) );
  NOR3_X1 U20492 ( .A1(n18114), .A2(n17259), .A3(n17338), .ZN(n17262) );
  OAI22_X1 U20493 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17262), .B1(n17261), .B2(
        n17260), .ZN(n17263) );
  NAND2_X1 U20494 ( .A1(n17264), .A2(n17263), .ZN(P3_U2734) );
  NOR2_X2 U20495 ( .A1(n18688), .A2(n17533), .ZN(n18729) );
  INV_X1 U20496 ( .A(n17265), .ZN(n17266) );
  NOR2_X4 U20497 ( .A1(n18729), .A2(n17284), .ZN(n17281) );
  AND2_X1 U20498 ( .A1(n17281), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20499 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20500 ( .A1(n18729), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17281), .ZN(n17267) );
  OAI21_X1 U20501 ( .B1(n17336), .B2(n17283), .A(n17267), .ZN(P3_U2737) );
  INV_X1 U20502 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U20503 ( .A1(n18729), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17268) );
  OAI21_X1 U20504 ( .B1(n17334), .B2(n17283), .A(n17268), .ZN(P3_U2738) );
  AOI22_X1 U20505 ( .A1(n18729), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17269) );
  OAI21_X1 U20506 ( .B1(n17332), .B2(n17283), .A(n17269), .ZN(P3_U2739) );
  INV_X1 U20507 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20508 ( .A1(n18729), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17270) );
  OAI21_X1 U20509 ( .B1(n17329), .B2(n17283), .A(n17270), .ZN(P3_U2740) );
  AOI22_X1 U20510 ( .A1(n18729), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17271) );
  OAI21_X1 U20511 ( .B1(n17327), .B2(n17283), .A(n17271), .ZN(P3_U2741) );
  INV_X1 U20512 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20513 ( .A1(n18729), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20514 ( .B1(n17325), .B2(n17283), .A(n17272), .ZN(P3_U2742) );
  INV_X1 U20515 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20516 ( .A1(n18729), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17273) );
  OAI21_X1 U20517 ( .B1(n17323), .B2(n17283), .A(n17273), .ZN(P3_U2743) );
  INV_X1 U20518 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17321) );
  AOI22_X1 U20519 ( .A1(n18729), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17274) );
  OAI21_X1 U20520 ( .B1(n17321), .B2(n17283), .A(n17274), .ZN(P3_U2744) );
  CLKBUF_X1 U20521 ( .A(n18729), .Z(n18574) );
  AOI22_X1 U20522 ( .A1(n18574), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17275) );
  OAI21_X1 U20523 ( .B1(n17319), .B2(n17283), .A(n17275), .ZN(P3_U2745) );
  AOI22_X1 U20524 ( .A1(n18574), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17276) );
  OAI21_X1 U20525 ( .B1(n17317), .B2(n17283), .A(n17276), .ZN(P3_U2746) );
  INV_X1 U20526 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20527 ( .A1(n18574), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17277) );
  OAI21_X1 U20528 ( .B1(n17315), .B2(n17283), .A(n17277), .ZN(P3_U2747) );
  AOI22_X1 U20529 ( .A1(n18574), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17278) );
  OAI21_X1 U20530 ( .B1(n17313), .B2(n17283), .A(n17278), .ZN(P3_U2748) );
  INV_X1 U20531 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17311) );
  AOI22_X1 U20532 ( .A1(n18574), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17279) );
  OAI21_X1 U20533 ( .B1(n17311), .B2(n17283), .A(n17279), .ZN(P3_U2749) );
  INV_X1 U20534 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20535 ( .A1(n18574), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17280) );
  OAI21_X1 U20536 ( .B1(n17309), .B2(n17283), .A(n17280), .ZN(P3_U2750) );
  INV_X1 U20537 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U20538 ( .A1(n18574), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17282) );
  OAI21_X1 U20539 ( .B1(n17307), .B2(n17283), .A(n17282), .ZN(P3_U2751) );
  AOI22_X1 U20540 ( .A1(n18574), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17285) );
  OAI21_X1 U20541 ( .B1(n17371), .B2(n17301), .A(n17285), .ZN(P3_U2752) );
  INV_X1 U20542 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20543 ( .A1(n18574), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17286) );
  OAI21_X1 U20544 ( .B1(n17367), .B2(n17301), .A(n17286), .ZN(P3_U2753) );
  INV_X1 U20545 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20546 ( .A1(n18574), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17287) );
  OAI21_X1 U20547 ( .B1(n17365), .B2(n17301), .A(n17287), .ZN(P3_U2754) );
  INV_X1 U20548 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U20549 ( .A1(n18574), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17288) );
  OAI21_X1 U20550 ( .B1(n17363), .B2(n17301), .A(n17288), .ZN(P3_U2755) );
  AOI22_X1 U20551 ( .A1(n18574), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17289) );
  OAI21_X1 U20552 ( .B1(n17361), .B2(n17301), .A(n17289), .ZN(P3_U2756) );
  INV_X1 U20553 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20554 ( .A1(n18574), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17290) );
  OAI21_X1 U20555 ( .B1(n17359), .B2(n17301), .A(n17290), .ZN(P3_U2757) );
  AOI22_X1 U20556 ( .A1(n18574), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17291) );
  OAI21_X1 U20557 ( .B1(n17357), .B2(n17301), .A(n17291), .ZN(P3_U2758) );
  INV_X1 U20558 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U20559 ( .A1(n18574), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17292) );
  OAI21_X1 U20560 ( .B1(n17355), .B2(n17301), .A(n17292), .ZN(P3_U2759) );
  INV_X1 U20561 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20562 ( .A1(n18574), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17293) );
  OAI21_X1 U20563 ( .B1(n17352), .B2(n17301), .A(n17293), .ZN(P3_U2760) );
  AOI22_X1 U20564 ( .A1(n18574), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17294) );
  OAI21_X1 U20565 ( .B1(n17350), .B2(n17301), .A(n17294), .ZN(P3_U2761) );
  INV_X1 U20566 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17348) );
  AOI22_X1 U20567 ( .A1(n18574), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17295) );
  OAI21_X1 U20568 ( .B1(n17348), .B2(n17301), .A(n17295), .ZN(P3_U2762) );
  AOI22_X1 U20569 ( .A1(n18574), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17296) );
  OAI21_X1 U20570 ( .B1(n17346), .B2(n17301), .A(n17296), .ZN(P3_U2763) );
  INV_X1 U20571 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U20572 ( .A1(n18574), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17297) );
  OAI21_X1 U20573 ( .B1(n17344), .B2(n17301), .A(n17297), .ZN(P3_U2764) );
  INV_X1 U20574 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20575 ( .A1(n18574), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17298) );
  OAI21_X1 U20576 ( .B1(n17342), .B2(n17301), .A(n17298), .ZN(P3_U2765) );
  AOI22_X1 U20577 ( .A1(n18574), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17299) );
  OAI21_X1 U20578 ( .B1(n17340), .B2(n17301), .A(n17299), .ZN(P3_U2766) );
  AOI22_X1 U20579 ( .A1(n18574), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17281), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17300) );
  OAI21_X1 U20580 ( .B1(n17338), .B2(n17301), .A(n17300), .ZN(P3_U2767) );
  OR2_X2 U20581 ( .A1(n17303), .A2(n18576), .ZN(n17370) );
  NOR4_X1 U20582 ( .A1(n18732), .A2(n18599), .A3(n17302), .A4(n17303), .ZN(
        n17330) );
  AOI21_X1 U20583 ( .B1(n18599), .B2(n18085), .A(n17303), .ZN(n17304) );
  AOI22_X1 U20584 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17353), .ZN(n17306) );
  OAI21_X1 U20585 ( .B1(n17307), .B2(n17370), .A(n17306), .ZN(P3_U2768) );
  AOI22_X1 U20586 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17353), .ZN(n17308) );
  OAI21_X1 U20587 ( .B1(n17309), .B2(n17370), .A(n17308), .ZN(P3_U2769) );
  AOI22_X1 U20588 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17353), .ZN(n17310) );
  OAI21_X1 U20589 ( .B1(n17311), .B2(n17370), .A(n17310), .ZN(P3_U2770) );
  AOI22_X1 U20590 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17353), .ZN(n17312) );
  OAI21_X1 U20591 ( .B1(n17313), .B2(n17370), .A(n17312), .ZN(P3_U2771) );
  AOI22_X1 U20592 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17353), .ZN(n17314) );
  OAI21_X1 U20593 ( .B1(n17315), .B2(n17370), .A(n17314), .ZN(P3_U2772) );
  AOI22_X1 U20594 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17353), .ZN(n17316) );
  OAI21_X1 U20595 ( .B1(n17317), .B2(n17370), .A(n17316), .ZN(P3_U2773) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17330), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17353), .ZN(n17318) );
  OAI21_X1 U20597 ( .B1(n17319), .B2(n17370), .A(n17318), .ZN(P3_U2774) );
  AOI22_X1 U20598 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17330), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17353), .ZN(n17320) );
  OAI21_X1 U20599 ( .B1(n17321), .B2(n17370), .A(n17320), .ZN(P3_U2775) );
  AOI22_X1 U20600 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17330), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17353), .ZN(n17322) );
  OAI21_X1 U20601 ( .B1(n17323), .B2(n17370), .A(n17322), .ZN(P3_U2776) );
  AOI22_X1 U20602 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17353), .ZN(n17324) );
  OAI21_X1 U20603 ( .B1(n17325), .B2(n17370), .A(n17324), .ZN(P3_U2777) );
  AOI22_X1 U20604 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17353), .ZN(n17326) );
  OAI21_X1 U20605 ( .B1(n17327), .B2(n17370), .A(n17326), .ZN(P3_U2778) );
  AOI22_X1 U20606 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17353), .ZN(n17328) );
  OAI21_X1 U20607 ( .B1(n17329), .B2(n17370), .A(n17328), .ZN(P3_U2779) );
  AOI22_X1 U20608 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17353), .ZN(n17331) );
  OAI21_X1 U20609 ( .B1(n17332), .B2(n17370), .A(n17331), .ZN(P3_U2780) );
  AOI22_X1 U20610 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17353), .ZN(n17333) );
  OAI21_X1 U20611 ( .B1(n17334), .B2(n17370), .A(n17333), .ZN(P3_U2781) );
  AOI22_X1 U20612 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17368), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17353), .ZN(n17335) );
  OAI21_X1 U20613 ( .B1(n17336), .B2(n17370), .A(n17335), .ZN(P3_U2782) );
  AOI22_X1 U20614 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17353), .ZN(n17337) );
  OAI21_X1 U20615 ( .B1(n17338), .B2(n17370), .A(n17337), .ZN(P3_U2783) );
  AOI22_X1 U20616 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17353), .ZN(n17339) );
  OAI21_X1 U20617 ( .B1(n17340), .B2(n17370), .A(n17339), .ZN(P3_U2784) );
  AOI22_X1 U20618 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17353), .ZN(n17341) );
  OAI21_X1 U20619 ( .B1(n17342), .B2(n17370), .A(n17341), .ZN(P3_U2785) );
  AOI22_X1 U20620 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17353), .ZN(n17343) );
  OAI21_X1 U20621 ( .B1(n17344), .B2(n17370), .A(n17343), .ZN(P3_U2786) );
  AOI22_X1 U20622 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17353), .ZN(n17345) );
  OAI21_X1 U20623 ( .B1(n17346), .B2(n17370), .A(n17345), .ZN(P3_U2787) );
  AOI22_X1 U20624 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17353), .ZN(n17347) );
  OAI21_X1 U20625 ( .B1(n17348), .B2(n17370), .A(n17347), .ZN(P3_U2788) );
  AOI22_X1 U20626 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17353), .ZN(n17349) );
  OAI21_X1 U20627 ( .B1(n17350), .B2(n17370), .A(n17349), .ZN(P3_U2789) );
  AOI22_X1 U20628 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17353), .ZN(n17351) );
  OAI21_X1 U20629 ( .B1(n17352), .B2(n17370), .A(n17351), .ZN(P3_U2790) );
  AOI22_X1 U20630 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17353), .ZN(n17354) );
  OAI21_X1 U20631 ( .B1(n17355), .B2(n17370), .A(n17354), .ZN(P3_U2791) );
  AOI22_X1 U20632 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17353), .ZN(n17356) );
  OAI21_X1 U20633 ( .B1(n17357), .B2(n17370), .A(n17356), .ZN(P3_U2792) );
  AOI22_X1 U20634 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17353), .ZN(n17358) );
  OAI21_X1 U20635 ( .B1(n17359), .B2(n17370), .A(n17358), .ZN(P3_U2793) );
  AOI22_X1 U20636 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17353), .ZN(n17360) );
  OAI21_X1 U20637 ( .B1(n17361), .B2(n17370), .A(n17360), .ZN(P3_U2794) );
  AOI22_X1 U20638 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17353), .ZN(n17362) );
  OAI21_X1 U20639 ( .B1(n17363), .B2(n17370), .A(n17362), .ZN(P3_U2795) );
  AOI22_X1 U20640 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17353), .ZN(n17364) );
  OAI21_X1 U20641 ( .B1(n17365), .B2(n17370), .A(n17364), .ZN(P3_U2796) );
  AOI22_X1 U20642 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17353), .ZN(n17366) );
  OAI21_X1 U20643 ( .B1(n17367), .B2(n17370), .A(n17366), .ZN(P3_U2797) );
  AOI22_X1 U20644 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17368), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17353), .ZN(n17369) );
  OAI21_X1 U20645 ( .B1(n17371), .B2(n17370), .A(n17369), .ZN(P3_U2798) );
  NOR3_X1 U20646 ( .A1(n17507), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17372), .ZN(n17381) );
  INV_X1 U20647 ( .A(n17374), .ZN(n17373) );
  NOR3_X1 U20648 ( .A1(n17507), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17373), .ZN(n17395) );
  INV_X1 U20649 ( .A(n17532), .ZN(n17698) );
  OAI21_X1 U20650 ( .B1(n17374), .B2(n17698), .A(n17745), .ZN(n17375) );
  AOI21_X1 U20651 ( .B1(n17574), .B2(n17376), .A(n17375), .ZN(n17408) );
  OAI21_X1 U20652 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17483), .A(
        n17408), .ZN(n17396) );
  OAI21_X1 U20653 ( .B1(n17395), .B2(n17396), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17378) );
  NAND2_X1 U20654 ( .A1(n18032), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17377) );
  OAI211_X1 U20655 ( .C1(n17576), .C2(n17379), .A(n17378), .B(n17377), .ZN(
        n17380) );
  AOI211_X1 U20656 ( .C1(n17382), .C2(n17527), .A(n17381), .B(n17380), .ZN(
        n17389) );
  NAND2_X1 U20657 ( .A1(n17750), .A2(n17649), .ZN(n17482) );
  AOI22_X1 U20658 ( .A1(n17738), .A2(n17755), .B1(n17570), .B2(n17383), .ZN(
        n17409) );
  NAND2_X1 U20659 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17409), .ZN(
        n17397) );
  NAND3_X1 U20660 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17482), .A3(
        n17397), .ZN(n17388) );
  OAI211_X1 U20661 ( .C1(n17386), .C2(n17385), .A(n17636), .B(n17384), .ZN(
        n17387) );
  NAND3_X1 U20662 ( .A1(n17389), .A2(n17388), .A3(n17387), .ZN(P3_U2802) );
  NOR2_X1 U20663 ( .A1(n17391), .A2(n17390), .ZN(n17392) );
  XOR2_X1 U20664 ( .A(n17392), .B(n9876), .Z(n17764) );
  OAI22_X1 U20665 ( .A1(n9637), .A2(n18662), .B1(n17576), .B2(n17393), .ZN(
        n17394) );
  AOI211_X1 U20666 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17396), .A(
        n17395), .B(n17394), .ZN(n17400) );
  OAI21_X1 U20667 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17398), .A(
        n17397), .ZN(n17399) );
  OAI211_X1 U20668 ( .C1(n17764), .C2(n17650), .A(n17400), .B(n17399), .ZN(
        P3_U2803) );
  AOI21_X1 U20669 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17402), .A(
        n17401), .ZN(n17770) );
  NAND3_X1 U20670 ( .A1(n18457), .A2(n17416), .A3(n17417), .ZN(n17406) );
  INV_X1 U20671 ( .A(n17483), .ZN(n17404) );
  OAI21_X1 U20672 ( .B1(n17597), .B2(n17404), .A(n17403), .ZN(n17405) );
  OAI221_X1 U20673 ( .B1(n17408), .B2(n17407), .C1(n17408), .C2(n17406), .A(
        n17405), .ZN(n17413) );
  INV_X1 U20674 ( .A(n17426), .ZN(n17765) );
  NOR2_X1 U20675 ( .A1(n17765), .A2(n17546), .ZN(n17411) );
  INV_X1 U20676 ( .A(n17409), .ZN(n17410) );
  MUX2_X1 U20677 ( .A(n17411), .B(n17410), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17412) );
  AOI211_X1 U20678 ( .C1(n18017), .C2(P3_REIP_REG_26__SCAN_IN), .A(n17413), 
        .B(n17412), .ZN(n17414) );
  OAI21_X1 U20679 ( .B1(n17770), .B2(n17650), .A(n17414), .ZN(P3_U2804) );
  NOR2_X1 U20680 ( .A1(n17757), .A2(n17883), .ZN(n17415) );
  OAI22_X1 U20681 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17415), .B1(
        n17765), .B2(n17883), .ZN(n17783) );
  NAND2_X1 U20682 ( .A1(n17416), .A2(n17588), .ZN(n17433) );
  AOI211_X1 U20683 ( .C1(n17432), .C2(n17422), .A(n17417), .B(n17433), .ZN(
        n17424) );
  AOI22_X1 U20684 ( .A1(n18457), .A2(n17419), .B1(n17574), .B2(n17418), .ZN(
        n17420) );
  NAND2_X1 U20685 ( .A1(n17420), .A2(n17745), .ZN(n17442) );
  AOI21_X1 U20686 ( .B1(n17574), .B2(n9952), .A(n17442), .ZN(n17431) );
  OAI22_X1 U20687 ( .A1(n17431), .A2(n17422), .B1(n17576), .B2(n17421), .ZN(
        n17423) );
  AOI211_X1 U20688 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n18032), .A(n17424), 
        .B(n17423), .ZN(n17430) );
  INV_X1 U20689 ( .A(n17757), .ZN(n17775) );
  AOI21_X1 U20690 ( .B1(n17775), .B2(n17884), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17425) );
  AOI21_X1 U20691 ( .B1(n17884), .B2(n17426), .A(n17425), .ZN(n17780) );
  AOI21_X1 U20692 ( .B1(n9870), .B2(n17648), .A(n17427), .ZN(n17428) );
  XOR2_X1 U20693 ( .A(n17428), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17779) );
  AOI22_X1 U20694 ( .A1(n17570), .A2(n17780), .B1(n17636), .B2(n17779), .ZN(
        n17429) );
  OAI211_X1 U20695 ( .C1(n17750), .C2(n17783), .A(n17430), .B(n17429), .ZN(
        P3_U2805) );
  NAND2_X1 U20696 ( .A1(n17555), .A2(n17436), .ZN(n17789) );
  NAND2_X1 U20697 ( .A1(n17436), .A2(n17884), .ZN(n17788) );
  AOI22_X1 U20698 ( .A1(n17738), .A2(n17789), .B1(n17570), .B2(n17788), .ZN(
        n17448) );
  NAND2_X1 U20699 ( .A1(n18032), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17795) );
  OAI221_X1 U20700 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17433), .C1(
        n17432), .C2(n17431), .A(n17795), .ZN(n17438) );
  AOI21_X1 U20701 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17435), .A(
        n17434), .ZN(n17786) );
  NAND2_X1 U20702 ( .A1(n17436), .A2(n9869), .ZN(n17785) );
  OAI22_X1 U20703 ( .A1(n17786), .A2(n17650), .B1(n17546), .B2(n17785), .ZN(
        n17437) );
  AOI211_X1 U20704 ( .C1(n17597), .C2(n17439), .A(n17438), .B(n17437), .ZN(
        n17440) );
  OAI21_X1 U20705 ( .B1(n17448), .B2(n9869), .A(n17440), .ZN(P3_U2806) );
  AOI22_X1 U20706 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17442), .B1(
        n17597), .B2(n17441), .ZN(n17454) );
  AOI22_X1 U20707 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17648), .B1(
        n17444), .B2(n17456), .ZN(n17445) );
  NAND2_X1 U20708 ( .A1(n17443), .A2(n17445), .ZN(n17447) );
  XOR2_X1 U20709 ( .A(n17447), .B(n17446), .Z(n17797) );
  NOR2_X1 U20710 ( .A1(n17851), .A2(n17457), .ZN(n17811) );
  NAND2_X1 U20711 ( .A1(n17527), .A2(n17811), .ZN(n17468) );
  NOR2_X1 U20712 ( .A1(n17820), .A2(n17468), .ZN(n17450) );
  INV_X1 U20713 ( .A(n17448), .ZN(n17449) );
  MUX2_X1 U20714 ( .A(n17450), .B(n17449), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17451) );
  AOI21_X1 U20715 ( .B1(n17636), .B2(n17797), .A(n17451), .ZN(n17453) );
  NAND2_X1 U20716 ( .A1(n18032), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17803) );
  AND2_X1 U20717 ( .A1(n17588), .A2(n9716), .ZN(n17473) );
  NAND3_X1 U20718 ( .A1(n17461), .A2(n17473), .A3(n9952), .ZN(n17452) );
  NAND4_X1 U20719 ( .A1(n17454), .A2(n17453), .A3(n17803), .A4(n17452), .ZN(
        P3_U2807) );
  INV_X1 U20720 ( .A(n17811), .ZN(n17805) );
  OAI22_X1 U20721 ( .A1(n17555), .A2(n17750), .B1(n17884), .B2(n17649), .ZN(
        n17543) );
  AOI21_X1 U20722 ( .B1(n17482), .B2(n17805), .A(n17543), .ZN(n17481) );
  INV_X1 U20723 ( .A(n17443), .ZN(n17455) );
  AOI221_X1 U20724 ( .B1(n17457), .B2(n17456), .C1(n17474), .C2(n17456), .A(
        n17455), .ZN(n17458) );
  XOR2_X1 U20725 ( .A(n17458), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n17817) );
  OAI21_X1 U20726 ( .B1(n9716), .B2(n17698), .A(n17745), .ZN(n17459) );
  AOI21_X1 U20727 ( .B1(n17574), .B2(n17460), .A(n17459), .ZN(n17484) );
  OAI21_X1 U20728 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17483), .A(
        n17484), .ZN(n17471) );
  AOI21_X1 U20729 ( .B1(n17472), .B2(n17462), .A(n17461), .ZN(n17463) );
  AOI22_X1 U20730 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17471), .B1(
        n17473), .B2(n17463), .ZN(n17464) );
  NAND2_X1 U20731 ( .A1(n18032), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17818) );
  OAI211_X1 U20732 ( .C1(n17576), .C2(n17465), .A(n17464), .B(n17818), .ZN(
        n17466) );
  AOI21_X1 U20733 ( .B1(n17636), .B2(n17817), .A(n17466), .ZN(n17467) );
  OAI221_X1 U20734 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17468), 
        .C1(n17820), .C2(n17481), .A(n17467), .ZN(P3_U2808) );
  OAI22_X1 U20735 ( .A1(n9637), .A2(n18650), .B1(n17576), .B2(n17469), .ZN(
        n17470) );
  AOI221_X1 U20736 ( .B1(n17473), .B2(n17472), .C1(n17471), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17470), .ZN(n17479) );
  INV_X1 U20737 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17518) );
  NOR3_X1 U20738 ( .A1(n17518), .A2(n17648), .A3(n17474), .ZN(n17500) );
  INV_X1 U20739 ( .A(n17475), .ZN(n17514) );
  AOI22_X1 U20740 ( .A1(n17823), .A2(n17500), .B1(n17514), .B2(n17476), .ZN(
        n17477) );
  XOR2_X1 U20741 ( .A(n17480), .B(n17477), .Z(n17828) );
  NOR2_X1 U20742 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17813), .ZN(
        n17827) );
  NOR2_X1 U20743 ( .A1(n17851), .A2(n17518), .ZN(n17821) );
  INV_X1 U20744 ( .A(n17821), .ZN(n17825) );
  NOR2_X1 U20745 ( .A1(n17546), .A2(n17825), .ZN(n17502) );
  AOI22_X1 U20746 ( .A1(n17636), .A2(n17828), .B1(n17827), .B2(n17502), .ZN(
        n17478) );
  OAI211_X1 U20747 ( .C1(n17481), .C2(n17480), .A(n17479), .B(n17478), .ZN(
        P3_U2809) );
  NAND2_X1 U20748 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17821), .ZN(
        n17834) );
  AOI21_X1 U20749 ( .B1(n17482), .B2(n17834), .A(n17543), .ZN(n17505) );
  INV_X1 U20750 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17841) );
  NAND2_X1 U20751 ( .A1(n18032), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17839) );
  INV_X1 U20752 ( .A(n17839), .ZN(n17488) );
  AOI221_X1 U20753 ( .B1(n18427), .B2(n17486), .C1(n17485), .C2(n17486), .A(
        n17484), .ZN(n17487) );
  AOI211_X1 U20754 ( .C1(n17489), .C2(n17737), .A(n17488), .B(n17487), .ZN(
        n17492) );
  OAI221_X1 U20755 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17513), 
        .C1(n17845), .C2(n17500), .A(n17443), .ZN(n17490) );
  XOR2_X1 U20756 ( .A(n17841), .B(n17490), .Z(n17838) );
  NOR2_X1 U20757 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17845), .ZN(
        n17837) );
  AOI22_X1 U20758 ( .A1(n17636), .A2(n17838), .B1(n17502), .B2(n17837), .ZN(
        n17491) );
  OAI211_X1 U20759 ( .C1(n17505), .C2(n17841), .A(n17492), .B(n17491), .ZN(
        P3_U2810) );
  INV_X1 U20760 ( .A(n17742), .ZN(n17670) );
  OAI21_X1 U20761 ( .B1(n17716), .B2(n17506), .A(n17670), .ZN(n17519) );
  OAI21_X1 U20762 ( .B1(n17493), .B2(n17533), .A(n17519), .ZN(n17510) );
  NOR2_X1 U20763 ( .A1(n9637), .A2(n18645), .ZN(n17844) );
  NOR2_X1 U20764 ( .A1(n17511), .A2(n17494), .ZN(n17498) );
  OAI211_X1 U20765 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17495), .B(n17588), .ZN(n17497) );
  OAI22_X1 U20766 ( .A1(n17498), .A2(n17497), .B1(n17496), .B2(n17576), .ZN(
        n17499) );
  AOI211_X1 U20767 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17510), .A(
        n17844), .B(n17499), .ZN(n17504) );
  AOI21_X1 U20768 ( .B1(n17513), .B2(n17514), .A(n17500), .ZN(n17501) );
  XOR2_X1 U20769 ( .A(n17845), .B(n17501), .Z(n17843) );
  AOI22_X1 U20770 ( .A1(n17636), .A2(n17843), .B1(n17502), .B2(n17845), .ZN(
        n17503) );
  OAI211_X1 U20771 ( .C1(n17505), .C2(n17845), .A(n17504), .B(n17503), .ZN(
        P3_U2811) );
  AOI21_X1 U20772 ( .B1(n17527), .B2(n17851), .A(n17543), .ZN(n17530) );
  NOR2_X1 U20773 ( .A1(n17507), .A2(n17506), .ZN(n17512) );
  OAI22_X1 U20774 ( .A1(n9637), .A2(n18643), .B1(n17576), .B2(n17508), .ZN(
        n17509) );
  AOI221_X1 U20775 ( .B1(n17512), .B2(n17511), .C1(n17510), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17509), .ZN(n17517) );
  AOI21_X1 U20776 ( .B1(n9876), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17513), .ZN(n17515) );
  XOR2_X1 U20777 ( .A(n17515), .B(n17514), .Z(n17860) );
  NOR2_X1 U20778 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17851), .ZN(
        n17859) );
  AOI22_X1 U20779 ( .A1(n17636), .A2(n17860), .B1(n17527), .B2(n17859), .ZN(
        n17516) );
  OAI211_X1 U20780 ( .C1(n17530), .C2(n17518), .A(n17517), .B(n17516), .ZN(
        P3_U2812) );
  NAND2_X1 U20781 ( .A1(n18032), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17867) );
  INV_X1 U20782 ( .A(n17867), .ZN(n17523) );
  AOI221_X1 U20783 ( .B1(n18427), .B2(n17521), .C1(n17520), .C2(n17521), .A(
        n17519), .ZN(n17522) );
  AOI211_X1 U20784 ( .C1(n17524), .C2(n17737), .A(n17523), .B(n17522), .ZN(
        n17529) );
  OAI21_X1 U20785 ( .B1(n17526), .B2(n17855), .A(n17525), .ZN(n17864) );
  NOR2_X1 U20786 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17877), .ZN(
        n17863) );
  AOI22_X1 U20787 ( .A1(n17636), .A2(n17864), .B1(n17527), .B2(n17863), .ZN(
        n17528) );
  OAI211_X1 U20788 ( .C1(n17530), .C2(n17855), .A(n17529), .B(n17528), .ZN(
        P3_U2813) );
  AOI21_X1 U20789 ( .B1(n17532), .B2(n17531), .A(n17716), .ZN(n17562) );
  OAI21_X1 U20790 ( .B1(n17534), .B2(n17533), .A(n17562), .ZN(n17554) );
  NAND2_X1 U20791 ( .A1(n17535), .A2(n17588), .ZN(n17552) );
  AOI221_X1 U20792 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C1(n17537), .C2(n17536), .A(
        n17552), .ZN(n17540) );
  OAI22_X1 U20793 ( .A1(n9637), .A2(n18639), .B1(n17576), .B2(n17538), .ZN(
        n17539) );
  AOI211_X1 U20794 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n17554), .A(
        n17540), .B(n17539), .ZN(n17545) );
  NOR2_X1 U20795 ( .A1(n17648), .A2(n17937), .ZN(n17628) );
  INV_X1 U20796 ( .A(n17628), .ZN(n17619) );
  OAI22_X1 U20797 ( .A1(n9876), .A2(n17541), .B1(n17619), .B2(n17858), .ZN(
        n17542) );
  XOR2_X1 U20798 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17542), .Z(
        n17879) );
  AOI22_X1 U20799 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17543), .B1(
        n17636), .B2(n17879), .ZN(n17544) );
  OAI211_X1 U20800 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17546), .A(
        n17545), .B(n17544), .ZN(P3_U2814) );
  NOR3_X1 U20801 ( .A1(n17595), .A2(n10040), .A3(n15598), .ZN(n17548) );
  AOI21_X1 U20802 ( .B1(n9681), .B2(n17548), .A(n17547), .ZN(n17549) );
  AOI221_X1 U20803 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17933), 
        .C1(n17648), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17549), .ZN(
        n17550) );
  XOR2_X1 U20804 ( .A(n15597), .B(n17550), .Z(n17890) );
  NOR2_X1 U20805 ( .A1(n9637), .A2(n18637), .ZN(n17893) );
  OAI22_X1 U20806 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17552), .B1(
        n17551), .B2(n17576), .ZN(n17553) );
  AOI211_X1 U20807 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17554), .A(
        n17893), .B(n17553), .ZN(n17559) );
  NOR2_X1 U20808 ( .A1(n17555), .A2(n17750), .ZN(n17557) );
  NAND2_X1 U20809 ( .A1(n17560), .A2(n15597), .ZN(n17882) );
  NOR2_X1 U20810 ( .A1(n17884), .A2(n17649), .ZN(n17556) );
  OR2_X1 U20811 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17567), .ZN(
        n17888) );
  AOI22_X1 U20812 ( .A1(n17557), .A2(n17882), .B1(n17556), .B2(n17888), .ZN(
        n17558) );
  OAI211_X1 U20813 ( .C1(n17650), .C2(n17890), .A(n17559), .B(n17558), .ZN(
        P3_U2815) );
  OAI21_X1 U20814 ( .B1(n17561), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17560), .ZN(n17911) );
  AOI221_X1 U20815 ( .B1(n17564), .B2(n17563), .C1(n18427), .C2(n17563), .A(
        n17562), .ZN(n17565) );
  NOR2_X1 U20816 ( .A1(n9637), .A2(n18635), .ZN(n17905) );
  AOI211_X1 U20817 ( .C1(n17566), .C2(n17737), .A(n17565), .B(n17905), .ZN(
        n17572) );
  AOI221_X1 U20818 ( .B1(n17937), .B2(n15598), .C1(n17903), .C2(n15598), .A(
        n17567), .ZN(n17907) );
  OAI21_X1 U20819 ( .B1(n17903), .B2(n17619), .A(n17568), .ZN(n17569) );
  XOR2_X1 U20820 ( .A(n17569), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n17906) );
  AOI22_X1 U20821 ( .A1(n17570), .A2(n17907), .B1(n17636), .B2(n17906), .ZN(
        n17571) );
  OAI211_X1 U20822 ( .C1(n17750), .C2(n17911), .A(n17572), .B(n17571), .ZN(
        P3_U2816) );
  NAND2_X1 U20823 ( .A1(n17915), .A2(n10040), .ZN(n17922) );
  AOI21_X1 U20824 ( .B1(n17574), .B2(n17573), .A(n17716), .ZN(n17575) );
  OAI21_X1 U20825 ( .B1(n17605), .B2(n17698), .A(n17575), .ZN(n17589) );
  NOR2_X1 U20826 ( .A1(n9637), .A2(n18633), .ZN(n17581) );
  OAI211_X1 U20827 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17605), .B(n17588), .ZN(n17578) );
  OAI22_X1 U20828 ( .A1(n17579), .A2(n17578), .B1(n17577), .B2(n17576), .ZN(
        n17580) );
  AOI211_X1 U20829 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17589), .A(
        n17581), .B(n17580), .ZN(n17587) );
  NOR2_X1 U20830 ( .A1(n17923), .A2(n17937), .ZN(n17582) );
  OAI22_X1 U20831 ( .A1(n17583), .A2(n17750), .B1(n17582), .B2(n17649), .ZN(
        n17594) );
  AOI22_X1 U20832 ( .A1(n9681), .A2(n17915), .B1(n17933), .B2(n17648), .ZN(
        n17584) );
  AOI21_X1 U20833 ( .B1(n17592), .B2(n17648), .A(n17584), .ZN(n17585) );
  XOR2_X1 U20834 ( .A(n17585), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n17912) );
  AOI22_X1 U20835 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17594), .B1(
        n17636), .B2(n17912), .ZN(n17586) );
  OAI211_X1 U20836 ( .C1(n17639), .C2(n17922), .A(n17587), .B(n17586), .ZN(
        P3_U2817) );
  AND2_X1 U20837 ( .A1(n17588), .A2(n17605), .ZN(n17591) );
  NOR2_X1 U20838 ( .A1(n9637), .A2(n18631), .ZN(n17930) );
  AOI221_X1 U20839 ( .B1(n17591), .B2(n17590), .C1(n17589), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17930), .ZN(n17601) );
  OAI21_X1 U20840 ( .B1(n17595), .B2(n17619), .A(n17592), .ZN(n17593) );
  XOR2_X1 U20841 ( .A(n17593), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17931) );
  AOI22_X1 U20842 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17594), .B1(
        n17636), .B2(n17931), .ZN(n17600) );
  INV_X1 U20843 ( .A(n17595), .ZN(n17925) );
  INV_X1 U20844 ( .A(n17639), .ZN(n17615) );
  NAND3_X1 U20845 ( .A1(n17925), .A2(n17933), .A3(n17615), .ZN(n17599) );
  NAND2_X1 U20846 ( .A1(n17597), .A2(n17596), .ZN(n17598) );
  NAND4_X1 U20847 ( .A1(n17601), .A2(n17600), .A3(n17599), .A4(n17598), .ZN(
        P3_U2818) );
  OAI22_X1 U20848 ( .A1(n17914), .A2(n17649), .B1(n17750), .B2(n17602), .ZN(
        n17626) );
  AOI21_X1 U20849 ( .B1(n17943), .B2(n17615), .A(n17626), .ZN(n17625) );
  INV_X1 U20850 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17631) );
  NAND4_X1 U20851 ( .A1(n18457), .A2(n17658), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A4(n17603), .ZN(n17632) );
  NOR2_X1 U20852 ( .A1(n17631), .A2(n17632), .ZN(n17630) );
  AOI22_X1 U20853 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17670), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17630), .ZN(n17604) );
  AOI21_X1 U20854 ( .B1(n17605), .B2(n18457), .A(n17604), .ZN(n17607) );
  NOR2_X1 U20855 ( .A1(n9637), .A2(n18629), .ZN(n17606) );
  AOI211_X1 U20856 ( .C1(n17608), .C2(n17737), .A(n17607), .B(n17606), .ZN(
        n17613) );
  AOI21_X1 U20857 ( .B1(n17610), .B2(n17628), .A(n17609), .ZN(n17611) );
  XOR2_X1 U20858 ( .A(n17614), .B(n17611), .Z(n17935) );
  NOR2_X1 U20859 ( .A1(n17943), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17934) );
  AOI22_X1 U20860 ( .A1(n17636), .A2(n17935), .B1(n17934), .B2(n17615), .ZN(
        n17612) );
  OAI211_X1 U20861 ( .C1(n17625), .C2(n17614), .A(n17613), .B(n17612), .ZN(
        P3_U2819) );
  AOI21_X1 U20862 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17615), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17624) );
  NOR2_X1 U20863 ( .A1(n17630), .A2(n17617), .ZN(n17616) );
  NOR2_X1 U20864 ( .A1(n9637), .A2(n18627), .ZN(n17950) );
  AOI221_X1 U20865 ( .B1(n17630), .B2(n17617), .C1(n17616), .C2(n17670), .A(
        n17950), .ZN(n17623) );
  OAI21_X1 U20866 ( .B1(n17962), .B2(n17619), .A(n17618), .ZN(n17620) );
  XOR2_X1 U20867 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n17620), .Z(
        n17951) );
  AOI22_X1 U20868 ( .A1(n17636), .A2(n17951), .B1(n17621), .B2(n17737), .ZN(
        n17622) );
  OAI211_X1 U20869 ( .C1(n17625), .C2(n17624), .A(n17623), .B(n17622), .ZN(
        P3_U2820) );
  INV_X1 U20870 ( .A(n17626), .ZN(n17638) );
  NOR2_X1 U20871 ( .A1(n17628), .A2(n17627), .ZN(n17629) );
  XOR2_X1 U20872 ( .A(n17629), .B(n17962), .Z(n17966) );
  AOI211_X1 U20873 ( .C1(n17632), .C2(n17631), .A(n17742), .B(n17630), .ZN(
        n17635) );
  NAND2_X1 U20874 ( .A1(n18032), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17968) );
  OAI21_X1 U20875 ( .B1(n17729), .B2(n17633), .A(n17968), .ZN(n17634) );
  AOI211_X1 U20876 ( .C1(n17636), .C2(n17966), .A(n17635), .B(n17634), .ZN(
        n17637) );
  OAI221_X1 U20877 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17639), .C1(
        n17962), .C2(n17638), .A(n17637), .ZN(P3_U2821) );
  OAI21_X1 U20878 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17641), .A(
        n17640), .ZN(n17988) );
  OAI21_X1 U20879 ( .B1(n17642), .B2(n17698), .A(n17745), .ZN(n17659) );
  OAI211_X1 U20880 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17644), .A(
        n18457), .B(n17643), .ZN(n17645) );
  NAND2_X1 U20881 ( .A1(n18032), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17979) );
  OAI211_X1 U20882 ( .C1(n17729), .C2(n17646), .A(n17645), .B(n17979), .ZN(
        n17652) );
  AOI21_X1 U20883 ( .B1(n17648), .B2(n17981), .A(n17647), .ZN(n17983) );
  OAI22_X1 U20884 ( .A1(n17983), .A2(n17650), .B1(n17649), .B2(n17981), .ZN(
        n17651) );
  AOI211_X1 U20885 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17659), .A(
        n17652), .B(n17651), .ZN(n17653) );
  OAI21_X1 U20886 ( .B1(n17750), .B2(n17988), .A(n17653), .ZN(P3_U2822) );
  OAI21_X1 U20887 ( .B1(n17656), .B2(n17655), .A(n17654), .ZN(n17657) );
  XOR2_X1 U20888 ( .A(n17657), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n17997) );
  NAND2_X1 U20889 ( .A1(n18457), .A2(n17658), .ZN(n17676) );
  NOR2_X1 U20890 ( .A1(n17675), .A2(n17676), .ZN(n17661) );
  NOR2_X1 U20891 ( .A1(n9637), .A2(n18621), .ZN(n17989) );
  AOI221_X1 U20892 ( .B1(n17661), .B2(n17660), .C1(n17659), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17989), .ZN(n17667) );
  AOI21_X1 U20893 ( .B1(n17664), .B2(n17663), .A(n17662), .ZN(n17994) );
  AOI22_X1 U20894 ( .A1(n17734), .A2(n17994), .B1(n17665), .B2(n17737), .ZN(
        n17666) );
  OAI211_X1 U20895 ( .C1(n17750), .C2(n17997), .A(n17667), .B(n17666), .ZN(
        P3_U2823) );
  OAI21_X1 U20896 ( .B1(n17669), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17668), .ZN(n18005) );
  NAND2_X1 U20897 ( .A1(n17670), .A2(n17676), .ZN(n17692) );
  AOI21_X1 U20898 ( .B1(n17673), .B2(n17672), .A(n17671), .ZN(n17998) );
  AOI22_X1 U20899 ( .A1(n17734), .A2(n17998), .B1(n18032), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17674) );
  OAI221_X1 U20900 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17676), .C1(
        n17675), .C2(n17692), .A(n17674), .ZN(n17677) );
  AOI21_X1 U20901 ( .B1(n17678), .B2(n17737), .A(n17677), .ZN(n17679) );
  OAI21_X1 U20902 ( .B1(n17750), .B2(n18005), .A(n17679), .ZN(P3_U2824) );
  INV_X1 U20903 ( .A(n17680), .ZN(n17681) );
  AOI21_X1 U20904 ( .B1(n17681), .B2(n17745), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17693) );
  OAI21_X1 U20905 ( .B1(n17684), .B2(n17683), .A(n17682), .ZN(n17685) );
  XNOR2_X1 U20906 ( .A(n17685), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18012) );
  NOR2_X1 U20907 ( .A1(n9637), .A2(n18618), .ZN(n18009) );
  OAI21_X1 U20908 ( .B1(n17688), .B2(n17687), .A(n17686), .ZN(n18006) );
  OAI22_X1 U20909 ( .A1(n17729), .A2(n17689), .B1(n17750), .B2(n18006), .ZN(
        n17690) );
  AOI211_X1 U20910 ( .C1(n17734), .C2(n18012), .A(n18009), .B(n17690), .ZN(
        n17691) );
  OAI21_X1 U20911 ( .B1(n17693), .B2(n17692), .A(n17691), .ZN(P3_U2825) );
  INV_X1 U20912 ( .A(n17694), .ZN(n17707) );
  AOI21_X1 U20913 ( .B1(n17697), .B2(n17696), .A(n17695), .ZN(n18016) );
  AOI22_X1 U20914 ( .A1(n17734), .A2(n18016), .B1(n18032), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n17706) );
  OAI21_X1 U20915 ( .B1(n9919), .B2(n17698), .A(n17745), .ZN(n17719) );
  OAI21_X1 U20916 ( .B1(n17701), .B2(n17700), .A(n17699), .ZN(n17702) );
  XOR2_X1 U20917 ( .A(n17702), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18025) );
  OAI22_X1 U20918 ( .A1(n17729), .A2(n17703), .B1(n17750), .B2(n18025), .ZN(
        n17704) );
  AOI21_X1 U20919 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17719), .A(
        n17704), .ZN(n17705) );
  OAI211_X1 U20920 ( .C1(n18427), .C2(n17707), .A(n17706), .B(n17705), .ZN(
        P3_U2826) );
  OAI21_X1 U20921 ( .B1(n17710), .B2(n17709), .A(n17708), .ZN(n18027) );
  OAI21_X1 U20922 ( .B1(n17713), .B2(n17712), .A(n17711), .ZN(n17714) );
  XOR2_X1 U20923 ( .A(n17714), .B(n10039), .Z(n18031) );
  AOI22_X1 U20924 ( .A1(n17734), .A2(n18031), .B1(n18032), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17721) );
  INV_X1 U20925 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17732) );
  OAI21_X1 U20926 ( .B1(n17716), .B2(n17732), .A(n17715), .ZN(n17718) );
  AOI22_X1 U20927 ( .A1(n17719), .A2(n17718), .B1(n17717), .B2(n17737), .ZN(
        n17720) );
  OAI211_X1 U20928 ( .C1(n17750), .C2(n18027), .A(n17721), .B(n17720), .ZN(
        P3_U2827) );
  AOI21_X1 U20929 ( .B1(n17724), .B2(n17723), .A(n17722), .ZN(n18040) );
  NOR2_X1 U20930 ( .A1(n9637), .A2(n18611), .ZN(n18049) );
  OAI21_X1 U20931 ( .B1(n17727), .B2(n17726), .A(n17725), .ZN(n18044) );
  OAI22_X1 U20932 ( .A1(n17729), .A2(n17728), .B1(n17750), .B2(n18044), .ZN(
        n17730) );
  AOI211_X1 U20933 ( .C1(n17734), .C2(n18040), .A(n18049), .B(n17730), .ZN(
        n17731) );
  OAI221_X1 U20934 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18427), .C1(
        n17732), .C2(n17745), .A(n17731), .ZN(P3_U2828) );
  AOI21_X1 U20935 ( .B1(n17735), .B2(n17743), .A(n17733), .ZN(n18056) );
  AOI22_X1 U20936 ( .A1(n17734), .A2(n18056), .B1(n18032), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17740) );
  NOR2_X1 U20937 ( .A1(n17744), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17736) );
  XNOR2_X1 U20938 ( .A(n17736), .B(n17735), .ZN(n18052) );
  AOI22_X1 U20939 ( .A1(n17738), .A2(n18052), .B1(n17741), .B2(n17737), .ZN(
        n17739) );
  OAI211_X1 U20940 ( .C1(n17742), .C2(n17741), .A(n17740), .B(n17739), .ZN(
        P3_U2829) );
  OAI21_X1 U20941 ( .B1(n17744), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17743), .ZN(n17749) );
  INV_X1 U20942 ( .A(n17749), .ZN(n18069) );
  OAI211_X1 U20943 ( .C1(P3_STATE2_REG_0__SCAN_IN), .C2(n18742), .A(n18688), 
        .B(n17745), .ZN(n17746) );
  AOI22_X1 U20944 ( .A1(n18017), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17746), .ZN(n17747) );
  OAI221_X1 U20945 ( .B1(n18069), .B2(n17750), .C1(n17749), .C2(n17748), .A(
        n17747), .ZN(P3_U2830) );
  AOI22_X1 U20946 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18058), .B1(
        n18032), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n17763) );
  NOR3_X1 U20947 ( .A1(n17799), .A2(n17751), .A3(n17765), .ZN(n17761) );
  AND2_X1 U20948 ( .A1(n17972), .A2(n17752), .ZN(n17754) );
  AOI211_X1 U20949 ( .C1(n18509), .C2(n17755), .A(n17754), .B(n17753), .ZN(
        n17758) );
  OAI21_X1 U20950 ( .B1(n18537), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17756), .ZN(n17852) );
  OAI21_X1 U20951 ( .B1(n17757), .B2(n17852), .A(n17972), .ZN(n17771) );
  OAI211_X1 U20952 ( .C1(n17759), .C2(n17913), .A(n17758), .B(n17771), .ZN(
        n17766) );
  OAI221_X1 U20953 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17761), 
        .C1(n17760), .C2(n17766), .A(n18019), .ZN(n17762) );
  OAI211_X1 U20954 ( .C1(n17764), .C2(n17982), .A(n17763), .B(n17762), .ZN(
        P3_U2835) );
  AOI22_X1 U20955 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18058), .B1(
        n18032), .B2(P3_REIP_REG_26__SCAN_IN), .ZN(n17769) );
  NOR2_X1 U20956 ( .A1(n17799), .A2(n17765), .ZN(n17767) );
  OAI211_X1 U20957 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17767), .A(
        n17766), .B(n18019), .ZN(n17768) );
  OAI211_X1 U20958 ( .C1(n17770), .C2(n17982), .A(n17769), .B(n17768), .ZN(
        P3_U2836) );
  NAND3_X1 U20959 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17772), .A3(
        n17771), .ZN(n17773) );
  OAI221_X1 U20960 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17775), 
        .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n17774), .A(n17773), .ZN(
        n17777) );
  OAI22_X1 U20961 ( .A1(n18065), .A2(n17777), .B1(n17776), .B2(n18035), .ZN(
        n17778) );
  AOI21_X1 U20962 ( .B1(n18017), .B2(P3_REIP_REG_25__SCAN_IN), .A(n17778), 
        .ZN(n17782) );
  AOI22_X1 U20963 ( .A1(n17908), .A2(n17780), .B1(n17967), .B2(n17779), .ZN(
        n17781) );
  OAI211_X1 U20964 ( .C1(n18068), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        P3_U2837) );
  INV_X1 U20965 ( .A(n17784), .ZN(n17826) );
  OAI22_X1 U20966 ( .A1(n17786), .A2(n17982), .B1(n17826), .B2(n17785), .ZN(
        n17787) );
  INV_X1 U20967 ( .A(n17787), .ZN(n17796) );
  INV_X1 U20968 ( .A(n18020), .ZN(n17992) );
  AOI22_X1 U20969 ( .A1(n18509), .A2(n17789), .B1(n17938), .B2(n17788), .ZN(
        n17791) );
  OAI21_X1 U20970 ( .B1(n17798), .B2(n17852), .A(n17972), .ZN(n17790) );
  NAND3_X1 U20971 ( .A1(n17791), .A2(n18035), .A3(n17790), .ZN(n17793) );
  AOI221_X1 U20972 ( .B1(n17798), .B2(n18548), .C1(n17850), .C2(n18548), .A(
        n17793), .ZN(n17792) );
  AOI21_X1 U20973 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17792), .A(
        n18032), .ZN(n17800) );
  OAI211_X1 U20974 ( .C1(n17992), .C2(n17793), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17800), .ZN(n17794) );
  NAND3_X1 U20975 ( .A1(n17796), .A2(n17795), .A3(n17794), .ZN(P3_U2838) );
  INV_X1 U20976 ( .A(n17797), .ZN(n17804) );
  NOR3_X1 U20977 ( .A1(n18058), .A2(n17799), .A3(n17798), .ZN(n17801) );
  OAI21_X1 U20978 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17801), .A(
        n17800), .ZN(n17802) );
  OAI211_X1 U20979 ( .C1(n17804), .C2(n17982), .A(n17803), .B(n17802), .ZN(
        P3_U2839) );
  OAI22_X1 U20980 ( .A1(n18065), .A2(n17820), .B1(n17826), .B2(n17805), .ZN(
        n17816) );
  OAI21_X1 U20981 ( .B1(n17850), .B2(n17825), .A(n18548), .ZN(n17809) );
  OAI21_X1 U20982 ( .B1(n17807), .B2(n17834), .A(n18539), .ZN(n17808) );
  NOR2_X1 U20983 ( .A1(n18509), .A2(n17938), .ZN(n17831) );
  OAI22_X1 U20984 ( .A1(n18552), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17811), .B2(n17831), .ZN(n17810) );
  NOR2_X1 U20985 ( .A1(n17832), .A2(n17810), .ZN(n17822) );
  AOI21_X1 U20986 ( .B1(n17871), .B2(n17811), .A(n18537), .ZN(n17812) );
  AOI211_X1 U20987 ( .C1(n18548), .C2(n17813), .A(n17812), .B(n17820), .ZN(
        n17814) );
  OAI211_X1 U20988 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n17954), .A(
        n17822), .B(n17814), .ZN(n17815) );
  AOI22_X1 U20989 ( .A1(n17967), .A2(n17817), .B1(n17816), .B2(n17815), .ZN(
        n17819) );
  OAI211_X1 U20990 ( .C1(n18035), .C2(n17820), .A(n17819), .B(n17818), .ZN(
        P3_U2840) );
  OAI221_X1 U20991 ( .B1(n18537), .B2(n17871), .C1(n18537), .C2(n17821), .A(
        n18019), .ZN(n17833) );
  NOR2_X1 U20992 ( .A1(n18548), .A2(n18524), .ZN(n18057) );
  OAI21_X1 U20993 ( .B1(n17823), .B2(n18057), .A(n17822), .ZN(n17824) );
  OAI21_X1 U20994 ( .B1(n17833), .B2(n17824), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17830) );
  NOR2_X1 U20995 ( .A1(n17826), .A2(n17825), .ZN(n17846) );
  AOI22_X1 U20996 ( .A1(n17967), .A2(n17828), .B1(n17827), .B2(n17846), .ZN(
        n17829) );
  OAI221_X1 U20997 ( .B1(n18017), .B2(n17830), .C1(n9637), .C2(n18650), .A(
        n17829), .ZN(P3_U2841) );
  NOR3_X1 U20998 ( .A1(n18057), .A2(n18742), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17836) );
  INV_X1 U20999 ( .A(n17831), .ZN(n17942) );
  NOR2_X1 U21000 ( .A1(n18032), .A2(n17835), .ZN(n17847) );
  NOR2_X1 U21001 ( .A1(n17836), .A2(n17847), .ZN(n17842) );
  AOI22_X1 U21002 ( .A1(n17967), .A2(n17838), .B1(n17837), .B2(n17846), .ZN(
        n17840) );
  OAI211_X1 U21003 ( .C1(n17842), .C2(n17841), .A(n17840), .B(n17839), .ZN(
        P3_U2842) );
  INV_X1 U21004 ( .A(n17843), .ZN(n17849) );
  AOI221_X1 U21005 ( .B1(n17847), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), 
        .C1(n17846), .C2(n17845), .A(n17844), .ZN(n17848) );
  OAI21_X1 U21006 ( .B1(n17849), .B2(n17982), .A(n17848), .ZN(P3_U2843) );
  AOI222_X1 U21007 ( .A1(n18548), .A2(n17851), .B1(n18548), .B2(n17850), .C1(
        n17851), .C2(n17942), .ZN(n17854) );
  OAI21_X1 U21008 ( .B1(n17877), .B2(n17852), .A(n17972), .ZN(n17853) );
  NAND4_X1 U21009 ( .A1(n17869), .A2(n18019), .A3(n17854), .A4(n17853), .ZN(
        n17865) );
  OAI221_X1 U21010 ( .B1(n17865), .B2(n17972), .C1(n17865), .C2(n17855), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17862) );
  OAI22_X1 U21011 ( .A1(n17973), .A2(n18039), .B1(n17971), .B2(n18036), .ZN(
        n18026) );
  AND2_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18026), .ZN(
        n17975) );
  NAND2_X1 U21013 ( .A1(n17856), .A2(n17975), .ZN(n17902) );
  NAND2_X1 U21014 ( .A1(n17857), .A2(n17902), .ZN(n17924) );
  NAND2_X1 U21015 ( .A1(n18019), .A2(n17924), .ZN(n17970) );
  NOR2_X1 U21016 ( .A1(n17858), .A2(n17970), .ZN(n17878) );
  AOI22_X1 U21017 ( .A1(n17967), .A2(n17860), .B1(n17878), .B2(n17859), .ZN(
        n17861) );
  OAI221_X1 U21018 ( .B1(n18017), .B2(n17862), .C1(n9637), .C2(n18643), .A(
        n17861), .ZN(P3_U2844) );
  AOI22_X1 U21019 ( .A1(n17967), .A2(n17864), .B1(n17878), .B2(n17863), .ZN(
        n17868) );
  NAND3_X1 U21020 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n9637), .A3(
        n17865), .ZN(n17866) );
  NAND3_X1 U21021 ( .A1(n17868), .A2(n17867), .A3(n17866), .ZN(P3_U2845) );
  NAND2_X1 U21022 ( .A1(n17869), .A2(n18019), .ZN(n17876) );
  OR2_X1 U21023 ( .A1(n18552), .A2(n17870), .ZN(n17952) );
  NAND2_X1 U21024 ( .A1(n18537), .A2(n17952), .ZN(n17960) );
  INV_X1 U21025 ( .A(n17871), .ZN(n17872) );
  OAI21_X1 U21026 ( .B1(n15597), .B2(n17960), .A(n17872), .ZN(n17874) );
  INV_X1 U21027 ( .A(n17873), .ZN(n17897) );
  NAND2_X1 U21028 ( .A1(n18548), .A2(n17897), .ZN(n17963) );
  OAI211_X1 U21029 ( .C1(n17875), .C2(n17954), .A(n17874), .B(n17963), .ZN(
        n17887) );
  OAI221_X1 U21030 ( .B1(n17876), .B2(n17992), .C1(n17876), .C2(n17887), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17881) );
  AOI22_X1 U21031 ( .A1(n17967), .A2(n17879), .B1(n17878), .B2(n17877), .ZN(
        n17880) );
  OAI221_X1 U21032 ( .B1(n18017), .B2(n17881), .C1(n9637), .C2(n18639), .A(
        n17880), .ZN(P3_U2846) );
  NAND3_X1 U21033 ( .A1(n17883), .A2(n18010), .A3(n17882), .ZN(n17895) );
  NOR2_X1 U21034 ( .A1(n17884), .A2(n17913), .ZN(n17889) );
  OAI21_X1 U21035 ( .B1(n17885), .B2(n17902), .A(n15597), .ZN(n17886) );
  AOI22_X1 U21036 ( .A1(n17889), .A2(n17888), .B1(n17887), .B2(n17886), .ZN(
        n17891) );
  OAI22_X1 U21037 ( .A1(n18065), .A2(n17891), .B1(n17890), .B2(n17982), .ZN(
        n17892) );
  AOI211_X1 U21038 ( .C1(n18058), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17893), .B(n17892), .ZN(n17894) );
  NAND2_X1 U21039 ( .A1(n17895), .A2(n17894), .ZN(P3_U2847) );
  INV_X1 U21040 ( .A(n17903), .ZN(n17896) );
  OAI22_X1 U21041 ( .A1(n18552), .A2(n17896), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18057), .ZN(n17900) );
  OAI21_X1 U21042 ( .B1(n17923), .B2(n17961), .A(n18524), .ZN(n17918) );
  OAI21_X1 U21043 ( .B1(n17923), .B2(n17897), .A(n18548), .ZN(n17898) );
  NAND4_X1 U21044 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17918), .A3(
        n17952), .A4(n17898), .ZN(n17899) );
  OAI21_X1 U21045 ( .B1(n17900), .B2(n17899), .A(n18019), .ZN(n17901) );
  AOI221_X1 U21046 ( .B1(n17903), .B2(n15598), .C1(n17902), .C2(n15598), .A(
        n17901), .ZN(n17904) );
  AOI211_X1 U21047 ( .C1(n18058), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17905), .B(n17904), .ZN(n17910) );
  AOI22_X1 U21048 ( .A1(n17908), .A2(n17907), .B1(n17967), .B2(n17906), .ZN(
        n17909) );
  OAI211_X1 U21049 ( .C1(n18068), .C2(n17911), .A(n17910), .B(n17909), .ZN(
        P3_U2848) );
  AOI22_X1 U21050 ( .A1(n18017), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17967), 
        .B2(n17912), .ZN(n17921) );
  AOI21_X1 U21051 ( .B1(n17915), .B2(n17914), .A(n17913), .ZN(n17916) );
  OAI211_X1 U21052 ( .C1(n17925), .C2(n17954), .A(n17952), .B(n17963), .ZN(
        n17945) );
  AOI211_X1 U21053 ( .C1(n18509), .C2(n17917), .A(n17916), .B(n17945), .ZN(
        n17928) );
  OAI211_X1 U21054 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17954), .A(
        n17928), .B(n17918), .ZN(n17919) );
  OAI211_X1 U21055 ( .C1(n18065), .C2(n17919), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n9637), .ZN(n17920) );
  OAI211_X1 U21056 ( .C1(n17970), .C2(n17922), .A(n17921), .B(n17920), .ZN(
        P3_U2849) );
  OAI22_X1 U21057 ( .A1(n18524), .A2(n17933), .B1(n17923), .B2(n17961), .ZN(
        n17927) );
  AOI21_X1 U21058 ( .B1(n17925), .B2(n17924), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17926) );
  AOI211_X1 U21059 ( .C1(n17928), .C2(n17927), .A(n18065), .B(n17926), .ZN(
        n17929) );
  AOI211_X1 U21060 ( .C1(n17967), .C2(n17931), .A(n17930), .B(n17929), .ZN(
        n17932) );
  OAI21_X1 U21061 ( .B1(n17933), .B2(n18035), .A(n17932), .ZN(P3_U2850) );
  INV_X1 U21062 ( .A(n17934), .ZN(n17948) );
  AOI22_X1 U21063 ( .A1(n18017), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17967), 
        .B2(n17935), .ZN(n17947) );
  OAI21_X1 U21064 ( .B1(n17962), .B2(n17961), .A(n18524), .ZN(n17936) );
  INV_X1 U21065 ( .A(n17936), .ZN(n17941) );
  AOI22_X1 U21066 ( .A1(n18509), .A2(n17939), .B1(n17938), .B2(n17937), .ZN(
        n17940) );
  NAND2_X1 U21067 ( .A1(n17940), .A2(n18019), .ZN(n17959) );
  AOI211_X1 U21068 ( .C1(n17943), .C2(n17942), .A(n17941), .B(n17959), .ZN(
        n17953) );
  OAI21_X1 U21069 ( .B1(n18537), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17953), .ZN(n17944) );
  OAI211_X1 U21070 ( .C1(n17945), .C2(n17944), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n9637), .ZN(n17946) );
  OAI211_X1 U21071 ( .C1(n17948), .C2(n17970), .A(n17947), .B(n17946), .ZN(
        P3_U2851) );
  NOR3_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17962), .A3(
        n17970), .ZN(n17949) );
  AOI211_X1 U21073 ( .C1(n17967), .C2(n17951), .A(n17950), .B(n17949), .ZN(
        n17958) );
  NAND2_X1 U21074 ( .A1(n17963), .A2(n17952), .ZN(n17956) );
  OAI21_X1 U21075 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17954), .A(
        n17953), .ZN(n17955) );
  OAI211_X1 U21076 ( .C1(n17956), .C2(n17955), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n9637), .ZN(n17957) );
  NAND2_X1 U21077 ( .A1(n17958), .A2(n17957), .ZN(P3_U2852) );
  AOI21_X1 U21078 ( .B1(n17961), .B2(n17960), .A(n17959), .ZN(n17964) );
  AOI211_X1 U21079 ( .C1(n17964), .C2(n17963), .A(n18017), .B(n17962), .ZN(
        n17965) );
  AOI21_X1 U21080 ( .B1(n17967), .B2(n17966), .A(n17965), .ZN(n17969) );
  OAI211_X1 U21081 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17970), .A(
        n17969), .B(n17968), .ZN(P3_U2853) );
  AOI22_X1 U21082 ( .A1(n18524), .A2(n18705), .B1(n17972), .B2(n17971), .ZN(
        n18037) );
  NAND2_X1 U21083 ( .A1(n18548), .A2(n17973), .ZN(n18043) );
  NAND3_X1 U21084 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18037), .A3(
        n18043), .ZN(n18018) );
  NOR2_X1 U21085 ( .A1(n17974), .A2(n18018), .ZN(n17991) );
  OAI21_X1 U21086 ( .B1(n17991), .B2(n18053), .A(n18035), .ZN(n17986) );
  INV_X1 U21087 ( .A(n17974), .ZN(n17977) );
  INV_X1 U21088 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17976) );
  NAND2_X1 U21089 ( .A1(n17975), .A2(n18019), .ZN(n18007) );
  INV_X1 U21090 ( .A(n18007), .ZN(n18021) );
  NAND3_X1 U21091 ( .A1(n17977), .A2(n17976), .A3(n18021), .ZN(n17978) );
  NAND2_X1 U21092 ( .A1(n17979), .A2(n17978), .ZN(n17985) );
  OAI22_X1 U21093 ( .A1(n17983), .A2(n17982), .B1(n17981), .B2(n17980), .ZN(
        n17984) );
  AOI211_X1 U21094 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n17986), .A(
        n17985), .B(n17984), .ZN(n17987) );
  OAI21_X1 U21095 ( .B1(n18068), .B2(n17988), .A(n17987), .ZN(P3_U2854) );
  AOI21_X1 U21096 ( .B1(n18058), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17989), .ZN(n17996) );
  NAND2_X1 U21097 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17999) );
  NOR2_X1 U21098 ( .A1(n17999), .A2(n18007), .ZN(n18002) );
  AOI22_X1 U21099 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18019), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18002), .ZN(n17990) );
  NOR2_X1 U21100 ( .A1(n17991), .A2(n17990), .ZN(n17993) );
  AOI22_X1 U21101 ( .A1(n17994), .A2(n18064), .B1(n17993), .B2(n17992), .ZN(
        n17995) );
  OAI211_X1 U21102 ( .C1(n18068), .C2(n17997), .A(n17996), .B(n17995), .ZN(
        P3_U2855) );
  AOI22_X1 U21103 ( .A1(n18017), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18064), 
        .B2(n17998), .ZN(n18004) );
  NOR2_X1 U21104 ( .A1(n18018), .A2(n17999), .ZN(n18000) );
  OAI21_X1 U21105 ( .B1(n18000), .B2(n18053), .A(n18035), .ZN(n18013) );
  AOI22_X1 U21106 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18013), .B1(
        n18002), .B2(n18001), .ZN(n18003) );
  OAI211_X1 U21107 ( .C1(n18068), .C2(n18005), .A(n18004), .B(n18003), .ZN(
        P3_U2856) );
  INV_X1 U21108 ( .A(n18006), .ZN(n18011) );
  NOR3_X1 U21109 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20898), .A3(
        n18007), .ZN(n18008) );
  AOI211_X1 U21110 ( .C1(n18011), .C2(n18010), .A(n18009), .B(n18008), .ZN(
        n18015) );
  AOI22_X1 U21111 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18013), .B1(
        n18064), .B2(n18012), .ZN(n18014) );
  NAND2_X1 U21112 ( .A1(n18015), .A2(n18014), .ZN(P3_U2857) );
  AOI22_X1 U21113 ( .A1(n18017), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18064), 
        .B2(n18016), .ZN(n18024) );
  NAND2_X1 U21114 ( .A1(n18019), .A2(n18018), .ZN(n18028) );
  OAI21_X1 U21115 ( .B1(n18020), .B2(n18028), .A(n18035), .ZN(n18022) );
  AOI22_X1 U21116 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18022), .B1(
        n18021), .B2(n20898), .ZN(n18023) );
  OAI211_X1 U21117 ( .C1(n18068), .C2(n18025), .A(n18024), .B(n18023), .ZN(
        P3_U2858) );
  NOR2_X1 U21118 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18026), .ZN(
        n18029) );
  OAI22_X1 U21119 ( .A1(n18029), .A2(n18028), .B1(n18068), .B2(n18027), .ZN(
        n18030) );
  AOI21_X1 U21120 ( .B1(n18064), .B2(n18031), .A(n18030), .ZN(n18034) );
  NAND2_X1 U21121 ( .A1(n18032), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18033) );
  OAI211_X1 U21122 ( .C1(n18035), .C2(n10039), .A(n18034), .B(n18033), .ZN(
        P3_U2859) );
  NOR2_X1 U21123 ( .A1(n18689), .A2(n18036), .ZN(n18048) );
  NAND2_X1 U21124 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18038) );
  OAI21_X1 U21125 ( .B1(n18039), .B2(n18038), .A(n18037), .ZN(n18047) );
  NAND2_X1 U21126 ( .A1(n18041), .A2(n18040), .ZN(n18042) );
  OAI211_X1 U21127 ( .C1(n18045), .C2(n18044), .A(n18043), .B(n18042), .ZN(
        n18046) );
  AOI221_X1 U21128 ( .B1(n18048), .B2(n15583), .C1(n18047), .C2(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n18046), .ZN(n18051) );
  AOI21_X1 U21129 ( .B1(n18058), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18049), .ZN(n18050) );
  OAI21_X1 U21130 ( .B1(n18065), .B2(n18051), .A(n18050), .ZN(P3_U2860) );
  INV_X1 U21131 ( .A(n18052), .ZN(n18061) );
  NOR2_X1 U21132 ( .A1(n9637), .A2(n18721), .ZN(n18055) );
  AOI211_X1 U21133 ( .C1(n18552), .C2(n18705), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18053), .ZN(n18054) );
  AOI211_X1 U21134 ( .C1(n18064), .C2(n18056), .A(n18055), .B(n18054), .ZN(
        n18060) );
  NOR3_X1 U21135 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18065), .A3(
        n18057), .ZN(n18062) );
  OAI21_X1 U21136 ( .B1(n18058), .B2(n18062), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18059) );
  OAI211_X1 U21137 ( .C1(n18061), .C2(n18068), .A(n18060), .B(n18059), .ZN(
        P3_U2861) );
  NOR2_X1 U21138 ( .A1(n9637), .A2(n18712), .ZN(n18063) );
  AOI211_X1 U21139 ( .C1(n18064), .C2(n18069), .A(n18063), .B(n18062), .ZN(
        n18067) );
  OAI211_X1 U21140 ( .C1(n18065), .C2(n18539), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n9637), .ZN(n18066) );
  OAI211_X1 U21141 ( .C1(n18069), .C2(n18068), .A(n18067), .B(n18066), .ZN(
        P3_U2862) );
  OAI211_X1 U21142 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18070), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18071)
         );
  INV_X1 U21143 ( .A(n18071), .ZN(n18578) );
  OAI21_X1 U21144 ( .B1(n18578), .B2(n18122), .A(n18076), .ZN(n18072) );
  OAI221_X1 U21145 ( .B1(n18540), .B2(n18726), .C1(n18540), .C2(n18076), .A(
        n18072), .ZN(P3_U2863) );
  NAND2_X1 U21146 ( .A1(n18561), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18347) );
  NAND2_X1 U21147 ( .A1(n18562), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18229) );
  NOR2_X1 U21148 ( .A1(n18369), .A2(n18255), .ZN(n18074) );
  OAI22_X1 U21149 ( .A1(n18075), .A2(n18562), .B1(n18074), .B2(n18073), .ZN(
        P3_U2866) );
  NOR2_X1 U21150 ( .A1(n18563), .A2(n18076), .ZN(P3_U2867) );
  NOR2_X1 U21151 ( .A1(n18427), .A2(n18077), .ZN(n18453) );
  NAND2_X1 U21152 ( .A1(n18540), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18230) );
  NAND2_X1 U21153 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18078) );
  NOR2_X2 U21154 ( .A1(n18230), .A2(n18078), .ZN(n18430) );
  AND2_X1 U21155 ( .A1(n18374), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18452) );
  NOR2_X1 U21156 ( .A1(n18562), .A2(n18253), .ZN(n18455) );
  NAND2_X1 U21157 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18455), .ZN(
        n18508) );
  NOR2_X1 U21158 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18544) );
  NAND2_X1 U21159 ( .A1(n18561), .A2(n18562), .ZN(n18163) );
  INV_X1 U21160 ( .A(n18163), .ZN(n18164) );
  NAND2_X1 U21161 ( .A1(n18544), .A2(n18164), .ZN(n18153) );
  NOR2_X1 U21162 ( .A1(n18159), .A2(n18181), .ZN(n18141) );
  NOR2_X1 U21163 ( .A1(n18571), .A2(n18141), .ZN(n18118) );
  AND2_X1 U21164 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18457), .ZN(n18458) );
  NOR2_X1 U21165 ( .A1(n18078), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18456) );
  NAND2_X1 U21166 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18456), .ZN(
        n18423) );
  INV_X1 U21167 ( .A(n18423), .ZN(n18502) );
  AOI22_X1 U21168 ( .A1(n18452), .A2(n18118), .B1(n18458), .B2(n18502), .ZN(
        n18084) );
  INV_X1 U21169 ( .A(n18230), .ZN(n18323) );
  NOR2_X1 U21170 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18540), .ZN(
        n18301) );
  NOR2_X1 U21171 ( .A1(n18323), .A2(n18301), .ZN(n18372) );
  NOR2_X1 U21172 ( .A1(n18372), .A2(n18078), .ZN(n18424) );
  AOI211_X1 U21173 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18141), .B(n18426), .ZN(
        n18079) );
  AOI21_X1 U21174 ( .B1(n18457), .B2(n18424), .A(n18079), .ZN(n18119) );
  NOR2_X1 U21175 ( .A1(n18081), .A2(n18080), .ZN(n18115) );
  NAND2_X1 U21176 ( .A1(n18082), .A2(n18115), .ZN(n18461) );
  INV_X1 U21177 ( .A(n18461), .ZN(n18397) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18119), .B1(
        n18181), .B2(n18397), .ZN(n18083) );
  OAI211_X1 U21179 ( .C1(n18400), .C2(n18450), .A(n18084), .B(n18083), .ZN(
        P3_U2868) );
  NAND2_X1 U21180 ( .A1(n18115), .A2(n18085), .ZN(n18467) );
  NOR2_X2 U21181 ( .A1(n18086), .A2(n18427), .ZN(n18463) );
  AND2_X1 U21182 ( .A1(n18374), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18462) );
  AOI22_X1 U21183 ( .A1(n18463), .A2(n18502), .B1(n18462), .B2(n18118), .ZN(
        n18088) );
  AND2_X1 U21184 ( .A1(n18457), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18464) );
  AOI22_X1 U21185 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18119), .B1(
        n18464), .B2(n18430), .ZN(n18087) );
  OAI211_X1 U21186 ( .C1(n18153), .C2(n18467), .A(n18088), .B(n18087), .ZN(
        P3_U2869) );
  NAND2_X1 U21187 ( .A1(n18089), .A2(n18115), .ZN(n18473) );
  NAND2_X1 U21188 ( .A1(n18457), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18286) );
  INV_X1 U21189 ( .A(n18286), .ZN(n18469) );
  NOR2_X2 U21190 ( .A1(n18426), .A2(n18090), .ZN(n18468) );
  AOI22_X1 U21191 ( .A1(n18469), .A2(n18430), .B1(n18468), .B2(n18118), .ZN(
        n18093) );
  NOR2_X2 U21192 ( .A1(n18091), .A2(n18427), .ZN(n18470) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18119), .B1(
        n18470), .B2(n18502), .ZN(n18092) );
  OAI211_X1 U21194 ( .C1(n18153), .C2(n18473), .A(n18093), .B(n18092), .ZN(
        P3_U2870) );
  NOR2_X1 U21195 ( .A1(n18427), .A2(n18094), .ZN(n18475) );
  INV_X1 U21196 ( .A(n18475), .ZN(n18408) );
  NOR2_X2 U21197 ( .A1(n20933), .A2(n18427), .ZN(n18476) );
  NOR2_X2 U21198 ( .A1(n18426), .A2(n18095), .ZN(n18474) );
  AOI22_X1 U21199 ( .A1(n18476), .A2(n18502), .B1(n18474), .B2(n18118), .ZN(
        n18098) );
  NAND2_X1 U21200 ( .A1(n18096), .A2(n18115), .ZN(n18479) );
  INV_X1 U21201 ( .A(n18479), .ZN(n18405) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18119), .B1(
        n18181), .B2(n18405), .ZN(n18097) );
  OAI211_X1 U21203 ( .C1(n18408), .C2(n18450), .A(n18098), .B(n18097), .ZN(
        P3_U2871) );
  NAND2_X1 U21204 ( .A1(n18099), .A2(n18115), .ZN(n18485) );
  INV_X1 U21205 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18100) );
  NOR2_X2 U21206 ( .A1(n18426), .A2(n18101), .ZN(n18480) );
  AOI22_X1 U21207 ( .A1(n18481), .A2(n18430), .B1(n18480), .B2(n18118), .ZN(
        n18103) );
  AND2_X1 U21208 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18457), .ZN(n18482) );
  AOI22_X1 U21209 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18119), .B1(
        n18482), .B2(n18502), .ZN(n18102) );
  OAI211_X1 U21210 ( .C1(n18153), .C2(n18485), .A(n18103), .B(n18102), .ZN(
        P3_U2872) );
  NAND2_X1 U21211 ( .A1(n18115), .A2(n18104), .ZN(n18491) );
  NOR2_X2 U21212 ( .A1(n18426), .A2(n18105), .ZN(n18487) );
  NOR2_X2 U21213 ( .A1(n18427), .A2(n18106), .ZN(n18486) );
  AOI22_X1 U21214 ( .A1(n18487), .A2(n18118), .B1(n18486), .B2(n18430), .ZN(
        n18108) );
  AND2_X1 U21215 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18457), .ZN(n18488) );
  AOI22_X1 U21216 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18119), .B1(
        n18488), .B2(n18502), .ZN(n18107) );
  OAI211_X1 U21217 ( .C1(n18153), .C2(n18491), .A(n18108), .B(n18107), .ZN(
        P3_U2873) );
  NAND2_X1 U21218 ( .A1(n18115), .A2(n18109), .ZN(n18497) );
  NOR2_X2 U21219 ( .A1(n18110), .A2(n18427), .ZN(n18493) );
  NOR2_X2 U21220 ( .A1(n18426), .A2(n18111), .ZN(n18492) );
  AOI22_X1 U21221 ( .A1(n18493), .A2(n18502), .B1(n18492), .B2(n18118), .ZN(
        n18113) );
  AND2_X1 U21222 ( .A1(n18457), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18494) );
  AOI22_X1 U21223 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18119), .B1(
        n18494), .B2(n18430), .ZN(n18112) );
  OAI211_X1 U21224 ( .C1(n18153), .C2(n18497), .A(n18113), .B(n18112), .ZN(
        P3_U2874) );
  NAND2_X1 U21225 ( .A1(n18115), .A2(n18114), .ZN(n18507) );
  NOR2_X2 U21226 ( .A1(n18427), .A2(n18116), .ZN(n18501) );
  NOR2_X2 U21227 ( .A1(n18117), .A2(n18426), .ZN(n18499) );
  AOI22_X1 U21228 ( .A1(n18501), .A2(n18502), .B1(n18499), .B2(n18118), .ZN(
        n18121) );
  AND2_X1 U21229 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18457), .ZN(n18503) );
  AOI22_X1 U21230 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18119), .B1(
        n18503), .B2(n18430), .ZN(n18120) );
  OAI211_X1 U21231 ( .C1(n18153), .C2(n18507), .A(n18121), .B(n18120), .ZN(
        P3_U2875) );
  NAND2_X1 U21232 ( .A1(n18164), .A2(n18301), .ZN(n18175) );
  NAND2_X1 U21233 ( .A1(n18541), .A2(n18451), .ZN(n18302) );
  NOR2_X1 U21234 ( .A1(n18163), .A2(n18302), .ZN(n18137) );
  AOI22_X1 U21235 ( .A1(n18159), .A2(n18453), .B1(n18452), .B2(n18137), .ZN(
        n18124) );
  NOR2_X1 U21236 ( .A1(n18426), .A2(n18122), .ZN(n18454) );
  AND2_X1 U21237 ( .A1(n18541), .A2(n18454), .ZN(n18208) );
  AOI22_X1 U21238 ( .A1(n18457), .A2(n18455), .B1(n18164), .B2(n18208), .ZN(
        n18138) );
  AOI22_X1 U21239 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18138), .B1(
        n18458), .B2(n18430), .ZN(n18123) );
  OAI211_X1 U21240 ( .C1(n18175), .C2(n18461), .A(n18124), .B(n18123), .ZN(
        P3_U2876) );
  AOI22_X1 U21241 ( .A1(n18463), .A2(n18430), .B1(n18462), .B2(n18137), .ZN(
        n18126) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18138), .B1(
        n18159), .B2(n18464), .ZN(n18125) );
  OAI211_X1 U21243 ( .C1(n18175), .C2(n18467), .A(n18126), .B(n18125), .ZN(
        P3_U2877) );
  AOI22_X1 U21244 ( .A1(n18468), .A2(n18137), .B1(n18470), .B2(n18430), .ZN(
        n18128) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18138), .B1(
        n18159), .B2(n18469), .ZN(n18127) );
  OAI211_X1 U21246 ( .C1(n18175), .C2(n18473), .A(n18128), .B(n18127), .ZN(
        P3_U2878) );
  AOI22_X1 U21247 ( .A1(n18159), .A2(n18475), .B1(n18474), .B2(n18137), .ZN(
        n18130) );
  AOI22_X1 U21248 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18138), .B1(
        n18476), .B2(n18430), .ZN(n18129) );
  OAI211_X1 U21249 ( .C1(n18175), .C2(n18479), .A(n18130), .B(n18129), .ZN(
        P3_U2879) );
  AOI22_X1 U21250 ( .A1(n18480), .A2(n18137), .B1(n18482), .B2(n18430), .ZN(
        n18132) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18138), .B1(
        n18159), .B2(n18481), .ZN(n18131) );
  OAI211_X1 U21252 ( .C1(n18175), .C2(n18485), .A(n18132), .B(n18131), .ZN(
        P3_U2880) );
  AOI22_X1 U21253 ( .A1(n18488), .A2(n18430), .B1(n18487), .B2(n18137), .ZN(
        n18134) );
  AOI22_X1 U21254 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18138), .B1(
        n18159), .B2(n18486), .ZN(n18133) );
  OAI211_X1 U21255 ( .C1(n18175), .C2(n18491), .A(n18134), .B(n18133), .ZN(
        P3_U2881) );
  AOI22_X1 U21256 ( .A1(n18493), .A2(n18430), .B1(n18492), .B2(n18137), .ZN(
        n18136) );
  AOI22_X1 U21257 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18138), .B1(
        n18159), .B2(n18494), .ZN(n18135) );
  OAI211_X1 U21258 ( .C1(n18175), .C2(n18497), .A(n18136), .B(n18135), .ZN(
        P3_U2882) );
  AOI22_X1 U21259 ( .A1(n18159), .A2(n18503), .B1(n18499), .B2(n18137), .ZN(
        n18140) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18138), .B1(
        n18501), .B2(n18430), .ZN(n18139) );
  OAI211_X1 U21261 ( .C1(n18175), .C2(n18507), .A(n18140), .B(n18139), .ZN(
        P3_U2883) );
  NOR2_X2 U21262 ( .A1(n18230), .A2(n18163), .ZN(n18225) );
  INV_X1 U21263 ( .A(n18225), .ZN(n18194) );
  AOI21_X1 U21264 ( .B1(n18194), .B2(n18175), .A(n18571), .ZN(n18158) );
  AOI22_X1 U21265 ( .A1(n18159), .A2(n18458), .B1(n18452), .B2(n18158), .ZN(
        n18144) );
  AOI221_X1 U21266 ( .B1(n18141), .B2(n18175), .C1(n18324), .C2(n18175), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18142) );
  OAI21_X1 U21267 ( .B1(n18225), .B2(n18142), .A(n18374), .ZN(n18160) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18160), .B1(
        n18225), .B2(n18397), .ZN(n18143) );
  OAI211_X1 U21269 ( .C1(n18153), .C2(n18400), .A(n18144), .B(n18143), .ZN(
        P3_U2884) );
  AOI22_X1 U21270 ( .A1(n18181), .A2(n18464), .B1(n18158), .B2(n18462), .ZN(
        n18146) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18160), .B1(
        n18159), .B2(n18463), .ZN(n18145) );
  OAI211_X1 U21272 ( .C1(n18194), .C2(n18467), .A(n18146), .B(n18145), .ZN(
        P3_U2885) );
  AOI22_X1 U21273 ( .A1(n18159), .A2(n18470), .B1(n18158), .B2(n18468), .ZN(
        n18148) );
  INV_X1 U21274 ( .A(n18473), .ZN(n18283) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18160), .B1(
        n18225), .B2(n18283), .ZN(n18147) );
  OAI211_X1 U21276 ( .C1(n18153), .C2(n18286), .A(n18148), .B(n18147), .ZN(
        P3_U2886) );
  AOI22_X1 U21277 ( .A1(n18159), .A2(n18476), .B1(n18158), .B2(n18474), .ZN(
        n18150) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18160), .B1(
        n18225), .B2(n18405), .ZN(n18149) );
  OAI211_X1 U21279 ( .C1(n18153), .C2(n18408), .A(n18150), .B(n18149), .ZN(
        P3_U2887) );
  INV_X1 U21280 ( .A(n18481), .ZN(n18413) );
  AOI22_X1 U21281 ( .A1(n18159), .A2(n18482), .B1(n18158), .B2(n18480), .ZN(
        n18152) );
  INV_X1 U21282 ( .A(n18485), .ZN(n18409) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18160), .B1(
        n18225), .B2(n18409), .ZN(n18151) );
  OAI211_X1 U21284 ( .C1(n18153), .C2(n18413), .A(n18152), .B(n18151), .ZN(
        P3_U2888) );
  AOI22_X1 U21285 ( .A1(n18181), .A2(n18486), .B1(n18158), .B2(n18487), .ZN(
        n18155) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18160), .B1(
        n18159), .B2(n18488), .ZN(n18154) );
  OAI211_X1 U21287 ( .C1(n18194), .C2(n18491), .A(n18155), .B(n18154), .ZN(
        P3_U2889) );
  AOI22_X1 U21288 ( .A1(n18181), .A2(n18494), .B1(n18158), .B2(n18492), .ZN(
        n18157) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18160), .B1(
        n18159), .B2(n18493), .ZN(n18156) );
  OAI211_X1 U21290 ( .C1(n18194), .C2(n18497), .A(n18157), .B(n18156), .ZN(
        P3_U2890) );
  AOI22_X1 U21291 ( .A1(n18181), .A2(n18503), .B1(n18158), .B2(n18499), .ZN(
        n18162) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18160), .B1(
        n18159), .B2(n18501), .ZN(n18161) );
  OAI211_X1 U21293 ( .C1(n18194), .C2(n18507), .A(n18162), .B(n18161), .ZN(
        P3_U2891) );
  NOR2_X1 U21294 ( .A1(n18541), .A2(n18163), .ZN(n18209) );
  NAND2_X1 U21295 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18209), .ZN(
        n18185) );
  AOI21_X1 U21296 ( .B1(n18541), .B2(n18324), .A(n18426), .ZN(n18254) );
  OAI211_X1 U21297 ( .C1(n18249), .C2(n18679), .A(n18164), .B(n18254), .ZN(
        n18182) );
  AND2_X1 U21298 ( .A1(n18451), .A2(n18209), .ZN(n18180) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18182), .B1(
        n18452), .B2(n18180), .ZN(n18166) );
  AOI22_X1 U21300 ( .A1(n18181), .A2(n18458), .B1(n18397), .B2(n18249), .ZN(
        n18165) );
  OAI211_X1 U21301 ( .C1(n18175), .C2(n18400), .A(n18166), .B(n18165), .ZN(
        P3_U2892) );
  AOI22_X1 U21302 ( .A1(n18181), .A2(n18463), .B1(n18462), .B2(n18180), .ZN(
        n18168) );
  INV_X1 U21303 ( .A(n18175), .ZN(n18204) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18182), .B1(
        n18204), .B2(n18464), .ZN(n18167) );
  OAI211_X1 U21305 ( .C1(n18467), .C2(n18185), .A(n18168), .B(n18167), .ZN(
        P3_U2893) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18182), .B1(
        n18468), .B2(n18180), .ZN(n18170) );
  AOI22_X1 U21307 ( .A1(n18181), .A2(n18470), .B1(n18283), .B2(n18249), .ZN(
        n18169) );
  OAI211_X1 U21308 ( .C1(n18175), .C2(n18286), .A(n18170), .B(n18169), .ZN(
        P3_U2894) );
  AOI22_X1 U21309 ( .A1(n18204), .A2(n18475), .B1(n18474), .B2(n18180), .ZN(
        n18172) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18182), .B1(
        n18181), .B2(n18476), .ZN(n18171) );
  OAI211_X1 U21311 ( .C1(n18479), .C2(n18185), .A(n18172), .B(n18171), .ZN(
        P3_U2895) );
  AOI22_X1 U21312 ( .A1(n18181), .A2(n18482), .B1(n18480), .B2(n18180), .ZN(
        n18174) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18182), .B1(
        n18409), .B2(n18249), .ZN(n18173) );
  OAI211_X1 U21314 ( .C1(n18175), .C2(n18413), .A(n18174), .B(n18173), .ZN(
        P3_U2896) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18182), .B1(
        n18487), .B2(n18180), .ZN(n18177) );
  AOI22_X1 U21316 ( .A1(n18204), .A2(n18486), .B1(n18181), .B2(n18488), .ZN(
        n18176) );
  OAI211_X1 U21317 ( .C1(n18491), .C2(n18185), .A(n18177), .B(n18176), .ZN(
        P3_U2897) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18182), .B1(
        n18492), .B2(n18180), .ZN(n18179) );
  AOI22_X1 U21319 ( .A1(n18204), .A2(n18494), .B1(n18181), .B2(n18493), .ZN(
        n18178) );
  OAI211_X1 U21320 ( .C1(n18497), .C2(n18185), .A(n18179), .B(n18178), .ZN(
        P3_U2898) );
  AOI22_X1 U21321 ( .A1(n18204), .A2(n18503), .B1(n18499), .B2(n18180), .ZN(
        n18184) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18182), .B1(
        n18181), .B2(n18501), .ZN(n18183) );
  OAI211_X1 U21323 ( .C1(n18507), .C2(n18185), .A(n18184), .B(n18183), .ZN(
        P3_U2899) );
  NAND2_X1 U21324 ( .A1(n18544), .A2(n18255), .ZN(n18239) );
  INV_X1 U21325 ( .A(n18239), .ZN(n18272) );
  NOR2_X1 U21326 ( .A1(n18272), .A2(n18249), .ZN(n18231) );
  NOR2_X1 U21327 ( .A1(n18571), .A2(n18231), .ZN(n18203) );
  AOI22_X1 U21328 ( .A1(n18204), .A2(n18458), .B1(n18452), .B2(n18203), .ZN(
        n18189) );
  NOR2_X1 U21329 ( .A1(n18225), .A2(n18204), .ZN(n18186) );
  OAI21_X1 U21330 ( .B1(n18186), .B2(n18324), .A(n18231), .ZN(n18187) );
  OAI211_X1 U21331 ( .C1(n18272), .C2(n18679), .A(n18374), .B(n18187), .ZN(
        n18205) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18205), .B1(
        n18397), .B2(n18272), .ZN(n18188) );
  OAI211_X1 U21333 ( .C1(n18194), .C2(n18400), .A(n18189), .B(n18188), .ZN(
        P3_U2900) );
  AOI22_X1 U21334 ( .A1(n18225), .A2(n18464), .B1(n18462), .B2(n18203), .ZN(
        n18191) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18205), .B1(
        n18204), .B2(n18463), .ZN(n18190) );
  OAI211_X1 U21336 ( .C1(n18467), .C2(n18239), .A(n18191), .B(n18190), .ZN(
        P3_U2901) );
  AOI22_X1 U21337 ( .A1(n18204), .A2(n18470), .B1(n18468), .B2(n18203), .ZN(
        n18193) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18205), .B1(
        n18283), .B2(n18272), .ZN(n18192) );
  OAI211_X1 U21339 ( .C1(n18194), .C2(n18286), .A(n18193), .B(n18192), .ZN(
        P3_U2902) );
  AOI22_X1 U21340 ( .A1(n18225), .A2(n18475), .B1(n18474), .B2(n18203), .ZN(
        n18196) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18205), .B1(
        n18204), .B2(n18476), .ZN(n18195) );
  OAI211_X1 U21342 ( .C1(n18479), .C2(n18239), .A(n18196), .B(n18195), .ZN(
        P3_U2903) );
  AOI22_X1 U21343 ( .A1(n18225), .A2(n18481), .B1(n18480), .B2(n18203), .ZN(
        n18198) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18205), .B1(
        n18204), .B2(n18482), .ZN(n18197) );
  OAI211_X1 U21345 ( .C1(n18485), .C2(n18239), .A(n18198), .B(n18197), .ZN(
        P3_U2904) );
  AOI22_X1 U21346 ( .A1(n18225), .A2(n18486), .B1(n18487), .B2(n18203), .ZN(
        n18200) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18205), .B1(
        n18204), .B2(n18488), .ZN(n18199) );
  OAI211_X1 U21348 ( .C1(n18491), .C2(n18239), .A(n18200), .B(n18199), .ZN(
        P3_U2905) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18205), .B1(
        n18492), .B2(n18203), .ZN(n18202) );
  AOI22_X1 U21350 ( .A1(n18225), .A2(n18494), .B1(n18204), .B2(n18493), .ZN(
        n18201) );
  OAI211_X1 U21351 ( .C1(n18497), .C2(n18239), .A(n18202), .B(n18201), .ZN(
        P3_U2906) );
  AOI22_X1 U21352 ( .A1(n18225), .A2(n18503), .B1(n18499), .B2(n18203), .ZN(
        n18207) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18205), .B1(
        n18204), .B2(n18501), .ZN(n18206) );
  OAI211_X1 U21354 ( .C1(n18507), .C2(n18239), .A(n18207), .B(n18206), .ZN(
        P3_U2907) );
  NAND2_X1 U21355 ( .A1(n18301), .A2(n18255), .ZN(n18266) );
  NOR2_X1 U21356 ( .A1(n18229), .A2(n18302), .ZN(n18224) );
  AOI22_X1 U21357 ( .A1(n18453), .A2(n18249), .B1(n18452), .B2(n18224), .ZN(
        n18211) );
  AOI22_X1 U21358 ( .A1(n18457), .A2(n18209), .B1(n18255), .B2(n18208), .ZN(
        n18226) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18226), .B1(
        n18225), .B2(n18458), .ZN(n18210) );
  OAI211_X1 U21360 ( .C1(n18461), .C2(n18266), .A(n18211), .B(n18210), .ZN(
        P3_U2908) );
  AOI22_X1 U21361 ( .A1(n18464), .A2(n18249), .B1(n18462), .B2(n18224), .ZN(
        n18213) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18226), .B1(
        n18225), .B2(n18463), .ZN(n18212) );
  OAI211_X1 U21363 ( .C1(n18467), .C2(n18266), .A(n18213), .B(n18212), .ZN(
        P3_U2909) );
  AOI22_X1 U21364 ( .A1(n18225), .A2(n18470), .B1(n18468), .B2(n18224), .ZN(
        n18215) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18226), .B1(
        n18469), .B2(n18249), .ZN(n18214) );
  OAI211_X1 U21366 ( .C1(n18473), .C2(n18266), .A(n18215), .B(n18214), .ZN(
        P3_U2910) );
  AOI22_X1 U21367 ( .A1(n18475), .A2(n18249), .B1(n18474), .B2(n18224), .ZN(
        n18217) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18226), .B1(
        n18225), .B2(n18476), .ZN(n18216) );
  OAI211_X1 U21369 ( .C1(n18479), .C2(n18266), .A(n18217), .B(n18216), .ZN(
        P3_U2911) );
  AOI22_X1 U21370 ( .A1(n18225), .A2(n18482), .B1(n18480), .B2(n18224), .ZN(
        n18219) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18226), .B1(
        n18481), .B2(n18249), .ZN(n18218) );
  OAI211_X1 U21372 ( .C1(n18485), .C2(n18266), .A(n18219), .B(n18218), .ZN(
        P3_U2912) );
  AOI22_X1 U21373 ( .A1(n18487), .A2(n18224), .B1(n18486), .B2(n18249), .ZN(
        n18221) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18226), .B1(
        n18225), .B2(n18488), .ZN(n18220) );
  OAI211_X1 U21375 ( .C1(n18491), .C2(n18266), .A(n18221), .B(n18220), .ZN(
        P3_U2913) );
  AOI22_X1 U21376 ( .A1(n18225), .A2(n18493), .B1(n18492), .B2(n18224), .ZN(
        n18223) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18226), .B1(
        n18494), .B2(n18249), .ZN(n18222) );
  OAI211_X1 U21378 ( .C1(n18497), .C2(n18266), .A(n18223), .B(n18222), .ZN(
        P3_U2914) );
  AOI22_X1 U21379 ( .A1(n18499), .A2(n18224), .B1(n18503), .B2(n18249), .ZN(
        n18228) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18226), .B1(
        n18225), .B2(n18501), .ZN(n18227) );
  OAI211_X1 U21381 ( .C1(n18507), .C2(n18266), .A(n18228), .B(n18227), .ZN(
        P3_U2915) );
  NOR2_X2 U21382 ( .A1(n18230), .A2(n18229), .ZN(n18319) );
  AOI21_X1 U21383 ( .B1(n18291), .B2(n18266), .A(n18571), .ZN(n18248) );
  AOI22_X1 U21384 ( .A1(n18452), .A2(n18248), .B1(n18458), .B2(n18249), .ZN(
        n18234) );
  AOI221_X1 U21385 ( .B1(n18231), .B2(n18266), .C1(n18324), .C2(n18266), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18232) );
  OAI21_X1 U21386 ( .B1(n18319), .B2(n18232), .A(n18374), .ZN(n18250) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18250), .B1(
        n18397), .B2(n18319), .ZN(n18233) );
  OAI211_X1 U21388 ( .C1(n18400), .C2(n18239), .A(n18234), .B(n18233), .ZN(
        P3_U2916) );
  AOI22_X1 U21389 ( .A1(n18463), .A2(n18249), .B1(n18462), .B2(n18248), .ZN(
        n18236) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18250), .B1(
        n18464), .B2(n18272), .ZN(n18235) );
  OAI211_X1 U21391 ( .C1(n18467), .C2(n18291), .A(n18236), .B(n18235), .ZN(
        P3_U2917) );
  AOI22_X1 U21392 ( .A1(n18468), .A2(n18248), .B1(n18470), .B2(n18249), .ZN(
        n18238) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18250), .B1(
        n18283), .B2(n18319), .ZN(n18237) );
  OAI211_X1 U21394 ( .C1(n18286), .C2(n18239), .A(n18238), .B(n18237), .ZN(
        P3_U2918) );
  AOI22_X1 U21395 ( .A1(n18475), .A2(n18272), .B1(n18474), .B2(n18248), .ZN(
        n18241) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18250), .B1(
        n18476), .B2(n18249), .ZN(n18240) );
  OAI211_X1 U21397 ( .C1(n18479), .C2(n18291), .A(n18241), .B(n18240), .ZN(
        P3_U2919) );
  AOI22_X1 U21398 ( .A1(n18481), .A2(n18272), .B1(n18480), .B2(n18248), .ZN(
        n18243) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18250), .B1(
        n18482), .B2(n18249), .ZN(n18242) );
  OAI211_X1 U21400 ( .C1(n18485), .C2(n18291), .A(n18243), .B(n18242), .ZN(
        P3_U2920) );
  AOI22_X1 U21401 ( .A1(n18488), .A2(n18249), .B1(n18487), .B2(n18248), .ZN(
        n18245) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18250), .B1(
        n18486), .B2(n18272), .ZN(n18244) );
  OAI211_X1 U21403 ( .C1(n18491), .C2(n18291), .A(n18245), .B(n18244), .ZN(
        P3_U2921) );
  AOI22_X1 U21404 ( .A1(n18493), .A2(n18249), .B1(n18492), .B2(n18248), .ZN(
        n18247) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18250), .B1(
        n18494), .B2(n18272), .ZN(n18246) );
  OAI211_X1 U21406 ( .C1(n18497), .C2(n18291), .A(n18247), .B(n18246), .ZN(
        P3_U2922) );
  AOI22_X1 U21407 ( .A1(n18501), .A2(n18249), .B1(n18499), .B2(n18248), .ZN(
        n18252) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18250), .B1(
        n18503), .B2(n18272), .ZN(n18251) );
  OAI211_X1 U21409 ( .C1(n18507), .C2(n18291), .A(n18252), .B(n18251), .ZN(
        P3_U2923) );
  NOR2_X1 U21410 ( .A1(n18253), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18303) );
  NAND2_X1 U21411 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18303), .ZN(
        n18276) );
  AND2_X1 U21412 ( .A1(n18451), .A2(n18303), .ZN(n18271) );
  AOI22_X1 U21413 ( .A1(n18453), .A2(n18298), .B1(n18452), .B2(n18271), .ZN(
        n18257) );
  OAI211_X1 U21414 ( .C1(n18343), .C2(n18679), .A(n18255), .B(n18254), .ZN(
        n18273) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18273), .B1(
        n18458), .B2(n18272), .ZN(n18256) );
  OAI211_X1 U21416 ( .C1(n18461), .C2(n18276), .A(n18257), .B(n18256), .ZN(
        P3_U2924) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18273), .B1(
        n18462), .B2(n18271), .ZN(n18259) );
  AOI22_X1 U21418 ( .A1(n18463), .A2(n18272), .B1(n18464), .B2(n18298), .ZN(
        n18258) );
  OAI211_X1 U21419 ( .C1(n18467), .C2(n18276), .A(n18259), .B(n18258), .ZN(
        P3_U2925) );
  AOI22_X1 U21420 ( .A1(n18469), .A2(n18298), .B1(n18468), .B2(n18271), .ZN(
        n18261) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18273), .B1(
        n18470), .B2(n18272), .ZN(n18260) );
  OAI211_X1 U21422 ( .C1(n18473), .C2(n18276), .A(n18261), .B(n18260), .ZN(
        P3_U2926) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18273), .B1(
        n18474), .B2(n18271), .ZN(n18263) );
  AOI22_X1 U21424 ( .A1(n18405), .A2(n18343), .B1(n18476), .B2(n18272), .ZN(
        n18262) );
  OAI211_X1 U21425 ( .C1(n18408), .C2(n18266), .A(n18263), .B(n18262), .ZN(
        P3_U2927) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18273), .B1(
        n18480), .B2(n18271), .ZN(n18265) );
  AOI22_X1 U21427 ( .A1(n18409), .A2(n18343), .B1(n18482), .B2(n18272), .ZN(
        n18264) );
  OAI211_X1 U21428 ( .C1(n18413), .C2(n18266), .A(n18265), .B(n18264), .ZN(
        P3_U2928) );
  AOI22_X1 U21429 ( .A1(n18487), .A2(n18271), .B1(n18486), .B2(n18298), .ZN(
        n18268) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18273), .B1(
        n18488), .B2(n18272), .ZN(n18267) );
  OAI211_X1 U21431 ( .C1(n18491), .C2(n18276), .A(n18268), .B(n18267), .ZN(
        P3_U2929) );
  AOI22_X1 U21432 ( .A1(n18494), .A2(n18298), .B1(n18492), .B2(n18271), .ZN(
        n18270) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18273), .B1(
        n18493), .B2(n18272), .ZN(n18269) );
  OAI211_X1 U21434 ( .C1(n18497), .C2(n18276), .A(n18270), .B(n18269), .ZN(
        P3_U2930) );
  AOI22_X1 U21435 ( .A1(n18499), .A2(n18271), .B1(n18503), .B2(n18298), .ZN(
        n18275) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18273), .B1(
        n18501), .B2(n18272), .ZN(n18274) );
  OAI211_X1 U21437 ( .C1(n18507), .C2(n18276), .A(n18275), .B(n18274), .ZN(
        P3_U2931) );
  NAND2_X1 U21438 ( .A1(n18544), .A2(n18369), .ZN(n18335) );
  NOR2_X1 U21439 ( .A1(n18319), .A2(n18298), .ZN(n18277) );
  NOR2_X1 U21440 ( .A1(n18365), .A2(n18343), .ZN(n18325) );
  OAI21_X1 U21441 ( .B1(n18277), .B2(n18324), .A(n18325), .ZN(n18278) );
  OAI211_X1 U21442 ( .C1(n18365), .C2(n18679), .A(n18374), .B(n18278), .ZN(
        n18297) );
  NOR2_X1 U21443 ( .A1(n18571), .A2(n18325), .ZN(n18296) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18297), .B1(
        n18452), .B2(n18296), .ZN(n18280) );
  AOI22_X1 U21445 ( .A1(n18397), .A2(n18365), .B1(n18458), .B2(n18298), .ZN(
        n18279) );
  OAI211_X1 U21446 ( .C1(n18400), .C2(n18291), .A(n18280), .B(n18279), .ZN(
        P3_U2932) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18297), .B1(
        n18462), .B2(n18296), .ZN(n18282) );
  AOI22_X1 U21448 ( .A1(n18463), .A2(n18298), .B1(n18464), .B2(n18319), .ZN(
        n18281) );
  OAI211_X1 U21449 ( .C1(n18467), .C2(n18335), .A(n18282), .B(n18281), .ZN(
        P3_U2933) );
  AOI22_X1 U21450 ( .A1(n18468), .A2(n18296), .B1(n18470), .B2(n18298), .ZN(
        n18285) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18297), .B1(
        n18283), .B2(n18365), .ZN(n18284) );
  OAI211_X1 U21452 ( .C1(n18286), .C2(n18291), .A(n18285), .B(n18284), .ZN(
        P3_U2934) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18297), .B1(
        n18474), .B2(n18296), .ZN(n18288) );
  AOI22_X1 U21454 ( .A1(n18405), .A2(n18365), .B1(n18476), .B2(n18298), .ZN(
        n18287) );
  OAI211_X1 U21455 ( .C1(n18408), .C2(n18291), .A(n18288), .B(n18287), .ZN(
        P3_U2935) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18297), .B1(
        n18480), .B2(n18296), .ZN(n18290) );
  AOI22_X1 U21457 ( .A1(n18409), .A2(n18365), .B1(n18482), .B2(n18298), .ZN(
        n18289) );
  OAI211_X1 U21458 ( .C1(n18413), .C2(n18291), .A(n18290), .B(n18289), .ZN(
        P3_U2936) );
  AOI22_X1 U21459 ( .A1(n18487), .A2(n18296), .B1(n18486), .B2(n18319), .ZN(
        n18293) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18297), .B1(
        n18488), .B2(n18298), .ZN(n18292) );
  OAI211_X1 U21461 ( .C1(n18491), .C2(n18335), .A(n18293), .B(n18292), .ZN(
        P3_U2937) );
  AOI22_X1 U21462 ( .A1(n18494), .A2(n18319), .B1(n18492), .B2(n18296), .ZN(
        n18295) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18297), .B1(
        n18493), .B2(n18298), .ZN(n18294) );
  OAI211_X1 U21464 ( .C1(n18497), .C2(n18335), .A(n18295), .B(n18294), .ZN(
        P3_U2938) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18297), .B1(
        n18499), .B2(n18296), .ZN(n18300) );
  AOI22_X1 U21466 ( .A1(n18501), .A2(n18298), .B1(n18503), .B2(n18319), .ZN(
        n18299) );
  OAI211_X1 U21467 ( .C1(n18507), .C2(n18335), .A(n18300), .B(n18299), .ZN(
        P3_U2939) );
  NAND2_X1 U21468 ( .A1(n18301), .A2(n18369), .ZN(n18348) );
  NOR2_X1 U21469 ( .A1(n18347), .A2(n18302), .ZN(n18318) );
  AOI22_X1 U21470 ( .A1(n18453), .A2(n18343), .B1(n18452), .B2(n18318), .ZN(
        n18305) );
  NOR2_X1 U21471 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18347), .ZN(
        n18349) );
  AOI22_X1 U21472 ( .A1(n18457), .A2(n18303), .B1(n18454), .B2(n18349), .ZN(
        n18320) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18320), .B1(
        n18458), .B2(n18319), .ZN(n18304) );
  OAI211_X1 U21474 ( .C1(n18461), .C2(n18348), .A(n18305), .B(n18304), .ZN(
        P3_U2940) );
  AOI22_X1 U21475 ( .A1(n18464), .A2(n18343), .B1(n18462), .B2(n18318), .ZN(
        n18307) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18320), .B1(
        n18463), .B2(n18319), .ZN(n18306) );
  OAI211_X1 U21477 ( .C1(n18467), .C2(n18348), .A(n18307), .B(n18306), .ZN(
        P3_U2941) );
  AOI22_X1 U21478 ( .A1(n18468), .A2(n18318), .B1(n18470), .B2(n18319), .ZN(
        n18309) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18320), .B1(
        n18469), .B2(n18343), .ZN(n18308) );
  OAI211_X1 U21480 ( .C1(n18473), .C2(n18348), .A(n18309), .B(n18308), .ZN(
        P3_U2942) );
  AOI22_X1 U21481 ( .A1(n18476), .A2(n18319), .B1(n18474), .B2(n18318), .ZN(
        n18311) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18320), .B1(
        n18475), .B2(n18343), .ZN(n18310) );
  OAI211_X1 U21483 ( .C1(n18479), .C2(n18348), .A(n18311), .B(n18310), .ZN(
        P3_U2943) );
  AOI22_X1 U21484 ( .A1(n18481), .A2(n18343), .B1(n18480), .B2(n18318), .ZN(
        n18313) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18320), .B1(
        n18482), .B2(n18319), .ZN(n18312) );
  OAI211_X1 U21486 ( .C1(n18485), .C2(n18348), .A(n18313), .B(n18312), .ZN(
        P3_U2944) );
  AOI22_X1 U21487 ( .A1(n18488), .A2(n18319), .B1(n18487), .B2(n18318), .ZN(
        n18315) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18320), .B1(
        n18486), .B2(n18343), .ZN(n18314) );
  OAI211_X1 U21489 ( .C1(n18491), .C2(n18348), .A(n18315), .B(n18314), .ZN(
        P3_U2945) );
  AOI22_X1 U21490 ( .A1(n18493), .A2(n18319), .B1(n18492), .B2(n18318), .ZN(
        n18317) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18320), .B1(
        n18494), .B2(n18343), .ZN(n18316) );
  OAI211_X1 U21492 ( .C1(n18497), .C2(n18348), .A(n18317), .B(n18316), .ZN(
        P3_U2946) );
  AOI22_X1 U21493 ( .A1(n18499), .A2(n18318), .B1(n18503), .B2(n18343), .ZN(
        n18322) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18320), .B1(
        n18501), .B2(n18319), .ZN(n18321) );
  OAI211_X1 U21495 ( .C1(n18507), .C2(n18348), .A(n18322), .B(n18321), .ZN(
        P3_U2947) );
  AOI22_X1 U21496 ( .A1(n18452), .A2(n18342), .B1(n18458), .B2(n18343), .ZN(
        n18328) );
  NAND2_X1 U21497 ( .A1(n18323), .A2(n18369), .ZN(n18383) );
  AOI221_X1 U21498 ( .B1(n18325), .B2(n18348), .C1(n18324), .C2(n18348), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18326) );
  OAI21_X1 U21499 ( .B1(n18419), .B2(n18326), .A(n18374), .ZN(n18344) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18344), .B1(
        n18397), .B2(n18419), .ZN(n18327) );
  OAI211_X1 U21501 ( .C1(n18400), .C2(n18335), .A(n18328), .B(n18327), .ZN(
        P3_U2948) );
  AOI22_X1 U21502 ( .A1(n18464), .A2(n18365), .B1(n18462), .B2(n18342), .ZN(
        n18330) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18344), .B1(
        n18463), .B2(n18343), .ZN(n18329) );
  OAI211_X1 U21504 ( .C1(n18467), .C2(n18383), .A(n18330), .B(n18329), .ZN(
        P3_U2949) );
  AOI22_X1 U21505 ( .A1(n18469), .A2(n18365), .B1(n18468), .B2(n18342), .ZN(
        n18332) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18344), .B1(
        n18470), .B2(n18343), .ZN(n18331) );
  OAI211_X1 U21507 ( .C1(n18473), .C2(n18383), .A(n18332), .B(n18331), .ZN(
        P3_U2950) );
  AOI22_X1 U21508 ( .A1(n18476), .A2(n18343), .B1(n18474), .B2(n18342), .ZN(
        n18334) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18344), .B1(
        n18405), .B2(n18419), .ZN(n18333) );
  OAI211_X1 U21510 ( .C1(n18408), .C2(n18335), .A(n18334), .B(n18333), .ZN(
        P3_U2951) );
  AOI22_X1 U21511 ( .A1(n18481), .A2(n18365), .B1(n18480), .B2(n18342), .ZN(
        n18337) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18344), .B1(
        n18482), .B2(n18343), .ZN(n18336) );
  OAI211_X1 U21513 ( .C1(n18485), .C2(n18383), .A(n18337), .B(n18336), .ZN(
        P3_U2952) );
  AOI22_X1 U21514 ( .A1(n18488), .A2(n18343), .B1(n18487), .B2(n18342), .ZN(
        n18339) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18344), .B1(
        n18486), .B2(n18365), .ZN(n18338) );
  OAI211_X1 U21516 ( .C1(n18491), .C2(n18383), .A(n18339), .B(n18338), .ZN(
        P3_U2953) );
  AOI22_X1 U21517 ( .A1(n18493), .A2(n18343), .B1(n18492), .B2(n18342), .ZN(
        n18341) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18344), .B1(
        n18494), .B2(n18365), .ZN(n18340) );
  OAI211_X1 U21519 ( .C1(n18497), .C2(n18383), .A(n18341), .B(n18340), .ZN(
        P3_U2954) );
  AOI22_X1 U21520 ( .A1(n18501), .A2(n18343), .B1(n18499), .B2(n18342), .ZN(
        n18346) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18344), .B1(
        n18503), .B2(n18365), .ZN(n18345) );
  OAI211_X1 U21522 ( .C1(n18507), .C2(n18383), .A(n18346), .B(n18345), .ZN(
        P3_U2955) );
  NOR2_X1 U21523 ( .A1(n18541), .A2(n18347), .ZN(n18396) );
  NAND2_X1 U21524 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18396), .ZN(
        n18412) );
  INV_X1 U21525 ( .A(n18348), .ZN(n18391) );
  AND2_X1 U21526 ( .A1(n18451), .A2(n18396), .ZN(n18364) );
  AOI22_X1 U21527 ( .A1(n18453), .A2(n18391), .B1(n18452), .B2(n18364), .ZN(
        n18351) );
  AOI22_X1 U21528 ( .A1(n18457), .A2(n18349), .B1(n18454), .B2(n18396), .ZN(
        n18366) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18366), .B1(
        n18458), .B2(n18365), .ZN(n18350) );
  OAI211_X1 U21530 ( .C1(n18461), .C2(n18412), .A(n18351), .B(n18350), .ZN(
        P3_U2956) );
  AOI22_X1 U21531 ( .A1(n18464), .A2(n18391), .B1(n18462), .B2(n18364), .ZN(
        n18353) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18366), .B1(
        n18463), .B2(n18365), .ZN(n18352) );
  OAI211_X1 U21533 ( .C1(n18467), .C2(n18412), .A(n18353), .B(n18352), .ZN(
        P3_U2957) );
  AOI22_X1 U21534 ( .A1(n18468), .A2(n18364), .B1(n18470), .B2(n18365), .ZN(
        n18355) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18366), .B1(
        n18469), .B2(n18391), .ZN(n18354) );
  OAI211_X1 U21536 ( .C1(n18473), .C2(n18412), .A(n18355), .B(n18354), .ZN(
        P3_U2958) );
  AOI22_X1 U21537 ( .A1(n18475), .A2(n18391), .B1(n18474), .B2(n18364), .ZN(
        n18357) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18366), .B1(
        n18476), .B2(n18365), .ZN(n18356) );
  OAI211_X1 U21539 ( .C1(n18479), .C2(n18412), .A(n18357), .B(n18356), .ZN(
        P3_U2959) );
  AOI22_X1 U21540 ( .A1(n18481), .A2(n18391), .B1(n18480), .B2(n18364), .ZN(
        n18359) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18366), .B1(
        n18482), .B2(n18365), .ZN(n18358) );
  OAI211_X1 U21542 ( .C1(n18485), .C2(n18412), .A(n18359), .B(n18358), .ZN(
        P3_U2960) );
  AOI22_X1 U21543 ( .A1(n18488), .A2(n18365), .B1(n18487), .B2(n18364), .ZN(
        n18361) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18366), .B1(
        n18486), .B2(n18391), .ZN(n18360) );
  OAI211_X1 U21545 ( .C1(n18491), .C2(n18412), .A(n18361), .B(n18360), .ZN(
        P3_U2961) );
  AOI22_X1 U21546 ( .A1(n18493), .A2(n18365), .B1(n18492), .B2(n18364), .ZN(
        n18363) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18366), .B1(
        n18494), .B2(n18391), .ZN(n18362) );
  OAI211_X1 U21548 ( .C1(n18497), .C2(n18412), .A(n18363), .B(n18362), .ZN(
        P3_U2962) );
  AOI22_X1 U21549 ( .A1(n18501), .A2(n18365), .B1(n18499), .B2(n18364), .ZN(
        n18368) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18366), .B1(
        n18503), .B2(n18391), .ZN(n18367) );
  OAI211_X1 U21551 ( .C1(n18507), .C2(n18412), .A(n18368), .B(n18367), .ZN(
        P3_U2963) );
  NAND2_X1 U21552 ( .A1(n18540), .A2(n18456), .ZN(n18395) );
  INV_X1 U21553 ( .A(n18395), .ZN(n18500) );
  NAND2_X1 U21554 ( .A1(n18370), .A2(n18369), .ZN(n18371) );
  NOR2_X1 U21555 ( .A1(n18446), .A2(n18500), .ZN(n18428) );
  OAI21_X1 U21556 ( .B1(n18372), .B2(n18371), .A(n18428), .ZN(n18373) );
  OAI211_X1 U21557 ( .C1(n18500), .C2(n18679), .A(n18374), .B(n18373), .ZN(
        n18392) );
  NOR2_X1 U21558 ( .A1(n18571), .A2(n18428), .ZN(n18390) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18392), .B1(
        n18452), .B2(n18390), .ZN(n18376) );
  AOI22_X1 U21560 ( .A1(n18397), .A2(n18500), .B1(n18458), .B2(n18391), .ZN(
        n18375) );
  OAI211_X1 U21561 ( .C1(n18400), .C2(n18383), .A(n18376), .B(n18375), .ZN(
        P3_U2964) );
  AOI22_X1 U21562 ( .A1(n18464), .A2(n18419), .B1(n18462), .B2(n18390), .ZN(
        n18378) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18392), .B1(
        n18463), .B2(n18391), .ZN(n18377) );
  OAI211_X1 U21564 ( .C1(n18467), .C2(n18395), .A(n18378), .B(n18377), .ZN(
        P3_U2965) );
  AOI22_X1 U21565 ( .A1(n18469), .A2(n18419), .B1(n18468), .B2(n18390), .ZN(
        n18380) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18392), .B1(
        n18470), .B2(n18391), .ZN(n18379) );
  OAI211_X1 U21567 ( .C1(n18473), .C2(n18395), .A(n18380), .B(n18379), .ZN(
        P3_U2966) );
  AOI22_X1 U21568 ( .A1(n18476), .A2(n18391), .B1(n18474), .B2(n18390), .ZN(
        n18382) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18392), .B1(
        n18405), .B2(n18500), .ZN(n18381) );
  OAI211_X1 U21570 ( .C1(n18408), .C2(n18383), .A(n18382), .B(n18381), .ZN(
        P3_U2967) );
  AOI22_X1 U21571 ( .A1(n18481), .A2(n18419), .B1(n18480), .B2(n18390), .ZN(
        n18385) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18392), .B1(
        n18482), .B2(n18391), .ZN(n18384) );
  OAI211_X1 U21573 ( .C1(n18485), .C2(n18395), .A(n18385), .B(n18384), .ZN(
        P3_U2968) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18392), .B1(
        n18487), .B2(n18390), .ZN(n18387) );
  AOI22_X1 U21575 ( .A1(n18488), .A2(n18391), .B1(n18486), .B2(n18419), .ZN(
        n18386) );
  OAI211_X1 U21576 ( .C1(n18491), .C2(n18395), .A(n18387), .B(n18386), .ZN(
        P3_U2969) );
  AOI22_X1 U21577 ( .A1(n18493), .A2(n18391), .B1(n18492), .B2(n18390), .ZN(
        n18389) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18392), .B1(
        n18494), .B2(n18419), .ZN(n18388) );
  OAI211_X1 U21579 ( .C1(n18497), .C2(n18395), .A(n18389), .B(n18388), .ZN(
        P3_U2970) );
  AOI22_X1 U21580 ( .A1(n18499), .A2(n18390), .B1(n18503), .B2(n18419), .ZN(
        n18394) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18392), .B1(
        n18501), .B2(n18391), .ZN(n18393) );
  OAI211_X1 U21582 ( .C1(n18507), .C2(n18395), .A(n18394), .B(n18393), .ZN(
        P3_U2971) );
  AND2_X1 U21583 ( .A1(n18451), .A2(n18456), .ZN(n18418) );
  AOI22_X1 U21584 ( .A1(n18452), .A2(n18418), .B1(n18458), .B2(n18419), .ZN(
        n18399) );
  AOI22_X1 U21585 ( .A1(n18457), .A2(n18396), .B1(n18456), .B2(n18454), .ZN(
        n18420) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18420), .B1(
        n18397), .B2(n18502), .ZN(n18398) );
  OAI211_X1 U21587 ( .C1(n18400), .C2(n18412), .A(n18399), .B(n18398), .ZN(
        P3_U2972) );
  AOI22_X1 U21588 ( .A1(n18464), .A2(n18446), .B1(n18462), .B2(n18418), .ZN(
        n18402) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18420), .B1(
        n18463), .B2(n18419), .ZN(n18401) );
  OAI211_X1 U21590 ( .C1(n18467), .C2(n18423), .A(n18402), .B(n18401), .ZN(
        P3_U2973) );
  AOI22_X1 U21591 ( .A1(n18469), .A2(n18446), .B1(n18468), .B2(n18418), .ZN(
        n18404) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18420), .B1(
        n18470), .B2(n18419), .ZN(n18403) );
  OAI211_X1 U21593 ( .C1(n18473), .C2(n18423), .A(n18404), .B(n18403), .ZN(
        P3_U2974) );
  AOI22_X1 U21594 ( .A1(n18476), .A2(n18419), .B1(n18474), .B2(n18418), .ZN(
        n18407) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18420), .B1(
        n18405), .B2(n18502), .ZN(n18406) );
  OAI211_X1 U21596 ( .C1(n18408), .C2(n18412), .A(n18407), .B(n18406), .ZN(
        P3_U2975) );
  AOI22_X1 U21597 ( .A1(n18480), .A2(n18418), .B1(n18482), .B2(n18419), .ZN(
        n18411) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18420), .B1(
        n18409), .B2(n18502), .ZN(n18410) );
  OAI211_X1 U21599 ( .C1(n18413), .C2(n18412), .A(n18411), .B(n18410), .ZN(
        P3_U2976) );
  AOI22_X1 U21600 ( .A1(n18488), .A2(n18419), .B1(n18487), .B2(n18418), .ZN(
        n18415) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18420), .B1(
        n18486), .B2(n18446), .ZN(n18414) );
  OAI211_X1 U21602 ( .C1(n18491), .C2(n18423), .A(n18415), .B(n18414), .ZN(
        P3_U2977) );
  AOI22_X1 U21603 ( .A1(n18494), .A2(n18446), .B1(n18492), .B2(n18418), .ZN(
        n18417) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18420), .B1(
        n18493), .B2(n18419), .ZN(n18416) );
  OAI211_X1 U21605 ( .C1(n18497), .C2(n18423), .A(n18417), .B(n18416), .ZN(
        P3_U2978) );
  AOI22_X1 U21606 ( .A1(n18501), .A2(n18419), .B1(n18499), .B2(n18418), .ZN(
        n18422) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18420), .B1(
        n18503), .B2(n18446), .ZN(n18421) );
  OAI211_X1 U21608 ( .C1(n18507), .C2(n18423), .A(n18422), .B(n18421), .ZN(
        P3_U2979) );
  INV_X1 U21609 ( .A(n18424), .ZN(n18425) );
  NOR2_X1 U21610 ( .A1(n18571), .A2(n18425), .ZN(n18445) );
  AOI22_X1 U21611 ( .A1(n18453), .A2(n18500), .B1(n18452), .B2(n18445), .ZN(
        n18432) );
  OAI22_X1 U21612 ( .A1(n18428), .A2(n18427), .B1(n18426), .B2(n18425), .ZN(
        n18429) );
  OAI21_X1 U21613 ( .B1(n18430), .B2(n18679), .A(n18429), .ZN(n18447) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18447), .B1(
        n18458), .B2(n18446), .ZN(n18431) );
  OAI211_X1 U21615 ( .C1(n18461), .C2(n18450), .A(n18432), .B(n18431), .ZN(
        P3_U2980) );
  AOI22_X1 U21616 ( .A1(n18464), .A2(n18500), .B1(n18462), .B2(n18445), .ZN(
        n18434) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18447), .B1(
        n18463), .B2(n18446), .ZN(n18433) );
  OAI211_X1 U21618 ( .C1(n18467), .C2(n18450), .A(n18434), .B(n18433), .ZN(
        P3_U2981) );
  AOI22_X1 U21619 ( .A1(n18469), .A2(n18500), .B1(n18468), .B2(n18445), .ZN(
        n18436) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18447), .B1(
        n18470), .B2(n18446), .ZN(n18435) );
  OAI211_X1 U21621 ( .C1(n18473), .C2(n18450), .A(n18436), .B(n18435), .ZN(
        P3_U2982) );
  AOI22_X1 U21622 ( .A1(n18475), .A2(n18500), .B1(n18474), .B2(n18445), .ZN(
        n18438) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18447), .B1(
        n18476), .B2(n18446), .ZN(n18437) );
  OAI211_X1 U21624 ( .C1(n18479), .C2(n18450), .A(n18438), .B(n18437), .ZN(
        P3_U2983) );
  AOI22_X1 U21625 ( .A1(n18481), .A2(n18500), .B1(n18480), .B2(n18445), .ZN(
        n18440) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18447), .B1(
        n18482), .B2(n18446), .ZN(n18439) );
  OAI211_X1 U21627 ( .C1(n18485), .C2(n18450), .A(n18440), .B(n18439), .ZN(
        P3_U2984) );
  AOI22_X1 U21628 ( .A1(n18487), .A2(n18445), .B1(n18486), .B2(n18500), .ZN(
        n18442) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18447), .B1(
        n18488), .B2(n18446), .ZN(n18441) );
  OAI211_X1 U21630 ( .C1(n18491), .C2(n18450), .A(n18442), .B(n18441), .ZN(
        P3_U2985) );
  AOI22_X1 U21631 ( .A1(n18494), .A2(n18500), .B1(n18492), .B2(n18445), .ZN(
        n18444) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18447), .B1(
        n18493), .B2(n18446), .ZN(n18443) );
  OAI211_X1 U21633 ( .C1(n18497), .C2(n18450), .A(n18444), .B(n18443), .ZN(
        P3_U2986) );
  AOI22_X1 U21634 ( .A1(n18499), .A2(n18445), .B1(n18503), .B2(n18500), .ZN(
        n18449) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18447), .B1(
        n18501), .B2(n18446), .ZN(n18448) );
  OAI211_X1 U21636 ( .C1(n18507), .C2(n18450), .A(n18449), .B(n18448), .ZN(
        P3_U2987) );
  AND2_X1 U21637 ( .A1(n18451), .A2(n18455), .ZN(n18498) );
  AOI22_X1 U21638 ( .A1(n18453), .A2(n18502), .B1(n18452), .B2(n18498), .ZN(
        n18460) );
  AOI22_X1 U21639 ( .A1(n18457), .A2(n18456), .B1(n18455), .B2(n18454), .ZN(
        n18504) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18504), .B1(
        n18458), .B2(n18500), .ZN(n18459) );
  OAI211_X1 U21641 ( .C1(n18508), .C2(n18461), .A(n18460), .B(n18459), .ZN(
        P3_U2988) );
  AOI22_X1 U21642 ( .A1(n18463), .A2(n18500), .B1(n18462), .B2(n18498), .ZN(
        n18466) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18504), .B1(
        n18464), .B2(n18502), .ZN(n18465) );
  OAI211_X1 U21644 ( .C1(n18508), .C2(n18467), .A(n18466), .B(n18465), .ZN(
        P3_U2989) );
  AOI22_X1 U21645 ( .A1(n18469), .A2(n18502), .B1(n18468), .B2(n18498), .ZN(
        n18472) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18504), .B1(
        n18470), .B2(n18500), .ZN(n18471) );
  OAI211_X1 U21647 ( .C1(n18508), .C2(n18473), .A(n18472), .B(n18471), .ZN(
        P3_U2990) );
  AOI22_X1 U21648 ( .A1(n18475), .A2(n18502), .B1(n18474), .B2(n18498), .ZN(
        n18478) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18504), .B1(
        n18476), .B2(n18500), .ZN(n18477) );
  OAI211_X1 U21650 ( .C1(n18508), .C2(n18479), .A(n18478), .B(n18477), .ZN(
        P3_U2991) );
  AOI22_X1 U21651 ( .A1(n18481), .A2(n18502), .B1(n18480), .B2(n18498), .ZN(
        n18484) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18504), .B1(
        n18482), .B2(n18500), .ZN(n18483) );
  OAI211_X1 U21653 ( .C1(n18508), .C2(n18485), .A(n18484), .B(n18483), .ZN(
        P3_U2992) );
  AOI22_X1 U21654 ( .A1(n18487), .A2(n18498), .B1(n18486), .B2(n18502), .ZN(
        n18490) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18504), .B1(
        n18488), .B2(n18500), .ZN(n18489) );
  OAI211_X1 U21656 ( .C1(n18508), .C2(n18491), .A(n18490), .B(n18489), .ZN(
        P3_U2993) );
  AOI22_X1 U21657 ( .A1(n18493), .A2(n18500), .B1(n18492), .B2(n18498), .ZN(
        n18496) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18504), .B1(
        n18494), .B2(n18502), .ZN(n18495) );
  OAI211_X1 U21659 ( .C1(n18508), .C2(n18497), .A(n18496), .B(n18495), .ZN(
        P3_U2994) );
  AOI22_X1 U21660 ( .A1(n18501), .A2(n18500), .B1(n18499), .B2(n18498), .ZN(
        n18506) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18504), .B1(
        n18503), .B2(n18502), .ZN(n18505) );
  OAI211_X1 U21662 ( .C1(n18508), .C2(n18507), .A(n18506), .B(n18505), .ZN(
        P3_U2995) );
  NOR2_X1 U21663 ( .A1(n18548), .A2(n18509), .ZN(n18511) );
  OAI222_X1 U21664 ( .A1(n18515), .A2(n18514), .B1(n18513), .B2(n18512), .C1(
        n18511), .C2(n18510), .ZN(n18724) );
  OAI21_X1 U21665 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18516), .ZN(n18517) );
  OAI211_X1 U21666 ( .C1(n18558), .C2(n18572), .A(n18518), .B(n18517), .ZN(
        n18569) );
  OAI21_X1 U21667 ( .B1(n18521), .B2(n18520), .A(n18519), .ZN(n18555) );
  AOI21_X1 U21668 ( .B1(n18702), .B2(n18522), .A(n18555), .ZN(n18534) );
  NAND2_X1 U21669 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18523), .ZN(
        n18533) );
  NAND2_X1 U21670 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18524), .ZN(
        n18525) );
  AOI211_X1 U21671 ( .C1(n18526), .C2(n18525), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18702), .ZN(n18527) );
  AOI21_X1 U21672 ( .B1(n18548), .B2(n18528), .A(n18527), .ZN(n18532) );
  OAI211_X1 U21673 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18530), .B(n18529), .ZN(
        n18531) );
  OAI211_X1 U21674 ( .C1(n18534), .C2(n18533), .A(n18532), .B(n18531), .ZN(
        n18693) );
  AOI22_X1 U21675 ( .A1(n18535), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18693), .B2(n18558), .ZN(n18547) );
  NAND2_X1 U21676 ( .A1(n18537), .A2(n18536), .ZN(n18538) );
  NAND2_X1 U21677 ( .A1(n18552), .A2(n18708), .ZN(n18549) );
  AOI22_X1 U21678 ( .A1(n18699), .A2(n18538), .B1(n18702), .B2(n18549), .ZN(
        n18696) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18539), .B1(
        n18538), .B2(n18708), .ZN(n18542) );
  INV_X1 U21680 ( .A(n18542), .ZN(n18704) );
  NOR3_X1 U21681 ( .A1(n18541), .A2(n18540), .A3(n18704), .ZN(n18543) );
  OAI22_X1 U21682 ( .A1(n18696), .A2(n18543), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18542), .ZN(n18545) );
  AOI21_X1 U21683 ( .B1(n18545), .B2(n18558), .A(n18544), .ZN(n18546) );
  AOI21_X1 U21684 ( .B1(n18547), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n18546), .ZN(n18559) );
  INV_X1 U21685 ( .A(n18547), .ZN(n18560) );
  AOI221_X1 U21686 ( .B1(n18559), .B2(n18563), .C1(n18562), .C2(n18563), .A(
        n18560), .ZN(n18567) );
  AOI22_X1 U21687 ( .A1(n18553), .A2(n18549), .B1(n18548), .B2(n18551), .ZN(
        n18550) );
  NOR2_X1 U21688 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18550), .ZN(
        n18681) );
  OAI21_X1 U21689 ( .B1(n18553), .B2(n18552), .A(n18551), .ZN(n18554) );
  AOI21_X1 U21690 ( .B1(n18556), .B2(n18555), .A(n18554), .ZN(n18682) );
  NAND2_X1 U21691 ( .A1(n18558), .A2(n18682), .ZN(n18557) );
  AOI22_X1 U21692 ( .A1(n18558), .A2(n18681), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18557), .ZN(n18566) );
  AOI21_X1 U21693 ( .B1(n18561), .B2(n18560), .A(n18559), .ZN(n18565) );
  NAND2_X1 U21694 ( .A1(n18563), .A2(n18562), .ZN(n18564) );
  OAI22_X1 U21695 ( .A1(n18567), .A2(n18566), .B1(n18565), .B2(n18564), .ZN(
        n18568) );
  NOR4_X1 U21696 ( .A1(n18570), .A2(n18724), .A3(n18569), .A4(n18568), .ZN(
        n18582) );
  NAND2_X1 U21697 ( .A1(n18688), .A2(n18571), .ZN(n18577) );
  INV_X1 U21698 ( .A(n18577), .ZN(n18573) );
  AOI22_X1 U21699 ( .A1(n18574), .A2(n18599), .B1(n18573), .B2(n18572), .ZN(
        n18579) );
  OAI211_X1 U21700 ( .C1(n18576), .C2(n18575), .A(n18727), .B(n18582), .ZN(
        n18678) );
  NAND2_X1 U21701 ( .A1(n18599), .A2(n18742), .ZN(n18583) );
  NAND4_X1 U21702 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18678), .A3(n18577), 
        .A4(n18583), .ZN(n18587) );
  OAI22_X1 U21703 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18579), .B1(n18578), 
        .B2(n18587), .ZN(n18580) );
  OAI21_X1 U21704 ( .B1(n18582), .B2(n18581), .A(n18580), .ZN(P3_U2996) );
  NOR3_X1 U21705 ( .A1(n18688), .A2(n18584), .A3(n18583), .ZN(n18589) );
  AOI211_X1 U21706 ( .C1(n18599), .C2(n18729), .A(n18585), .B(n18589), .ZN(
        n18586) );
  OAI21_X1 U21707 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18587), .A(n18586), 
        .ZN(P3_U2997) );
  NOR2_X1 U21708 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18735) );
  NOR4_X1 U21709 ( .A1(n18735), .A2(n18590), .A3(n18589), .A4(n18588), .ZN(
        P3_U2998) );
  AND2_X1 U21710 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18591), .ZN(
        P3_U2999) );
  AND2_X1 U21711 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18591), .ZN(
        P3_U3000) );
  AND2_X1 U21712 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18591), .ZN(
        P3_U3001) );
  AND2_X1 U21713 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18591), .ZN(
        P3_U3002) );
  AND2_X1 U21714 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18591), .ZN(
        P3_U3003) );
  AND2_X1 U21715 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18591), .ZN(
        P3_U3004) );
  AND2_X1 U21716 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18591), .ZN(
        P3_U3005) );
  AND2_X1 U21717 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18591), .ZN(
        P3_U3006) );
  AND2_X1 U21718 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18591), .ZN(
        P3_U3007) );
  AND2_X1 U21719 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18591), .ZN(
        P3_U3008) );
  AND2_X1 U21720 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18591), .ZN(
        P3_U3009) );
  AND2_X1 U21721 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18591), .ZN(
        P3_U3010) );
  AND2_X1 U21722 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18591), .ZN(
        P3_U3011) );
  AND2_X1 U21723 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18591), .ZN(
        P3_U3012) );
  AND2_X1 U21724 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18591), .ZN(
        P3_U3013) );
  AND2_X1 U21725 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18591), .ZN(
        P3_U3014) );
  AND2_X1 U21726 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18591), .ZN(
        P3_U3015) );
  AND2_X1 U21727 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18591), .ZN(
        P3_U3016) );
  AND2_X1 U21728 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18591), .ZN(
        P3_U3017) );
  AND2_X1 U21729 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18591), .ZN(
        P3_U3018) );
  AND2_X1 U21730 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18591), .ZN(
        P3_U3019) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18591), .ZN(
        P3_U3020) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18591), .ZN(P3_U3021) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18591), .ZN(P3_U3022) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18591), .ZN(P3_U3023) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18591), .ZN(P3_U3024) );
  INV_X1 U21736 ( .A(P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20807) );
  NOR2_X1 U21737 ( .A1(n20807), .A2(n18676), .ZN(P3_U3025) );
  AND2_X1 U21738 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18591), .ZN(P3_U3026) );
  AND2_X1 U21739 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18591), .ZN(P3_U3027) );
  AND2_X1 U21740 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18591), .ZN(P3_U3028) );
  OAI21_X1 U21741 ( .B1(n18592), .B2(n20660), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18593) );
  AOI22_X1 U21742 ( .A1(n18607), .A2(n18609), .B1(n18740), .B2(n18593), .ZN(
        n18595) );
  INV_X1 U21743 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18594) );
  NAND3_X1 U21744 ( .A1(NA), .A2(n18607), .A3(n18594), .ZN(n18602) );
  OAI211_X1 U21745 ( .C1(n18733), .C2(n18596), .A(n18595), .B(n18602), .ZN(
        P3_U3029) );
  NOR2_X1 U21746 ( .A1(n18609), .A2(n20660), .ZN(n18605) );
  INV_X1 U21747 ( .A(n18605), .ZN(n18598) );
  INV_X1 U21748 ( .A(n18596), .ZN(n18597) );
  AOI22_X1 U21749 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18598), .B1(HOLD), 
        .B2(n18597), .ZN(n18600) );
  NAND2_X1 U21750 ( .A1(n18599), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18603) );
  OAI211_X1 U21751 ( .C1(n18600), .C2(n18607), .A(n18603), .B(n18730), .ZN(
        P3_U3030) );
  INV_X1 U21752 ( .A(n18603), .ZN(n18601) );
  AOI21_X1 U21753 ( .B1(n18607), .B2(n18602), .A(n18601), .ZN(n18608) );
  OAI22_X1 U21754 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18603), .ZN(n18604) );
  OAI22_X1 U21755 ( .A1(n18605), .A2(n18604), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18606) );
  OAI22_X1 U21756 ( .A1(n18608), .A2(n18609), .B1(n18607), .B2(n18606), .ZN(
        P3_U3031) );
  OAI222_X1 U21757 ( .A1(n18721), .A2(n18672), .B1(n18610), .B2(n18669), .C1(
        n18611), .C2(n18657), .ZN(P3_U3032) );
  OAI222_X1 U21758 ( .A1(n18657), .A2(n18613), .B1(n18612), .B2(n18669), .C1(
        n18611), .C2(n18672), .ZN(P3_U3033) );
  OAI222_X1 U21759 ( .A1(n18657), .A2(n18615), .B1(n18614), .B2(n18669), .C1(
        n18613), .C2(n18672), .ZN(P3_U3034) );
  OAI222_X1 U21760 ( .A1(n18657), .A2(n18618), .B1(n18616), .B2(n18669), .C1(
        n18615), .C2(n18672), .ZN(P3_U3035) );
  OAI222_X1 U21761 ( .A1(n18618), .A2(n18672), .B1(n18617), .B2(n18669), .C1(
        n18619), .C2(n18657), .ZN(P3_U3036) );
  OAI222_X1 U21762 ( .A1(n18657), .A2(n18621), .B1(n18620), .B2(n18669), .C1(
        n18619), .C2(n18672), .ZN(P3_U3037) );
  OAI222_X1 U21763 ( .A1(n18657), .A2(n18624), .B1(n18622), .B2(n18669), .C1(
        n18621), .C2(n18672), .ZN(P3_U3038) );
  OAI222_X1 U21764 ( .A1(n18624), .A2(n18672), .B1(n18623), .B2(n18669), .C1(
        n18625), .C2(n18657), .ZN(P3_U3039) );
  OAI222_X1 U21765 ( .A1(n18657), .A2(n18627), .B1(n18626), .B2(n18669), .C1(
        n18625), .C2(n18672), .ZN(P3_U3040) );
  OAI222_X1 U21766 ( .A1(n18657), .A2(n18629), .B1(n18628), .B2(n18669), .C1(
        n18627), .C2(n18672), .ZN(P3_U3041) );
  INV_X1 U21767 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18630) );
  OAI222_X1 U21768 ( .A1(n18657), .A2(n18631), .B1(n18630), .B2(n18669), .C1(
        n18629), .C2(n18672), .ZN(P3_U3042) );
  OAI222_X1 U21769 ( .A1(n18657), .A2(n18633), .B1(n18632), .B2(n18669), .C1(
        n18631), .C2(n18672), .ZN(P3_U3043) );
  OAI222_X1 U21770 ( .A1(n18657), .A2(n18635), .B1(n18634), .B2(n18669), .C1(
        n18633), .C2(n18672), .ZN(P3_U3044) );
  OAI222_X1 U21771 ( .A1(n18657), .A2(n18637), .B1(n18636), .B2(n18669), .C1(
        n18635), .C2(n18672), .ZN(P3_U3045) );
  OAI222_X1 U21772 ( .A1(n18657), .A2(n18639), .B1(n18638), .B2(n18669), .C1(
        n18637), .C2(n18672), .ZN(P3_U3046) );
  OAI222_X1 U21773 ( .A1(n18657), .A2(n18641), .B1(n18640), .B2(n18669), .C1(
        n18639), .C2(n18672), .ZN(P3_U3047) );
  OAI222_X1 U21774 ( .A1(n18657), .A2(n18643), .B1(n18642), .B2(n18669), .C1(
        n18641), .C2(n18672), .ZN(P3_U3048) );
  OAI222_X1 U21775 ( .A1(n18657), .A2(n18645), .B1(n18644), .B2(n18669), .C1(
        n18643), .C2(n18672), .ZN(P3_U3049) );
  OAI222_X1 U21776 ( .A1(n18657), .A2(n18647), .B1(n18646), .B2(n18669), .C1(
        n18645), .C2(n18672), .ZN(P3_U3050) );
  OAI222_X1 U21777 ( .A1(n18657), .A2(n18650), .B1(n18648), .B2(n18669), .C1(
        n18647), .C2(n18672), .ZN(P3_U3051) );
  INV_X1 U21778 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18651) );
  OAI222_X1 U21779 ( .A1(n18650), .A2(n18672), .B1(n18649), .B2(n18669), .C1(
        n18651), .C2(n18657), .ZN(P3_U3052) );
  OAI222_X1 U21780 ( .A1(n18657), .A2(n18654), .B1(n18652), .B2(n18669), .C1(
        n18651), .C2(n18672), .ZN(P3_U3053) );
  OAI222_X1 U21781 ( .A1(n18654), .A2(n18672), .B1(n18653), .B2(n18669), .C1(
        n18655), .C2(n18657), .ZN(P3_U3054) );
  OAI222_X1 U21782 ( .A1(n18657), .A2(n18658), .B1(n18656), .B2(n18669), .C1(
        n18655), .C2(n18672), .ZN(P3_U3055) );
  INV_X1 U21783 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18660) );
  OAI222_X1 U21784 ( .A1(n18657), .A2(n18660), .B1(n18659), .B2(n18669), .C1(
        n18658), .C2(n18672), .ZN(P3_U3056) );
  OAI222_X1 U21785 ( .A1(n18657), .A2(n18662), .B1(n18661), .B2(n18669), .C1(
        n18660), .C2(n18672), .ZN(P3_U3057) );
  INV_X1 U21786 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18664) );
  OAI222_X1 U21787 ( .A1(n18657), .A2(n18664), .B1(n18663), .B2(n18669), .C1(
        n18662), .C2(n18672), .ZN(P3_U3058) );
  OAI222_X1 U21788 ( .A1(n18657), .A2(n18666), .B1(n18665), .B2(n18669), .C1(
        n18664), .C2(n18672), .ZN(P3_U3059) );
  OAI222_X1 U21789 ( .A1(n18657), .A2(n18671), .B1(n18667), .B2(n18669), .C1(
        n18666), .C2(n18672), .ZN(P3_U3060) );
  OAI222_X1 U21790 ( .A1(n18672), .A2(n18671), .B1(n18670), .B2(n18669), .C1(
        n18668), .C2(n18657), .ZN(P3_U3061) );
  MUX2_X1 U21791 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .B(P3_BE_N_REG_3__SCAN_IN), .S(n18740), .Z(P3_U3274) );
  MUX2_X1 U21792 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n18740), .Z(P3_U3275) );
  MUX2_X1 U21793 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .B(P3_BE_N_REG_1__SCAN_IN), .S(n18740), .Z(P3_U3276) );
  MUX2_X1 U21794 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .B(P3_BE_N_REG_0__SCAN_IN), .S(n18740), .Z(P3_U3277) );
  OAI21_X1 U21795 ( .B1(n18676), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18674), 
        .ZN(n18673) );
  INV_X1 U21796 ( .A(n18673), .ZN(P3_U3280) );
  INV_X1 U21797 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18675) );
  OAI21_X1 U21798 ( .B1(n18676), .B2(n18675), .A(n18674), .ZN(P3_U3281) );
  OAI221_X1 U21799 ( .B1(n18679), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18679), 
        .C2(n18678), .A(n18677), .ZN(P3_U3282) );
  INV_X1 U21800 ( .A(n18683), .ZN(n18743) );
  AOI22_X1 U21801 ( .A1(n18743), .A2(n18681), .B1(n18703), .B2(n18680), .ZN(
        n18687) );
  OAI21_X1 U21802 ( .B1(n18683), .B2(n18682), .A(n18706), .ZN(n18684) );
  INV_X1 U21803 ( .A(n18684), .ZN(n18686) );
  OAI22_X1 U21804 ( .A1(n18709), .A2(n18687), .B1(n18686), .B2(n18685), .ZN(
        P3_U3285) );
  NOR2_X1 U21805 ( .A1(n18688), .A2(n18705), .ZN(n18697) );
  OAI22_X1 U21806 ( .A1(n18690), .A2(n18689), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18698) );
  INV_X1 U21807 ( .A(n18698), .ZN(n18692) );
  AOI222_X1 U21808 ( .A1(n18693), .A2(n18743), .B1(n18697), .B2(n18692), .C1(
        n18703), .C2(n18691), .ZN(n18694) );
  AOI22_X1 U21809 ( .A1(n18709), .A2(n18695), .B1(n18694), .B2(n18706), .ZN(
        P3_U3288) );
  INV_X1 U21810 ( .A(n18696), .ZN(n18700) );
  AOI222_X1 U21811 ( .A1(n18700), .A2(n18743), .B1(n18703), .B2(n18699), .C1(
        n18698), .C2(n18697), .ZN(n18701) );
  AOI22_X1 U21812 ( .A1(n18709), .A2(n18702), .B1(n18701), .B2(n18706), .ZN(
        P3_U3289) );
  AOI222_X1 U21813 ( .A1(n18705), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18743), 
        .B2(n18704), .C1(n18708), .C2(n18703), .ZN(n18707) );
  AOI22_X1 U21814 ( .A1(n18709), .A2(n18708), .B1(n18707), .B2(n18706), .ZN(
        P3_U3290) );
  NOR2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18711) );
  AOI211_X1 U21816 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(n18712), .A(n18711), 
        .B(n18710), .ZN(n18716) );
  NOR2_X1 U21817 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n18721), .ZN(n18714) );
  INV_X1 U21818 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18713) );
  MUX2_X1 U21819 ( .A(n18714), .B(n18713), .S(n18720), .Z(n18715) );
  NOR2_X1 U21820 ( .A1(n18716), .A2(n18715), .ZN(P3_U3292) );
  OAI21_X1 U21821 ( .B1(n18718), .B2(P3_BYTEENABLE_REG_0__SCAN_IN), .A(n18717), 
        .ZN(n18719) );
  OAI21_X1 U21822 ( .B1(n18721), .B2(n18720), .A(n18719), .ZN(P3_U3293) );
  INV_X1 U21823 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n20924) );
  OAI22_X1 U21824 ( .A1(n18740), .A2(n20924), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18669), .ZN(n18722) );
  INV_X1 U21825 ( .A(n18722), .ZN(P3_U3294) );
  MUX2_X1 U21826 ( .A(P3_MORE_REG_SCAN_IN), .B(n18724), .S(n18723), .Z(
        P3_U3295) );
  OAI21_X1 U21827 ( .B1(n18727), .B2(n18726), .A(n18725), .ZN(n18728) );
  AOI21_X1 U21828 ( .B1(n18729), .B2(n18733), .A(n18728), .ZN(n18739) );
  AOI21_X1 U21829 ( .B1(n18732), .B2(n18731), .A(n18730), .ZN(n18734) );
  OAI211_X1 U21830 ( .C1(n18744), .C2(n18734), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18733), .ZN(n18736) );
  AOI21_X1 U21831 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18736), .A(n18735), 
        .ZN(n18738) );
  NAND2_X1 U21832 ( .A1(n18739), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18737) );
  OAI21_X1 U21833 ( .B1(n18739), .B2(n18738), .A(n18737), .ZN(P3_U3296) );
  OAI22_X1 U21834 ( .A1(n18740), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18669), .ZN(n18741) );
  INV_X1 U21835 ( .A(n18741), .ZN(P3_U3297) );
  AOI21_X1 U21836 ( .B1(n18743), .B2(n18742), .A(n18746), .ZN(n18749) );
  INV_X1 U21837 ( .A(n18744), .ZN(n18745) );
  AOI22_X1 U21838 ( .A1(n18749), .A2(n20924), .B1(n18746), .B2(n18745), .ZN(
        P3_U3298) );
  INV_X1 U21839 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18748) );
  AOI21_X1 U21840 ( .B1(n18749), .B2(n18748), .A(n18747), .ZN(P3_U3299) );
  INV_X1 U21841 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19614) );
  NAND2_X1 U21842 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19619), .ZN(n19608) );
  NAND2_X1 U21843 ( .A1(n19614), .A2(n19601), .ZN(n19605) );
  OAI21_X1 U21844 ( .B1(n19614), .B2(n19608), .A(n19605), .ZN(n19678) );
  AOI21_X1 U21845 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19678), .ZN(n18750) );
  INV_X1 U21846 ( .A(n18750), .ZN(P2_U2815) );
  INV_X1 U21847 ( .A(n18751), .ZN(n19727) );
  AOI22_X1 U21848 ( .A1(P2_CODEFETCH_REG_SCAN_IN), .A2(n19727), .B1(n18752), 
        .B2(n19733), .ZN(n18753) );
  INV_X1 U21849 ( .A(n18753), .ZN(P2_U2816) );
  INV_X2 U21850 ( .A(n19745), .ZN(n19744) );
  AOI21_X1 U21851 ( .B1(n19614), .B2(n19619), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18754) );
  AOI22_X1 U21852 ( .A1(n19744), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18754), 
        .B2(n19745), .ZN(P2_U2817) );
  OAI21_X1 U21853 ( .B1(n19612), .B2(BS16), .A(n19678), .ZN(n19676) );
  OAI21_X1 U21854 ( .B1(n19678), .B2(n19736), .A(n19676), .ZN(P2_U2818) );
  NOR2_X1 U21855 ( .A1(n18756), .A2(n18755), .ZN(n19717) );
  OAI21_X1 U21856 ( .B1(n19717), .B2(n18758), .A(n18757), .ZN(P2_U2819) );
  NOR4_X1 U21857 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n18768) );
  NOR4_X1 U21858 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18767) );
  NOR4_X1 U21859 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n18759) );
  INV_X1 U21860 ( .A(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(n19598) );
  INV_X1 U21861 ( .A(P2_DATAWIDTH_REG_20__SCAN_IN), .ZN(n20774) );
  NAND3_X1 U21862 ( .A1(n18759), .A2(n19598), .A3(n20774), .ZN(n18765) );
  NOR4_X1 U21863 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18763) );
  NOR4_X1 U21864 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n18762) );
  NOR4_X1 U21865 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18761) );
  NOR4_X1 U21866 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18760) );
  NAND4_X1 U21867 ( .A1(n18763), .A2(n18762), .A3(n18761), .A4(n18760), .ZN(
        n18764) );
  AOI211_X1 U21868 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n18765), .B(n18764), .ZN(n18766) );
  NAND3_X1 U21869 ( .A1(n18768), .A2(n18767), .A3(n18766), .ZN(n18771) );
  NOR2_X1 U21870 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18771), .ZN(n18770) );
  INV_X1 U21871 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18769) );
  AOI22_X1 U21872 ( .A1(n18770), .A2(n18919), .B1(n18771), .B2(n18769), .ZN(
        P2_U2820) );
  INV_X1 U21873 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20949) );
  OR4_X1 U21874 ( .A1(n18771), .A2(P2_REIP_REG_0__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A4(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18775) );
  OAI221_X1 U21875 ( .B1(n18770), .B2(n20949), .C1(n18770), .C2(n18771), .A(
        n18775), .ZN(P2_U2821) );
  INV_X1 U21876 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19677) );
  NAND2_X1 U21877 ( .A1(n18770), .A2(n19677), .ZN(n18774) );
  INV_X1 U21878 ( .A(n18771), .ZN(n18777) );
  OAI21_X1 U21879 ( .B1(n19620), .B2(n18919), .A(n18777), .ZN(n18772) );
  OAI21_X1 U21880 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18777), .A(n18772), 
        .ZN(n18773) );
  OAI221_X1 U21881 ( .B1(n18774), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18774), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18773), .ZN(P2_U2822) );
  INV_X1 U21882 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18776) );
  OAI211_X1 U21883 ( .C1(n18777), .C2(n18776), .A(n18775), .B(n18774), .ZN(
        P2_U2823) );
  INV_X1 U21884 ( .A(n18778), .ZN(n18779) );
  OAI22_X1 U21885 ( .A1(n18780), .A2(n18878), .B1(n18779), .B2(n18916), .ZN(
        n18781) );
  INV_X1 U21886 ( .A(n18781), .ZN(n18790) );
  AOI211_X1 U21887 ( .C1(n18784), .C2(n18783), .A(n18782), .B(n18883), .ZN(
        n18788) );
  AOI22_X1 U21888 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n18917), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18829), .ZN(n18785) );
  OAI21_X1 U21889 ( .B1(n18786), .B2(n18925), .A(n18785), .ZN(n18787) );
  AOI211_X1 U21890 ( .C1(n18906), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n18788), .B(n18787), .ZN(n18789) );
  NAND2_X1 U21891 ( .A1(n18790), .A2(n18789), .ZN(P2_U2834) );
  INV_X1 U21892 ( .A(n18791), .ZN(n18792) );
  AOI22_X1 U21893 ( .A1(n18793), .A2(n18927), .B1(n18792), .B2(n18922), .ZN(
        n18802) );
  AOI211_X1 U21894 ( .C1(n18796), .C2(n18795), .A(n18794), .B(n18883), .ZN(
        n18800) );
  AOI22_X1 U21895 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18906), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18829), .ZN(n18797) );
  OAI21_X1 U21896 ( .B1(n18798), .B2(n18925), .A(n18797), .ZN(n18799) );
  AOI211_X1 U21897 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n18917), .A(n18800), .B(
        n18799), .ZN(n18801) );
  NAND2_X1 U21898 ( .A1(n18802), .A2(n18801), .ZN(P2_U2835) );
  INV_X1 U21899 ( .A(n18803), .ZN(n18812) );
  AOI22_X1 U21900 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n18917), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18906), .ZN(n18805) );
  AOI21_X1 U21901 ( .B1(P2_REIP_REG_19__SCAN_IN), .B2(n18829), .A(n15058), 
        .ZN(n18804) );
  OAI211_X1 U21902 ( .C1(n18878), .C2(n18806), .A(n18805), .B(n18804), .ZN(
        n18811) );
  AOI211_X1 U21903 ( .C1(n18809), .C2(n18808), .A(n18883), .B(n18807), .ZN(
        n18810) );
  AOI211_X1 U21904 ( .C1(n18901), .C2(n18812), .A(n18811), .B(n18810), .ZN(
        n18813) );
  OAI21_X1 U21905 ( .B1(n18814), .B2(n18916), .A(n18813), .ZN(P2_U2836) );
  AOI211_X1 U21906 ( .C1(n18817), .C2(n18816), .A(n18815), .B(n18936), .ZN(
        n18820) );
  AOI22_X1 U21907 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n18917), .B1(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18906), .ZN(n18818) );
  OAI211_X1 U21908 ( .C1(n19644), .C2(n18918), .A(n18818), .B(n18900), .ZN(
        n18819) );
  AOI211_X1 U21909 ( .C1(n18901), .C2(n18821), .A(n18820), .B(n18819), .ZN(
        n18825) );
  AOI22_X1 U21910 ( .A1(n18823), .A2(n18927), .B1(n18922), .B2(n18822), .ZN(
        n18824) );
  OAI211_X1 U21911 ( .C1(n18826), .C2(n18930), .A(n18825), .B(n18824), .ZN(
        P2_U2838) );
  INV_X1 U21912 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20927) );
  OAI22_X1 U21913 ( .A1(n18887), .A2(n13663), .B1(n18827), .B2(n18925), .ZN(
        n18828) );
  AOI211_X1 U21914 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18829), .A(n15058), 
        .B(n18828), .ZN(n18838) );
  NOR2_X1 U21915 ( .A1(n18891), .A2(n18830), .ZN(n18831) );
  XNOR2_X1 U21916 ( .A(n18832), .B(n18831), .ZN(n18836) );
  OAI22_X1 U21917 ( .A1(n18834), .A2(n18878), .B1(n18916), .B2(n18833), .ZN(
        n18835) );
  AOI21_X1 U21918 ( .B1(n18836), .B2(n18912), .A(n18835), .ZN(n18837) );
  OAI211_X1 U21919 ( .C1(n20927), .C2(n18931), .A(n18838), .B(n18837), .ZN(
        P2_U2839) );
  NAND2_X1 U21920 ( .A1(n9642), .A2(n18839), .ZN(n18841) );
  XOR2_X1 U21921 ( .A(n18841), .B(n18840), .Z(n18850) );
  AOI22_X1 U21922 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n18917), .B1(n18842), 
        .B2(n18901), .ZN(n18843) );
  OAI211_X1 U21923 ( .C1(n10781), .C2(n18918), .A(n18843), .B(n18885), .ZN(
        n18848) );
  INV_X1 U21924 ( .A(n18844), .ZN(n18846) );
  OAI22_X1 U21925 ( .A1(n18846), .A2(n18878), .B1(n18916), .B2(n18845), .ZN(
        n18847) );
  AOI211_X1 U21926 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18906), .A(
        n18848), .B(n18847), .ZN(n18849) );
  OAI21_X1 U21927 ( .B1(n18850), .B2(n18883), .A(n18849), .ZN(P2_U2844) );
  OAI21_X1 U21928 ( .B1(n19634), .B2(n18918), .A(n18900), .ZN(n18853) );
  OAI22_X1 U21929 ( .A1(n18887), .A2(n10499), .B1(n18851), .B2(n18925), .ZN(
        n18852) );
  AOI211_X1 U21930 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18906), .A(
        n18853), .B(n18852), .ZN(n18860) );
  NOR2_X1 U21931 ( .A1(n18891), .A2(n18854), .ZN(n18856) );
  XNOR2_X1 U21932 ( .A(n18856), .B(n18855), .ZN(n18858) );
  AOI22_X1 U21933 ( .A1(n18858), .A2(n18912), .B1(n18927), .B2(n18857), .ZN(
        n18859) );
  OAI211_X1 U21934 ( .C1(n18952), .C2(n18916), .A(n18860), .B(n18859), .ZN(
        P2_U2845) );
  NAND2_X1 U21935 ( .A1(n9642), .A2(n18861), .ZN(n18863) );
  XOR2_X1 U21936 ( .A(n18863), .B(n18862), .Z(n18871) );
  AOI22_X1 U21937 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18906), .B1(
        n18901), .B2(n18864), .ZN(n18865) );
  OAI211_X1 U21938 ( .C1(n10755), .C2(n18918), .A(n18865), .B(n18885), .ZN(
        n18869) );
  OAI22_X1 U21939 ( .A1(n18867), .A2(n18878), .B1(n18916), .B2(n18866), .ZN(
        n18868) );
  AOI211_X1 U21940 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n18917), .A(n18869), .B(
        n18868), .ZN(n18870) );
  OAI21_X1 U21941 ( .B1(n18871), .B2(n18883), .A(n18870), .ZN(P2_U2846) );
  NAND2_X1 U21942 ( .A1(n9642), .A2(n18872), .ZN(n18874) );
  XOR2_X1 U21943 ( .A(n18874), .B(n18873), .Z(n18884) );
  AOI22_X1 U21944 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18906), .B1(
        n18875), .B2(n18901), .ZN(n18876) );
  OAI211_X1 U21945 ( .C1(n19630), .C2(n18918), .A(n18876), .B(n18885), .ZN(
        n18881) );
  OAI22_X1 U21946 ( .A1(n18879), .A2(n18916), .B1(n18878), .B2(n18877), .ZN(
        n18880) );
  AOI211_X1 U21947 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n18917), .A(n18881), .B(
        n18880), .ZN(n18882) );
  OAI21_X1 U21948 ( .B1(n18884), .B2(n18883), .A(n18882), .ZN(P2_U2848) );
  OAI21_X1 U21949 ( .B1(n19628), .B2(n18918), .A(n18885), .ZN(n18889) );
  OAI22_X1 U21950 ( .A1(n18887), .A2(n10482), .B1(n18886), .B2(n18925), .ZN(
        n18888) );
  AOI211_X1 U21951 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18906), .A(
        n18889), .B(n18888), .ZN(n18898) );
  NOR2_X1 U21952 ( .A1(n18891), .A2(n18890), .ZN(n18893) );
  XNOR2_X1 U21953 ( .A(n18893), .B(n18892), .ZN(n18896) );
  INV_X1 U21954 ( .A(n18894), .ZN(n18895) );
  AOI22_X1 U21955 ( .A1(n18896), .A2(n18912), .B1(n18927), .B2(n18895), .ZN(
        n18897) );
  OAI211_X1 U21956 ( .C1(n18916), .C2(n18899), .A(n18898), .B(n18897), .ZN(
        P2_U2849) );
  OAI21_X1 U21957 ( .B1(n10703), .B2(n18918), .A(n18900), .ZN(n18905) );
  AOI22_X1 U21958 ( .A1(n18917), .A2(P2_EBX_REG_5__SCAN_IN), .B1(n18902), .B2(
        n18901), .ZN(n18903) );
  INV_X1 U21959 ( .A(n18903), .ZN(n18904) );
  AOI211_X1 U21960 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18906), .A(
        n18905), .B(n18904), .ZN(n18915) );
  NAND2_X1 U21961 ( .A1(n9642), .A2(n18907), .ZN(n18909) );
  XNOR2_X1 U21962 ( .A(n18910), .B(n18909), .ZN(n18913) );
  AOI22_X1 U21963 ( .A1(n18913), .A2(n18912), .B1(n18927), .B2(n18911), .ZN(
        n18914) );
  OAI211_X1 U21964 ( .C1(n18916), .C2(n18963), .A(n18915), .B(n18914), .ZN(
        P2_U2850) );
  OAI22_X1 U21965 ( .A1(n18887), .A2(n18920), .B1(n18919), .B2(n18918), .ZN(
        n18921) );
  AOI21_X1 U21966 ( .B1(n18922), .B2(n18988), .A(n18921), .ZN(n18923) );
  OAI21_X1 U21967 ( .B1(n18925), .B2(n18924), .A(n18923), .ZN(n18926) );
  AOI21_X1 U21968 ( .B1(n18928), .B2(n18927), .A(n18926), .ZN(n18935) );
  INV_X1 U21969 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18929) );
  AOI21_X1 U21970 ( .B1(n18931), .B2(n18930), .A(n18929), .ZN(n18932) );
  AOI21_X1 U21971 ( .B1(n18933), .B2(n18989), .A(n18932), .ZN(n18934) );
  OAI211_X1 U21972 ( .C1(n18937), .C2(n18936), .A(n18935), .B(n18934), .ZN(
        P2_U2855) );
  AOI22_X1 U21973 ( .A1(n18939), .A2(n18984), .B1(n18938), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n18942) );
  AOI22_X1 U21974 ( .A1(n18940), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18983), .ZN(n18941) );
  NAND2_X1 U21975 ( .A1(n18942), .A2(n18941), .ZN(P2_U2888) );
  INV_X1 U21976 ( .A(n18943), .ZN(n18945) );
  AOI22_X1 U21977 ( .A1(n18958), .A2(n19032), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n18983), .ZN(n18944) );
  OAI21_X1 U21978 ( .B1(n18964), .B2(n18945), .A(n18944), .ZN(P2_U2905) );
  INV_X1 U21979 ( .A(n18946), .ZN(n18949) );
  AOI22_X1 U21980 ( .A1(n18958), .A2(n18947), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n18983), .ZN(n18948) );
  OAI21_X1 U21981 ( .B1(n18964), .B2(n18949), .A(n18948), .ZN(P2_U2907) );
  AOI22_X1 U21982 ( .A1(n18958), .A2(n18950), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n18983), .ZN(n18951) );
  OAI21_X1 U21983 ( .B1(n18964), .B2(n18952), .A(n18951), .ZN(P2_U2909) );
  INV_X1 U21984 ( .A(n18953), .ZN(n18956) );
  AOI22_X1 U21985 ( .A1(n18958), .A2(n18954), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n18983), .ZN(n18955) );
  OAI21_X1 U21986 ( .B1(n18964), .B2(n18956), .A(n18955), .ZN(P2_U2911) );
  AOI22_X1 U21987 ( .A1(n18958), .A2(n18957), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n18983), .ZN(n18962) );
  OR3_X1 U21988 ( .A1(n18960), .A2(n18959), .A3(n18978), .ZN(n18961) );
  OAI211_X1 U21989 ( .C1(n18964), .C2(n18963), .A(n18962), .B(n18961), .ZN(
        P2_U2914) );
  INV_X1 U21990 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18965) );
  OAI22_X1 U21991 ( .A1(n19686), .A2(n18967), .B1(n18966), .B2(n18965), .ZN(
        n18968) );
  INV_X1 U21992 ( .A(n18968), .ZN(n18974) );
  AOI21_X1 U21993 ( .B1(n18971), .B2(n18970), .A(n18969), .ZN(n18972) );
  OR2_X1 U21994 ( .A1(n18972), .A2(n18978), .ZN(n18973) );
  OAI211_X1 U21995 ( .C1(n18975), .C2(n18992), .A(n18974), .B(n18973), .ZN(
        P2_U2916) );
  AOI22_X1 U21996 ( .A1(n18984), .A2(n19703), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n18983), .ZN(n18981) );
  AOI21_X1 U21997 ( .B1(n18985), .B2(n18977), .A(n18976), .ZN(n18979) );
  OR2_X1 U21998 ( .A1(n18979), .A2(n18978), .ZN(n18980) );
  OAI211_X1 U21999 ( .C1(n18982), .C2(n18992), .A(n18981), .B(n18980), .ZN(
        P2_U2918) );
  AOI22_X1 U22000 ( .A1(n18984), .A2(n18988), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n18983), .ZN(n18991) );
  INV_X1 U22001 ( .A(n18985), .ZN(n18987) );
  OAI211_X1 U22002 ( .C1(n18989), .C2(n18988), .A(n18987), .B(n18986), .ZN(
        n18990) );
  OAI211_X1 U22003 ( .C1(n18993), .C2(n18992), .A(n18991), .B(n18990), .ZN(
        P2_U2919) );
  NOR2_X1 U22004 ( .A1(n18998), .A2(n18994), .ZN(P2_U2920) );
  INV_X1 U22005 ( .A(n18995), .ZN(n18996) );
  AOI22_X1 U22006 ( .A1(n18996), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19025), .ZN(n18997) );
  OAI21_X1 U22007 ( .B1(n18999), .B2(n18998), .A(n18997), .ZN(P2_U2921) );
  AOI22_X1 U22008 ( .A1(n19025), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19000) );
  OAI21_X1 U22009 ( .B1(n12672), .B2(n19030), .A(n19000), .ZN(P2_U2936) );
  INV_X1 U22010 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19002) );
  AOI22_X1 U22011 ( .A1(n19025), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19001) );
  OAI21_X1 U22012 ( .B1(n19002), .B2(n19030), .A(n19001), .ZN(P2_U2937) );
  AOI22_X1 U22013 ( .A1(n19025), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19003) );
  OAI21_X1 U22014 ( .B1(n19004), .B2(n19030), .A(n19003), .ZN(P2_U2938) );
  AOI22_X1 U22015 ( .A1(n19025), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19005) );
  OAI21_X1 U22016 ( .B1(n19006), .B2(n19030), .A(n19005), .ZN(P2_U2939) );
  AOI22_X1 U22017 ( .A1(n19025), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19007) );
  OAI21_X1 U22018 ( .B1(n19008), .B2(n19030), .A(n19007), .ZN(P2_U2940) );
  AOI22_X1 U22019 ( .A1(n19025), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19009) );
  OAI21_X1 U22020 ( .B1(n10766), .B2(n19030), .A(n19009), .ZN(P2_U2941) );
  AOI22_X1 U22021 ( .A1(n19025), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19010) );
  OAI21_X1 U22022 ( .B1(n19011), .B2(n19030), .A(n19010), .ZN(P2_U2942) );
  AOI22_X1 U22023 ( .A1(n19025), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19012) );
  OAI21_X1 U22024 ( .B1(n19013), .B2(n19030), .A(n19012), .ZN(P2_U2943) );
  AOI22_X1 U22025 ( .A1(n19025), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19014) );
  OAI21_X1 U22026 ( .B1(n19015), .B2(n19030), .A(n19014), .ZN(P2_U2944) );
  AOI22_X1 U22027 ( .A1(n19025), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19016) );
  OAI21_X1 U22028 ( .B1(n19017), .B2(n19030), .A(n19016), .ZN(P2_U2945) );
  INV_X1 U22029 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19019) );
  AOI22_X1 U22030 ( .A1(n19025), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19018) );
  OAI21_X1 U22031 ( .B1(n19019), .B2(n19030), .A(n19018), .ZN(P2_U2946) );
  INV_X1 U22032 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19021) );
  AOI22_X1 U22033 ( .A1(n19025), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19020) );
  OAI21_X1 U22034 ( .B1(n19021), .B2(n19030), .A(n19020), .ZN(P2_U2947) );
  AOI22_X1 U22035 ( .A1(n19025), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19022) );
  OAI21_X1 U22036 ( .B1(n18965), .B2(n19030), .A(n19022), .ZN(P2_U2948) );
  INV_X1 U22037 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19024) );
  AOI22_X1 U22038 ( .A1(n19025), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19023) );
  OAI21_X1 U22039 ( .B1(n19024), .B2(n19030), .A(n19023), .ZN(P2_U2949) );
  INV_X1 U22040 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19027) );
  AOI22_X1 U22041 ( .A1(n19025), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19026) );
  OAI21_X1 U22042 ( .B1(n19027), .B2(n19030), .A(n19026), .ZN(P2_U2950) );
  INV_X1 U22043 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19031) );
  AOI22_X1 U22044 ( .A1(n19025), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19028), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19029) );
  OAI21_X1 U22045 ( .B1(n19031), .B2(n19030), .A(n19029), .ZN(P2_U2951) );
  AOI22_X1 U22046 ( .A1(n19036), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19035), .ZN(n19034) );
  NAND2_X1 U22047 ( .A1(n19033), .A2(n19032), .ZN(n19037) );
  NAND2_X1 U22048 ( .A1(n19034), .A2(n19037), .ZN(P2_U2966) );
  AOI22_X1 U22049 ( .A1(n19036), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19035), .ZN(n19038) );
  NAND2_X1 U22050 ( .A1(n19038), .A2(n19037), .ZN(P2_U2981) );
  AOI22_X1 U22051 ( .A1(n19039), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n15397), .ZN(n19050) );
  NAND2_X1 U22052 ( .A1(n19041), .A2(n19040), .ZN(n19045) );
  NAND2_X1 U22053 ( .A1(n19043), .A2(n19042), .ZN(n19044) );
  OAI211_X1 U22054 ( .C1(n19047), .C2(n19046), .A(n19045), .B(n19044), .ZN(
        n19048) );
  INV_X1 U22055 ( .A(n19048), .ZN(n19049) );
  OAI211_X1 U22056 ( .C1(n19052), .C2(n19051), .A(n19050), .B(n19049), .ZN(
        P2_U3010) );
  AOI211_X1 U22057 ( .C1(n19056), .C2(n19055), .A(n19054), .B(n19053), .ZN(
        n19073) );
  INV_X1 U22058 ( .A(n19063), .ZN(n19058) );
  OAI21_X1 U22059 ( .B1(n19059), .B2(n19058), .A(n19057), .ZN(n19060) );
  NAND2_X1 U22060 ( .A1(n19060), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19061) );
  OAI21_X1 U22061 ( .B1(n19063), .B2(n19062), .A(n19061), .ZN(n19064) );
  AOI21_X1 U22062 ( .B1(n19066), .B2(n19065), .A(n19064), .ZN(n19069) );
  NAND2_X1 U22063 ( .A1(n11911), .A2(n19067), .ZN(n19068) );
  OAI211_X1 U22064 ( .C1(n19692), .C2(n19070), .A(n19069), .B(n19068), .ZN(
        n19071) );
  INV_X1 U22065 ( .A(n19071), .ZN(n19072) );
  OAI211_X1 U22066 ( .C1(n19075), .C2(n19074), .A(n19073), .B(n19072), .ZN(
        P2_U3044) );
  NAND3_X1 U22067 ( .A1(n19078), .A2(n19682), .A3(n19147), .ZN(n19079) );
  NAND2_X1 U22068 ( .A1(n19682), .A2(n19736), .ZN(n19681) );
  NAND2_X1 U22069 ( .A1(n19079), .A2(n19681), .ZN(n19088) );
  NAND2_X1 U22070 ( .A1(n19088), .A2(n19080), .ZN(n19083) );
  AOI21_X1 U22071 ( .B1(n19081), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19082) );
  NAND2_X1 U22072 ( .A1(n19083), .A2(n19082), .ZN(n19086) );
  NAND2_X1 U22073 ( .A1(n19690), .A2(n12319), .ZN(n19195) );
  INV_X1 U22074 ( .A(n19195), .ZN(n19084) );
  NAND2_X1 U22075 ( .A1(n19084), .A2(n19705), .ZN(n19121) );
  NOR2_X1 U22076 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19121), .ZN(
        n19110) );
  INV_X1 U22077 ( .A(n19110), .ZN(n19085) );
  NAND2_X1 U22078 ( .A1(n19086), .A2(n19085), .ZN(n19087) );
  INV_X1 U22079 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19093) );
  AOI22_X1 U22080 ( .A1(n19591), .A2(n19512), .B1(n19511), .B2(n19110), .ZN(
        n19092) );
  OAI21_X1 U22081 ( .B1(n19587), .B2(n19110), .A(n19088), .ZN(n19090) );
  OAI21_X1 U22082 ( .B1(n11965), .B2(n19110), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19089) );
  NAND2_X1 U22083 ( .A1(n19090), .A2(n19089), .ZN(n19111) );
  AOI22_X1 U22084 ( .A1(n19467), .A2(n19111), .B1(n19156), .B2(n19519), .ZN(
        n19091) );
  OAI211_X1 U22085 ( .C1(n19107), .C2(n19093), .A(n19092), .B(n19091), .ZN(
        P2_U3048) );
  INV_X1 U22086 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19096) );
  AOI22_X1 U22087 ( .A1(n19591), .A2(n19554), .B1(n19551), .B2(n19110), .ZN(
        n19095) );
  AOI22_X1 U22088 ( .A1(n19552), .A2(n19111), .B1(n19156), .B2(n19553), .ZN(
        n19094) );
  OAI211_X1 U22089 ( .C1(n19107), .C2(n19096), .A(n19095), .B(n19094), .ZN(
        P2_U3049) );
  AOI22_X1 U22090 ( .A1(n19591), .A2(n19561), .B1(n19558), .B2(n19110), .ZN(
        n19098) );
  AOI22_X1 U22091 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19112), .B1(
        n19559), .B2(n19111), .ZN(n19097) );
  OAI211_X1 U22092 ( .C1(n19484), .C2(n19147), .A(n19098), .B(n19097), .ZN(
        P2_U3050) );
  AOI22_X1 U22093 ( .A1(n19591), .A2(n19530), .B1(n19529), .B2(n19110), .ZN(
        n19100) );
  AOI22_X1 U22094 ( .A1(n19485), .A2(n19111), .B1(n19156), .B2(n19531), .ZN(
        n19099) );
  OAI211_X1 U22095 ( .C1(n19107), .C2(n19101), .A(n19100), .B(n19099), .ZN(
        P2_U3051) );
  AOI22_X1 U22096 ( .A1(n19591), .A2(n19567), .B1(n19565), .B2(n19110), .ZN(
        n19103) );
  AOI22_X1 U22097 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19112), .B1(
        n19566), .B2(n19111), .ZN(n19102) );
  OAI211_X1 U22098 ( .C1(n19491), .C2(n19147), .A(n19103), .B(n19102), .ZN(
        P2_U3052) );
  AOI22_X1 U22099 ( .A1(n19591), .A2(n19574), .B1(n19572), .B2(n19110), .ZN(
        n19105) );
  AOI22_X1 U22100 ( .A1(n19573), .A2(n19111), .B1(n19156), .B2(n19575), .ZN(
        n19104) );
  OAI211_X1 U22101 ( .C1(n19107), .C2(n19106), .A(n19105), .B(n19104), .ZN(
        P2_U3053) );
  AOI22_X1 U22102 ( .A1(n19591), .A2(n19582), .B1(n19579), .B2(n19110), .ZN(
        n19109) );
  AOI22_X1 U22103 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19112), .B1(
        n19580), .B2(n19111), .ZN(n19108) );
  OAI211_X1 U22104 ( .C1(n19498), .C2(n19147), .A(n19109), .B(n19108), .ZN(
        P2_U3054) );
  AOI22_X1 U22105 ( .A1(n19591), .A2(n19592), .B1(n19586), .B2(n19110), .ZN(
        n19114) );
  AOI22_X1 U22106 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19112), .B1(
        n19588), .B2(n19111), .ZN(n19113) );
  OAI211_X1 U22107 ( .C1(n19505), .C2(n19147), .A(n19114), .B(n19113), .ZN(
        P2_U3055) );
  NOR2_X1 U22108 ( .A1(n19356), .A2(n19195), .ZN(n19124) );
  INV_X1 U22109 ( .A(n19124), .ZN(n19152) );
  NAND2_X1 U22110 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19152), .ZN(n19115) );
  NOR2_X1 U22111 ( .A1(n11936), .A2(n19115), .ZN(n19120) );
  INV_X1 U22112 ( .A(n19121), .ZN(n19116) );
  AOI21_X1 U22113 ( .B1(n19731), .B2(n19116), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19117) );
  OAI22_X1 U22114 ( .A1(n19154), .A2(n19522), .B1(n19118), .B2(n19152), .ZN(
        n19119) );
  INV_X1 U22115 ( .A(n19119), .ZN(n19126) );
  NAND2_X1 U22116 ( .A1(n19298), .A2(n19361), .ZN(n19122) );
  AOI21_X1 U22117 ( .B1(n19122), .B2(n19121), .A(n19120), .ZN(n19123) );
  OAI211_X1 U22118 ( .C1(n19124), .C2(n19731), .A(n19123), .B(n19516), .ZN(
        n19157) );
  AOI22_X1 U22119 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19157), .B1(
        n19189), .B2(n19519), .ZN(n19125) );
  OAI211_X1 U22120 ( .C1(n19478), .C2(n19147), .A(n19126), .B(n19125), .ZN(
        P2_U3056) );
  INV_X1 U22121 ( .A(n19189), .ZN(n19160) );
  INV_X1 U22122 ( .A(n19551), .ZN(n19127) );
  OAI22_X1 U22123 ( .A1(n19154), .A2(n19525), .B1(n19127), .B2(n19152), .ZN(
        n19128) );
  INV_X1 U22124 ( .A(n19128), .ZN(n19130) );
  AOI22_X1 U22125 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19157), .B1(
        n19156), .B2(n19554), .ZN(n19129) );
  OAI211_X1 U22126 ( .C1(n19481), .C2(n19160), .A(n19130), .B(n19129), .ZN(
        P2_U3057) );
  INV_X1 U22127 ( .A(n19558), .ZN(n19131) );
  OAI22_X1 U22128 ( .A1(n19154), .A2(n19528), .B1(n19152), .B2(n19131), .ZN(
        n19132) );
  INV_X1 U22129 ( .A(n19132), .ZN(n19134) );
  AOI22_X1 U22130 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19157), .B1(
        n19156), .B2(n19561), .ZN(n19133) );
  OAI211_X1 U22131 ( .C1(n19484), .C2(n19160), .A(n19134), .B(n19133), .ZN(
        P2_U3058) );
  OAI22_X1 U22132 ( .A1(n19154), .A2(n19534), .B1(n19135), .B2(n19152), .ZN(
        n19136) );
  INV_X1 U22133 ( .A(n19136), .ZN(n19138) );
  AOI22_X1 U22134 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19157), .B1(
        n19189), .B2(n19531), .ZN(n19137) );
  OAI211_X1 U22135 ( .C1(n19488), .C2(n19147), .A(n19138), .B(n19137), .ZN(
        P2_U3059) );
  INV_X1 U22136 ( .A(n19565), .ZN(n19139) );
  OAI22_X1 U22137 ( .A1(n19154), .A2(n19537), .B1(n19152), .B2(n19139), .ZN(
        n19140) );
  INV_X1 U22138 ( .A(n19140), .ZN(n19142) );
  AOI22_X1 U22139 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19157), .B1(
        n19189), .B2(n19568), .ZN(n19141) );
  OAI211_X1 U22140 ( .C1(n19452), .C2(n19147), .A(n19142), .B(n19141), .ZN(
        P2_U3060) );
  INV_X1 U22141 ( .A(n19572), .ZN(n19143) );
  OAI22_X1 U22142 ( .A1(n19154), .A2(n19540), .B1(n19143), .B2(n19152), .ZN(
        n19144) );
  INV_X1 U22143 ( .A(n19144), .ZN(n19146) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19157), .B1(
        n19189), .B2(n19575), .ZN(n19145) );
  OAI211_X1 U22145 ( .C1(n19495), .C2(n19147), .A(n19146), .B(n19145), .ZN(
        P2_U3061) );
  INV_X1 U22146 ( .A(n19579), .ZN(n19148) );
  OAI22_X1 U22147 ( .A1(n19154), .A2(n19543), .B1(n19152), .B2(n19148), .ZN(
        n19149) );
  INV_X1 U22148 ( .A(n19149), .ZN(n19151) );
  AOI22_X1 U22149 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19157), .B1(
        n19156), .B2(n19582), .ZN(n19150) );
  OAI211_X1 U22150 ( .C1(n19498), .C2(n19160), .A(n19151), .B(n19150), .ZN(
        P2_U3062) );
  INV_X1 U22151 ( .A(n19586), .ZN(n19153) );
  OAI22_X1 U22152 ( .A1(n19154), .A2(n19549), .B1(n19153), .B2(n19152), .ZN(
        n19155) );
  INV_X1 U22153 ( .A(n19155), .ZN(n19159) );
  AOI22_X1 U22154 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19157), .B1(
        n19156), .B2(n19592), .ZN(n19158) );
  OAI211_X1 U22155 ( .C1(n19505), .C2(n19160), .A(n19159), .B(n19158), .ZN(
        P2_U3063) );
  NOR2_X1 U22156 ( .A1(n19389), .A2(n19195), .ZN(n19161) );
  AOI221_X1 U22157 ( .B1(n19189), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19224), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19161), .ZN(n19165) );
  INV_X1 U22158 ( .A(n11958), .ZN(n19162) );
  AOI21_X1 U22159 ( .B1(n19162), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19163) );
  NOR2_X1 U22160 ( .A1(n19387), .A2(n19195), .ZN(n19187) );
  OAI21_X1 U22161 ( .B1(n19163), .B2(n19187), .A(n19516), .ZN(n19164) );
  INV_X1 U22162 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n20896) );
  OAI21_X1 U22163 ( .B1(n11958), .B2(n19187), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19166) );
  OAI21_X1 U22164 ( .B1(n19195), .B2(n19389), .A(n19166), .ZN(n19188) );
  AOI22_X1 U22165 ( .A1(n19188), .A2(n19467), .B1(n19511), .B2(n19187), .ZN(
        n19168) );
  AOI22_X1 U22166 ( .A1(n19224), .A2(n19519), .B1(n19189), .B2(n19512), .ZN(
        n19167) );
  OAI211_X1 U22167 ( .C1(n19193), .C2(n20896), .A(n19168), .B(n19167), .ZN(
        P2_U3064) );
  INV_X1 U22168 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n19171) );
  AOI22_X1 U22169 ( .A1(n19188), .A2(n19552), .B1(n19551), .B2(n19187), .ZN(
        n19170) );
  AOI22_X1 U22170 ( .A1(n19189), .A2(n19554), .B1(n19224), .B2(n19553), .ZN(
        n19169) );
  OAI211_X1 U22171 ( .C1(n19193), .C2(n19171), .A(n19170), .B(n19169), .ZN(
        P2_U3065) );
  INV_X1 U22172 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n19174) );
  AOI22_X1 U22173 ( .A1(n19188), .A2(n19559), .B1(n19187), .B2(n19558), .ZN(
        n19173) );
  AOI22_X1 U22174 ( .A1(n19189), .A2(n19561), .B1(n19224), .B2(n19560), .ZN(
        n19172) );
  OAI211_X1 U22175 ( .C1(n19193), .C2(n19174), .A(n19173), .B(n19172), .ZN(
        P2_U3066) );
  INV_X1 U22176 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n19177) );
  AOI22_X1 U22177 ( .A1(n19188), .A2(n19485), .B1(n19529), .B2(n19187), .ZN(
        n19176) );
  AOI22_X1 U22178 ( .A1(n19224), .A2(n19531), .B1(n19189), .B2(n19530), .ZN(
        n19175) );
  OAI211_X1 U22179 ( .C1(n19193), .C2(n19177), .A(n19176), .B(n19175), .ZN(
        P2_U3067) );
  INV_X1 U22180 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n19180) );
  AOI22_X1 U22181 ( .A1(n19188), .A2(n19566), .B1(n19187), .B2(n19565), .ZN(
        n19179) );
  AOI22_X1 U22182 ( .A1(n19224), .A2(n19568), .B1(n19189), .B2(n19567), .ZN(
        n19178) );
  OAI211_X1 U22183 ( .C1(n19193), .C2(n19180), .A(n19179), .B(n19178), .ZN(
        P2_U3068) );
  INV_X1 U22184 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n19183) );
  AOI22_X1 U22185 ( .A1(n19188), .A2(n19573), .B1(n19572), .B2(n19187), .ZN(
        n19182) );
  AOI22_X1 U22186 ( .A1(n19224), .A2(n19575), .B1(n19189), .B2(n19574), .ZN(
        n19181) );
  OAI211_X1 U22187 ( .C1(n19193), .C2(n19183), .A(n19182), .B(n19181), .ZN(
        P2_U3069) );
  INV_X1 U22188 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n19186) );
  AOI22_X1 U22189 ( .A1(n19188), .A2(n19580), .B1(n19187), .B2(n19579), .ZN(
        n19185) );
  AOI22_X1 U22190 ( .A1(n19189), .A2(n19582), .B1(n19224), .B2(n19581), .ZN(
        n19184) );
  OAI211_X1 U22191 ( .C1(n19193), .C2(n19186), .A(n19185), .B(n19184), .ZN(
        P2_U3070) );
  INV_X1 U22192 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19192) );
  AOI22_X1 U22193 ( .A1(n19188), .A2(n19588), .B1(n19586), .B2(n19187), .ZN(
        n19191) );
  AOI22_X1 U22194 ( .A1(n19189), .A2(n19592), .B1(n19224), .B2(n19590), .ZN(
        n19190) );
  OAI211_X1 U22195 ( .C1(n19193), .C2(n19192), .A(n19191), .B(n19190), .ZN(
        P2_U3071) );
  NOR2_X1 U22196 ( .A1(n19705), .A2(n19195), .ZN(n19203) );
  INV_X1 U22197 ( .A(n19203), .ZN(n19194) );
  NOR2_X1 U22198 ( .A1(n19194), .A2(n19684), .ZN(n19200) );
  INV_X1 U22199 ( .A(n19201), .ZN(n19198) );
  NOR2_X1 U22200 ( .A1(n19196), .A2(n19195), .ZN(n19223) );
  INV_X1 U22201 ( .A(n19223), .ZN(n19197) );
  AOI21_X1 U22202 ( .B1(n19198), .B2(n19197), .A(n19733), .ZN(n19199) );
  AOI22_X1 U22203 ( .A1(n19224), .A2(n19512), .B1(n19511), .B2(n19223), .ZN(
        n19210) );
  AOI21_X1 U22204 ( .B1(n19201), .B2(n19731), .A(n19223), .ZN(n19206) );
  INV_X1 U22205 ( .A(n19298), .ZN(n19202) );
  NOR2_X1 U22206 ( .A1(n19202), .A2(n19208), .ZN(n19204) );
  NOR2_X1 U22207 ( .A1(n19204), .A2(n19203), .ZN(n19205) );
  MUX2_X1 U22208 ( .A(n19206), .B(n19205), .S(n19682), .Z(n19207) );
  AOI22_X1 U22209 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19225), .B1(
        n19259), .B2(n19519), .ZN(n19209) );
  OAI211_X1 U22210 ( .C1(n19228), .C2(n19522), .A(n19210), .B(n19209), .ZN(
        P2_U3072) );
  AOI22_X1 U22211 ( .A1(n19224), .A2(n19554), .B1(n19551), .B2(n19223), .ZN(
        n19212) );
  AOI22_X1 U22212 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19225), .B1(
        n19259), .B2(n19553), .ZN(n19211) );
  OAI211_X1 U22213 ( .C1(n19228), .C2(n19525), .A(n19212), .B(n19211), .ZN(
        P2_U3073) );
  AOI22_X1 U22214 ( .A1(n19259), .A2(n19560), .B1(n19558), .B2(n19223), .ZN(
        n19214) );
  AOI22_X1 U22215 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19225), .B1(
        n19224), .B2(n19561), .ZN(n19213) );
  OAI211_X1 U22216 ( .C1(n19228), .C2(n19528), .A(n19214), .B(n19213), .ZN(
        P2_U3074) );
  AOI22_X1 U22217 ( .A1(n19259), .A2(n19531), .B1(n19529), .B2(n19223), .ZN(
        n19216) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19225), .B1(
        n19224), .B2(n19530), .ZN(n19215) );
  OAI211_X1 U22219 ( .C1(n19228), .C2(n19534), .A(n19216), .B(n19215), .ZN(
        P2_U3075) );
  AOI22_X1 U22220 ( .A1(n19259), .A2(n19568), .B1(n19565), .B2(n19223), .ZN(
        n19218) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19225), .B1(
        n19224), .B2(n19567), .ZN(n19217) );
  OAI211_X1 U22222 ( .C1(n19228), .C2(n19537), .A(n19218), .B(n19217), .ZN(
        P2_U3076) );
  AOI22_X1 U22223 ( .A1(n19224), .A2(n19574), .B1(n19572), .B2(n19223), .ZN(
        n19220) );
  AOI22_X1 U22224 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19225), .B1(
        n19259), .B2(n19575), .ZN(n19219) );
  OAI211_X1 U22225 ( .C1(n19228), .C2(n19540), .A(n19220), .B(n19219), .ZN(
        P2_U3077) );
  AOI22_X1 U22226 ( .A1(n19224), .A2(n19582), .B1(n19579), .B2(n19223), .ZN(
        n19222) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19225), .B1(
        n19259), .B2(n19581), .ZN(n19221) );
  OAI211_X1 U22228 ( .C1(n19228), .C2(n19543), .A(n19222), .B(n19221), .ZN(
        P2_U3078) );
  AOI22_X1 U22229 ( .A1(n19259), .A2(n19590), .B1(n19586), .B2(n19223), .ZN(
        n19227) );
  AOI22_X1 U22230 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19225), .B1(
        n19224), .B2(n19592), .ZN(n19226) );
  OAI211_X1 U22231 ( .C1(n19228), .C2(n19549), .A(n19227), .B(n19226), .ZN(
        P2_U3079) );
  INV_X1 U22232 ( .A(n19229), .ZN(n19436) );
  NAND2_X1 U22233 ( .A1(n19690), .A2(n19436), .ZN(n19237) );
  INV_X1 U22234 ( .A(n19230), .ZN(n19233) );
  NOR2_X1 U22235 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19231), .ZN(
        n19257) );
  OAI21_X1 U22236 ( .B1(n11973), .B2(n19257), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19232) );
  OAI21_X1 U22237 ( .B1(n19237), .B2(n19233), .A(n19232), .ZN(n19258) );
  AOI22_X1 U22238 ( .A1(n19258), .A2(n19467), .B1(n19511), .B2(n19257), .ZN(
        n19242) );
  INV_X1 U22239 ( .A(n19257), .ZN(n19234) );
  OAI211_X1 U22240 ( .C1(n19235), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19234), 
        .B(n19684), .ZN(n19240) );
  INV_X1 U22241 ( .A(n19437), .ZN(n19238) );
  OAI21_X1 U22242 ( .B1(n19259), .B2(n19251), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19236) );
  OAI21_X1 U22243 ( .B1(n19238), .B2(n19237), .A(n19236), .ZN(n19239) );
  NAND3_X1 U22244 ( .A1(n19240), .A2(n19516), .A3(n19239), .ZN(n19260) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19260), .B1(
        n19251), .B2(n19519), .ZN(n19241) );
  OAI211_X1 U22246 ( .C1(n19478), .C2(n19254), .A(n19242), .B(n19241), .ZN(
        P2_U3080) );
  INV_X1 U22247 ( .A(n19251), .ZN(n19263) );
  AOI22_X1 U22248 ( .A1(n19258), .A2(n19552), .B1(n19551), .B2(n19257), .ZN(
        n19244) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19260), .B1(
        n19259), .B2(n19554), .ZN(n19243) );
  OAI211_X1 U22250 ( .C1(n19481), .C2(n19263), .A(n19244), .B(n19243), .ZN(
        P2_U3081) );
  AOI22_X1 U22251 ( .A1(n19258), .A2(n19559), .B1(n19257), .B2(n19558), .ZN(
        n19246) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19260), .B1(
        n19259), .B2(n19561), .ZN(n19245) );
  OAI211_X1 U22253 ( .C1(n19484), .C2(n19263), .A(n19246), .B(n19245), .ZN(
        P2_U3082) );
  AOI22_X1 U22254 ( .A1(n19258), .A2(n19485), .B1(n19529), .B2(n19257), .ZN(
        n19248) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19260), .B1(
        n19251), .B2(n19531), .ZN(n19247) );
  OAI211_X1 U22256 ( .C1(n19488), .C2(n19254), .A(n19248), .B(n19247), .ZN(
        P2_U3083) );
  AOI22_X1 U22257 ( .A1(n19258), .A2(n19566), .B1(n19257), .B2(n19565), .ZN(
        n19250) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19260), .B1(
        n19251), .B2(n19568), .ZN(n19249) );
  OAI211_X1 U22259 ( .C1(n19452), .C2(n19254), .A(n19250), .B(n19249), .ZN(
        P2_U3084) );
  AOI22_X1 U22260 ( .A1(n19258), .A2(n19573), .B1(n19572), .B2(n19257), .ZN(
        n19253) );
  AOI22_X1 U22261 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19260), .B1(
        n19251), .B2(n19575), .ZN(n19252) );
  OAI211_X1 U22262 ( .C1(n19495), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        P2_U3085) );
  AOI22_X1 U22263 ( .A1(n19258), .A2(n19580), .B1(n19257), .B2(n19579), .ZN(
        n19256) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19260), .B1(
        n19259), .B2(n19582), .ZN(n19255) );
  OAI211_X1 U22265 ( .C1(n19498), .C2(n19263), .A(n19256), .B(n19255), .ZN(
        P2_U3086) );
  AOI22_X1 U22266 ( .A1(n19258), .A2(n19588), .B1(n19586), .B2(n19257), .ZN(
        n19262) );
  AOI22_X1 U22267 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19260), .B1(
        n19259), .B2(n19592), .ZN(n19261) );
  OAI211_X1 U22268 ( .C1(n19505), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U3087) );
  INV_X1 U22269 ( .A(n19290), .ZN(n19285) );
  NOR2_X1 U22270 ( .A1(n19387), .A2(n19268), .ZN(n19288) );
  OAI21_X1 U22271 ( .B1(n19268), .B2(n19389), .A(n19264), .ZN(n19289) );
  AOI22_X1 U22272 ( .A1(n19289), .A2(n19467), .B1(n19511), .B2(n19288), .ZN(
        n19274) );
  OAI21_X1 U22273 ( .B1(n19290), .B2(n19321), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19267) );
  OAI21_X1 U22274 ( .B1(n19436), .B2(n19268), .A(n19267), .ZN(n19272) );
  INV_X1 U22275 ( .A(n19288), .ZN(n19269) );
  OAI211_X1 U22276 ( .C1(n19270), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19269), 
        .B(n19684), .ZN(n19271) );
  NAND3_X1 U22277 ( .A1(n19272), .A2(n19516), .A3(n19271), .ZN(n19291) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19291), .B1(
        n19321), .B2(n19519), .ZN(n19273) );
  OAI211_X1 U22279 ( .C1(n19478), .C2(n19285), .A(n19274), .B(n19273), .ZN(
        P2_U3096) );
  AOI22_X1 U22280 ( .A1(n19289), .A2(n19552), .B1(n19551), .B2(n19288), .ZN(
        n19276) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19554), .ZN(n19275) );
  OAI211_X1 U22282 ( .C1(n19481), .C2(n19317), .A(n19276), .B(n19275), .ZN(
        P2_U3097) );
  AOI22_X1 U22283 ( .A1(n19289), .A2(n19559), .B1(n19288), .B2(n19558), .ZN(
        n19278) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19561), .ZN(n19277) );
  OAI211_X1 U22285 ( .C1(n19484), .C2(n19317), .A(n19278), .B(n19277), .ZN(
        P2_U3098) );
  AOI22_X1 U22286 ( .A1(n19289), .A2(n19485), .B1(n19529), .B2(n19288), .ZN(
        n19280) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19291), .B1(
        n19321), .B2(n19531), .ZN(n19279) );
  OAI211_X1 U22288 ( .C1(n19488), .C2(n19285), .A(n19280), .B(n19279), .ZN(
        P2_U3099) );
  AOI22_X1 U22289 ( .A1(n19289), .A2(n19566), .B1(n19288), .B2(n19565), .ZN(
        n19282) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19567), .ZN(n19281) );
  OAI211_X1 U22291 ( .C1(n19491), .C2(n19317), .A(n19282), .B(n19281), .ZN(
        P2_U3100) );
  AOI22_X1 U22292 ( .A1(n19289), .A2(n19573), .B1(n19572), .B2(n19288), .ZN(
        n19284) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19291), .B1(
        n19321), .B2(n19575), .ZN(n19283) );
  OAI211_X1 U22294 ( .C1(n19495), .C2(n19285), .A(n19284), .B(n19283), .ZN(
        P2_U3101) );
  AOI22_X1 U22295 ( .A1(n19289), .A2(n19580), .B1(n19288), .B2(n19579), .ZN(
        n19287) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19582), .ZN(n19286) );
  OAI211_X1 U22297 ( .C1(n19498), .C2(n19317), .A(n19287), .B(n19286), .ZN(
        P2_U3102) );
  AOI22_X1 U22298 ( .A1(n19289), .A2(n19588), .B1(n19586), .B2(n19288), .ZN(
        n19293) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19291), .B1(
        n19290), .B2(n19592), .ZN(n19292) );
  OAI211_X1 U22300 ( .C1(n19505), .C2(n19317), .A(n19293), .B(n19292), .ZN(
        P2_U3103) );
  NAND2_X1 U22301 ( .A1(n19295), .A2(n19294), .ZN(n19327) );
  NAND3_X1 U22302 ( .A1(n11968), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19327), 
        .ZN(n19301) );
  NAND2_X1 U22303 ( .A1(n19296), .A2(n19690), .ZN(n19299) );
  OAI21_X1 U22304 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19299), .A(n19733), 
        .ZN(n19297) );
  AND2_X1 U22305 ( .A1(n19301), .A2(n19297), .ZN(n19320) );
  INV_X1 U22306 ( .A(n19327), .ZN(n19330) );
  AOI22_X1 U22307 ( .A1(n19320), .A2(n19467), .B1(n19511), .B2(n19330), .ZN(
        n19306) );
  NAND2_X1 U22308 ( .A1(n19303), .A2(n19298), .ZN(n19685) );
  AOI22_X1 U22309 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19327), .B1(n19685), 
        .B2(n19299), .ZN(n19300) );
  NAND3_X1 U22310 ( .A1(n19301), .A2(n19300), .A3(n19516), .ZN(n19322) );
  INV_X1 U22311 ( .A(n19302), .ZN(n19304) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19322), .B1(
        n19349), .B2(n19519), .ZN(n19305) );
  OAI211_X1 U22313 ( .C1(n19478), .C2(n19317), .A(n19306), .B(n19305), .ZN(
        P2_U3104) );
  AOI22_X1 U22314 ( .A1(n19320), .A2(n19552), .B1(n19551), .B2(n19330), .ZN(
        n19308) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19322), .B1(
        n19321), .B2(n19554), .ZN(n19307) );
  OAI211_X1 U22316 ( .C1(n19481), .C2(n19345), .A(n19308), .B(n19307), .ZN(
        P2_U3105) );
  AOI22_X1 U22317 ( .A1(n19320), .A2(n19559), .B1(n19330), .B2(n19558), .ZN(
        n19310) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19322), .B1(
        n19321), .B2(n19561), .ZN(n19309) );
  OAI211_X1 U22319 ( .C1(n19484), .C2(n19345), .A(n19310), .B(n19309), .ZN(
        P2_U3106) );
  AOI22_X1 U22320 ( .A1(n19320), .A2(n19485), .B1(n19529), .B2(n19330), .ZN(
        n19312) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19322), .B1(
        n19349), .B2(n19531), .ZN(n19311) );
  OAI211_X1 U22322 ( .C1(n19488), .C2(n19317), .A(n19312), .B(n19311), .ZN(
        P2_U3107) );
  AOI22_X1 U22323 ( .A1(n19320), .A2(n19566), .B1(n19330), .B2(n19565), .ZN(
        n19314) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19322), .B1(
        n19321), .B2(n19567), .ZN(n19313) );
  OAI211_X1 U22325 ( .C1(n19491), .C2(n19345), .A(n19314), .B(n19313), .ZN(
        P2_U3108) );
  AOI22_X1 U22326 ( .A1(n19320), .A2(n19573), .B1(n19572), .B2(n19330), .ZN(
        n19316) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19322), .B1(
        n19349), .B2(n19575), .ZN(n19315) );
  OAI211_X1 U22328 ( .C1(n19495), .C2(n19317), .A(n19316), .B(n19315), .ZN(
        P2_U3109) );
  AOI22_X1 U22329 ( .A1(n19320), .A2(n19580), .B1(n19330), .B2(n19579), .ZN(
        n19319) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19322), .B1(
        n19321), .B2(n19582), .ZN(n19318) );
  OAI211_X1 U22331 ( .C1(n19498), .C2(n19345), .A(n19319), .B(n19318), .ZN(
        P2_U3110) );
  AOI22_X1 U22332 ( .A1(n19320), .A2(n19588), .B1(n19586), .B2(n19330), .ZN(
        n19324) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19322), .B1(
        n19321), .B2(n19592), .ZN(n19323) );
  OAI211_X1 U22334 ( .C1(n19505), .C2(n19345), .A(n19324), .B(n19323), .ZN(
        P2_U3111) );
  NOR2_X1 U22335 ( .A1(n19390), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19355) );
  AND2_X1 U22336 ( .A1(n19714), .A2(n19355), .ZN(n19348) );
  AOI22_X1 U22337 ( .A1(n19382), .A2(n19519), .B1(n19511), .B2(n19348), .ZN(
        n19334) );
  NAND2_X1 U22338 ( .A1(n19345), .A2(n19354), .ZN(n19325) );
  AOI21_X1 U22339 ( .B1(n19325), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19684), 
        .ZN(n19329) );
  AOI21_X1 U22340 ( .B1(n11960), .B2(n19731), .A(n19682), .ZN(n19326) );
  AOI21_X1 U22341 ( .B1(n19329), .B2(n19327), .A(n19326), .ZN(n19328) );
  OAI21_X1 U22342 ( .B1(n19348), .B2(n19328), .A(n19516), .ZN(n19351) );
  OAI21_X1 U22343 ( .B1(n19330), .B2(n19348), .A(n19329), .ZN(n19332) );
  OAI21_X1 U22344 ( .B1(n11960), .B2(n19348), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19331) );
  NAND2_X1 U22345 ( .A1(n19332), .A2(n19331), .ZN(n19350) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19351), .B1(
        n19467), .B2(n19350), .ZN(n19333) );
  OAI211_X1 U22347 ( .C1(n19478), .C2(n19345), .A(n19334), .B(n19333), .ZN(
        P2_U3112) );
  AOI22_X1 U22348 ( .A1(n19349), .A2(n19554), .B1(n19551), .B2(n19348), .ZN(
        n19336) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19552), .ZN(n19335) );
  OAI211_X1 U22350 ( .C1(n19481), .C2(n19354), .A(n19336), .B(n19335), .ZN(
        P2_U3113) );
  AOI22_X1 U22351 ( .A1(n19349), .A2(n19561), .B1(n19558), .B2(n19348), .ZN(
        n19338) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19559), .ZN(n19337) );
  OAI211_X1 U22353 ( .C1(n19484), .C2(n19354), .A(n19338), .B(n19337), .ZN(
        P2_U3114) );
  AOI22_X1 U22354 ( .A1(n19382), .A2(n19531), .B1(n19529), .B2(n19348), .ZN(
        n19340) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19485), .ZN(n19339) );
  OAI211_X1 U22356 ( .C1(n19488), .C2(n19345), .A(n19340), .B(n19339), .ZN(
        P2_U3115) );
  AOI22_X1 U22357 ( .A1(n19382), .A2(n19568), .B1(n19565), .B2(n19348), .ZN(
        n19342) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19566), .ZN(n19341) );
  OAI211_X1 U22359 ( .C1(n19452), .C2(n19345), .A(n19342), .B(n19341), .ZN(
        P2_U3116) );
  AOI22_X1 U22360 ( .A1(n19382), .A2(n19575), .B1(n19572), .B2(n19348), .ZN(
        n19344) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19573), .ZN(n19343) );
  OAI211_X1 U22362 ( .C1(n19495), .C2(n19345), .A(n19344), .B(n19343), .ZN(
        P2_U3117) );
  AOI22_X1 U22363 ( .A1(n19349), .A2(n19582), .B1(n19579), .B2(n19348), .ZN(
        n19347) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19580), .ZN(n19346) );
  OAI211_X1 U22365 ( .C1(n19498), .C2(n19354), .A(n19347), .B(n19346), .ZN(
        P2_U3118) );
  AOI22_X1 U22366 ( .A1(n19349), .A2(n19592), .B1(n19586), .B2(n19348), .ZN(
        n19353) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19351), .B1(
        n19350), .B2(n19588), .ZN(n19352) );
  OAI211_X1 U22368 ( .C1(n19505), .C2(n19354), .A(n19353), .B(n19352), .ZN(
        P2_U3119) );
  INV_X1 U22369 ( .A(n19355), .ZN(n19362) );
  NOR2_X1 U22370 ( .A1(n19684), .A2(n19362), .ZN(n19358) );
  NOR2_X1 U22371 ( .A1(n19356), .A2(n19390), .ZN(n19391) );
  INV_X1 U22372 ( .A(n19391), .ZN(n19359) );
  AOI21_X1 U22373 ( .B1(n19360), .B2(n19359), .A(n19733), .ZN(n19357) );
  NOR2_X1 U22374 ( .A1(n19358), .A2(n19357), .ZN(n19386) );
  AOI22_X1 U22375 ( .A1(n19382), .A2(n19512), .B1(n19511), .B2(n19391), .ZN(
        n19369) );
  OAI21_X1 U22376 ( .B1(n19360), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19359), 
        .ZN(n19365) );
  NAND2_X1 U22377 ( .A1(n19471), .A2(n19361), .ZN(n19363) );
  NAND2_X1 U22378 ( .A1(n19363), .A2(n19362), .ZN(n19364) );
  MUX2_X1 U22379 ( .A(n19365), .B(n19364), .S(n19682), .Z(n19366) );
  NAND2_X1 U22380 ( .A1(n19366), .A2(n19516), .ZN(n19383) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19383), .B1(
        n19412), .B2(n19519), .ZN(n19368) );
  OAI211_X1 U22382 ( .C1(n19386), .C2(n19522), .A(n19369), .B(n19368), .ZN(
        P2_U3120) );
  AOI22_X1 U22383 ( .A1(n19412), .A2(n19553), .B1(n19551), .B2(n19391), .ZN(
        n19371) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19554), .ZN(n19370) );
  OAI211_X1 U22385 ( .C1(n19386), .C2(n19525), .A(n19371), .B(n19370), .ZN(
        P2_U3121) );
  AOI22_X1 U22386 ( .A1(n19412), .A2(n19560), .B1(n19558), .B2(n19391), .ZN(
        n19373) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19561), .ZN(n19372) );
  OAI211_X1 U22388 ( .C1(n19386), .C2(n19528), .A(n19373), .B(n19372), .ZN(
        P2_U3122) );
  AOI22_X1 U22389 ( .A1(n19412), .A2(n19531), .B1(n19529), .B2(n19391), .ZN(
        n19375) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19530), .ZN(n19374) );
  OAI211_X1 U22391 ( .C1(n19386), .C2(n19534), .A(n19375), .B(n19374), .ZN(
        P2_U3123) );
  AOI22_X1 U22392 ( .A1(n19382), .A2(n19567), .B1(n19565), .B2(n19391), .ZN(
        n19377) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19383), .B1(
        n19412), .B2(n19568), .ZN(n19376) );
  OAI211_X1 U22394 ( .C1(n19386), .C2(n19537), .A(n19377), .B(n19376), .ZN(
        P2_U3124) );
  AOI22_X1 U22395 ( .A1(n19412), .A2(n19575), .B1(n19572), .B2(n19391), .ZN(
        n19379) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19383), .B1(
        n19382), .B2(n19574), .ZN(n19378) );
  OAI211_X1 U22397 ( .C1(n19386), .C2(n19540), .A(n19379), .B(n19378), .ZN(
        P2_U3125) );
  AOI22_X1 U22398 ( .A1(n19382), .A2(n19582), .B1(n19579), .B2(n19391), .ZN(
        n19381) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19383), .B1(
        n19412), .B2(n19581), .ZN(n19380) );
  OAI211_X1 U22400 ( .C1(n19386), .C2(n19543), .A(n19381), .B(n19380), .ZN(
        P2_U3126) );
  AOI22_X1 U22401 ( .A1(n19382), .A2(n19592), .B1(n19586), .B2(n19391), .ZN(
        n19385) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19383), .B1(
        n19412), .B2(n19590), .ZN(n19384) );
  OAI211_X1 U22403 ( .C1(n19386), .C2(n19549), .A(n19385), .B(n19384), .ZN(
        P2_U3127) );
  NOR2_X1 U22404 ( .A1(n19387), .A2(n19390), .ZN(n19410) );
  OAI21_X1 U22405 ( .B1(n11959), .B2(n19410), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19388) );
  OAI21_X1 U22406 ( .B1(n19390), .B2(n19389), .A(n19388), .ZN(n19411) );
  AOI22_X1 U22407 ( .A1(n19411), .A2(n19467), .B1(n19511), .B2(n19410), .ZN(
        n19396) );
  INV_X1 U22408 ( .A(n11959), .ZN(n19393) );
  AOI221_X1 U22409 ( .B1(n19429), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19412), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19391), .ZN(n19392) );
  AOI211_X1 U22410 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19393), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19392), .ZN(n19394) );
  OAI21_X1 U22411 ( .B1(n19394), .B2(n19410), .A(n19516), .ZN(n19413) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19413), .B1(
        n19429), .B2(n19519), .ZN(n19395) );
  OAI211_X1 U22413 ( .C1(n19478), .C2(n19407), .A(n19396), .B(n19395), .ZN(
        P2_U3128) );
  AOI22_X1 U22414 ( .A1(n19411), .A2(n19552), .B1(n19551), .B2(n19410), .ZN(
        n19398) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19413), .B1(
        n19412), .B2(n19554), .ZN(n19397) );
  OAI211_X1 U22416 ( .C1(n19481), .C2(n19424), .A(n19398), .B(n19397), .ZN(
        P2_U3129) );
  AOI22_X1 U22417 ( .A1(n19411), .A2(n19559), .B1(n19410), .B2(n19558), .ZN(
        n19400) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19413), .B1(
        n19412), .B2(n19561), .ZN(n19399) );
  OAI211_X1 U22419 ( .C1(n19484), .C2(n19424), .A(n19400), .B(n19399), .ZN(
        P2_U3130) );
  AOI22_X1 U22420 ( .A1(n19411), .A2(n19485), .B1(n19529), .B2(n19410), .ZN(
        n19402) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19413), .B1(
        n19429), .B2(n19531), .ZN(n19401) );
  OAI211_X1 U22422 ( .C1(n19488), .C2(n19407), .A(n19402), .B(n19401), .ZN(
        P2_U3131) );
  AOI22_X1 U22423 ( .A1(n19411), .A2(n19566), .B1(n19410), .B2(n19565), .ZN(
        n19404) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19413), .B1(
        n19429), .B2(n19568), .ZN(n19403) );
  OAI211_X1 U22425 ( .C1(n19452), .C2(n19407), .A(n19404), .B(n19403), .ZN(
        P2_U3132) );
  AOI22_X1 U22426 ( .A1(n19411), .A2(n19573), .B1(n19572), .B2(n19410), .ZN(
        n19406) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19413), .B1(
        n19429), .B2(n19575), .ZN(n19405) );
  OAI211_X1 U22428 ( .C1(n19495), .C2(n19407), .A(n19406), .B(n19405), .ZN(
        P2_U3133) );
  AOI22_X1 U22429 ( .A1(n19411), .A2(n19580), .B1(n19410), .B2(n19579), .ZN(
        n19409) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19413), .B1(
        n19412), .B2(n19582), .ZN(n19408) );
  OAI211_X1 U22431 ( .C1(n19498), .C2(n19424), .A(n19409), .B(n19408), .ZN(
        P2_U3134) );
  AOI22_X1 U22432 ( .A1(n19411), .A2(n19588), .B1(n19586), .B2(n19410), .ZN(
        n19415) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19413), .B1(
        n19412), .B2(n19592), .ZN(n19414) );
  OAI211_X1 U22434 ( .C1(n19505), .C2(n19424), .A(n19415), .B(n19414), .ZN(
        P2_U3135) );
  AOI22_X1 U22435 ( .A1(n19428), .A2(n19552), .B1(n19551), .B2(n19427), .ZN(
        n19417) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19554), .ZN(n19416) );
  OAI211_X1 U22437 ( .C1(n19481), .C2(n19455), .A(n19417), .B(n19416), .ZN(
        P2_U3137) );
  AOI22_X1 U22438 ( .A1(n19428), .A2(n19559), .B1(n19427), .B2(n19558), .ZN(
        n19419) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19561), .ZN(n19418) );
  OAI211_X1 U22440 ( .C1(n19484), .C2(n19455), .A(n19419), .B(n19418), .ZN(
        P2_U3138) );
  AOI22_X1 U22441 ( .A1(n19428), .A2(n19566), .B1(n19427), .B2(n19565), .ZN(
        n19421) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19430), .B1(
        n19460), .B2(n19568), .ZN(n19420) );
  OAI211_X1 U22443 ( .C1(n19452), .C2(n19424), .A(n19421), .B(n19420), .ZN(
        P2_U3140) );
  AOI22_X1 U22444 ( .A1(n19428), .A2(n19573), .B1(n19572), .B2(n19427), .ZN(
        n19423) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19430), .B1(
        n19460), .B2(n19575), .ZN(n19422) );
  OAI211_X1 U22446 ( .C1(n19495), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U3141) );
  AOI22_X1 U22447 ( .A1(n19428), .A2(n19580), .B1(n19427), .B2(n19579), .ZN(
        n19426) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19582), .ZN(n19425) );
  OAI211_X1 U22449 ( .C1(n19498), .C2(n19455), .A(n19426), .B(n19425), .ZN(
        P2_U3142) );
  AOI22_X1 U22450 ( .A1(n19428), .A2(n19588), .B1(n19586), .B2(n19427), .ZN(
        n19432) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19430), .B1(
        n19429), .B2(n19592), .ZN(n19431) );
  OAI211_X1 U22452 ( .C1(n19505), .C2(n19455), .A(n19432), .B(n19431), .ZN(
        P2_U3143) );
  NAND4_X1 U22453 ( .A1(n19437), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19436), .A4(n19731), .ZN(n19434) );
  NAND3_X1 U22454 ( .A1(n19705), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19465) );
  NOR2_X1 U22455 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19465), .ZN(
        n19458) );
  NOR3_X1 U22456 ( .A1(n19433), .A2(n19458), .A3(n19733), .ZN(n19438) );
  AOI21_X1 U22457 ( .B1(n19733), .B2(n19434), .A(n19438), .ZN(n19459) );
  AOI22_X1 U22458 ( .A1(n19459), .A2(n19467), .B1(n19511), .B2(n19458), .ZN(
        n19443) );
  OAI21_X1 U22459 ( .B1(n19460), .B2(n19501), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19440) );
  NAND3_X1 U22460 ( .A1(n19437), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19436), .ZN(n19439) );
  AOI211_X1 U22461 ( .C1(n19440), .C2(n19439), .A(n19469), .B(n19438), .ZN(
        n19441) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19461), .B1(
        n19501), .B2(n19519), .ZN(n19442) );
  OAI211_X1 U22463 ( .C1(n19478), .C2(n19455), .A(n19443), .B(n19442), .ZN(
        P2_U3144) );
  AOI22_X1 U22464 ( .A1(n19459), .A2(n19552), .B1(n19551), .B2(n19458), .ZN(
        n19445) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19461), .B1(
        n19460), .B2(n19554), .ZN(n19444) );
  OAI211_X1 U22466 ( .C1(n19481), .C2(n19494), .A(n19445), .B(n19444), .ZN(
        P2_U3145) );
  AOI22_X1 U22467 ( .A1(n19459), .A2(n19559), .B1(n19458), .B2(n19558), .ZN(
        n19447) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19461), .B1(
        n19460), .B2(n19561), .ZN(n19446) );
  OAI211_X1 U22469 ( .C1(n19484), .C2(n19494), .A(n19447), .B(n19446), .ZN(
        P2_U3146) );
  AOI22_X1 U22470 ( .A1(n19459), .A2(n19485), .B1(n19529), .B2(n19458), .ZN(
        n19449) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19461), .B1(
        n19501), .B2(n19531), .ZN(n19448) );
  OAI211_X1 U22472 ( .C1(n19488), .C2(n19455), .A(n19449), .B(n19448), .ZN(
        P2_U3147) );
  AOI22_X1 U22473 ( .A1(n19459), .A2(n19566), .B1(n19458), .B2(n19565), .ZN(
        n19451) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19461), .B1(
        n19501), .B2(n19568), .ZN(n19450) );
  OAI211_X1 U22475 ( .C1(n19452), .C2(n19455), .A(n19451), .B(n19450), .ZN(
        P2_U3148) );
  AOI22_X1 U22476 ( .A1(n19459), .A2(n19573), .B1(n19572), .B2(n19458), .ZN(
        n19454) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19461), .B1(
        n19501), .B2(n19575), .ZN(n19453) );
  OAI211_X1 U22478 ( .C1(n19495), .C2(n19455), .A(n19454), .B(n19453), .ZN(
        P2_U3149) );
  AOI22_X1 U22479 ( .A1(n19459), .A2(n19580), .B1(n19458), .B2(n19579), .ZN(
        n19457) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19461), .B1(
        n19460), .B2(n19582), .ZN(n19456) );
  OAI211_X1 U22481 ( .C1(n19498), .C2(n19494), .A(n19457), .B(n19456), .ZN(
        P2_U3150) );
  AOI22_X1 U22482 ( .A1(n19459), .A2(n19588), .B1(n19586), .B2(n19458), .ZN(
        n19463) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19461), .B1(
        n19460), .B2(n19592), .ZN(n19462) );
  OAI211_X1 U22484 ( .C1(n19505), .C2(n19494), .A(n19463), .B(n19462), .ZN(
        P2_U3151) );
  NOR2_X1 U22485 ( .A1(n19714), .A2(n19465), .ZN(n19499) );
  NOR3_X1 U22486 ( .A1(n19464), .A2(n19499), .A3(n19733), .ZN(n19468) );
  INV_X1 U22487 ( .A(n19465), .ZN(n19473) );
  AOI21_X1 U22488 ( .B1(n19731), .B2(n19473), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19466) );
  NOR2_X1 U22489 ( .A1(n19468), .A2(n19466), .ZN(n19500) );
  AOI22_X1 U22490 ( .A1(n19500), .A2(n19467), .B1(n19511), .B2(n19499), .ZN(
        n19477) );
  INV_X1 U22491 ( .A(n19499), .ZN(n19509) );
  AOI211_X1 U22492 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19509), .A(n19469), 
        .B(n19468), .ZN(n19470) );
  OAI221_X1 U22493 ( .B1(n19473), .B2(n19472), .C1(n19473), .C2(n19471), .A(
        n19470), .ZN(n19502) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19502), .B1(
        n19545), .B2(n19519), .ZN(n19476) );
  OAI211_X1 U22495 ( .C1(n19478), .C2(n19494), .A(n19477), .B(n19476), .ZN(
        P2_U3152) );
  AOI22_X1 U22496 ( .A1(n19500), .A2(n19552), .B1(n19551), .B2(n19499), .ZN(
        n19480) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19502), .B1(
        n19501), .B2(n19554), .ZN(n19479) );
  OAI211_X1 U22498 ( .C1(n19481), .C2(n19506), .A(n19480), .B(n19479), .ZN(
        P2_U3153) );
  AOI22_X1 U22499 ( .A1(n19500), .A2(n19559), .B1(n19499), .B2(n19558), .ZN(
        n19483) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19502), .B1(
        n19501), .B2(n19561), .ZN(n19482) );
  OAI211_X1 U22501 ( .C1(n19484), .C2(n19506), .A(n19483), .B(n19482), .ZN(
        P2_U3154) );
  AOI22_X1 U22502 ( .A1(n19500), .A2(n19485), .B1(n19529), .B2(n19499), .ZN(
        n19487) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19502), .B1(
        n19545), .B2(n19531), .ZN(n19486) );
  OAI211_X1 U22504 ( .C1(n19488), .C2(n19494), .A(n19487), .B(n19486), .ZN(
        P2_U3155) );
  AOI22_X1 U22505 ( .A1(n19500), .A2(n19566), .B1(n19499), .B2(n19565), .ZN(
        n19490) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19502), .B1(
        n19501), .B2(n19567), .ZN(n19489) );
  OAI211_X1 U22507 ( .C1(n19491), .C2(n19506), .A(n19490), .B(n19489), .ZN(
        P2_U3156) );
  AOI22_X1 U22508 ( .A1(n19500), .A2(n19573), .B1(n19572), .B2(n19499), .ZN(
        n19493) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19502), .B1(
        n19545), .B2(n19575), .ZN(n19492) );
  OAI211_X1 U22510 ( .C1(n19495), .C2(n19494), .A(n19493), .B(n19492), .ZN(
        P2_U3157) );
  AOI22_X1 U22511 ( .A1(n19500), .A2(n19580), .B1(n19499), .B2(n19579), .ZN(
        n19497) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19502), .B1(
        n19501), .B2(n19582), .ZN(n19496) );
  OAI211_X1 U22513 ( .C1(n19498), .C2(n19506), .A(n19497), .B(n19496), .ZN(
        P2_U3158) );
  AOI22_X1 U22514 ( .A1(n19500), .A2(n19588), .B1(n19586), .B2(n19499), .ZN(
        n19504) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19502), .B1(
        n19501), .B2(n19592), .ZN(n19503) );
  OAI211_X1 U22516 ( .C1(n19505), .C2(n19506), .A(n19504), .B(n19503), .ZN(
        P2_U3159) );
  NAND2_X1 U22517 ( .A1(n19506), .A2(n19682), .ZN(n19507) );
  OAI21_X1 U22518 ( .B1(n19507), .B2(n19593), .A(n19681), .ZN(n19513) );
  NOR3_X2 U22519 ( .A1(n19690), .A2(n19508), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19544) );
  INV_X1 U22520 ( .A(n19544), .ZN(n19514) );
  NAND2_X1 U22521 ( .A1(n19514), .A2(n19509), .ZN(n19517) );
  AOI21_X1 U22522 ( .B1(n11943), .B2(n19514), .A(n19733), .ZN(n19510) );
  AOI22_X1 U22523 ( .A1(n19545), .A2(n19512), .B1(n19511), .B2(n19544), .ZN(
        n19521) );
  INV_X1 U22524 ( .A(n19513), .ZN(n19518) );
  OAI211_X1 U22525 ( .C1(n11943), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19514), 
        .B(n19684), .ZN(n19515) );
  OAI211_X1 U22526 ( .C1(n19518), .C2(n19517), .A(n19516), .B(n19515), .ZN(
        n19546) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19546), .B1(
        n19593), .B2(n19519), .ZN(n19520) );
  OAI211_X1 U22528 ( .C1(n19550), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P2_U3160) );
  AOI22_X1 U22529 ( .A1(n19545), .A2(n19554), .B1(n19551), .B2(n19544), .ZN(
        n19524) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19546), .B1(
        n19593), .B2(n19553), .ZN(n19523) );
  OAI211_X1 U22531 ( .C1(n19550), .C2(n19525), .A(n19524), .B(n19523), .ZN(
        P2_U3161) );
  AOI22_X1 U22532 ( .A1(n19593), .A2(n19560), .B1(n19558), .B2(n19544), .ZN(
        n19527) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19561), .ZN(n19526) );
  OAI211_X1 U22534 ( .C1(n19550), .C2(n19528), .A(n19527), .B(n19526), .ZN(
        P2_U3162) );
  AOI22_X1 U22535 ( .A1(n19545), .A2(n19530), .B1(n19529), .B2(n19544), .ZN(
        n19533) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19546), .B1(
        n19593), .B2(n19531), .ZN(n19532) );
  OAI211_X1 U22537 ( .C1(n19550), .C2(n19534), .A(n19533), .B(n19532), .ZN(
        P2_U3163) );
  AOI22_X1 U22538 ( .A1(n19593), .A2(n19568), .B1(n19565), .B2(n19544), .ZN(
        n19536) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19567), .ZN(n19535) );
  OAI211_X1 U22540 ( .C1(n19550), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P2_U3164) );
  AOI22_X1 U22541 ( .A1(n19545), .A2(n19574), .B1(n19572), .B2(n19544), .ZN(
        n19539) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19546), .B1(
        n19593), .B2(n19575), .ZN(n19538) );
  OAI211_X1 U22543 ( .C1(n19550), .C2(n19540), .A(n19539), .B(n19538), .ZN(
        P2_U3165) );
  AOI22_X1 U22544 ( .A1(n19593), .A2(n19581), .B1(n19579), .B2(n19544), .ZN(
        n19542) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19546), .B1(
        n19545), .B2(n19582), .ZN(n19541) );
  OAI211_X1 U22546 ( .C1(n19550), .C2(n19543), .A(n19542), .B(n19541), .ZN(
        P2_U3166) );
  AOI22_X1 U22547 ( .A1(n19545), .A2(n19592), .B1(n19586), .B2(n19544), .ZN(
        n19548) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19546), .B1(
        n19593), .B2(n19590), .ZN(n19547) );
  OAI211_X1 U22549 ( .C1(n19550), .C2(n19549), .A(n19548), .B(n19547), .ZN(
        P2_U3167) );
  INV_X1 U22550 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n19557) );
  AOI22_X1 U22551 ( .A1(n19589), .A2(n19552), .B1(n19587), .B2(n19551), .ZN(
        n19556) );
  AOI22_X1 U22552 ( .A1(n19593), .A2(n19554), .B1(n19591), .B2(n19553), .ZN(
        n19555) );
  OAI211_X1 U22553 ( .C1(n19597), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P2_U3169) );
  INV_X1 U22554 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n19564) );
  AOI22_X1 U22555 ( .A1(n19589), .A2(n19559), .B1(n19587), .B2(n19558), .ZN(
        n19563) );
  AOI22_X1 U22556 ( .A1(n19593), .A2(n19561), .B1(n19591), .B2(n19560), .ZN(
        n19562) );
  OAI211_X1 U22557 ( .C1(n19597), .C2(n19564), .A(n19563), .B(n19562), .ZN(
        P2_U3170) );
  INV_X1 U22558 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n19571) );
  AOI22_X1 U22559 ( .A1(n19589), .A2(n19566), .B1(n19587), .B2(n19565), .ZN(
        n19570) );
  AOI22_X1 U22560 ( .A1(n19591), .A2(n19568), .B1(n19593), .B2(n19567), .ZN(
        n19569) );
  OAI211_X1 U22561 ( .C1(n19597), .C2(n19571), .A(n19570), .B(n19569), .ZN(
        P2_U3172) );
  INV_X1 U22562 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n19578) );
  AOI22_X1 U22563 ( .A1(n19589), .A2(n19573), .B1(n19587), .B2(n19572), .ZN(
        n19577) );
  AOI22_X1 U22564 ( .A1(n19591), .A2(n19575), .B1(n19593), .B2(n19574), .ZN(
        n19576) );
  OAI211_X1 U22565 ( .C1(n19597), .C2(n19578), .A(n19577), .B(n19576), .ZN(
        P2_U3173) );
  AOI22_X1 U22566 ( .A1(n19589), .A2(n19580), .B1(n19587), .B2(n19579), .ZN(
        n19584) );
  AOI22_X1 U22567 ( .A1(n19593), .A2(n19582), .B1(n19591), .B2(n19581), .ZN(
        n19583) );
  OAI211_X1 U22568 ( .C1(n19597), .C2(n19585), .A(n19584), .B(n19583), .ZN(
        P2_U3174) );
  INV_X1 U22569 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19596) );
  AOI22_X1 U22570 ( .A1(n19589), .A2(n19588), .B1(n19587), .B2(n19586), .ZN(
        n19595) );
  AOI22_X1 U22571 ( .A1(n19593), .A2(n19592), .B1(n19591), .B2(n19590), .ZN(
        n19594) );
  OAI211_X1 U22572 ( .C1(n19597), .C2(n19596), .A(n19595), .B(n19594), .ZN(
        P2_U3175) );
  AND2_X1 U22573 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19599), .ZN(
        P2_U3179) );
  AND2_X1 U22574 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19599), .ZN(
        P2_U3180) );
  AND2_X1 U22575 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19599), .ZN(
        P2_U3181) );
  NOR2_X1 U22576 ( .A1(n19598), .A2(n19678), .ZN(P2_U3182) );
  AND2_X1 U22577 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19599), .ZN(
        P2_U3183) );
  AND2_X1 U22578 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19599), .ZN(
        P2_U3184) );
  AND2_X1 U22579 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19599), .ZN(
        P2_U3185) );
  AND2_X1 U22580 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19599), .ZN(
        P2_U3186) );
  AND2_X1 U22581 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19599), .ZN(
        P2_U3187) );
  AND2_X1 U22582 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19599), .ZN(
        P2_U3188) );
  AND2_X1 U22583 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19599), .ZN(
        P2_U3189) );
  NOR2_X1 U22584 ( .A1(n20774), .A2(n19678), .ZN(P2_U3190) );
  AND2_X1 U22585 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19599), .ZN(
        P2_U3191) );
  AND2_X1 U22586 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19599), .ZN(
        P2_U3192) );
  AND2_X1 U22587 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19599), .ZN(
        P2_U3193) );
  AND2_X1 U22588 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19599), .ZN(
        P2_U3194) );
  AND2_X1 U22589 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19599), .ZN(
        P2_U3195) );
  AND2_X1 U22590 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19599), .ZN(
        P2_U3196) );
  AND2_X1 U22591 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19599), .ZN(
        P2_U3197) );
  AND2_X1 U22592 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19599), .ZN(
        P2_U3198) );
  AND2_X1 U22593 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19599), .ZN(
        P2_U3199) );
  AND2_X1 U22594 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19599), .ZN(
        P2_U3200) );
  AND2_X1 U22595 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19599), .ZN(P2_U3201) );
  AND2_X1 U22596 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19599), .ZN(P2_U3202) );
  AND2_X1 U22597 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19599), .ZN(P2_U3203) );
  AND2_X1 U22598 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19599), .ZN(P2_U3204) );
  AND2_X1 U22599 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19599), .ZN(P2_U3205) );
  AND2_X1 U22600 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19599), .ZN(P2_U3206) );
  AND2_X1 U22601 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19599), .ZN(P2_U3207) );
  AND2_X1 U22602 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19599), .ZN(P2_U3208) );
  NOR2_X1 U22603 ( .A1(n19601), .A2(n19600), .ZN(n19611) );
  INV_X1 U22604 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19743) );
  OR3_X1 U22605 ( .A1(n19611), .A2(n19743), .A3(n19614), .ZN(n19603) );
  AOI211_X1 U22606 ( .C1(n20660), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19612), .B(n19744), .ZN(n19602) );
  INV_X1 U22607 ( .A(NA), .ZN(n20658) );
  NOR2_X1 U22608 ( .A1(n20658), .A2(n19605), .ZN(n19618) );
  AOI211_X1 U22609 ( .C1(n19619), .C2(n19603), .A(n19602), .B(n19618), .ZN(
        n19604) );
  INV_X1 U22610 ( .A(n19604), .ZN(P2_U3209) );
  AOI21_X1 U22611 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20660), .A(n19619), 
        .ZN(n19609) );
  NOR2_X1 U22612 ( .A1(n19743), .A2(n19609), .ZN(n19606) );
  AOI21_X1 U22613 ( .B1(n19606), .B2(n19605), .A(n19611), .ZN(n19607) );
  OAI211_X1 U22614 ( .C1(n20660), .C2(n19608), .A(n19607), .B(n19735), .ZN(
        P2_U3210) );
  AOI21_X1 U22615 ( .B1(n19734), .B2(n19610), .A(n19609), .ZN(n19617) );
  AOI22_X1 U22616 ( .A1(n19743), .A2(n19612), .B1(n20658), .B2(n19611), .ZN(
        n19613) );
  AOI211_X1 U22617 ( .C1(n19743), .C2(n20660), .A(n19614), .B(n19613), .ZN(
        n19615) );
  INV_X1 U22618 ( .A(n19615), .ZN(n19616) );
  OAI21_X1 U22619 ( .B1(n19618), .B2(n19617), .A(n19616), .ZN(P2_U3211) );
  OAI222_X1 U22620 ( .A1(n19668), .A2(n19622), .B1(n19621), .B2(n19744), .C1(
        n19620), .C2(n19669), .ZN(P2_U3212) );
  OAI222_X1 U22621 ( .A1(n19668), .A2(n10675), .B1(n19623), .B2(n19744), .C1(
        n19622), .C2(n19669), .ZN(P2_U3213) );
  OAI222_X1 U22622 ( .A1(n19668), .A2(n19625), .B1(n19624), .B2(n19744), .C1(
        n10675), .C2(n19669), .ZN(P2_U3214) );
  OAI222_X1 U22623 ( .A1(n19668), .A2(n10703), .B1(n19626), .B2(n19744), .C1(
        n19625), .C2(n19669), .ZN(P2_U3215) );
  OAI222_X1 U22624 ( .A1(n19668), .A2(n19628), .B1(n19627), .B2(n19744), .C1(
        n10703), .C2(n19669), .ZN(P2_U3216) );
  OAI222_X1 U22625 ( .A1(n19668), .A2(n19630), .B1(n19629), .B2(n19744), .C1(
        n19628), .C2(n19669), .ZN(P2_U3217) );
  OAI222_X1 U22626 ( .A1(n19668), .A2(n13116), .B1(n19631), .B2(n19744), .C1(
        n19630), .C2(n19669), .ZN(P2_U3218) );
  OAI222_X1 U22627 ( .A1(n19668), .A2(n10755), .B1(n19632), .B2(n19744), .C1(
        n13116), .C2(n19669), .ZN(P2_U3219) );
  OAI222_X1 U22628 ( .A1(n19668), .A2(n19634), .B1(n19633), .B2(n19744), .C1(
        n10755), .C2(n19669), .ZN(P2_U3220) );
  OAI222_X1 U22629 ( .A1(n19668), .A2(n10781), .B1(n19635), .B2(n19744), .C1(
        n19634), .C2(n19669), .ZN(P2_U3221) );
  INV_X1 U22630 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19637) );
  INV_X1 U22631 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19636) );
  OAI222_X1 U22632 ( .A1(n19668), .A2(n19637), .B1(n19636), .B2(n19744), .C1(
        n10781), .C2(n19669), .ZN(P2_U3222) );
  OAI222_X1 U22633 ( .A1(n19668), .A2(n20932), .B1(n19638), .B2(n19744), .C1(
        n19637), .C2(n19669), .ZN(P2_U3223) );
  OAI222_X1 U22634 ( .A1(n19668), .A2(n13619), .B1(n19639), .B2(n19744), .C1(
        n20932), .C2(n19669), .ZN(P2_U3224) );
  OAI222_X1 U22635 ( .A1(n19668), .A2(n19641), .B1(n19640), .B2(n19744), .C1(
        n13619), .C2(n19669), .ZN(P2_U3225) );
  OAI222_X1 U22636 ( .A1(n19668), .A2(n10833), .B1(n19642), .B2(n19744), .C1(
        n19641), .C2(n19669), .ZN(P2_U3226) );
  OAI222_X1 U22637 ( .A1(n19668), .A2(n19644), .B1(n19643), .B2(n19744), .C1(
        n10833), .C2(n19669), .ZN(P2_U3227) );
  OAI222_X1 U22638 ( .A1(n19668), .A2(n19646), .B1(n19645), .B2(n19744), .C1(
        n19644), .C2(n19669), .ZN(P2_U3228) );
  OAI222_X1 U22639 ( .A1(n19668), .A2(n19648), .B1(n19647), .B2(n19744), .C1(
        n19646), .C2(n19669), .ZN(P2_U3229) );
  OAI222_X1 U22640 ( .A1(n19668), .A2(n15128), .B1(n19649), .B2(n19744), .C1(
        n19648), .C2(n19669), .ZN(P2_U3230) );
  OAI222_X1 U22641 ( .A1(n19668), .A2(n19651), .B1(n19650), .B2(n19744), .C1(
        n15128), .C2(n19669), .ZN(P2_U3231) );
  OAI222_X1 U22642 ( .A1(n19668), .A2(n10842), .B1(n19652), .B2(n19744), .C1(
        n19651), .C2(n19669), .ZN(P2_U3232) );
  OAI222_X1 U22643 ( .A1(n19668), .A2(n19654), .B1(n19653), .B2(n19744), .C1(
        n10842), .C2(n19669), .ZN(P2_U3233) );
  OAI222_X1 U22644 ( .A1(n19668), .A2(n19656), .B1(n19655), .B2(n19744), .C1(
        n19654), .C2(n19669), .ZN(P2_U3234) );
  OAI222_X1 U22645 ( .A1(n19668), .A2(n19658), .B1(n19657), .B2(n19744), .C1(
        n19656), .C2(n19669), .ZN(P2_U3235) );
  OAI222_X1 U22646 ( .A1(n19668), .A2(n19660), .B1(n19659), .B2(n19744), .C1(
        n19658), .C2(n19669), .ZN(P2_U3236) );
  OAI222_X1 U22647 ( .A1(n19668), .A2(n19663), .B1(n19661), .B2(n19744), .C1(
        n19660), .C2(n19669), .ZN(P2_U3237) );
  INV_X1 U22648 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19664) );
  OAI222_X1 U22649 ( .A1(n19669), .A2(n19663), .B1(n19662), .B2(n19744), .C1(
        n19664), .C2(n19668), .ZN(P2_U3238) );
  OAI222_X1 U22650 ( .A1(n19668), .A2(n19666), .B1(n19665), .B2(n19744), .C1(
        n19664), .C2(n19669), .ZN(P2_U3239) );
  OAI222_X1 U22651 ( .A1(n19668), .A2(n15026), .B1(n19667), .B2(n19744), .C1(
        n19666), .C2(n19669), .ZN(P2_U3240) );
  OAI222_X1 U22652 ( .A1(n19668), .A2(n19671), .B1(n19670), .B2(n19744), .C1(
        n15026), .C2(n19669), .ZN(P2_U3241) );
  OAI22_X1 U22653 ( .A1(n19745), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19744), .ZN(n19672) );
  INV_X1 U22654 ( .A(n19672), .ZN(P2_U3585) );
  MUX2_X1 U22655 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19745), .Z(P2_U3586) );
  OAI22_X1 U22656 ( .A1(n19745), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19744), .ZN(n19673) );
  INV_X1 U22657 ( .A(n19673), .ZN(P2_U3587) );
  OAI22_X1 U22658 ( .A1(n19745), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19744), .ZN(n19674) );
  INV_X1 U22659 ( .A(n19674), .ZN(P2_U3588) );
  OAI21_X1 U22660 ( .B1(n19678), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19676), 
        .ZN(n19675) );
  INV_X1 U22661 ( .A(n19675), .ZN(P2_U3591) );
  OAI21_X1 U22662 ( .B1(n19678), .B2(n19677), .A(n19676), .ZN(P2_U3592) );
  NOR2_X1 U22663 ( .A1(n19684), .A2(n19736), .ZN(n19700) );
  NAND2_X1 U22664 ( .A1(n19679), .A2(n19700), .ZN(n19693) );
  NAND2_X1 U22665 ( .A1(n19681), .A2(n19680), .ZN(n19701) );
  AOI21_X1 U22666 ( .B1(n19699), .B2(n19682), .A(n19701), .ZN(n19691) );
  AOI21_X1 U22667 ( .B1(n19693), .B2(n19691), .A(n19683), .ZN(n19688) );
  OAI22_X1 U22668 ( .A1(n19686), .A2(n19731), .B1(n19685), .B2(n19684), .ZN(
        n19687) );
  NOR2_X1 U22669 ( .A1(n19688), .A2(n19687), .ZN(n19689) );
  AOI22_X1 U22670 ( .A1(n19715), .A2(n19690), .B1(n19689), .B2(n19712), .ZN(
        P2_U3602) );
  INV_X1 U22671 ( .A(n19691), .ZN(n19696) );
  NOR2_X1 U22672 ( .A1(n19692), .A2(n19731), .ZN(n19695) );
  INV_X1 U22673 ( .A(n19693), .ZN(n19694) );
  AOI211_X1 U22674 ( .C1(n19697), .C2(n19696), .A(n19695), .B(n19694), .ZN(
        n19698) );
  AOI22_X1 U22675 ( .A1(n19715), .A2(n12319), .B1(n19698), .B2(n19712), .ZN(
        P2_U3603) );
  MUX2_X1 U22676 ( .A(n19701), .B(n19700), .S(n19699), .Z(n19702) );
  AOI21_X1 U22677 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19703), .A(n19702), 
        .ZN(n19704) );
  AOI22_X1 U22678 ( .A1(n19715), .A2(n19705), .B1(n19704), .B2(n19712), .ZN(
        P2_U3604) );
  INV_X1 U22679 ( .A(n19706), .ZN(n19707) );
  OAI22_X1 U22680 ( .A1(n19708), .A2(n19707), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19731), .ZN(n19709) );
  AOI21_X1 U22681 ( .B1(n19711), .B2(n19710), .A(n19709), .ZN(n19713) );
  AOI22_X1 U22682 ( .A1(n19715), .A2(n19714), .B1(n19713), .B2(n19712), .ZN(
        P2_U3605) );
  INV_X1 U22683 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19716) );
  AOI22_X1 U22684 ( .A1(n19744), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19716), 
        .B2(n19745), .ZN(P2_U3608) );
  INV_X1 U22685 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19726) );
  INV_X1 U22686 ( .A(n19717), .ZN(n19725) );
  AOI22_X1 U22687 ( .A1(n19721), .A2(n19720), .B1(n19719), .B2(n19718), .ZN(
        n19724) );
  NOR2_X1 U22688 ( .A1(n19725), .A2(n19722), .ZN(n19723) );
  AOI22_X1 U22689 ( .A1(n19726), .A2(n19725), .B1(n19724), .B2(n19723), .ZN(
        P2_U3609) );
  OAI21_X1 U22690 ( .B1(n19734), .B2(n19728), .A(n19727), .ZN(n19729) );
  AOI21_X1 U22691 ( .B1(n19731), .B2(n19730), .A(n19729), .ZN(n19742) );
  OAI21_X1 U22692 ( .B1(n19734), .B2(n19733), .A(n19732), .ZN(n19741) );
  AOI21_X1 U22693 ( .B1(n19737), .B2(n19736), .A(n19735), .ZN(n19738) );
  NOR3_X1 U22694 ( .A1(n12275), .A2(n19738), .A3(n13371), .ZN(n19739) );
  NOR2_X1 U22695 ( .A1(n19742), .A2(n19739), .ZN(n19740) );
  AOI22_X1 U22696 ( .A1(n19743), .A2(n19742), .B1(n19741), .B2(n19740), .ZN(
        P2_U3610) );
  OAI22_X1 U22697 ( .A1(n19745), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19744), .ZN(n19746) );
  INV_X1 U22698 ( .A(n19746), .ZN(P2_U3611) );
  NOR2_X1 U22699 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n19747), .ZN(n20662) );
  NOR2_X1 U22700 ( .A1(n20662), .A2(n20659), .ZN(n19755) );
  INV_X1 U22701 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19748) );
  AOI21_X1 U22702 ( .B1(n19755), .B2(n19748), .A(n20749), .ZN(P1_U2802) );
  INV_X1 U22703 ( .A(n19749), .ZN(n19751) );
  OAI21_X1 U22704 ( .B1(n19751), .B2(n19750), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19752) );
  OAI21_X1 U22705 ( .B1(n19753), .B2(n20759), .A(n19752), .ZN(P1_U2803) );
  INV_X1 U22706 ( .A(n20749), .ZN(n20747) );
  NOR2_X1 U22707 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20653) );
  INV_X1 U22708 ( .A(n20749), .ZN(n20770) );
  OAI21_X1 U22709 ( .B1(n20653), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20770), .ZN(
        n19754) );
  OAI21_X1 U22710 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20747), .A(n19754), 
        .ZN(P1_U2804) );
  NOR2_X1 U22711 ( .A1(n20749), .A2(n19755), .ZN(n20717) );
  OAI21_X1 U22712 ( .B1(BS16), .B2(n20653), .A(n20717), .ZN(n20715) );
  OAI21_X1 U22713 ( .B1(n20717), .B2(n20757), .A(n20715), .ZN(P1_U2805) );
  AOI21_X1 U22714 ( .B1(n19756), .B2(P1_FLUSH_REG_SCAN_IN), .A(n19939), .ZN(
        n19757) );
  INV_X1 U22715 ( .A(n19757), .ZN(P1_U2806) );
  NOR4_X1 U22716 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19761) );
  NOR4_X1 U22717 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19760) );
  NOR4_X1 U22718 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19759) );
  NOR4_X1 U22719 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19758) );
  NAND4_X1 U22720 ( .A1(n19761), .A2(n19760), .A3(n19759), .A4(n19758), .ZN(
        n19767) );
  NOR4_X1 U22721 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19765) );
  AOI211_X1 U22722 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19764) );
  NOR4_X1 U22723 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19763) );
  NOR4_X1 U22724 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19762) );
  NAND4_X1 U22725 ( .A1(n19765), .A2(n19764), .A3(n19763), .A4(n19762), .ZN(
        n19766) );
  NOR2_X1 U22726 ( .A1(n19767), .A2(n19766), .ZN(n20742) );
  INV_X1 U22727 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19769) );
  NOR3_X1 U22728 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19770) );
  OAI21_X1 U22729 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19770), .A(n20742), .ZN(
        n19768) );
  OAI21_X1 U22730 ( .B1(n20742), .B2(n19769), .A(n19768), .ZN(P1_U2807) );
  INV_X1 U22731 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20716) );
  AOI21_X1 U22732 ( .B1(n14390), .B2(n20716), .A(n19770), .ZN(n19772) );
  INV_X1 U22733 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19771) );
  INV_X1 U22734 ( .A(n20742), .ZN(n20745) );
  AOI22_X1 U22735 ( .A1(n20742), .A2(n19772), .B1(n19771), .B2(n20745), .ZN(
        P1_U2808) );
  OAI22_X1 U22736 ( .A1(n19774), .A2(n19819), .B1(n19865), .B2(n19773), .ZN(
        n19775) );
  AOI211_X1 U22737 ( .C1(n19849), .C2(P1_EBX_REG_9__SCAN_IN), .A(n19776), .B(
        n19775), .ZN(n19784) );
  INV_X1 U22738 ( .A(n19777), .ZN(n19779) );
  AOI22_X1 U22739 ( .A1(n19779), .A2(n19797), .B1(n19850), .B2(n19778), .ZN(
        n19783) );
  OAI21_X1 U22740 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n19781), .A(n19780), .ZN(
        n19782) );
  NAND3_X1 U22741 ( .A1(n19784), .A2(n19783), .A3(n19782), .ZN(P1_U2831) );
  OAI21_X1 U22742 ( .B1(n19819), .B2(n20945), .A(n19817), .ZN(n19788) );
  NAND2_X1 U22743 ( .A1(n19837), .A2(n19789), .ZN(n19786) );
  OAI22_X1 U22744 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19786), .B1(n19865), 
        .B2(n19785), .ZN(n19787) );
  AOI211_X1 U22745 ( .C1(P1_EBX_REG_7__SCAN_IN), .C2(n19849), .A(n19788), .B(
        n19787), .ZN(n19792) );
  OAI21_X1 U22746 ( .B1(n19826), .B2(n19789), .A(n19827), .ZN(n19802) );
  AOI22_X1 U22747 ( .A1(n19790), .A2(n19797), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19802), .ZN(n19791) );
  OAI211_X1 U22748 ( .C1(n19793), .C2(n19833), .A(n19792), .B(n19791), .ZN(
        P1_U2833) );
  AOI22_X1 U22749 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19853), .B1(
        n19834), .B2(n19794), .ZN(n19795) );
  OAI211_X1 U22750 ( .C1(n19847), .C2(n20895), .A(n19795), .B(n19817), .ZN(
        n19796) );
  AOI21_X1 U22751 ( .B1(n19798), .B2(n19797), .A(n19796), .ZN(n19804) );
  INV_X1 U22752 ( .A(n19799), .ZN(n19825) );
  NAND2_X1 U22753 ( .A1(n19827), .A2(n19825), .ZN(n19800) );
  AOI21_X1 U22754 ( .B1(n19801), .B2(n19800), .A(n20669), .ZN(n19806) );
  OAI21_X1 U22755 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n19806), .A(n19802), .ZN(
        n19803) );
  OAI211_X1 U22756 ( .C1(n19833), .C2(n19805), .A(n19804), .B(n19803), .ZN(
        P1_U2834) );
  NAND2_X1 U22757 ( .A1(n19837), .A2(n19825), .ZN(n19807) );
  AOI21_X1 U22758 ( .B1(n20669), .B2(n19807), .A(n19806), .ZN(n19811) );
  AOI22_X1 U22759 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n19849), .B1(n19834), .B2(
        n19866), .ZN(n19808) );
  OAI211_X1 U22760 ( .C1(n19819), .C2(n19809), .A(n19808), .B(n19817), .ZN(
        n19810) );
  AOI211_X1 U22761 ( .C1(n19867), .C2(n19830), .A(n19811), .B(n19810), .ZN(
        n19812) );
  OAI21_X1 U22762 ( .B1(n19813), .B2(n19833), .A(n19812), .ZN(P1_U2835) );
  AOI21_X1 U22763 ( .B1(n19816), .B2(n19815), .A(n19814), .ZN(n19945) );
  OAI21_X1 U22764 ( .B1(n19819), .B2(n19818), .A(n19817), .ZN(n19823) );
  OAI22_X1 U22765 ( .A1(n19872), .A2(n19847), .B1(n19821), .B2(n19820), .ZN(
        n19822) );
  AOI211_X1 U22766 ( .C1(n19834), .C2(n19945), .A(n19823), .B(n19822), .ZN(
        n19832) );
  NAND3_X1 U22767 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19824) );
  INV_X1 U22768 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20671) );
  AOI22_X1 U22769 ( .A1(n19827), .A2(n19825), .B1(n19824), .B2(n20671), .ZN(
        n19829) );
  OAI21_X1 U22770 ( .B1(n20671), .B2(n19827), .A(n19826), .ZN(n19828) );
  AOI22_X1 U22771 ( .A1(n19937), .A2(n19830), .B1(n19829), .B2(n19828), .ZN(
        n19831) );
  OAI211_X1 U22772 ( .C1(n19942), .C2(n19833), .A(n19832), .B(n19831), .ZN(
        P1_U2836) );
  AOI22_X1 U22773 ( .A1(n19835), .A2(n19850), .B1(n19834), .B2(n19955), .ZN(
        n19846) );
  AOI21_X1 U22774 ( .B1(n19837), .B2(n14390), .A(n19836), .ZN(n19857) );
  NOR2_X1 U22775 ( .A1(n19839), .A2(n19854), .ZN(n19838) );
  NAND2_X1 U22776 ( .A1(n19837), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19852) );
  AOI211_X1 U22777 ( .C1(n19839), .C2(n19854), .A(n19838), .B(n19852), .ZN(
        n19840) );
  AOI21_X1 U22778 ( .B1(n19853), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n19840), .ZN(n19841) );
  OAI21_X1 U22779 ( .B1(n19839), .B2(n19857), .A(n19841), .ZN(n19844) );
  NOR2_X1 U22780 ( .A1(n19842), .A2(n19858), .ZN(n19843) );
  AOI211_X1 U22781 ( .C1(n19862), .C2(n20727), .A(n19844), .B(n19843), .ZN(
        n19845) );
  OAI211_X1 U22782 ( .C1(n19848), .C2(n19847), .A(n19846), .B(n19845), .ZN(
        P1_U2837) );
  AOI22_X1 U22783 ( .A1(n19851), .A2(n19850), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n19849), .ZN(n19864) );
  INV_X1 U22784 ( .A(n12915), .ZN(n20003) );
  INV_X1 U22785 ( .A(n19852), .ZN(n19855) );
  AOI22_X1 U22786 ( .A1(n19855), .A2(n19854), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19853), .ZN(n19856) );
  OAI21_X1 U22787 ( .B1(n19857), .B2(n19854), .A(n19856), .ZN(n19861) );
  NOR2_X1 U22788 ( .A1(n19859), .A2(n19858), .ZN(n19860) );
  AOI211_X1 U22789 ( .C1(n19862), .C2(n20003), .A(n19861), .B(n19860), .ZN(
        n19863) );
  OAI211_X1 U22790 ( .C1(n19865), .C2(n19964), .A(n19864), .B(n19863), .ZN(
        P1_U2838) );
  INV_X1 U22791 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20795) );
  AOI22_X1 U22792 ( .A1(n19867), .A2(n19870), .B1(n19869), .B2(n19866), .ZN(
        n19868) );
  OAI21_X1 U22793 ( .B1(n19873), .B2(n20795), .A(n19868), .ZN(P1_U2867) );
  AOI22_X1 U22794 ( .A1(n19937), .A2(n19870), .B1(n19869), .B2(n19945), .ZN(
        n19871) );
  OAI21_X1 U22795 ( .B1(n19873), .B2(n19872), .A(n19871), .ZN(P1_U2868) );
  AOI22_X1 U22796 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19877), .B1(n15733), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U22797 ( .B1(n19876), .B2(n19875), .A(n19874), .ZN(P1_U2921) );
  INV_X1 U22798 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U22799 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U22800 ( .B1(n19879), .B2(n19903), .A(n19878), .ZN(P1_U2922) );
  AOI22_X1 U22801 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U22802 ( .B1(n14501), .B2(n19903), .A(n19880), .ZN(P1_U2923) );
  AOI22_X1 U22803 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19881) );
  OAI21_X1 U22804 ( .B1(n14506), .B2(n19903), .A(n19881), .ZN(P1_U2924) );
  INV_X1 U22805 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U22806 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19882) );
  OAI21_X1 U22807 ( .B1(n19883), .B2(n19903), .A(n19882), .ZN(P1_U2925) );
  INV_X1 U22808 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U22809 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19884) );
  OAI21_X1 U22810 ( .B1(n19885), .B2(n19903), .A(n19884), .ZN(P1_U2926) );
  INV_X1 U22811 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U22812 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19886) );
  OAI21_X1 U22813 ( .B1(n19887), .B2(n19903), .A(n19886), .ZN(P1_U2927) );
  AOI22_X1 U22814 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19888) );
  OAI21_X1 U22815 ( .B1(n19889), .B2(n19903), .A(n19888), .ZN(P1_U2928) );
  AOI22_X1 U22816 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19890) );
  OAI21_X1 U22817 ( .B1(n13536), .B2(n19903), .A(n19890), .ZN(P1_U2929) );
  AOI22_X1 U22818 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19891) );
  OAI21_X1 U22819 ( .B1(n11411), .B2(n19903), .A(n19891), .ZN(P1_U2930) );
  AOI22_X1 U22820 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19892) );
  OAI21_X1 U22821 ( .B1(n13339), .B2(n19903), .A(n19892), .ZN(P1_U2931) );
  AOI22_X1 U22822 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19893) );
  OAI21_X1 U22823 ( .B1(n19894), .B2(n19903), .A(n19893), .ZN(P1_U2932) );
  AOI22_X1 U22824 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19895) );
  OAI21_X1 U22825 ( .B1(n19896), .B2(n19903), .A(n19895), .ZN(P1_U2933) );
  AOI22_X1 U22826 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19897) );
  OAI21_X1 U22827 ( .B1(n19898), .B2(n19903), .A(n19897), .ZN(P1_U2934) );
  AOI22_X1 U22828 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19899) );
  OAI21_X1 U22829 ( .B1(n19900), .B2(n19903), .A(n19899), .ZN(P1_U2935) );
  AOI22_X1 U22830 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19901), .B1(n15733), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19902) );
  OAI21_X1 U22831 ( .B1(n19904), .B2(n19903), .A(n19902), .ZN(P1_U2936) );
  AOI22_X1 U22832 ( .A1(n19929), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n19926), .ZN(n19906) );
  NAND2_X1 U22833 ( .A1(n19916), .A2(n19905), .ZN(n19918) );
  NAND2_X1 U22834 ( .A1(n19906), .A2(n19918), .ZN(P1_U2946) );
  AOI22_X1 U22835 ( .A1(n19929), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n19926), .ZN(n19908) );
  NAND2_X1 U22836 ( .A1(n19916), .A2(n19907), .ZN(n19920) );
  NAND2_X1 U22837 ( .A1(n19908), .A2(n19920), .ZN(P1_U2947) );
  AOI22_X1 U22838 ( .A1(n19929), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n19926), .ZN(n19910) );
  NAND2_X1 U22839 ( .A1(n19916), .A2(n19909), .ZN(n19922) );
  NAND2_X1 U22840 ( .A1(n19910), .A2(n19922), .ZN(P1_U2948) );
  AOI22_X1 U22841 ( .A1(n19929), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n19926), .ZN(n19912) );
  NAND2_X1 U22842 ( .A1(n19916), .A2(n19911), .ZN(n19924) );
  NAND2_X1 U22843 ( .A1(n19912), .A2(n19924), .ZN(P1_U2949) );
  AOI22_X1 U22844 ( .A1(n19929), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n19926), .ZN(n19914) );
  NAND2_X1 U22845 ( .A1(n19916), .A2(n19913), .ZN(n19927) );
  NAND2_X1 U22846 ( .A1(n19914), .A2(n19927), .ZN(P1_U2950) );
  AOI22_X1 U22847 ( .A1(n19929), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19926), .ZN(n19917) );
  NAND2_X1 U22848 ( .A1(n19916), .A2(n19915), .ZN(n19930) );
  NAND2_X1 U22849 ( .A1(n19917), .A2(n19930), .ZN(P1_U2951) );
  AOI22_X1 U22850 ( .A1(n19929), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19926), .ZN(n19919) );
  NAND2_X1 U22851 ( .A1(n19919), .A2(n19918), .ZN(P1_U2961) );
  AOI22_X1 U22852 ( .A1(n19929), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19926), .ZN(n19921) );
  NAND2_X1 U22853 ( .A1(n19921), .A2(n19920), .ZN(P1_U2962) );
  AOI22_X1 U22854 ( .A1(n19929), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19926), .ZN(n19923) );
  NAND2_X1 U22855 ( .A1(n19923), .A2(n19922), .ZN(P1_U2963) );
  AOI22_X1 U22856 ( .A1(n19929), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19926), .ZN(n19925) );
  NAND2_X1 U22857 ( .A1(n19925), .A2(n19924), .ZN(P1_U2964) );
  AOI22_X1 U22858 ( .A1(n19929), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19926), .ZN(n19928) );
  NAND2_X1 U22859 ( .A1(n19928), .A2(n19927), .ZN(P1_U2965) );
  AOI22_X1 U22860 ( .A1(n19929), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19926), .ZN(n19931) );
  NAND2_X1 U22861 ( .A1(n19931), .A2(n19930), .ZN(P1_U2966) );
  AOI22_X1 U22862 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19944), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19941) );
  OAI21_X1 U22863 ( .B1(n19935), .B2(n19934), .A(n19933), .ZN(n19936) );
  INV_X1 U22864 ( .A(n19936), .ZN(n19948) );
  AOI22_X1 U22865 ( .A1(n19948), .A2(n19939), .B1(n19938), .B2(n19937), .ZN(
        n19940) );
  OAI211_X1 U22866 ( .C1(n19943), .C2(n19942), .A(n19941), .B(n19940), .ZN(
        P1_U2995) );
  AOI22_X1 U22867 ( .A1(n19945), .A2(n19974), .B1(n19944), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n19952) );
  NAND2_X1 U22868 ( .A1(n19962), .A2(n19946), .ZN(n19968) );
  NAND3_X1 U22869 ( .A1(n19977), .A2(n19947), .A3(n19968), .ZN(n19956) );
  AOI22_X1 U22870 ( .A1(n19948), .A2(n19988), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19956), .ZN(n19951) );
  OAI211_X1 U22871 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n19953), .B(n19949), .ZN(n19950) );
  NAND3_X1 U22872 ( .A1(n19952), .A2(n19951), .A3(n19950), .ZN(P1_U3027) );
  INV_X1 U22873 ( .A(n19953), .ZN(n19960) );
  AOI21_X1 U22874 ( .B1(n19955), .B2(n19974), .A(n19954), .ZN(n19959) );
  AOI22_X1 U22875 ( .A1(n19957), .A2(n19988), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n19956), .ZN(n19958) );
  OAI211_X1 U22876 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n19960), .A(
        n19959), .B(n19958), .ZN(P1_U3028) );
  NOR2_X1 U22877 ( .A1(n13034), .A2(n19984), .ZN(n19963) );
  AOI22_X1 U22878 ( .A1(n19963), .A2(n19962), .B1(n19984), .B2(n19961), .ZN(
        n19976) );
  INV_X1 U22879 ( .A(n19964), .ZN(n19973) );
  OR3_X1 U22880 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19984), .A3(
        n19965), .ZN(n19966) );
  NAND3_X1 U22881 ( .A1(n19968), .A2(n19967), .A3(n19966), .ZN(n19972) );
  AND3_X1 U22882 ( .A1(n19970), .A2(n19969), .A3(n19988), .ZN(n19971) );
  AOI211_X1 U22883 ( .C1(n19974), .C2(n19973), .A(n19972), .B(n19971), .ZN(
        n19975) );
  OAI221_X1 U22884 ( .B1(n19978), .B2(n19977), .C1(n19978), .C2(n19976), .A(
        n19975), .ZN(P1_U3029) );
  OAI21_X1 U22885 ( .B1(n19981), .B2(n19980), .A(n19979), .ZN(n19982) );
  INV_X1 U22886 ( .A(n19982), .ZN(n19994) );
  INV_X1 U22887 ( .A(n19983), .ZN(n19989) );
  AND2_X1 U22888 ( .A1(n19985), .A2(n19984), .ZN(n19987) );
  AOI22_X1 U22889 ( .A1(n19989), .A2(n19988), .B1(n19987), .B2(n19986), .ZN(
        n19993) );
  OAI21_X1 U22890 ( .B1(n19991), .B2(n19990), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19992) );
  NAND3_X1 U22891 ( .A1(n19994), .A2(n19993), .A3(n19992), .ZN(P1_U3030) );
  NOR2_X1 U22892 ( .A1(n19995), .A2(n20738), .ZN(P1_U3032) );
  AOI22_X1 U22893 ( .A1(DATAI_16_), .A2(n20038), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20037), .ZN(n20477) );
  AOI22_X1 U22894 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20037), .B1(DATAI_24_), 
        .B2(n20038), .ZN(n20526) );
  INV_X1 U22895 ( .A(n20526), .ZN(n20584) );
  NAND2_X1 U22896 ( .A1(n20040), .A2(n9956), .ZN(n20582) );
  NOR3_X1 U22897 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20051) );
  INV_X1 U22898 ( .A(n20051), .ZN(n20048) );
  NOR2_X1 U22899 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20048), .ZN(
        n20041) );
  AOI22_X1 U22900 ( .A1(n20644), .A2(n20584), .B1(n20514), .B2(n20041), .ZN(
        n20013) );
  OR2_X1 U22901 ( .A1(n20008), .A2(n20750), .ZN(n20512) );
  INV_X1 U22902 ( .A(n20512), .ZN(n20001) );
  INV_X1 U22903 ( .A(n20068), .ZN(n20071) );
  NOR3_X1 U22904 ( .A1(n20644), .A2(n20071), .A3(n20573), .ZN(n20002) );
  NAND2_X1 U22905 ( .A1(n20757), .A2(n20576), .ZN(n20431) );
  INV_X1 U22906 ( .A(n20431), .ZN(n20729) );
  NOR2_X1 U22907 ( .A1(n20002), .A2(n20729), .ZN(n20011) );
  INV_X1 U22908 ( .A(n20011), .ZN(n20005) );
  NAND2_X1 U22909 ( .A1(n9741), .A2(n20433), .ZN(n20010) );
  INV_X1 U22910 ( .A(n20004), .ZN(n20296) );
  NAND2_X1 U22911 ( .A1(n20296), .A2(n20354), .ZN(n20150) );
  AOI22_X1 U22912 ( .A1(n20005), .A2(n20010), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20150), .ZN(n20006) );
  INV_X1 U22913 ( .A(n20008), .ZN(n20009) );
  NOR2_X1 U22914 ( .A1(n20009), .A2(n20750), .ZN(n20155) );
  INV_X1 U22915 ( .A(n20155), .ZN(n20358) );
  AOI22_X1 U22916 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20044), .B1(
        n20513), .B2(n20043), .ZN(n20012) );
  OAI211_X1 U22917 ( .C1(n20477), .C2(n20068), .A(n20013), .B(n20012), .ZN(
        P1_U3033) );
  AOI22_X1 U22918 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20037), .B1(DATAI_17_), 
        .B2(n20038), .ZN(n20481) );
  AOI22_X1 U22919 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20037), .B1(DATAI_25_), 
        .B2(n20038), .ZN(n20531) );
  INV_X1 U22920 ( .A(n20531), .ZN(n20592) );
  NAND2_X1 U22921 ( .A1(n20040), .A2(n20014), .ZN(n20589) );
  AOI22_X1 U22922 ( .A1(n20644), .A2(n20592), .B1(n20528), .B2(n20041), .ZN(
        n20017) );
  AOI22_X1 U22923 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20044), .B1(
        n20527), .B2(n20043), .ZN(n20016) );
  OAI211_X1 U22924 ( .C1(n20481), .C2(n20068), .A(n20017), .B(n20016), .ZN(
        P1_U3034) );
  AOI22_X1 U22925 ( .A1(DATAI_18_), .A2(n20038), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20037), .ZN(n20485) );
  INV_X1 U22926 ( .A(n20536), .ZN(n20600) );
  NAND2_X1 U22927 ( .A1(n20040), .A2(n20018), .ZN(n20597) );
  AOI22_X1 U22928 ( .A1(n20644), .A2(n20600), .B1(n20533), .B2(n20041), .ZN(
        n20021) );
  AOI22_X1 U22929 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20044), .B1(
        n20532), .B2(n20043), .ZN(n20020) );
  OAI211_X1 U22930 ( .C1(n20485), .C2(n20068), .A(n20021), .B(n20020), .ZN(
        P1_U3035) );
  AOI22_X1 U22931 ( .A1(DATAI_19_), .A2(n20038), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20037), .ZN(n20489) );
  INV_X1 U22932 ( .A(n20541), .ZN(n20607) );
  NAND2_X1 U22933 ( .A1(n20040), .A2(n20022), .ZN(n20605) );
  AOI22_X1 U22934 ( .A1(n20644), .A2(n20607), .B1(n20538), .B2(n20041), .ZN(
        n20025) );
  AOI22_X1 U22935 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20044), .B1(
        n20537), .B2(n20043), .ZN(n20024) );
  OAI211_X1 U22936 ( .C1(n20489), .C2(n20068), .A(n20025), .B(n20024), .ZN(
        P1_U3036) );
  AOI22_X1 U22937 ( .A1(DATAI_20_), .A2(n20038), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20037), .ZN(n20493) );
  INV_X1 U22938 ( .A(n20546), .ZN(n20615) );
  NAND2_X1 U22939 ( .A1(n20040), .A2(n11112), .ZN(n20613) );
  AOI22_X1 U22940 ( .A1(n20644), .A2(n20615), .B1(n20041), .B2(n20543), .ZN(
        n20028) );
  AOI22_X1 U22941 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20044), .B1(
        n20542), .B2(n20043), .ZN(n20027) );
  OAI211_X1 U22942 ( .C1(n20493), .C2(n20068), .A(n20028), .B(n20027), .ZN(
        P1_U3037) );
  AOI22_X1 U22943 ( .A1(DATAI_21_), .A2(n20038), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20037), .ZN(n20497) );
  AOI22_X2 U22944 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20037), .B1(DATAI_29_), 
        .B2(n20038), .ZN(n20551) );
  INV_X1 U22945 ( .A(n20551), .ZN(n20623) );
  NAND2_X1 U22946 ( .A1(n20040), .A2(n20029), .ZN(n20621) );
  AOI22_X1 U22947 ( .A1(n20644), .A2(n20623), .B1(n20548), .B2(n20041), .ZN(
        n20032) );
  AOI22_X1 U22948 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20044), .B1(
        n20547), .B2(n20043), .ZN(n20031) );
  OAI211_X1 U22949 ( .C1(n20497), .C2(n20068), .A(n20032), .B(n20031), .ZN(
        P1_U3038) );
  AOI22_X1 U22950 ( .A1(DATAI_22_), .A2(n20038), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20037), .ZN(n20501) );
  AOI22_X1 U22951 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20037), .B1(DATAI_30_), 
        .B2(n20038), .ZN(n20556) );
  INV_X1 U22952 ( .A(n20556), .ZN(n20631) );
  NAND2_X1 U22953 ( .A1(n20040), .A2(n20033), .ZN(n20629) );
  AOI22_X1 U22954 ( .A1(n20644), .A2(n20631), .B1(n20553), .B2(n20041), .ZN(
        n20036) );
  AOI22_X1 U22955 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20044), .B1(
        n20552), .B2(n20043), .ZN(n20035) );
  OAI211_X1 U22956 ( .C1(n20501), .C2(n20068), .A(n20036), .B(n20035), .ZN(
        P1_U3039) );
  AOI22_X1 U22957 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20037), .B1(DATAI_23_), 
        .B2(n20038), .ZN(n20509) );
  AOI22_X1 U22958 ( .A1(DATAI_31_), .A2(n20038), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20037), .ZN(n20565) );
  INV_X1 U22959 ( .A(n20565), .ZN(n20641) );
  NAND2_X1 U22960 ( .A1(n20040), .A2(n20039), .ZN(n20639) );
  AOI22_X1 U22961 ( .A1(n20644), .A2(n20641), .B1(n20560), .B2(n20041), .ZN(
        n20046) );
  AOI22_X1 U22962 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20044), .B1(
        n20558), .B2(n20043), .ZN(n20045) );
  OAI211_X1 U22963 ( .C1(n20509), .C2(n20068), .A(n20046), .B(n20045), .ZN(
        P1_U3040) );
  NOR2_X1 U22964 ( .A1(n20464), .A2(n20048), .ZN(n20070) );
  INV_X1 U22965 ( .A(n20047), .ZN(n20465) );
  AOI21_X1 U22966 ( .B1(n9741), .B2(n20465), .A(n20070), .ZN(n20049) );
  OAI22_X1 U22967 ( .A1(n20049), .A2(n20573), .B1(n20048), .B2(n20750), .ZN(
        n20069) );
  AOI22_X1 U22968 ( .A1(n20514), .A2(n20070), .B1(n20513), .B2(n20069), .ZN(
        n20054) );
  INV_X1 U22969 ( .A(n20725), .ZN(n20395) );
  NOR2_X1 U22970 ( .A1(n9654), .A2(n20395), .ZN(n20471) );
  INV_X1 U22971 ( .A(n20471), .ZN(n20050) );
  NOR2_X1 U22972 ( .A1(n20115), .A2(n20050), .ZN(n20052) );
  OAI21_X1 U22973 ( .B1(n20052), .B2(n20051), .A(n20472), .ZN(n20072) );
  INV_X1 U22974 ( .A(n20477), .ZN(n20585) );
  AOI22_X1 U22975 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20072), .B1(
        n20065), .B2(n20585), .ZN(n20053) );
  OAI211_X1 U22976 ( .C1(n20526), .C2(n20068), .A(n20054), .B(n20053), .ZN(
        P1_U3041) );
  AOI22_X1 U22977 ( .A1(n20528), .A2(n20070), .B1(n20527), .B2(n20069), .ZN(
        n20056) );
  INV_X1 U22978 ( .A(n20481), .ZN(n20591) );
  AOI22_X1 U22979 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20072), .B1(
        n20065), .B2(n20591), .ZN(n20055) );
  OAI211_X1 U22980 ( .C1(n20531), .C2(n20068), .A(n20056), .B(n20055), .ZN(
        P1_U3042) );
  AOI22_X1 U22981 ( .A1(n20533), .A2(n20070), .B1(n20532), .B2(n20069), .ZN(
        n20058) );
  INV_X1 U22982 ( .A(n20485), .ZN(n20599) );
  AOI22_X1 U22983 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20072), .B1(
        n20065), .B2(n20599), .ZN(n20057) );
  OAI211_X1 U22984 ( .C1(n20536), .C2(n20068), .A(n20058), .B(n20057), .ZN(
        P1_U3043) );
  AOI22_X1 U22985 ( .A1(n20538), .A2(n20070), .B1(n20537), .B2(n20069), .ZN(
        n20060) );
  INV_X1 U22986 ( .A(n20489), .ZN(n20608) );
  AOI22_X1 U22987 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20072), .B1(
        n20065), .B2(n20608), .ZN(n20059) );
  OAI211_X1 U22988 ( .C1(n20541), .C2(n20068), .A(n20060), .B(n20059), .ZN(
        P1_U3044) );
  AOI22_X1 U22989 ( .A1(n20543), .A2(n20070), .B1(n20542), .B2(n20069), .ZN(
        n20062) );
  INV_X1 U22990 ( .A(n20493), .ZN(n20616) );
  AOI22_X1 U22991 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20072), .B1(
        n20065), .B2(n20616), .ZN(n20061) );
  OAI211_X1 U22992 ( .C1(n20546), .C2(n20068), .A(n20062), .B(n20061), .ZN(
        P1_U3045) );
  AOI22_X1 U22993 ( .A1(n20548), .A2(n20070), .B1(n20547), .B2(n20069), .ZN(
        n20064) );
  INV_X1 U22994 ( .A(n20497), .ZN(n20624) );
  AOI22_X1 U22995 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20072), .B1(
        n20065), .B2(n20624), .ZN(n20063) );
  OAI211_X1 U22996 ( .C1(n20551), .C2(n20068), .A(n20064), .B(n20063), .ZN(
        P1_U3046) );
  AOI22_X1 U22997 ( .A1(n20553), .A2(n20070), .B1(n20552), .B2(n20069), .ZN(
        n20067) );
  INV_X1 U22998 ( .A(n20501), .ZN(n20632) );
  AOI22_X1 U22999 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20072), .B1(
        n20065), .B2(n20632), .ZN(n20066) );
  OAI211_X1 U23000 ( .C1(n20556), .C2(n20068), .A(n20067), .B(n20066), .ZN(
        P1_U3047) );
  AOI22_X1 U23001 ( .A1(n20560), .A2(n20070), .B1(n20558), .B2(n20069), .ZN(
        n20074) );
  AOI22_X1 U23002 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20072), .B1(
        n20071), .B2(n20641), .ZN(n20073) );
  OAI211_X1 U23003 ( .C1(n20509), .C2(n20107), .A(n20074), .B(n20073), .ZN(
        P1_U3048) );
  NAND2_X1 U23004 ( .A1(n9654), .A2(n9650), .ZN(n20515) );
  NAND3_X1 U23005 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20737), .A3(
        n20428), .ZN(n20118) );
  OR2_X1 U23006 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20118), .ZN(
        n20101) );
  OAI22_X1 U23007 ( .A1(n20147), .A2(n20477), .B1(n20582), .B2(n20101), .ZN(
        n20075) );
  INV_X1 U23008 ( .A(n20075), .ZN(n20082) );
  NAND3_X1 U23009 ( .A1(n20107), .A2(n20576), .A3(n20147), .ZN(n20076) );
  NAND2_X1 U23010 ( .A1(n20076), .A2(n20431), .ZN(n20078) );
  INV_X1 U23011 ( .A(n20433), .ZN(n20519) );
  NAND2_X1 U23012 ( .A1(n9741), .A2(n20519), .ZN(n20079) );
  AOI22_X1 U23013 ( .A1(n20078), .A2(n20079), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20101), .ZN(n20077) );
  OAI21_X1 U23014 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20354), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20218) );
  NAND3_X1 U23015 ( .A1(n20356), .A2(n20077), .A3(n20218), .ZN(n20104) );
  INV_X1 U23016 ( .A(n20078), .ZN(n20080) );
  INV_X1 U23017 ( .A(n20354), .ZN(n20295) );
  NAND2_X1 U23018 ( .A1(n20295), .A2(n20737), .ZN(n20221) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20104), .B1(
        n20513), .B2(n20103), .ZN(n20081) );
  OAI211_X1 U23020 ( .C1(n20526), .C2(n20107), .A(n20082), .B(n20081), .ZN(
        P1_U3049) );
  OAI22_X1 U23021 ( .A1(n20107), .A2(n20531), .B1(n20589), .B2(n20101), .ZN(
        n20083) );
  INV_X1 U23022 ( .A(n20083), .ZN(n20085) );
  AOI22_X1 U23023 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20104), .B1(
        n20527), .B2(n20103), .ZN(n20084) );
  OAI211_X1 U23024 ( .C1(n20481), .C2(n20147), .A(n20085), .B(n20084), .ZN(
        P1_U3050) );
  OAI22_X1 U23025 ( .A1(n20107), .A2(n20536), .B1(n20597), .B2(n20101), .ZN(
        n20086) );
  INV_X1 U23026 ( .A(n20086), .ZN(n20088) );
  AOI22_X1 U23027 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20104), .B1(
        n20532), .B2(n20103), .ZN(n20087) );
  OAI211_X1 U23028 ( .C1(n20485), .C2(n20147), .A(n20088), .B(n20087), .ZN(
        P1_U3051) );
  OAI22_X1 U23029 ( .A1(n20147), .A2(n20489), .B1(n20605), .B2(n20101), .ZN(
        n20089) );
  INV_X1 U23030 ( .A(n20089), .ZN(n20091) );
  AOI22_X1 U23031 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20104), .B1(
        n20537), .B2(n20103), .ZN(n20090) );
  OAI211_X1 U23032 ( .C1(n20541), .C2(n20107), .A(n20091), .B(n20090), .ZN(
        P1_U3052) );
  OAI22_X1 U23033 ( .A1(n20147), .A2(n20493), .B1(n20101), .B2(n20613), .ZN(
        n20092) );
  INV_X1 U23034 ( .A(n20092), .ZN(n20094) );
  AOI22_X1 U23035 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20104), .B1(
        n20542), .B2(n20103), .ZN(n20093) );
  OAI211_X1 U23036 ( .C1(n20546), .C2(n20107), .A(n20094), .B(n20093), .ZN(
        P1_U3053) );
  OAI22_X1 U23037 ( .A1(n20147), .A2(n20497), .B1(n20621), .B2(n20101), .ZN(
        n20095) );
  INV_X1 U23038 ( .A(n20095), .ZN(n20097) );
  AOI22_X1 U23039 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20104), .B1(
        n20547), .B2(n20103), .ZN(n20096) );
  OAI211_X1 U23040 ( .C1(n20551), .C2(n20107), .A(n20097), .B(n20096), .ZN(
        P1_U3054) );
  OAI22_X1 U23041 ( .A1(n20147), .A2(n20501), .B1(n20629), .B2(n20101), .ZN(
        n20098) );
  INV_X1 U23042 ( .A(n20098), .ZN(n20100) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20104), .B1(
        n20552), .B2(n20103), .ZN(n20099) );
  OAI211_X1 U23044 ( .C1(n20556), .C2(n20107), .A(n20100), .B(n20099), .ZN(
        P1_U3055) );
  OAI22_X1 U23045 ( .A1(n20147), .A2(n20509), .B1(n20639), .B2(n20101), .ZN(
        n20102) );
  INV_X1 U23046 ( .A(n20102), .ZN(n20106) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20104), .B1(
        n20558), .B2(n20103), .ZN(n20105) );
  OAI211_X1 U23048 ( .C1(n20565), .C2(n20107), .A(n20106), .B(n20105), .ZN(
        P1_U3056) );
  OR2_X1 U23049 ( .A1(n20388), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20141) );
  OAI22_X1 U23050 ( .A1(n20177), .A2(n20477), .B1(n20582), .B2(n20141), .ZN(
        n20109) );
  INV_X1 U23051 ( .A(n20109), .ZN(n20122) );
  NAND2_X1 U23052 ( .A1(n20111), .A2(n20110), .ZN(n20389) );
  INV_X1 U23053 ( .A(n20141), .ZN(n20112) );
  AOI21_X1 U23054 ( .B1(n9741), .B2(n20567), .A(n20112), .ZN(n20120) );
  INV_X1 U23055 ( .A(n20113), .ZN(n20114) );
  AOI21_X1 U23056 ( .B1(n20115), .B2(n20576), .A(n20114), .ZN(n20119) );
  INV_X1 U23057 ( .A(n20119), .ZN(n20116) );
  AOI22_X1 U23058 ( .A1(n20120), .A2(n20116), .B1(n20573), .B2(n20118), .ZN(
        n20117) );
  NAND2_X1 U23059 ( .A1(n20472), .A2(n20117), .ZN(n20144) );
  OAI22_X1 U23060 ( .A1(n20120), .A2(n20119), .B1(n20750), .B2(n20118), .ZN(
        n20143) );
  AOI22_X1 U23061 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20144), .B1(
        n20513), .B2(n20143), .ZN(n20121) );
  OAI211_X1 U23062 ( .C1(n20526), .C2(n20147), .A(n20122), .B(n20121), .ZN(
        P1_U3057) );
  OAI22_X1 U23063 ( .A1(n20177), .A2(n20481), .B1(n20589), .B2(n20141), .ZN(
        n20123) );
  INV_X1 U23064 ( .A(n20123), .ZN(n20125) );
  AOI22_X1 U23065 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20144), .B1(
        n20527), .B2(n20143), .ZN(n20124) );
  OAI211_X1 U23066 ( .C1(n20531), .C2(n20147), .A(n20125), .B(n20124), .ZN(
        P1_U3058) );
  OAI22_X1 U23067 ( .A1(n20147), .A2(n20536), .B1(n20597), .B2(n20141), .ZN(
        n20126) );
  INV_X1 U23068 ( .A(n20126), .ZN(n20128) );
  AOI22_X1 U23069 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20144), .B1(
        n20532), .B2(n20143), .ZN(n20127) );
  OAI211_X1 U23070 ( .C1(n20485), .C2(n20177), .A(n20128), .B(n20127), .ZN(
        P1_U3059) );
  OAI22_X1 U23071 ( .A1(n20177), .A2(n20489), .B1(n20605), .B2(n20141), .ZN(
        n20129) );
  INV_X1 U23072 ( .A(n20129), .ZN(n20131) );
  AOI22_X1 U23073 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20144), .B1(
        n20537), .B2(n20143), .ZN(n20130) );
  OAI211_X1 U23074 ( .C1(n20541), .C2(n20147), .A(n20131), .B(n20130), .ZN(
        P1_U3060) );
  OAI22_X1 U23075 ( .A1(n20147), .A2(n20546), .B1(n20141), .B2(n20613), .ZN(
        n20132) );
  INV_X1 U23076 ( .A(n20132), .ZN(n20134) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20144), .B1(
        n20542), .B2(n20143), .ZN(n20133) );
  OAI211_X1 U23078 ( .C1(n20493), .C2(n20177), .A(n20134), .B(n20133), .ZN(
        P1_U3061) );
  OAI22_X1 U23079 ( .A1(n20177), .A2(n20497), .B1(n20621), .B2(n20141), .ZN(
        n20135) );
  INV_X1 U23080 ( .A(n20135), .ZN(n20137) );
  AOI22_X1 U23081 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20144), .B1(
        n20547), .B2(n20143), .ZN(n20136) );
  OAI211_X1 U23082 ( .C1(n20551), .C2(n20147), .A(n20137), .B(n20136), .ZN(
        P1_U3062) );
  OAI22_X1 U23083 ( .A1(n20177), .A2(n20501), .B1(n20629), .B2(n20141), .ZN(
        n20138) );
  INV_X1 U23084 ( .A(n20138), .ZN(n20140) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20144), .B1(
        n20552), .B2(n20143), .ZN(n20139) );
  OAI211_X1 U23086 ( .C1(n20556), .C2(n20147), .A(n20140), .B(n20139), .ZN(
        P1_U3063) );
  OAI22_X1 U23087 ( .A1(n20177), .A2(n20509), .B1(n20639), .B2(n20141), .ZN(
        n20142) );
  INV_X1 U23088 ( .A(n20142), .ZN(n20146) );
  AOI22_X1 U23089 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20144), .B1(
        n20558), .B2(n20143), .ZN(n20145) );
  OAI211_X1 U23090 ( .C1(n20565), .C2(n20147), .A(n20146), .B(n20145), .ZN(
        P1_U3064) );
  NOR3_X1 U23091 ( .A1(n20428), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20186) );
  INV_X1 U23092 ( .A(n20186), .ZN(n20178) );
  NOR2_X1 U23093 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20178), .ZN(
        n20173) );
  NOR2_X1 U23094 ( .A1(n12915), .A2(n20148), .ZN(n20251) );
  NAND3_X1 U23095 ( .A1(n20251), .A2(n20576), .A3(n20433), .ZN(n20149) );
  OAI21_X1 U23096 ( .B1(n20150), .B2(n20512), .A(n20149), .ZN(n20172) );
  AOI22_X1 U23097 ( .A1(n20514), .A2(n20173), .B1(n20513), .B2(n20172), .ZN(
        n20158) );
  AOI21_X1 U23098 ( .B1(n20177), .B2(n20215), .A(n20757), .ZN(n20152) );
  AOI21_X1 U23099 ( .B1(n20251), .B2(n20433), .A(n20152), .ZN(n20153) );
  NOR2_X1 U23100 ( .A1(n20153), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20156) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20174), .B1(
        n20187), .B2(n20585), .ZN(n20157) );
  OAI211_X1 U23102 ( .C1(n20526), .C2(n20177), .A(n20158), .B(n20157), .ZN(
        P1_U3065) );
  AOI22_X1 U23103 ( .A1(n20528), .A2(n20173), .B1(n20527), .B2(n20172), .ZN(
        n20160) );
  INV_X1 U23104 ( .A(n20177), .ZN(n20161) );
  AOI22_X1 U23105 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20174), .B1(
        n20161), .B2(n20592), .ZN(n20159) );
  OAI211_X1 U23106 ( .C1(n20481), .C2(n20215), .A(n20160), .B(n20159), .ZN(
        P1_U3066) );
  AOI22_X1 U23107 ( .A1(n20533), .A2(n20173), .B1(n20532), .B2(n20172), .ZN(
        n20163) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20174), .B1(
        n20161), .B2(n20600), .ZN(n20162) );
  OAI211_X1 U23109 ( .C1(n20485), .C2(n20215), .A(n20163), .B(n20162), .ZN(
        P1_U3067) );
  AOI22_X1 U23110 ( .A1(n20538), .A2(n20173), .B1(n20537), .B2(n20172), .ZN(
        n20165) );
  AOI22_X1 U23111 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20174), .B1(
        n20187), .B2(n20608), .ZN(n20164) );
  OAI211_X1 U23112 ( .C1(n20541), .C2(n20177), .A(n20165), .B(n20164), .ZN(
        P1_U3068) );
  AOI22_X1 U23113 ( .A1(n20543), .A2(n20173), .B1(n20542), .B2(n20172), .ZN(
        n20167) );
  AOI22_X1 U23114 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20174), .B1(
        n20187), .B2(n20616), .ZN(n20166) );
  OAI211_X1 U23115 ( .C1(n20546), .C2(n20177), .A(n20167), .B(n20166), .ZN(
        P1_U3069) );
  AOI22_X1 U23116 ( .A1(n20548), .A2(n20173), .B1(n20547), .B2(n20172), .ZN(
        n20169) );
  AOI22_X1 U23117 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20174), .B1(
        n20187), .B2(n20624), .ZN(n20168) );
  OAI211_X1 U23118 ( .C1(n20551), .C2(n20177), .A(n20169), .B(n20168), .ZN(
        P1_U3070) );
  AOI22_X1 U23119 ( .A1(n20553), .A2(n20173), .B1(n20552), .B2(n20172), .ZN(
        n20171) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20174), .B1(
        n20187), .B2(n20632), .ZN(n20170) );
  OAI211_X1 U23121 ( .C1(n20556), .C2(n20177), .A(n20171), .B(n20170), .ZN(
        P1_U3071) );
  AOI22_X1 U23122 ( .A1(n20560), .A2(n20173), .B1(n20558), .B2(n20172), .ZN(
        n20176) );
  INV_X1 U23123 ( .A(n20509), .ZN(n20643) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20174), .B1(
        n20187), .B2(n20643), .ZN(n20175) );
  OAI211_X1 U23125 ( .C1(n20565), .C2(n20177), .A(n20176), .B(n20175), .ZN(
        P1_U3072) );
  OR2_X1 U23126 ( .A1(n20464), .A2(n20178), .ZN(n20209) );
  NAND2_X1 U23127 ( .A1(n20251), .A2(n20465), .ZN(n20179) );
  NAND2_X1 U23128 ( .A1(n20179), .A2(n20209), .ZN(n20183) );
  NAND2_X1 U23129 ( .A1(n20183), .A2(n20576), .ZN(n20181) );
  NAND2_X1 U23130 ( .A1(n20186), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20180) );
  INV_X1 U23131 ( .A(n20513), .ZN(n20581) );
  OAI22_X1 U23132 ( .A1(n20582), .A2(n20209), .B1(n20208), .B2(n20581), .ZN(
        n20182) );
  INV_X1 U23133 ( .A(n20182), .ZN(n20189) );
  INV_X1 U23134 ( .A(n20183), .ZN(n20184) );
  OAI21_X1 U23135 ( .B1(n20259), .B2(n20757), .A(n20184), .ZN(n20185) );
  OAI221_X1 U23136 ( .B1(n20576), .B2(n20186), .C1(n20573), .C2(n20185), .A(
        n20472), .ZN(n20212) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20212), .B1(
        n20187), .B2(n20584), .ZN(n20188) );
  OAI211_X1 U23138 ( .C1(n20477), .C2(n20250), .A(n20189), .B(n20188), .ZN(
        P1_U3073) );
  INV_X1 U23139 ( .A(n20527), .ZN(n20588) );
  OAI22_X1 U23140 ( .A1(n20589), .A2(n20209), .B1(n20208), .B2(n20588), .ZN(
        n20190) );
  INV_X1 U23141 ( .A(n20190), .ZN(n20192) );
  AOI22_X1 U23142 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20212), .B1(
        n20211), .B2(n20591), .ZN(n20191) );
  OAI211_X1 U23143 ( .C1(n20531), .C2(n20215), .A(n20192), .B(n20191), .ZN(
        P1_U3074) );
  INV_X1 U23144 ( .A(n20532), .ZN(n20596) );
  OAI22_X1 U23145 ( .A1(n20597), .A2(n20209), .B1(n20208), .B2(n20596), .ZN(
        n20193) );
  INV_X1 U23146 ( .A(n20193), .ZN(n20195) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20212), .B1(
        n20211), .B2(n20599), .ZN(n20194) );
  OAI211_X1 U23148 ( .C1(n20536), .C2(n20215), .A(n20195), .B(n20194), .ZN(
        P1_U3075) );
  INV_X1 U23149 ( .A(n20537), .ZN(n20604) );
  OAI22_X1 U23150 ( .A1(n20605), .A2(n20209), .B1(n20208), .B2(n20604), .ZN(
        n20196) );
  INV_X1 U23151 ( .A(n20196), .ZN(n20198) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20212), .B1(
        n20211), .B2(n20608), .ZN(n20197) );
  OAI211_X1 U23153 ( .C1(n20541), .C2(n20215), .A(n20198), .B(n20197), .ZN(
        P1_U3076) );
  INV_X1 U23154 ( .A(n20542), .ZN(n20612) );
  OAI22_X1 U23155 ( .A1(n20613), .A2(n20209), .B1(n20208), .B2(n20612), .ZN(
        n20199) );
  INV_X1 U23156 ( .A(n20199), .ZN(n20201) );
  AOI22_X1 U23157 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20212), .B1(
        n20211), .B2(n20616), .ZN(n20200) );
  OAI211_X1 U23158 ( .C1(n20546), .C2(n20215), .A(n20201), .B(n20200), .ZN(
        P1_U3077) );
  INV_X1 U23159 ( .A(n20547), .ZN(n20620) );
  OAI22_X1 U23160 ( .A1(n20621), .A2(n20209), .B1(n20208), .B2(n20620), .ZN(
        n20202) );
  INV_X1 U23161 ( .A(n20202), .ZN(n20204) );
  AOI22_X1 U23162 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20212), .B1(
        n20211), .B2(n20624), .ZN(n20203) );
  OAI211_X1 U23163 ( .C1(n20551), .C2(n20215), .A(n20204), .B(n20203), .ZN(
        P1_U3078) );
  INV_X1 U23164 ( .A(n20552), .ZN(n20628) );
  OAI22_X1 U23165 ( .A1(n20629), .A2(n20209), .B1(n20208), .B2(n20628), .ZN(
        n20205) );
  INV_X1 U23166 ( .A(n20205), .ZN(n20207) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20212), .B1(
        n20211), .B2(n20632), .ZN(n20206) );
  OAI211_X1 U23168 ( .C1(n20556), .C2(n20215), .A(n20207), .B(n20206), .ZN(
        P1_U3079) );
  INV_X1 U23169 ( .A(n20558), .ZN(n20636) );
  OAI22_X1 U23170 ( .A1(n20639), .A2(n20209), .B1(n20208), .B2(n20636), .ZN(
        n20210) );
  INV_X1 U23171 ( .A(n20210), .ZN(n20214) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20212), .B1(
        n20211), .B2(n20643), .ZN(n20213) );
  OAI211_X1 U23173 ( .C1(n20565), .C2(n20215), .A(n20214), .B(n20213), .ZN(
        P1_U3080) );
  OR2_X1 U23174 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20260), .ZN(
        n20244) );
  OAI22_X1 U23175 ( .A1(n20250), .A2(n20526), .B1(n20582), .B2(n20244), .ZN(
        n20216) );
  INV_X1 U23176 ( .A(n20216), .ZN(n20225) );
  NAND3_X1 U23177 ( .A1(n20250), .A2(n20576), .A3(n20291), .ZN(n20217) );
  NAND2_X1 U23178 ( .A1(n20217), .A2(n20431), .ZN(n20220) );
  NAND2_X1 U23179 ( .A1(n20251), .A2(n20519), .ZN(n20222) );
  AOI22_X1 U23180 ( .A1(n20220), .A2(n20222), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20244), .ZN(n20219) );
  NAND3_X1 U23181 ( .A1(n20522), .A2(n20219), .A3(n20218), .ZN(n20247) );
  INV_X1 U23182 ( .A(n20220), .ZN(n20223) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20247), .B1(
        n20513), .B2(n20246), .ZN(n20224) );
  OAI211_X1 U23184 ( .C1(n20477), .C2(n20291), .A(n20225), .B(n20224), .ZN(
        P1_U3081) );
  OAI22_X1 U23185 ( .A1(n20589), .A2(n20244), .B1(n20291), .B2(n20481), .ZN(
        n20226) );
  INV_X1 U23186 ( .A(n20226), .ZN(n20228) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20247), .B1(
        n20527), .B2(n20246), .ZN(n20227) );
  OAI211_X1 U23188 ( .C1(n20531), .C2(n20250), .A(n20228), .B(n20227), .ZN(
        P1_U3082) );
  OAI22_X1 U23189 ( .A1(n20597), .A2(n20244), .B1(n20291), .B2(n20485), .ZN(
        n20229) );
  INV_X1 U23190 ( .A(n20229), .ZN(n20231) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20247), .B1(
        n20532), .B2(n20246), .ZN(n20230) );
  OAI211_X1 U23192 ( .C1(n20536), .C2(n20250), .A(n20231), .B(n20230), .ZN(
        P1_U3083) );
  OAI22_X1 U23193 ( .A1(n20605), .A2(n20244), .B1(n20291), .B2(n20489), .ZN(
        n20232) );
  INV_X1 U23194 ( .A(n20232), .ZN(n20234) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20247), .B1(
        n20537), .B2(n20246), .ZN(n20233) );
  OAI211_X1 U23196 ( .C1(n20541), .C2(n20250), .A(n20234), .B(n20233), .ZN(
        P1_U3084) );
  OAI22_X1 U23197 ( .A1(n20250), .A2(n20546), .B1(n20613), .B2(n20244), .ZN(
        n20235) );
  INV_X1 U23198 ( .A(n20235), .ZN(n20237) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20247), .B1(
        n20542), .B2(n20246), .ZN(n20236) );
  OAI211_X1 U23200 ( .C1(n20493), .C2(n20291), .A(n20237), .B(n20236), .ZN(
        P1_U3085) );
  OAI22_X1 U23201 ( .A1(n20250), .A2(n20551), .B1(n20621), .B2(n20244), .ZN(
        n20238) );
  INV_X1 U23202 ( .A(n20238), .ZN(n20240) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20247), .B1(
        n20547), .B2(n20246), .ZN(n20239) );
  OAI211_X1 U23204 ( .C1(n20497), .C2(n20291), .A(n20240), .B(n20239), .ZN(
        P1_U3086) );
  OAI22_X1 U23205 ( .A1(n20250), .A2(n20556), .B1(n20629), .B2(n20244), .ZN(
        n20241) );
  INV_X1 U23206 ( .A(n20241), .ZN(n20243) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20247), .B1(
        n20552), .B2(n20246), .ZN(n20242) );
  OAI211_X1 U23208 ( .C1(n20501), .C2(n20291), .A(n20243), .B(n20242), .ZN(
        P1_U3087) );
  OAI22_X1 U23209 ( .A1(n20639), .A2(n20244), .B1(n20291), .B2(n20509), .ZN(
        n20245) );
  INV_X1 U23210 ( .A(n20245), .ZN(n20249) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20247), .B1(
        n20558), .B2(n20246), .ZN(n20248) );
  OAI211_X1 U23212 ( .C1(n20565), .C2(n20250), .A(n20249), .B(n20248), .ZN(
        P1_U3088) );
  NAND2_X1 U23213 ( .A1(n20251), .A2(n20567), .ZN(n20252) );
  NAND2_X1 U23214 ( .A1(n20252), .A2(n20286), .ZN(n20253) );
  NAND2_X1 U23215 ( .A1(n20253), .A2(n20576), .ZN(n20256) );
  NAND2_X1 U23216 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20254), .ZN(n20255) );
  AND2_X1 U23217 ( .A1(n20256), .A2(n20255), .ZN(n20285) );
  OAI22_X1 U23218 ( .A1(n20582), .A2(n20286), .B1(n20285), .B2(n20581), .ZN(
        n20257) );
  INV_X1 U23219 ( .A(n20257), .ZN(n20264) );
  OR2_X1 U23220 ( .A1(n20259), .A2(n20258), .ZN(n20732) );
  INV_X1 U23221 ( .A(n20472), .ZN(n20572) );
  AOI21_X1 U23222 ( .B1(n20260), .B2(n20732), .A(n20572), .ZN(n20261) );
  NAND2_X1 U23223 ( .A1(n20262), .A2(n9654), .ZN(n20284) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20288), .B1(
        n20318), .B2(n20585), .ZN(n20263) );
  OAI211_X1 U23225 ( .C1(n20526), .C2(n20291), .A(n20264), .B(n20263), .ZN(
        P1_U3089) );
  OAI22_X1 U23226 ( .A1(n20589), .A2(n20286), .B1(n20285), .B2(n20588), .ZN(
        n20265) );
  INV_X1 U23227 ( .A(n20265), .ZN(n20267) );
  INV_X1 U23228 ( .A(n20291), .ZN(n20281) );
  AOI22_X1 U23229 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20288), .B1(
        n20281), .B2(n20592), .ZN(n20266) );
  OAI211_X1 U23230 ( .C1(n20481), .C2(n20284), .A(n20267), .B(n20266), .ZN(
        P1_U3090) );
  OAI22_X1 U23231 ( .A1(n20597), .A2(n20286), .B1(n20285), .B2(n20596), .ZN(
        n20268) );
  INV_X1 U23232 ( .A(n20268), .ZN(n20270) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20288), .B1(
        n20318), .B2(n20599), .ZN(n20269) );
  OAI211_X1 U23234 ( .C1(n20536), .C2(n20291), .A(n20270), .B(n20269), .ZN(
        P1_U3091) );
  OAI22_X1 U23235 ( .A1(n20605), .A2(n20286), .B1(n20285), .B2(n20604), .ZN(
        n20271) );
  INV_X1 U23236 ( .A(n20271), .ZN(n20273) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20288), .B1(
        n20281), .B2(n20607), .ZN(n20272) );
  OAI211_X1 U23238 ( .C1(n20489), .C2(n20284), .A(n20273), .B(n20272), .ZN(
        P1_U3092) );
  OAI22_X1 U23239 ( .A1(n20613), .A2(n20286), .B1(n20285), .B2(n20612), .ZN(
        n20274) );
  INV_X1 U23240 ( .A(n20274), .ZN(n20276) );
  AOI22_X1 U23241 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20288), .B1(
        n20281), .B2(n20615), .ZN(n20275) );
  OAI211_X1 U23242 ( .C1(n20493), .C2(n20284), .A(n20276), .B(n20275), .ZN(
        P1_U3093) );
  OAI22_X1 U23243 ( .A1(n20621), .A2(n20286), .B1(n20285), .B2(n20620), .ZN(
        n20277) );
  INV_X1 U23244 ( .A(n20277), .ZN(n20279) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20288), .B1(
        n20318), .B2(n20624), .ZN(n20278) );
  OAI211_X1 U23246 ( .C1(n20551), .C2(n20291), .A(n20279), .B(n20278), .ZN(
        P1_U3094) );
  OAI22_X1 U23247 ( .A1(n20629), .A2(n20286), .B1(n20285), .B2(n20628), .ZN(
        n20280) );
  INV_X1 U23248 ( .A(n20280), .ZN(n20283) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20288), .B1(
        n20281), .B2(n20631), .ZN(n20282) );
  OAI211_X1 U23250 ( .C1(n20501), .C2(n20284), .A(n20283), .B(n20282), .ZN(
        P1_U3095) );
  OAI22_X1 U23251 ( .A1(n20639), .A2(n20286), .B1(n20285), .B2(n20636), .ZN(
        n20287) );
  INV_X1 U23252 ( .A(n20287), .ZN(n20290) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20288), .B1(
        n20318), .B2(n20643), .ZN(n20289) );
  OAI211_X1 U23254 ( .C1(n20565), .C2(n20291), .A(n20290), .B(n20289), .ZN(
        P1_U3096) );
  INV_X1 U23255 ( .A(n20292), .ZN(n20293) );
  NOR3_X1 U23256 ( .A1(n20737), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20327) );
  INV_X1 U23257 ( .A(n20327), .ZN(n20323) );
  NOR2_X1 U23258 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20323), .ZN(
        n20317) );
  NAND2_X1 U23259 ( .A1(n20727), .A2(n12915), .ZN(n20390) );
  INV_X1 U23260 ( .A(n20390), .ZN(n20322) );
  AOI21_X1 U23261 ( .B1(n20322), .B2(n20433), .A(n20317), .ZN(n20298) );
  NOR2_X1 U23262 ( .A1(n20296), .A2(n20295), .ZN(n20436) );
  INV_X1 U23263 ( .A(n20436), .ZN(n20438) );
  OAI22_X1 U23264 ( .A1(n20298), .A2(n20573), .B1(n20358), .B2(n20438), .ZN(
        n20316) );
  AOI22_X1 U23265 ( .A1(n20514), .A2(n20317), .B1(n20513), .B2(n20316), .ZN(
        n20303) );
  INV_X1 U23266 ( .A(n20349), .ZN(n20297) );
  OAI21_X1 U23267 ( .B1(n20318), .B2(n20297), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20299) );
  NAND2_X1 U23268 ( .A1(n20299), .A2(n20298), .ZN(n20300) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20584), .ZN(n20302) );
  OAI211_X1 U23270 ( .C1(n20477), .C2(n20349), .A(n20303), .B(n20302), .ZN(
        P1_U3097) );
  AOI22_X1 U23271 ( .A1(n20528), .A2(n20317), .B1(n20527), .B2(n20316), .ZN(
        n20305) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20592), .ZN(n20304) );
  OAI211_X1 U23273 ( .C1(n20481), .C2(n20349), .A(n20305), .B(n20304), .ZN(
        P1_U3098) );
  AOI22_X1 U23274 ( .A1(n20533), .A2(n20317), .B1(n20532), .B2(n20316), .ZN(
        n20307) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20600), .ZN(n20306) );
  OAI211_X1 U23276 ( .C1(n20485), .C2(n20349), .A(n20307), .B(n20306), .ZN(
        P1_U3099) );
  AOI22_X1 U23277 ( .A1(n20538), .A2(n20317), .B1(n20537), .B2(n20316), .ZN(
        n20309) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20607), .ZN(n20308) );
  OAI211_X1 U23279 ( .C1(n20489), .C2(n20349), .A(n20309), .B(n20308), .ZN(
        P1_U3100) );
  AOI22_X1 U23280 ( .A1(n20543), .A2(n20317), .B1(n20542), .B2(n20316), .ZN(
        n20311) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20615), .ZN(n20310) );
  OAI211_X1 U23282 ( .C1(n20493), .C2(n20349), .A(n20311), .B(n20310), .ZN(
        P1_U3101) );
  AOI22_X1 U23283 ( .A1(n20548), .A2(n20317), .B1(n20547), .B2(n20316), .ZN(
        n20313) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20623), .ZN(n20312) );
  OAI211_X1 U23285 ( .C1(n20497), .C2(n20349), .A(n20313), .B(n20312), .ZN(
        P1_U3102) );
  AOI22_X1 U23286 ( .A1(n20553), .A2(n20317), .B1(n20552), .B2(n20316), .ZN(
        n20315) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20631), .ZN(n20314) );
  OAI211_X1 U23288 ( .C1(n20501), .C2(n20349), .A(n20315), .B(n20314), .ZN(
        P1_U3103) );
  AOI22_X1 U23289 ( .A1(n20560), .A2(n20317), .B1(n20558), .B2(n20316), .ZN(
        n20321) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20319), .B1(
        n20318), .B2(n20641), .ZN(n20320) );
  OAI211_X1 U23291 ( .C1(n20509), .C2(n20349), .A(n20321), .B(n20320), .ZN(
        P1_U3104) );
  NOR2_X1 U23292 ( .A1(n20464), .A2(n20323), .ZN(n20344) );
  AOI21_X1 U23293 ( .B1(n20322), .B2(n20465), .A(n20344), .ZN(n20324) );
  OAI22_X1 U23294 ( .A1(n20324), .A2(n20573), .B1(n20323), .B2(n20750), .ZN(
        n20343) );
  AOI22_X1 U23295 ( .A1(n20514), .A2(n20344), .B1(n20513), .B2(n20343), .ZN(
        n20330) );
  INV_X1 U23296 ( .A(n20726), .ZN(n20325) );
  OAI21_X1 U23297 ( .B1(n20325), .B2(n20757), .A(n20324), .ZN(n20326) );
  OAI221_X1 U23298 ( .B1(n20576), .B2(n20327), .C1(n20573), .C2(n20326), .A(
        n20472), .ZN(n20346) );
  NOR2_X1 U23299 ( .A1(n9654), .A2(n9650), .ZN(n20328) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20585), .ZN(n20329) );
  OAI211_X1 U23301 ( .C1(n20526), .C2(n20349), .A(n20330), .B(n20329), .ZN(
        P1_U3105) );
  AOI22_X1 U23302 ( .A1(n20528), .A2(n20344), .B1(n20527), .B2(n20343), .ZN(
        n20332) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20591), .ZN(n20331) );
  OAI211_X1 U23304 ( .C1(n20531), .C2(n20349), .A(n20332), .B(n20331), .ZN(
        P1_U3106) );
  AOI22_X1 U23305 ( .A1(n20533), .A2(n20344), .B1(n20532), .B2(n20343), .ZN(
        n20334) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20599), .ZN(n20333) );
  OAI211_X1 U23307 ( .C1(n20536), .C2(n20349), .A(n20334), .B(n20333), .ZN(
        P1_U3107) );
  AOI22_X1 U23308 ( .A1(n20538), .A2(n20344), .B1(n20537), .B2(n20343), .ZN(
        n20336) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20608), .ZN(n20335) );
  OAI211_X1 U23310 ( .C1(n20541), .C2(n20349), .A(n20336), .B(n20335), .ZN(
        P1_U3108) );
  AOI22_X1 U23311 ( .A1(n20543), .A2(n20344), .B1(n20542), .B2(n20343), .ZN(
        n20338) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20616), .ZN(n20337) );
  OAI211_X1 U23313 ( .C1(n20546), .C2(n20349), .A(n20338), .B(n20337), .ZN(
        P1_U3109) );
  AOI22_X1 U23314 ( .A1(n20548), .A2(n20344), .B1(n20547), .B2(n20343), .ZN(
        n20340) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20624), .ZN(n20339) );
  OAI211_X1 U23316 ( .C1(n20551), .C2(n20349), .A(n20340), .B(n20339), .ZN(
        P1_U3110) );
  AOI22_X1 U23317 ( .A1(n20553), .A2(n20344), .B1(n20552), .B2(n20343), .ZN(
        n20342) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20632), .ZN(n20341) );
  OAI211_X1 U23319 ( .C1(n20556), .C2(n20349), .A(n20342), .B(n20341), .ZN(
        P1_U3111) );
  AOI22_X1 U23320 ( .A1(n20560), .A2(n20344), .B1(n20558), .B2(n20343), .ZN(
        n20348) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20643), .ZN(n20347) );
  OAI211_X1 U23322 ( .C1(n20565), .C2(n20349), .A(n20348), .B(n20347), .ZN(
        P1_U3112) );
  NAND2_X1 U23323 ( .A1(n20726), .A2(n9654), .ZN(n20396) );
  NOR3_X1 U23324 ( .A1(n20737), .A2(n20351), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20397) );
  NAND2_X1 U23325 ( .A1(n20464), .A2(n20397), .ZN(n20381) );
  OAI22_X1 U23326 ( .A1(n20417), .A2(n20477), .B1(n20582), .B2(n20381), .ZN(
        n20352) );
  INV_X1 U23327 ( .A(n20352), .ZN(n20362) );
  AOI21_X1 U23328 ( .B1(n20417), .B2(n20387), .A(n20757), .ZN(n20353) );
  NOR2_X1 U23329 ( .A1(n20353), .A2(n20573), .ZN(n20357) );
  OR2_X1 U23330 ( .A1(n20390), .A2(n20433), .ZN(n20359) );
  AOI22_X1 U23331 ( .A1(n20357), .A2(n20359), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20381), .ZN(n20355) );
  OR2_X1 U23332 ( .A1(n20354), .A2(n20737), .ZN(n20511) );
  NAND2_X1 U23333 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20511), .ZN(n20521) );
  NAND3_X1 U23334 ( .A1(n20356), .A2(n20355), .A3(n20521), .ZN(n20384) );
  INV_X1 U23335 ( .A(n20357), .ZN(n20360) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20384), .B1(
        n20513), .B2(n20383), .ZN(n20361) );
  OAI211_X1 U23337 ( .C1(n20526), .C2(n20387), .A(n20362), .B(n20361), .ZN(
        P1_U3113) );
  OAI22_X1 U23338 ( .A1(n20417), .A2(n20481), .B1(n20381), .B2(n20589), .ZN(
        n20363) );
  INV_X1 U23339 ( .A(n20363), .ZN(n20365) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20384), .B1(
        n20527), .B2(n20383), .ZN(n20364) );
  OAI211_X1 U23341 ( .C1(n20531), .C2(n20387), .A(n20365), .B(n20364), .ZN(
        P1_U3114) );
  OAI22_X1 U23342 ( .A1(n20417), .A2(n20485), .B1(n20381), .B2(n20597), .ZN(
        n20366) );
  INV_X1 U23343 ( .A(n20366), .ZN(n20368) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20384), .B1(
        n20532), .B2(n20383), .ZN(n20367) );
  OAI211_X1 U23345 ( .C1(n20536), .C2(n20387), .A(n20368), .B(n20367), .ZN(
        P1_U3115) );
  OAI22_X1 U23346 ( .A1(n20417), .A2(n20489), .B1(n20381), .B2(n20605), .ZN(
        n20369) );
  INV_X1 U23347 ( .A(n20369), .ZN(n20371) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20384), .B1(
        n20537), .B2(n20383), .ZN(n20370) );
  OAI211_X1 U23349 ( .C1(n20541), .C2(n20387), .A(n20371), .B(n20370), .ZN(
        P1_U3116) );
  OAI22_X1 U23350 ( .A1(n20387), .A2(n20546), .B1(n20381), .B2(n20613), .ZN(
        n20372) );
  INV_X1 U23351 ( .A(n20372), .ZN(n20374) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20384), .B1(
        n20542), .B2(n20383), .ZN(n20373) );
  OAI211_X1 U23353 ( .C1(n20493), .C2(n20417), .A(n20374), .B(n20373), .ZN(
        P1_U3117) );
  OAI22_X1 U23354 ( .A1(n20417), .A2(n20497), .B1(n20381), .B2(n20621), .ZN(
        n20375) );
  INV_X1 U23355 ( .A(n20375), .ZN(n20377) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20384), .B1(
        n20547), .B2(n20383), .ZN(n20376) );
  OAI211_X1 U23357 ( .C1(n20551), .C2(n20387), .A(n20377), .B(n20376), .ZN(
        P1_U3118) );
  OAI22_X1 U23358 ( .A1(n20417), .A2(n20501), .B1(n20381), .B2(n20629), .ZN(
        n20378) );
  INV_X1 U23359 ( .A(n20378), .ZN(n20380) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20384), .B1(
        n20552), .B2(n20383), .ZN(n20379) );
  OAI211_X1 U23361 ( .C1(n20556), .C2(n20387), .A(n20380), .B(n20379), .ZN(
        P1_U3119) );
  OAI22_X1 U23362 ( .A1(n20417), .A2(n20509), .B1(n20381), .B2(n20639), .ZN(
        n20382) );
  INV_X1 U23363 ( .A(n20382), .ZN(n20386) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20384), .B1(
        n20558), .B2(n20383), .ZN(n20385) );
  OAI211_X1 U23365 ( .C1(n20565), .C2(n20387), .A(n20386), .B(n20385), .ZN(
        P1_U3120) );
  OR2_X1 U23366 ( .A1(n20388), .A2(n20737), .ZN(n20422) );
  OAI21_X1 U23367 ( .B1(n20390), .B2(n20389), .A(n20422), .ZN(n20391) );
  NAND2_X1 U23368 ( .A1(n20391), .A2(n20576), .ZN(n20393) );
  NAND2_X1 U23369 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20397), .ZN(n20392) );
  OAI22_X1 U23370 ( .A1(n20582), .A2(n20422), .B1(n20421), .B2(n20581), .ZN(
        n20394) );
  INV_X1 U23371 ( .A(n20394), .ZN(n20400) );
  NOR2_X1 U23372 ( .A1(n20396), .A2(n20395), .ZN(n20398) );
  INV_X1 U23373 ( .A(n20417), .ZN(n20424) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20584), .ZN(n20399) );
  OAI211_X1 U23375 ( .C1(n20477), .C2(n20460), .A(n20400), .B(n20399), .ZN(
        P1_U3121) );
  OAI22_X1 U23376 ( .A1(n20589), .A2(n20422), .B1(n20421), .B2(n20588), .ZN(
        n20401) );
  INV_X1 U23377 ( .A(n20401), .ZN(n20403) );
  INV_X1 U23378 ( .A(n20460), .ZN(n20414) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20425), .B1(
        n20414), .B2(n20591), .ZN(n20402) );
  OAI211_X1 U23380 ( .C1(n20531), .C2(n20417), .A(n20403), .B(n20402), .ZN(
        P1_U3122) );
  OAI22_X1 U23381 ( .A1(n20597), .A2(n20422), .B1(n20421), .B2(n20596), .ZN(
        n20404) );
  INV_X1 U23382 ( .A(n20404), .ZN(n20406) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20425), .B1(
        n20414), .B2(n20599), .ZN(n20405) );
  OAI211_X1 U23384 ( .C1(n20536), .C2(n20417), .A(n20406), .B(n20405), .ZN(
        P1_U3123) );
  OAI22_X1 U23385 ( .A1(n20605), .A2(n20422), .B1(n20421), .B2(n20604), .ZN(
        n20407) );
  INV_X1 U23386 ( .A(n20407), .ZN(n20409) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20425), .B1(
        n20414), .B2(n20608), .ZN(n20408) );
  OAI211_X1 U23388 ( .C1(n20541), .C2(n20417), .A(n20409), .B(n20408), .ZN(
        P1_U3124) );
  OAI22_X1 U23389 ( .A1(n20613), .A2(n20422), .B1(n20421), .B2(n20612), .ZN(
        n20410) );
  INV_X1 U23390 ( .A(n20410), .ZN(n20412) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20425), .B1(
        n20414), .B2(n20616), .ZN(n20411) );
  OAI211_X1 U23392 ( .C1(n20546), .C2(n20417), .A(n20412), .B(n20411), .ZN(
        P1_U3125) );
  OAI22_X1 U23393 ( .A1(n20621), .A2(n20422), .B1(n20421), .B2(n20620), .ZN(
        n20413) );
  INV_X1 U23394 ( .A(n20413), .ZN(n20416) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20425), .B1(
        n20414), .B2(n20624), .ZN(n20415) );
  OAI211_X1 U23396 ( .C1(n20551), .C2(n20417), .A(n20416), .B(n20415), .ZN(
        P1_U3126) );
  OAI22_X1 U23397 ( .A1(n20629), .A2(n20422), .B1(n20421), .B2(n20628), .ZN(
        n20418) );
  INV_X1 U23398 ( .A(n20418), .ZN(n20420) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20631), .ZN(n20419) );
  OAI211_X1 U23400 ( .C1(n20501), .C2(n20460), .A(n20420), .B(n20419), .ZN(
        P1_U3127) );
  OAI22_X1 U23401 ( .A1(n20639), .A2(n20422), .B1(n20421), .B2(n20636), .ZN(
        n20423) );
  INV_X1 U23402 ( .A(n20423), .ZN(n20427) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20641), .ZN(n20426) );
  OAI211_X1 U23404 ( .C1(n20509), .C2(n20460), .A(n20427), .B(n20426), .ZN(
        P1_U3128) );
  NOR3_X1 U23405 ( .A1(n20428), .A2(n20737), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20473) );
  NAND2_X1 U23406 ( .A1(n20464), .A2(n20473), .ZN(n20434) );
  INV_X1 U23407 ( .A(n20434), .ZN(n20455) );
  AOI22_X1 U23408 ( .A1(n20514), .A2(n20455), .B1(n20505), .B2(n20585), .ZN(
        n20442) );
  INV_X1 U23409 ( .A(n20505), .ZN(n20430) );
  NAND3_X1 U23410 ( .A1(n20460), .A2(n20576), .A3(n20430), .ZN(n20432) );
  NAND2_X1 U23411 ( .A1(n20432), .A2(n20431), .ZN(n20437) );
  NOR2_X1 U23412 ( .A1(n12915), .A2(n9812), .ZN(n20568) );
  NAND2_X1 U23413 ( .A1(n20568), .A2(n20433), .ZN(n20439) );
  AOI22_X1 U23414 ( .A1(n20437), .A2(n20439), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20434), .ZN(n20435) );
  OAI211_X1 U23415 ( .C1(n20436), .C2(n20750), .A(n20522), .B(n20435), .ZN(
        n20457) );
  INV_X1 U23416 ( .A(n20437), .ZN(n20440) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20457), .B1(
        n20513), .B2(n20456), .ZN(n20441) );
  OAI211_X1 U23418 ( .C1(n20526), .C2(n20460), .A(n20442), .B(n20441), .ZN(
        P1_U3129) );
  AOI22_X1 U23419 ( .A1(n20528), .A2(n20455), .B1(n20505), .B2(n20591), .ZN(
        n20444) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20457), .B1(
        n20527), .B2(n20456), .ZN(n20443) );
  OAI211_X1 U23421 ( .C1(n20531), .C2(n20460), .A(n20444), .B(n20443), .ZN(
        P1_U3130) );
  AOI22_X1 U23422 ( .A1(n20533), .A2(n20455), .B1(n20505), .B2(n20599), .ZN(
        n20446) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20457), .B1(
        n20532), .B2(n20456), .ZN(n20445) );
  OAI211_X1 U23424 ( .C1(n20536), .C2(n20460), .A(n20446), .B(n20445), .ZN(
        P1_U3131) );
  AOI22_X1 U23425 ( .A1(n20538), .A2(n20455), .B1(n20505), .B2(n20608), .ZN(
        n20448) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20457), .B1(
        n20537), .B2(n20456), .ZN(n20447) );
  OAI211_X1 U23427 ( .C1(n20541), .C2(n20460), .A(n20448), .B(n20447), .ZN(
        P1_U3132) );
  AOI22_X1 U23428 ( .A1(n20543), .A2(n20455), .B1(n20505), .B2(n20616), .ZN(
        n20450) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20457), .B1(
        n20542), .B2(n20456), .ZN(n20449) );
  OAI211_X1 U23430 ( .C1(n20546), .C2(n20460), .A(n20450), .B(n20449), .ZN(
        P1_U3133) );
  AOI22_X1 U23431 ( .A1(n20548), .A2(n20455), .B1(n20505), .B2(n20624), .ZN(
        n20452) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20457), .B1(
        n20547), .B2(n20456), .ZN(n20451) );
  OAI211_X1 U23433 ( .C1(n20551), .C2(n20460), .A(n20452), .B(n20451), .ZN(
        P1_U3134) );
  AOI22_X1 U23434 ( .A1(n20553), .A2(n20455), .B1(n20505), .B2(n20632), .ZN(
        n20454) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20457), .B1(
        n20552), .B2(n20456), .ZN(n20453) );
  OAI211_X1 U23436 ( .C1(n20556), .C2(n20460), .A(n20454), .B(n20453), .ZN(
        P1_U3135) );
  AOI22_X1 U23437 ( .A1(n20560), .A2(n20455), .B1(n20505), .B2(n20643), .ZN(
        n20459) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20457), .B1(
        n20558), .B2(n20456), .ZN(n20458) );
  OAI211_X1 U23439 ( .C1(n20565), .C2(n20460), .A(n20459), .B(n20458), .ZN(
        P1_U3136) );
  INV_X1 U23440 ( .A(n20473), .ZN(n20463) );
  OR2_X1 U23441 ( .A1(n20464), .A2(n20463), .ZN(n20503) );
  NAND2_X1 U23442 ( .A1(n20568), .A2(n20465), .ZN(n20466) );
  NAND2_X1 U23443 ( .A1(n20466), .A2(n20503), .ZN(n20467) );
  NAND2_X1 U23444 ( .A1(n20467), .A2(n20576), .ZN(n20469) );
  NAND2_X1 U23445 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20473), .ZN(n20468) );
  AND2_X1 U23446 ( .A1(n20469), .A2(n20468), .ZN(n20502) );
  OAI22_X1 U23447 ( .A1(n20582), .A2(n20503), .B1(n20502), .B2(n20581), .ZN(
        n20470) );
  INV_X1 U23448 ( .A(n20470), .ZN(n20476) );
  NAND2_X1 U23449 ( .A1(n20571), .A2(n20471), .ZN(n20731) );
  INV_X1 U23450 ( .A(n20731), .ZN(n20474) );
  OAI21_X1 U23451 ( .B1(n20474), .B2(n20473), .A(n20472), .ZN(n20506) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20506), .B1(
        n20505), .B2(n20584), .ZN(n20475) );
  OAI211_X1 U23453 ( .C1(n20477), .C2(n20564), .A(n20476), .B(n20475), .ZN(
        P1_U3137) );
  OAI22_X1 U23454 ( .A1(n20589), .A2(n20503), .B1(n20502), .B2(n20588), .ZN(
        n20478) );
  INV_X1 U23455 ( .A(n20478), .ZN(n20480) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20506), .B1(
        n20505), .B2(n20592), .ZN(n20479) );
  OAI211_X1 U23457 ( .C1(n20481), .C2(n20564), .A(n20480), .B(n20479), .ZN(
        P1_U3138) );
  OAI22_X1 U23458 ( .A1(n20597), .A2(n20503), .B1(n20502), .B2(n20596), .ZN(
        n20482) );
  INV_X1 U23459 ( .A(n20482), .ZN(n20484) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20506), .B1(
        n20505), .B2(n20600), .ZN(n20483) );
  OAI211_X1 U23461 ( .C1(n20485), .C2(n20564), .A(n20484), .B(n20483), .ZN(
        P1_U3139) );
  OAI22_X1 U23462 ( .A1(n20605), .A2(n20503), .B1(n20502), .B2(n20604), .ZN(
        n20486) );
  INV_X1 U23463 ( .A(n20486), .ZN(n20488) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20506), .B1(
        n20505), .B2(n20607), .ZN(n20487) );
  OAI211_X1 U23465 ( .C1(n20489), .C2(n20564), .A(n20488), .B(n20487), .ZN(
        P1_U3140) );
  OAI22_X1 U23466 ( .A1(n20613), .A2(n20503), .B1(n20502), .B2(n20612), .ZN(
        n20490) );
  INV_X1 U23467 ( .A(n20490), .ZN(n20492) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20506), .B1(
        n20505), .B2(n20615), .ZN(n20491) );
  OAI211_X1 U23469 ( .C1(n20493), .C2(n20564), .A(n20492), .B(n20491), .ZN(
        P1_U3141) );
  OAI22_X1 U23470 ( .A1(n20621), .A2(n20503), .B1(n20502), .B2(n20620), .ZN(
        n20494) );
  INV_X1 U23471 ( .A(n20494), .ZN(n20496) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20506), .B1(
        n20505), .B2(n20623), .ZN(n20495) );
  OAI211_X1 U23473 ( .C1(n20497), .C2(n20564), .A(n20496), .B(n20495), .ZN(
        P1_U3142) );
  OAI22_X1 U23474 ( .A1(n20629), .A2(n20503), .B1(n20502), .B2(n20628), .ZN(
        n20498) );
  INV_X1 U23475 ( .A(n20498), .ZN(n20500) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20506), .B1(
        n20505), .B2(n20631), .ZN(n20499) );
  OAI211_X1 U23477 ( .C1(n20501), .C2(n20564), .A(n20500), .B(n20499), .ZN(
        P1_U3143) );
  OAI22_X1 U23478 ( .A1(n20639), .A2(n20503), .B1(n20502), .B2(n20636), .ZN(
        n20504) );
  INV_X1 U23479 ( .A(n20504), .ZN(n20508) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20506), .B1(
        n20505), .B2(n20641), .ZN(n20507) );
  OAI211_X1 U23481 ( .C1(n20509), .C2(n20564), .A(n20508), .B(n20507), .ZN(
        P1_U3144) );
  NOR2_X1 U23482 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20574), .ZN(
        n20559) );
  NAND3_X1 U23483 ( .A1(n20568), .A2(n20519), .A3(n20576), .ZN(n20510) );
  OAI21_X1 U23484 ( .B1(n20512), .B2(n20511), .A(n20510), .ZN(n20557) );
  AOI22_X1 U23485 ( .A1(n20514), .A2(n20559), .B1(n20513), .B2(n20557), .ZN(
        n20525) );
  INV_X1 U23486 ( .A(n20515), .ZN(n20516) );
  INV_X1 U23487 ( .A(n20642), .ZN(n20517) );
  AOI21_X1 U23488 ( .B1(n20517), .B2(n20564), .A(n20757), .ZN(n20518) );
  AOI21_X1 U23489 ( .B1(n20568), .B2(n20519), .A(n20518), .ZN(n20520) );
  NOR2_X1 U23490 ( .A1(n20520), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20523) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20561), .B1(
        n20642), .B2(n20585), .ZN(n20524) );
  OAI211_X1 U23492 ( .C1(n20526), .C2(n20564), .A(n20525), .B(n20524), .ZN(
        P1_U3145) );
  AOI22_X1 U23493 ( .A1(n20528), .A2(n20559), .B1(n20527), .B2(n20557), .ZN(
        n20530) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20561), .B1(
        n20642), .B2(n20591), .ZN(n20529) );
  OAI211_X1 U23495 ( .C1(n20531), .C2(n20564), .A(n20530), .B(n20529), .ZN(
        P1_U3146) );
  AOI22_X1 U23496 ( .A1(n20533), .A2(n20559), .B1(n20532), .B2(n20557), .ZN(
        n20535) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20561), .B1(
        n20642), .B2(n20599), .ZN(n20534) );
  OAI211_X1 U23498 ( .C1(n20536), .C2(n20564), .A(n20535), .B(n20534), .ZN(
        P1_U3147) );
  AOI22_X1 U23499 ( .A1(n20538), .A2(n20559), .B1(n20537), .B2(n20557), .ZN(
        n20540) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20561), .B1(
        n20642), .B2(n20608), .ZN(n20539) );
  OAI211_X1 U23501 ( .C1(n20541), .C2(n20564), .A(n20540), .B(n20539), .ZN(
        P1_U3148) );
  AOI22_X1 U23502 ( .A1(n20543), .A2(n20559), .B1(n20542), .B2(n20557), .ZN(
        n20545) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20561), .B1(
        n20642), .B2(n20616), .ZN(n20544) );
  OAI211_X1 U23504 ( .C1(n20546), .C2(n20564), .A(n20545), .B(n20544), .ZN(
        P1_U3149) );
  AOI22_X1 U23505 ( .A1(n20548), .A2(n20559), .B1(n20547), .B2(n20557), .ZN(
        n20550) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20561), .B1(
        n20642), .B2(n20624), .ZN(n20549) );
  OAI211_X1 U23507 ( .C1(n20551), .C2(n20564), .A(n20550), .B(n20549), .ZN(
        P1_U3150) );
  AOI22_X1 U23508 ( .A1(n20553), .A2(n20559), .B1(n20552), .B2(n20557), .ZN(
        n20555) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20561), .B1(
        n20642), .B2(n20632), .ZN(n20554) );
  OAI211_X1 U23510 ( .C1(n20556), .C2(n20564), .A(n20555), .B(n20554), .ZN(
        P1_U3151) );
  AOI22_X1 U23511 ( .A1(n20560), .A2(n20559), .B1(n20558), .B2(n20557), .ZN(
        n20563) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20561), .B1(
        n20642), .B2(n20643), .ZN(n20562) );
  OAI211_X1 U23513 ( .C1(n20565), .C2(n20564), .A(n20563), .B(n20562), .ZN(
        P1_U3152) );
  INV_X1 U23514 ( .A(n20566), .ZN(n20570) );
  NAND2_X1 U23515 ( .A1(n20568), .A2(n20567), .ZN(n20569) );
  NAND2_X1 U23516 ( .A1(n20569), .A2(n20638), .ZN(n20577) );
  AOI21_X1 U23517 ( .B1(n20571), .B2(n20570), .A(n20577), .ZN(n20575) );
  AOI221_X2 U23518 ( .B1(n20575), .B2(n20576), .C1(n20574), .C2(n20573), .A(
        n20572), .ZN(n20648) );
  INV_X1 U23519 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20915) );
  NAND2_X1 U23520 ( .A1(n20577), .A2(n20576), .ZN(n20580) );
  NAND2_X1 U23521 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20578), .ZN(n20579) );
  OAI22_X1 U23522 ( .A1(n20582), .A2(n20638), .B1(n20637), .B2(n20581), .ZN(
        n20583) );
  INV_X1 U23523 ( .A(n20583), .ZN(n20587) );
  AOI22_X1 U23524 ( .A1(n20644), .A2(n20585), .B1(n20642), .B2(n20584), .ZN(
        n20586) );
  OAI211_X1 U23525 ( .C1(n20648), .C2(n20915), .A(n20587), .B(n20586), .ZN(
        P1_U3153) );
  INV_X1 U23526 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20595) );
  OAI22_X1 U23527 ( .A1(n20589), .A2(n20638), .B1(n20637), .B2(n20588), .ZN(
        n20590) );
  INV_X1 U23528 ( .A(n20590), .ZN(n20594) );
  AOI22_X1 U23529 ( .A1(n20642), .A2(n20592), .B1(n20644), .B2(n20591), .ZN(
        n20593) );
  OAI211_X1 U23530 ( .C1(n20648), .C2(n20595), .A(n20594), .B(n20593), .ZN(
        P1_U3154) );
  INV_X1 U23531 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20603) );
  OAI22_X1 U23532 ( .A1(n20597), .A2(n20638), .B1(n20637), .B2(n20596), .ZN(
        n20598) );
  INV_X1 U23533 ( .A(n20598), .ZN(n20602) );
  AOI22_X1 U23534 ( .A1(n20642), .A2(n20600), .B1(n20644), .B2(n20599), .ZN(
        n20601) );
  OAI211_X1 U23535 ( .C1(n20648), .C2(n20603), .A(n20602), .B(n20601), .ZN(
        P1_U3155) );
  INV_X1 U23536 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20611) );
  OAI22_X1 U23537 ( .A1(n20605), .A2(n20638), .B1(n20637), .B2(n20604), .ZN(
        n20606) );
  INV_X1 U23538 ( .A(n20606), .ZN(n20610) );
  AOI22_X1 U23539 ( .A1(n20644), .A2(n20608), .B1(n20642), .B2(n20607), .ZN(
        n20609) );
  OAI211_X1 U23540 ( .C1(n20648), .C2(n20611), .A(n20610), .B(n20609), .ZN(
        P1_U3156) );
  INV_X1 U23541 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20619) );
  OAI22_X1 U23542 ( .A1(n20613), .A2(n20638), .B1(n20637), .B2(n20612), .ZN(
        n20614) );
  INV_X1 U23543 ( .A(n20614), .ZN(n20618) );
  AOI22_X1 U23544 ( .A1(n20644), .A2(n20616), .B1(n20642), .B2(n20615), .ZN(
        n20617) );
  OAI211_X1 U23545 ( .C1(n20648), .C2(n20619), .A(n20618), .B(n20617), .ZN(
        P1_U3157) );
  INV_X1 U23546 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20627) );
  OAI22_X1 U23547 ( .A1(n20621), .A2(n20638), .B1(n20637), .B2(n20620), .ZN(
        n20622) );
  INV_X1 U23548 ( .A(n20622), .ZN(n20626) );
  AOI22_X1 U23549 ( .A1(n20644), .A2(n20624), .B1(n20642), .B2(n20623), .ZN(
        n20625) );
  OAI211_X1 U23550 ( .C1(n20648), .C2(n20627), .A(n20626), .B(n20625), .ZN(
        P1_U3158) );
  INV_X1 U23551 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20635) );
  OAI22_X1 U23552 ( .A1(n20629), .A2(n20638), .B1(n20637), .B2(n20628), .ZN(
        n20630) );
  INV_X1 U23553 ( .A(n20630), .ZN(n20634) );
  AOI22_X1 U23554 ( .A1(n20644), .A2(n20632), .B1(n20642), .B2(n20631), .ZN(
        n20633) );
  OAI211_X1 U23555 ( .C1(n20648), .C2(n20635), .A(n20634), .B(n20633), .ZN(
        P1_U3159) );
  INV_X1 U23556 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20647) );
  OAI22_X1 U23557 ( .A1(n20639), .A2(n20638), .B1(n20637), .B2(n20636), .ZN(
        n20640) );
  INV_X1 U23558 ( .A(n20640), .ZN(n20646) );
  AOI22_X1 U23559 ( .A1(n20644), .A2(n20643), .B1(n20642), .B2(n20641), .ZN(
        n20645) );
  OAI211_X1 U23560 ( .C1(n20648), .C2(n20647), .A(n20646), .B(n20645), .ZN(
        P1_U3160) );
  NAND3_X1 U23561 ( .A1(n20650), .A2(n20649), .A3(n10231), .ZN(P1_U3163) );
  AND2_X1 U23562 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20651), .ZN(
        P1_U3164) );
  AND2_X1 U23563 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20651), .ZN(
        P1_U3165) );
  AND2_X1 U23564 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20651), .ZN(
        P1_U3166) );
  AND2_X1 U23565 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20651), .ZN(
        P1_U3167) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20651), .ZN(
        P1_U3168) );
  AND2_X1 U23567 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20651), .ZN(
        P1_U3169) );
  AND2_X1 U23568 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20651), .ZN(
        P1_U3170) );
  AND2_X1 U23569 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20651), .ZN(
        P1_U3171) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20651), .ZN(
        P1_U3172) );
  AND2_X1 U23571 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20651), .ZN(
        P1_U3173) );
  AND2_X1 U23572 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20651), .ZN(
        P1_U3174) );
  AND2_X1 U23573 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20651), .ZN(
        P1_U3175) );
  AND2_X1 U23574 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20651), .ZN(
        P1_U3176) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20651), .ZN(
        P1_U3177) );
  AND2_X1 U23576 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20651), .ZN(
        P1_U3178) );
  AND2_X1 U23577 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20651), .ZN(
        P1_U3179) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20651), .ZN(
        P1_U3180) );
  AND2_X1 U23579 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20651), .ZN(
        P1_U3181) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20651), .ZN(
        P1_U3182) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20651), .ZN(
        P1_U3183) );
  AND2_X1 U23582 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20651), .ZN(
        P1_U3184) );
  AND2_X1 U23583 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20651), .ZN(
        P1_U3185) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20651), .ZN(P1_U3186) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20651), .ZN(P1_U3187) );
  AND2_X1 U23586 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20651), .ZN(P1_U3188) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20651), .ZN(P1_U3189) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20651), .ZN(P1_U3190) );
  AND2_X1 U23589 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20651), .ZN(P1_U3191) );
  AND2_X1 U23590 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20651), .ZN(P1_U3192) );
  AND2_X1 U23591 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20651), .ZN(P1_U3193) );
  AOI211_X1 U23592 ( .C1(NA), .C2(n20659), .A(n20652), .B(n20769), .ZN(n20656)
         );
  NAND2_X1 U23593 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n20655) );
  AOI21_X1 U23594 ( .B1(n20662), .B2(n20751), .A(n20653), .ZN(n20654) );
  OAI221_X1 U23595 ( .B1(n20749), .B2(n20656), .C1(n20749), .C2(n20655), .A(
        n20654), .ZN(P1_U3194) );
  AOI21_X1 U23596 ( .B1(n20657), .B2(n20658), .A(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20666) );
  AOI22_X1 U23597 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20751), .B1(n20659), 
        .B2(n20658), .ZN(n20665) );
  AOI221_X1 U23598 ( .B1(NA), .B2(n20662), .C1(n20661), .C2(n20662), .A(n20660), .ZN(n20663) );
  OAI211_X1 U23599 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20769), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n20663), .ZN(n20664) );
  OAI211_X1 U23600 ( .C1(n20666), .C2(n20665), .A(n20704), .B(n20664), .ZN(
        P1_U3196) );
  INV_X1 U23601 ( .A(n20702), .ZN(n20708) );
  INV_X1 U23602 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20784) );
  OAI222_X1 U23603 ( .A1(n20708), .A2(n19854), .B1(n20784), .B2(n20749), .C1(
        n14390), .C2(n20704), .ZN(P1_U3197) );
  INV_X1 U23604 ( .A(n20667), .ZN(P1_U3198) );
  INV_X1 U23605 ( .A(n20668), .ZN(P1_U3199) );
  OAI222_X1 U23606 ( .A1(n20704), .A2(n20671), .B1(n20670), .B2(n20749), .C1(
        n20669), .C2(n20708), .ZN(P1_U3200) );
  AOI222_X1 U23607 ( .A1(n20702), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20706), .ZN(n20672) );
  INV_X1 U23608 ( .A(n20672), .ZN(P1_U3201) );
  AOI22_X1 U23609 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20702), .ZN(n20673) );
  OAI21_X1 U23610 ( .B1(n20674), .B2(n20704), .A(n20673), .ZN(P1_U3202) );
  AOI22_X1 U23611 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20706), .ZN(n20675) );
  OAI21_X1 U23612 ( .B1(n20677), .B2(n20708), .A(n20675), .ZN(P1_U3203) );
  AOI22_X1 U23613 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20702), .ZN(n20676) );
  OAI21_X1 U23614 ( .B1(n20677), .B2(n20704), .A(n20676), .ZN(P1_U3204) );
  AOI22_X1 U23615 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20706), .ZN(n20678) );
  OAI21_X1 U23616 ( .B1(n14229), .B2(n20708), .A(n20678), .ZN(P1_U3205) );
  AOI222_X1 U23617 ( .A1(n20702), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20706), .ZN(n20679) );
  INV_X1 U23618 ( .A(n20679), .ZN(P1_U3206) );
  INV_X1 U23619 ( .A(n20680), .ZN(P1_U3207) );
  INV_X1 U23620 ( .A(n20681), .ZN(P1_U3208) );
  AOI22_X1 U23621 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20702), .ZN(n20682) );
  OAI21_X1 U23622 ( .B1(n14643), .B2(n20704), .A(n20682), .ZN(P1_U3209) );
  AOI22_X1 U23623 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20706), .ZN(n20683) );
  OAI21_X1 U23624 ( .B1(n20684), .B2(n20708), .A(n20683), .ZN(P1_U3210) );
  INV_X1 U23625 ( .A(n20685), .ZN(P1_U3211) );
  INV_X1 U23626 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20772) );
  OAI222_X1 U23627 ( .A1(n20704), .A2(n15921), .B1(n20772), .B2(n20749), .C1(
        n20687), .C2(n20708), .ZN(P1_U3212) );
  AOI22_X1 U23628 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20702), .ZN(n20686) );
  OAI21_X1 U23629 ( .B1(n20687), .B2(n20704), .A(n20686), .ZN(P1_U3213) );
  AOI22_X1 U23630 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20706), .ZN(n20688) );
  OAI21_X1 U23631 ( .B1(n20689), .B2(n20708), .A(n20688), .ZN(P1_U3214) );
  AOI222_X1 U23632 ( .A1(n20702), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20706), .ZN(n20690) );
  INV_X1 U23633 ( .A(n20690), .ZN(P1_U3215) );
  AOI222_X1 U23634 ( .A1(n20706), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20770), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20702), .ZN(n20691) );
  INV_X1 U23635 ( .A(n20691), .ZN(P1_U3216) );
  AOI222_X1 U23636 ( .A1(n20702), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20706), .ZN(n20692) );
  INV_X1 U23637 ( .A(n20692), .ZN(P1_U3217) );
  AOI22_X1 U23638 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20702), .ZN(n20693) );
  OAI21_X1 U23639 ( .B1(n20694), .B2(n20704), .A(n20693), .ZN(P1_U3218) );
  AOI22_X1 U23640 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20770), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20706), .ZN(n20695) );
  OAI21_X1 U23641 ( .B1(n20696), .B2(n20708), .A(n20695), .ZN(P1_U3219) );
  AOI222_X1 U23642 ( .A1(n20706), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20702), .ZN(n20697) );
  INV_X1 U23643 ( .A(n20697), .ZN(P1_U3220) );
  AOI222_X1 U23644 ( .A1(n20706), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20702), .ZN(n20698) );
  INV_X1 U23645 ( .A(n20698), .ZN(P1_U3221) );
  AOI222_X1 U23646 ( .A1(n20706), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20702), .ZN(n20699) );
  INV_X1 U23647 ( .A(n20699), .ZN(P1_U3222) );
  AOI222_X1 U23648 ( .A1(n20706), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20702), .ZN(n20700) );
  INV_X1 U23649 ( .A(n20700), .ZN(P1_U3223) );
  AOI222_X1 U23650 ( .A1(n20706), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20702), .ZN(n20701) );
  INV_X1 U23651 ( .A(n20701), .ZN(P1_U3224) );
  AOI22_X1 U23652 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20702), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20747), .ZN(n20703) );
  OAI21_X1 U23653 ( .B1(n20705), .B2(n20704), .A(n20703), .ZN(P1_U3225) );
  AOI22_X1 U23654 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20706), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20747), .ZN(n20707) );
  OAI21_X1 U23655 ( .B1(n20709), .B2(n20708), .A(n20707), .ZN(P1_U3226) );
  OAI22_X1 U23656 ( .A1(n20770), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20749), .ZN(n20710) );
  INV_X1 U23657 ( .A(n20710), .ZN(P1_U3458) );
  OAI22_X1 U23658 ( .A1(n20747), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20749), .ZN(n20711) );
  INV_X1 U23659 ( .A(n20711), .ZN(P1_U3459) );
  OAI22_X1 U23660 ( .A1(n20747), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20749), .ZN(n20712) );
  INV_X1 U23661 ( .A(n20712), .ZN(P1_U3460) );
  OAI22_X1 U23662 ( .A1(n20747), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20749), .ZN(n20713) );
  INV_X1 U23663 ( .A(n20713), .ZN(P1_U3461) );
  OAI21_X1 U23664 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20717), .A(n20715), 
        .ZN(n20714) );
  INV_X1 U23665 ( .A(n20714), .ZN(P1_U3464) );
  OAI21_X1 U23666 ( .B1(n20717), .B2(n20716), .A(n20715), .ZN(P1_U3465) );
  AOI22_X1 U23667 ( .A1(n20721), .A2(n20720), .B1(n20719), .B2(n20718), .ZN(
        n20722) );
  INV_X1 U23668 ( .A(n20722), .ZN(n20724) );
  MUX2_X1 U23669 ( .A(n20724), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20723), .Z(P1_U3469) );
  NAND2_X1 U23670 ( .A1(n20726), .A2(n20725), .ZN(n20734) );
  AOI22_X1 U23671 ( .A1(n20730), .A2(n20729), .B1(n20728), .B2(n20727), .ZN(
        n20733) );
  NAND4_X1 U23672 ( .A1(n20734), .A2(n20733), .A3(n20732), .A4(n20731), .ZN(
        n20735) );
  NAND2_X1 U23673 ( .A1(n20738), .A2(n20735), .ZN(n20736) );
  OAI21_X1 U23674 ( .B1(n20738), .B2(n20737), .A(n20736), .ZN(P1_U3475) );
  AOI21_X1 U23675 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20739) );
  AOI22_X1 U23676 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20739), .B2(n14390), .ZN(n20741) );
  INV_X1 U23677 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20740) );
  AOI22_X1 U23678 ( .A1(n20742), .A2(n20741), .B1(n20740), .B2(n20745), .ZN(
        P1_U3481) );
  INV_X1 U23679 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20746) );
  INV_X1 U23680 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20744) );
  NOR2_X1 U23681 ( .A1(n20745), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20743) );
  AOI22_X1 U23682 ( .A1(n20746), .A2(n20745), .B1(n20744), .B2(n20743), .ZN(
        P1_U3482) );
  AOI22_X1 U23683 ( .A1(n20749), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20748), 
        .B2(n20747), .ZN(P1_U3483) );
  NOR2_X1 U23684 ( .A1(n20751), .A2(n20750), .ZN(n20760) );
  AOI211_X1 U23685 ( .C1(n20754), .C2(n20760), .A(n20753), .B(n20752), .ZN(
        n20768) );
  INV_X1 U23686 ( .A(n20755), .ZN(n20764) );
  OAI21_X1 U23687 ( .B1(n20758), .B2(n20757), .A(n20756), .ZN(n20761) );
  AOI21_X1 U23688 ( .B1(n20761), .B2(n20760), .A(n20759), .ZN(n20762) );
  AOI21_X1 U23689 ( .B1(n20764), .B2(n20763), .A(n20762), .ZN(n20767) );
  NOR2_X1 U23690 ( .A1(n20768), .A2(n20765), .ZN(n20766) );
  AOI22_X1 U23691 ( .A1(n20769), .A2(n20768), .B1(n20767), .B2(n20766), .ZN(
        P1_U3485) );
  MUX2_X1 U23692 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20770), .Z(P1_U3486) );
  AOI22_X1 U23693 ( .A1(n10842), .A2(keyinput103), .B1(keyinput107), .B2(
        n20772), .ZN(n20771) );
  OAI221_X1 U23694 ( .B1(n10842), .B2(keyinput103), .C1(n20772), .C2(
        keyinput107), .A(n20771), .ZN(n20782) );
  INV_X1 U23695 ( .A(DATAI_21_), .ZN(n20911) );
  AOI22_X1 U23696 ( .A1(n20911), .A2(keyinput116), .B1(keyinput88), .B2(n20774), .ZN(n20773) );
  OAI221_X1 U23697 ( .B1(n20911), .B2(keyinput116), .C1(n20774), .C2(
        keyinput88), .A(n20773), .ZN(n20781) );
  AOI22_X1 U23698 ( .A1(n20777), .A2(keyinput106), .B1(n20776), .B2(keyinput93), .ZN(n20775) );
  OAI221_X1 U23699 ( .B1(n20777), .B2(keyinput106), .C1(n20776), .C2(
        keyinput93), .A(n20775), .ZN(n20780) );
  AOI22_X1 U23700 ( .A1(n10490), .A2(keyinput125), .B1(keyinput117), .B2(
        n20913), .ZN(n20778) );
  OAI221_X1 U23701 ( .B1(n10490), .B2(keyinput125), .C1(n20913), .C2(
        keyinput117), .A(n20778), .ZN(n20779) );
  NOR4_X1 U23702 ( .A1(n20782), .A2(n20781), .A3(n20780), .A4(n20779), .ZN(
        n20819) );
  AOI22_X1 U23703 ( .A1(n20898), .A2(keyinput112), .B1(n20784), .B2(keyinput76), .ZN(n20783) );
  OAI221_X1 U23704 ( .B1(n20898), .B2(keyinput112), .C1(n20784), .C2(
        keyinput76), .A(n20783), .ZN(n20793) );
  AOI22_X1 U23705 ( .A1(n20786), .A2(keyinput109), .B1(n20910), .B2(keyinput73), .ZN(n20785) );
  OAI221_X1 U23706 ( .B1(n20786), .B2(keyinput109), .C1(n20910), .C2(
        keyinput73), .A(n20785), .ZN(n20792) );
  INV_X1 U23707 ( .A(P3_LWORD_REG_10__SCAN_IN), .ZN(n20788) );
  AOI22_X1 U23708 ( .A1(n20788), .A2(keyinput111), .B1(n20915), .B2(
        keyinput127), .ZN(n20787) );
  OAI221_X1 U23709 ( .B1(n20788), .B2(keyinput111), .C1(n20915), .C2(
        keyinput127), .A(n20787), .ZN(n20791) );
  AOI22_X1 U23710 ( .A1(n20945), .A2(keyinput120), .B1(keyinput87), .B2(n20895), .ZN(n20789) );
  OAI221_X1 U23711 ( .B1(n20945), .B2(keyinput120), .C1(n20895), .C2(
        keyinput87), .A(n20789), .ZN(n20790) );
  NOR4_X1 U23712 ( .A1(n20793), .A2(n20792), .A3(n20791), .A4(n20790), .ZN(
        n20818) );
  AOI22_X1 U23713 ( .A1(n20795), .A2(keyinput75), .B1(n20927), .B2(keyinput118), .ZN(n20794) );
  OAI221_X1 U23714 ( .B1(n20795), .B2(keyinput75), .C1(n20927), .C2(
        keyinput118), .A(n20794), .ZN(n20803) );
  AOI22_X1 U23715 ( .A1(n10755), .A2(keyinput79), .B1(n12103), .B2(keyinput69), 
        .ZN(n20796) );
  OAI221_X1 U23716 ( .B1(n10755), .B2(keyinput79), .C1(n12103), .C2(keyinput69), .A(n20796), .ZN(n20802) );
  INV_X1 U23717 ( .A(DATAI_6_), .ZN(n20948) );
  AOI22_X1 U23718 ( .A1(n20948), .A2(keyinput66), .B1(n20899), .B2(keyinput96), 
        .ZN(n20797) );
  OAI221_X1 U23719 ( .B1(n20948), .B2(keyinput66), .C1(n20899), .C2(keyinput96), .A(n20797), .ZN(n20801) );
  INV_X1 U23720 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n20799) );
  AOI22_X1 U23721 ( .A1(n20943), .A2(keyinput86), .B1(keyinput68), .B2(n20799), 
        .ZN(n20798) );
  OAI221_X1 U23722 ( .B1(n20943), .B2(keyinput86), .C1(n20799), .C2(keyinput68), .A(n20798), .ZN(n20800) );
  NOR4_X1 U23723 ( .A1(n20803), .A2(n20802), .A3(n20801), .A4(n20800), .ZN(
        n20817) );
  AOI22_X1 U23724 ( .A1(n20946), .A2(keyinput83), .B1(keyinput85), .B2(n13663), 
        .ZN(n20804) );
  OAI221_X1 U23725 ( .B1(n20946), .B2(keyinput83), .C1(n13663), .C2(keyinput85), .A(n20804), .ZN(n20815) );
  INV_X1 U23726 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n20806) );
  AOI22_X1 U23727 ( .A1(n20807), .A2(keyinput84), .B1(n20806), .B2(keyinput77), 
        .ZN(n20805) );
  OAI221_X1 U23728 ( .B1(n20807), .B2(keyinput84), .C1(n20806), .C2(keyinput77), .A(n20805), .ZN(n20814) );
  AOI22_X1 U23729 ( .A1(n20903), .A2(keyinput92), .B1(keyinput104), .B2(n20809), .ZN(n20808) );
  OAI221_X1 U23730 ( .B1(n20903), .B2(keyinput92), .C1(n20809), .C2(
        keyinput104), .A(n20808), .ZN(n20813) );
  AOI22_X1 U23731 ( .A1(n20949), .A2(keyinput114), .B1(n20811), .B2(
        keyinput123), .ZN(n20810) );
  OAI221_X1 U23732 ( .B1(n20949), .B2(keyinput114), .C1(n20811), .C2(
        keyinput123), .A(n20810), .ZN(n20812) );
  NOR4_X1 U23733 ( .A1(n20815), .A2(n20814), .A3(n20813), .A4(n20812), .ZN(
        n20816) );
  AND4_X1 U23734 ( .A1(n20819), .A2(n20818), .A3(n20817), .A4(n20816), .ZN(
        n20961) );
  OAI22_X1 U23735 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(keyinput119), 
        .B1(keyinput110), .B2(P3_REIP_REG_0__SCAN_IN), .ZN(n20820) );
  AOI221_X1 U23736 ( .B1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B2(keyinput119), 
        .C1(P3_REIP_REG_0__SCAN_IN), .C2(keyinput110), .A(n20820), .ZN(n20827)
         );
  OAI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(keyinput124), 
        .B1(BUF1_REG_2__SCAN_IN), .B2(keyinput102), .ZN(n20821) );
  AOI221_X1 U23738 ( .B1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B2(keyinput124), 
        .C1(keyinput102), .C2(BUF1_REG_2__SCAN_IN), .A(n20821), .ZN(n20826) );
  OAI22_X1 U23739 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(keyinput121), .B1(
        P3_READREQUEST_REG_SCAN_IN), .B2(keyinput65), .ZN(n20822) );
  AOI221_X1 U23740 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(keyinput121), .C1(
        keyinput65), .C2(P3_READREQUEST_REG_SCAN_IN), .A(n20822), .ZN(n20825)
         );
  OAI22_X1 U23741 ( .A1(BUF2_REG_30__SCAN_IN), .A2(keyinput80), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(keyinput94), .ZN(n20823) );
  AOI221_X1 U23742 ( .B1(BUF2_REG_30__SCAN_IN), .B2(keyinput80), .C1(
        keyinput94), .C2(P1_REIP_REG_5__SCAN_IN), .A(n20823), .ZN(n20824) );
  NAND4_X1 U23743 ( .A1(n20827), .A2(n20826), .A3(n20825), .A4(n20824), .ZN(
        n20857) );
  OAI22_X1 U23744 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput108), 
        .B1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput99), .ZN(n20828) );
  AOI221_X1 U23745 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput108), 
        .C1(keyinput99), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(n20828), 
        .ZN(n20835) );
  OAI22_X1 U23746 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(keyinput74), 
        .B1(keyinput78), .B2(P3_UWORD_REG_4__SCAN_IN), .ZN(n20829) );
  AOI221_X1 U23747 ( .B1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput74), 
        .C1(P3_UWORD_REG_4__SCAN_IN), .C2(keyinput78), .A(n20829), .ZN(n20834)
         );
  OAI22_X1 U23748 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(keyinput113), .B1(
        keyinput98), .B2(BUF2_REG_6__SCAN_IN), .ZN(n20830) );
  AOI221_X1 U23749 ( .B1(P2_EAX_REG_29__SCAN_IN), .B2(keyinput113), .C1(
        BUF2_REG_6__SCAN_IN), .C2(keyinput98), .A(n20830), .ZN(n20833) );
  OAI22_X1 U23750 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(keyinput89), .B1(
        BUF2_REG_16__SCAN_IN), .B2(keyinput70), .ZN(n20831) );
  AOI221_X1 U23751 ( .B1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B2(keyinput89), 
        .C1(keyinput70), .C2(BUF2_REG_16__SCAN_IN), .A(n20831), .ZN(n20832) );
  NAND4_X1 U23752 ( .A1(n20835), .A2(n20834), .A3(n20833), .A4(n20832), .ZN(
        n20856) );
  OAI22_X1 U23753 ( .A1(n20925), .A2(keyinput81), .B1(n20940), .B2(keyinput95), 
        .ZN(n20836) );
  AOI221_X1 U23754 ( .B1(n20925), .B2(keyinput81), .C1(keyinput95), .C2(n20940), .A(n20836), .ZN(n20844) );
  OAI22_X1 U23755 ( .A1(n20932), .A2(keyinput90), .B1(n13571), .B2(keyinput64), 
        .ZN(n20837) );
  AOI221_X1 U23756 ( .B1(n20932), .B2(keyinput90), .C1(keyinput64), .C2(n13571), .A(n20837), .ZN(n20843) );
  OAI22_X1 U23757 ( .A1(n12008), .A2(keyinput82), .B1(n20839), .B2(keyinput71), 
        .ZN(n20838) );
  AOI221_X1 U23758 ( .B1(n12008), .B2(keyinput82), .C1(keyinput71), .C2(n20839), .A(n20838), .ZN(n20842) );
  INV_X1 U23759 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n20904) );
  OAI22_X1 U23760 ( .A1(n20933), .A2(keyinput115), .B1(n20904), .B2(
        keyinput126), .ZN(n20840) );
  AOI221_X1 U23761 ( .B1(n20933), .B2(keyinput115), .C1(keyinput126), .C2(
        n20904), .A(n20840), .ZN(n20841) );
  NAND4_X1 U23762 ( .A1(n20844), .A2(n20843), .A3(n20842), .A4(n20841), .ZN(
        n20855) );
  OAI22_X1 U23763 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(keyinput67), 
        .B1(keyinput122), .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n20845) );
  AOI221_X1 U23764 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput67), 
        .C1(P2_UWORD_REG_8__SCAN_IN), .C2(keyinput122), .A(n20845), .ZN(n20853) );
  OAI22_X1 U23765 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(keyinput100), 
        .B1(keyinput91), .B2(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(n20846) );
  AOI221_X1 U23766 ( .B1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput100), 
        .C1(P2_DATAWIDTH_REG_28__SCAN_IN), .C2(keyinput91), .A(n20846), .ZN(
        n20852) );
  OAI22_X1 U23767 ( .A1(n20848), .A2(keyinput105), .B1(keyinput97), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20847) );
  AOI221_X1 U23768 ( .B1(n20848), .B2(keyinput105), .C1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .C2(keyinput97), .A(n20847), .ZN(
        n20851) );
  OAI22_X1 U23769 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput101), 
        .B1(BUF2_REG_18__SCAN_IN), .B2(keyinput72), .ZN(n20849) );
  AOI221_X1 U23770 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput101), 
        .C1(keyinput72), .C2(BUF2_REG_18__SCAN_IN), .A(n20849), .ZN(n20850) );
  NAND4_X1 U23771 ( .A1(n20853), .A2(n20852), .A3(n20851), .A4(n20850), .ZN(
        n20854) );
  NOR4_X1 U23772 ( .A1(n20857), .A2(n20856), .A3(n20855), .A4(n20854), .ZN(
        n20960) );
  AOI22_X1 U23773 ( .A1(P3_LWORD_REG_10__SCAN_IN), .A2(keyinput47), .B1(
        P1_INSTQUEUE_REG_3__1__SCAN_IN), .B2(keyinput60), .ZN(n20858) );
  OAI221_X1 U23774 ( .B1(P3_LWORD_REG_10__SCAN_IN), .B2(keyinput47), .C1(
        P1_INSTQUEUE_REG_3__1__SCAN_IN), .C2(keyinput60), .A(n20858), .ZN(
        n20865) );
  AOI22_X1 U23775 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(keyinput59), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(keyinput11), .ZN(n20859) );
  OAI221_X1 U23776 ( .B1(P1_EBX_REG_31__SCAN_IN), .B2(keyinput59), .C1(
        P1_EBX_REG_5__SCAN_IN), .C2(keyinput11), .A(n20859), .ZN(n20864) );
  AOI22_X1 U23777 ( .A1(P3_UWORD_REG_4__SCAN_IN), .A2(keyinput14), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(keyinput40), .ZN(n20860) );
  OAI221_X1 U23778 ( .B1(P3_UWORD_REG_4__SCAN_IN), .B2(keyinput14), .C1(
        P3_EBX_REG_21__SCAN_IN), .C2(keyinput40), .A(n20860), .ZN(n20863) );
  AOI22_X1 U23779 ( .A1(BUF2_REG_6__SCAN_IN), .A2(keyinput34), .B1(
        P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(keyinput18), .ZN(n20861) );
  OAI221_X1 U23780 ( .B1(BUF2_REG_6__SCAN_IN), .B2(keyinput34), .C1(
        P2_INSTQUEUE_REG_4__6__SCAN_IN), .C2(keyinput18), .A(n20861), .ZN(
        n20862) );
  NOR4_X1 U23781 ( .A1(n20865), .A2(n20864), .A3(n20863), .A4(n20862), .ZN(
        n20893) );
  AOI22_X1 U23782 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(keyinput45), .B1(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput37), .ZN(n20866) );
  OAI221_X1 U23783 ( .B1(P2_DATAO_REG_4__SCAN_IN), .B2(keyinput45), .C1(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput37), .A(n20866), .ZN(
        n20873) );
  AOI22_X1 U23784 ( .A1(BUF2_REG_18__SCAN_IN), .A2(keyinput8), .B1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput3), .ZN(n20867) );
  OAI221_X1 U23785 ( .B1(BUF2_REG_18__SCAN_IN), .B2(keyinput8), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(keyinput3), .A(n20867), .ZN(
        n20872) );
  AOI22_X1 U23786 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(keyinput12), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(keyinput49), .ZN(n20868) );
  OAI221_X1 U23787 ( .B1(P1_ADDRESS_REG_0__SCAN_IN), .B2(keyinput12), .C1(
        P2_EAX_REG_29__SCAN_IN), .C2(keyinput49), .A(n20868), .ZN(n20871) );
  AOI22_X1 U23788 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(keyinput20), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput44), .ZN(n20869) );
  OAI221_X1 U23789 ( .B1(P3_DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput20), .C1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(keyinput44), .A(n20869), .ZN(
        n20870) );
  NOR4_X1 U23790 ( .A1(n20873), .A2(n20872), .A3(n20871), .A4(n20870), .ZN(
        n20892) );
  AOI22_X1 U23791 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(keyinput27), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(keyinput46), .ZN(n20874) );
  OAI221_X1 U23792 ( .B1(P2_DATAWIDTH_REG_28__SCAN_IN), .B2(keyinput27), .C1(
        P3_REIP_REG_0__SCAN_IN), .C2(keyinput46), .A(n20874), .ZN(n20881) );
  AOI22_X1 U23793 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput24), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(keyinput39), .ZN(n20875) );
  OAI221_X1 U23794 ( .B1(P2_DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput24), .C1(
        P2_REIP_REG_22__SCAN_IN), .C2(keyinput39), .A(n20875), .ZN(n20880) );
  AOI22_X1 U23795 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(keyinput4), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(keyinput43), .ZN(n20876) );
  OAI221_X1 U23796 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(keyinput4), .C1(
        P1_ADDRESS_REG_15__SCAN_IN), .C2(keyinput43), .A(n20876), .ZN(n20879)
         );
  AOI22_X1 U23797 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput41), .B1(
        BUF2_REG_30__SCAN_IN), .B2(keyinput16), .ZN(n20877) );
  OAI221_X1 U23798 ( .B1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput41), 
        .C1(BUF2_REG_30__SCAN_IN), .C2(keyinput16), .A(n20877), .ZN(n20878) );
  NOR4_X1 U23799 ( .A1(n20881), .A2(n20880), .A3(n20879), .A4(n20878), .ZN(
        n20891) );
  AOI22_X1 U23800 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(keyinput42), .B1(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput13), .ZN(n20882) );
  OAI221_X1 U23801 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(keyinput42), .C1(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput13), .A(n20882), .ZN(
        n20889) );
  AOI22_X1 U23802 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(keyinput0), .B1(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput5), .ZN(n20883) );
  OAI221_X1 U23803 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(keyinput0), .C1(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(keyinput5), .A(n20883), .ZN(
        n20888) );
  AOI22_X1 U23804 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(keyinput30), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput7), .ZN(n20884) );
  OAI221_X1 U23805 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(keyinput30), .C1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(keyinput7), .A(n20884), .ZN(
        n20887) );
  AOI22_X1 U23806 ( .A1(BUF2_REG_16__SCAN_IN), .A2(keyinput6), .B1(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput29), .ZN(n20885) );
  OAI221_X1 U23807 ( .B1(BUF2_REG_16__SCAN_IN), .B2(keyinput6), .C1(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(keyinput29), .A(n20885), .ZN(
        n20886) );
  NOR4_X1 U23808 ( .A1(n20889), .A2(n20888), .A3(n20887), .A4(n20886), .ZN(
        n20890) );
  NAND4_X1 U23809 ( .A1(n20893), .A2(n20892), .A3(n20891), .A4(n20890), .ZN(
        n20959) );
  AOI22_X1 U23810 ( .A1(n20896), .A2(keyinput25), .B1(keyinput23), .B2(n20895), 
        .ZN(n20894) );
  OAI221_X1 U23811 ( .B1(n20896), .B2(keyinput25), .C1(n20895), .C2(keyinput23), .A(n20894), .ZN(n20908) );
  AOI22_X1 U23812 ( .A1(n20899), .A2(keyinput32), .B1(keyinput48), .B2(n20898), 
        .ZN(n20897) );
  OAI221_X1 U23813 ( .B1(n20899), .B2(keyinput32), .C1(n20898), .C2(keyinput48), .A(n20897), .ZN(n20907) );
  INV_X1 U23814 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20901) );
  AOI22_X1 U23815 ( .A1(n14229), .A2(keyinput57), .B1(keyinput35), .B2(n20901), 
        .ZN(n20900) );
  OAI221_X1 U23816 ( .B1(n14229), .B2(keyinput57), .C1(n20901), .C2(keyinput35), .A(n20900), .ZN(n20906) );
  AOI22_X1 U23817 ( .A1(n20904), .A2(keyinput62), .B1(n20903), .B2(keyinput28), 
        .ZN(n20902) );
  OAI221_X1 U23818 ( .B1(n20904), .B2(keyinput62), .C1(n20903), .C2(keyinput28), .A(n20902), .ZN(n20905) );
  NOR4_X1 U23819 ( .A1(n20908), .A2(n20907), .A3(n20906), .A4(n20905), .ZN(
        n20957) );
  AOI22_X1 U23820 ( .A1(n20911), .A2(keyinput52), .B1(n20910), .B2(keyinput9), 
        .ZN(n20909) );
  OAI221_X1 U23821 ( .B1(n20911), .B2(keyinput52), .C1(n20910), .C2(keyinput9), 
        .A(n20909), .ZN(n20922) );
  AOI22_X1 U23822 ( .A1(n10755), .A2(keyinput15), .B1(keyinput53), .B2(n20913), 
        .ZN(n20912) );
  OAI221_X1 U23823 ( .B1(n10755), .B2(keyinput15), .C1(n20913), .C2(keyinput53), .A(n20912), .ZN(n20921) );
  AOI22_X1 U23824 ( .A1(n20915), .A2(keyinput63), .B1(n13663), .B2(keyinput21), 
        .ZN(n20914) );
  OAI221_X1 U23825 ( .B1(n20915), .B2(keyinput63), .C1(n13663), .C2(keyinput21), .A(n20914), .ZN(n20920) );
  XOR2_X1 U23826 ( .A(n20916), .B(keyinput38), .Z(n20918) );
  XNOR2_X1 U23827 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B(keyinput33), .ZN(
        n20917) );
  NAND2_X1 U23828 ( .A1(n20918), .A2(n20917), .ZN(n20919) );
  NOR4_X1 U23829 ( .A1(n20922), .A2(n20921), .A3(n20920), .A4(n20919), .ZN(
        n20956) );
  AOI22_X1 U23830 ( .A1(n20925), .A2(keyinput17), .B1(keyinput1), .B2(n20924), 
        .ZN(n20923) );
  OAI221_X1 U23831 ( .B1(n20925), .B2(keyinput17), .C1(n20924), .C2(keyinput1), 
        .A(n20923), .ZN(n20937) );
  AOI22_X1 U23832 ( .A1(n20927), .A2(keyinput54), .B1(n10490), .B2(keyinput61), 
        .ZN(n20926) );
  OAI221_X1 U23833 ( .B1(n20927), .B2(keyinput54), .C1(n10490), .C2(keyinput61), .A(n20926), .ZN(n20936) );
  INV_X1 U23834 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20930) );
  AOI22_X1 U23835 ( .A1(n20930), .A2(keyinput55), .B1(keyinput36), .B2(n20929), 
        .ZN(n20928) );
  OAI221_X1 U23836 ( .B1(n20930), .B2(keyinput55), .C1(n20929), .C2(keyinput36), .A(n20928), .ZN(n20935) );
  AOI22_X1 U23837 ( .A1(n20933), .A2(keyinput51), .B1(n20932), .B2(keyinput26), 
        .ZN(n20931) );
  OAI221_X1 U23838 ( .B1(n20933), .B2(keyinput51), .C1(n20932), .C2(keyinput26), .A(n20931), .ZN(n20934) );
  NOR4_X1 U23839 ( .A1(n20937), .A2(n20936), .A3(n20935), .A4(n20934), .ZN(
        n20955) );
  INV_X1 U23840 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n20942) );
  AOI22_X1 U23841 ( .A1(n20943), .A2(keyinput22), .B1(keyinput58), .B2(n20942), 
        .ZN(n20941) );
  OAI221_X1 U23842 ( .B1(n20943), .B2(keyinput22), .C1(n20942), .C2(keyinput58), .A(n20941), .ZN(n20952) );
  AOI22_X1 U23843 ( .A1(n20946), .A2(keyinput19), .B1(keyinput56), .B2(n20945), 
        .ZN(n20944) );
  OAI221_X1 U23844 ( .B1(n20946), .B2(keyinput19), .C1(n20945), .C2(keyinput56), .A(n20944), .ZN(n20951) );
  AOI22_X1 U23845 ( .A1(n20949), .A2(keyinput50), .B1(n20948), .B2(keyinput2), 
        .ZN(n20947) );
  OAI221_X1 U23846 ( .B1(n20949), .B2(keyinput50), .C1(n20948), .C2(keyinput2), 
        .A(n20947), .ZN(n20950) );
  NOR4_X1 U23847 ( .A1(n20953), .A2(n20952), .A3(n20951), .A4(n20950), .ZN(
        n20954) );
  NAND4_X1 U23848 ( .A1(n20957), .A2(n20956), .A3(n20955), .A4(n20954), .ZN(
        n20958) );
  AOI211_X1 U23849 ( .C1(n20961), .C2(n20960), .A(n20959), .B(n20958), .ZN(
        n20965) );
  AOI22_X1 U23850 ( .A1(n20963), .A2(P3_ADDRESS_REG_10__SCAN_IN), .B1(
        P2_ADDRESS_REG_10__SCAN_IN), .B2(n20962), .ZN(n20964) );
  XNOR2_X1 U23851 ( .A(n20965), .B(n20964), .ZN(U375) );
  INV_X2 U11097 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18695) );
  BUF_X1 U11090 ( .A(n10646), .Z(n12413) );
  CLKBUF_X2 U11367 ( .A(n14087), .Z(n17044) );
  NOR2_X1 U12736 ( .A1(n11915), .A2(n15462), .ZN(n10004) );
  AOI222_X1 U11075 ( .A1(n20706), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20702), .ZN(n20685) );
  AOI222_X1 U11076 ( .A1(n20706), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20702), .ZN(n20681) );
  AOI222_X1 U11077 ( .A1(n20706), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20702), .ZN(n20680) );
  AOI222_X1 U11078 ( .A1(n20706), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20702), .ZN(n20668) );
  AOI222_X1 U11102 ( .A1(n20706), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20747), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20702), .ZN(n20667) );
  NOR2_X4 U11103 ( .A1(n11003), .A2(n20770), .ZN(n20706) );
  NOR2_X4 U11104 ( .A1(n20747), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20702) );
  CLKBUF_X1 U11136 ( .A(n10568), .Z(n13070) );
  CLKBUF_X1 U11148 ( .A(n10930), .Z(n11752) );
  CLKBUF_X3 U11149 ( .A(n10339), .Z(n9644) );
  AND4_X1 U11165 ( .A1(n10928), .A2(n10927), .A3(n10926), .A4(n10925), .ZN(
        n10243) );
  CLKBUF_X1 U11376 ( .A(n11884), .Z(n11897) );
  INV_X1 U11416 ( .A(n10615), .ZN(n10587) );
  CLKBUF_X1 U11507 ( .A(n12998), .Z(n14168) );
  CLKBUF_X1 U11866 ( .A(n14593), .Z(n14617) );
  CLKBUF_X1 U12435 ( .A(n14833), .Z(n9654) );
  CLKBUF_X1 U12478 ( .A(n16235), .Z(n18457) );
  XNOR2_X1 U12511 ( .A(n14104), .B(n14103), .ZN(n14666) );
  CLKBUF_X1 U13447 ( .A(n16941), .Z(n9643) );
  CLKBUF_X1 U15046 ( .A(n16387), .Z(n16395) );
endmodule

