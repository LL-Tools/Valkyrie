

module b17_C_AntiSAT_k_256_7 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9798, n9799, n9800, n9801, n9802, n9803,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136;

  NOR2_X1 U11227 ( .A1(n15083), .A2(n15069), .ZN(n14845) );
  NOR3_X1 U11228 ( .A1(n16289), .A2(n16298), .A3(n15647), .ZN(n15714) );
  AND2_X1 U11229 ( .A1(n16301), .A2(n16289), .ZN(n17366) );
  NAND2_X1 U11231 ( .A1(n9933), .A2(n9934), .ZN(n13527) );
  AND2_X1 U11232 ( .A1(n13702), .A2(n13701), .ZN(n13027) );
  AND3_X1 U11233 ( .A1(n9783), .A2(n13291), .A3(n10036), .ZN(n10218) );
  OR3_X1 U11234 ( .A1(n13251), .A2(n15400), .A3(n13252), .ZN(n19389) );
  OR2_X1 U11235 ( .A1(n13247), .A2(n13245), .ZN(n19212) );
  OR2_X1 U11236 ( .A1(n13244), .A2(n13245), .ZN(n19327) );
  CLKBUF_X2 U11237 ( .A(n13239), .Z(n13263) );
  INV_X2 U11238 ( .A(n13626), .ZN(n13621) );
  INV_X2 U11239 ( .A(n12150), .ZN(n13626) );
  AND2_X1 U11240 ( .A1(n10250), .A2(n10247), .ZN(n12489) );
  OR2_X1 U11241 ( .A1(n10506), .A2(n10505), .ZN(n10517) );
  NOR2_X2 U11242 ( .A1(n15532), .A2(n17219), .ZN(n15545) );
  NAND2_X1 U11243 ( .A1(n10554), .A2(n10553), .ZN(n11207) );
  CLKBUF_X2 U11244 ( .A(n10409), .Z(n10788) );
  INV_X1 U11245 ( .A(n10510), .ZN(n10524) );
  CLKBUF_X1 U11246 ( .A(n11566), .Z(n9790) );
  CLKBUF_X3 U11247 ( .A(n15492), .Z(n15546) );
  INV_X2 U11249 ( .A(n16842), .ZN(n17021) );
  AND2_X1 U11250 ( .A1(n9786), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13837) );
  MUX2_X1 U11252 ( .A(n12096), .B(n12103), .S(n12105), .Z(n11929) );
  INV_X1 U11253 ( .A(n15485), .ZN(n16929) );
  INV_X1 U11254 ( .A(n17018), .ZN(n16954) );
  INV_X2 U11255 ( .A(n11575), .ZN(n15486) );
  CLKBUF_X2 U11256 ( .A(n11950), .Z(n14030) );
  INV_X1 U11257 ( .A(n20729), .ZN(n11889) );
  INV_X1 U11258 ( .A(n11769), .ZN(n11907) );
  NAND2_X2 U11259 ( .A1(n11599), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11499) );
  INV_X2 U11260 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18665) );
  CLKBUF_X2 U11261 ( .A(n10408), .Z(n11076) );
  CLKBUF_X2 U11262 ( .A(n10493), .Z(n10458) );
  CLKBUF_X2 U11263 ( .A(n10913), .Z(n11077) );
  INV_X1 U11264 ( .A(n12325), .ZN(n20083) );
  NAND2_X2 U11265 ( .A1(n11742), .A2(n11741), .ZN(n13271) );
  CLKBUF_X2 U11266 ( .A(n10430), .Z(n12325) );
  CLKBUF_X2 U11267 ( .A(n10997), .Z(n10979) );
  AND2_X1 U11269 ( .A1(n10324), .A2(n12376), .ZN(n10349) );
  AND2_X1 U11270 ( .A1(n12383), .A2(n14516), .ZN(n10415) );
  AND2_X1 U11271 ( .A1(n10256), .A2(n10323), .ZN(n10416) );
  AND2_X1 U11272 ( .A1(n10324), .A2(n10323), .ZN(n10913) );
  AND2_X2 U11273 ( .A1(n11947), .A2(n11628), .ZN(n11946) );
  INV_X2 U11274 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10276) );
  CLKBUF_X2 U11275 ( .A(n10488), .Z(n10459) );
  CLKBUF_X2 U11276 ( .A(n10349), .Z(n9799) );
  AND4_X1 U11277 ( .A1(n11703), .A2(n11702), .A3(n11701), .A4(n11700), .ZN(
        n11704) );
  NOR2_X2 U11278 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12681) );
  NAND2_X1 U11279 ( .A1(n9953), .A2(n10430), .ZN(n10438) );
  AND2_X1 U11280 ( .A1(n14035), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U11281 ( .A1(n9926), .A2(n9925), .ZN(n15704) );
  INV_X2 U11283 ( .A(n9841), .ZN(n17036) );
  INV_X1 U11284 ( .A(n17038), .ZN(n16899) );
  OR2_X2 U11285 ( .A1(n10370), .A2(n10369), .ZN(n20074) );
  OAI21_X1 U11286 ( .B1(n15704), .B2(n11187), .A(n11189), .ZN(n14331) );
  NAND2_X1 U11287 ( .A1(n10567), .A2(n10566), .ZN(n12590) );
  AND2_X1 U11288 ( .A1(n13429), .A2(n13428), .ZN(n13449) );
  AND2_X1 U11289 ( .A1(n14601), .A2(n14602), .ZN(n14600) );
  NAND2_X1 U11290 ( .A1(n12082), .A2(n15433), .ZN(n12721) );
  OR2_X2 U11291 ( .A1(n14993), .A2(n14975), .ZN(n14973) );
  AND2_X1 U11292 ( .A1(n14992), .A2(n15203), .ZN(n15248) );
  NAND2_X1 U11293 ( .A1(n11707), .A2(n11918), .ZN(n15479) );
  INV_X1 U11294 ( .A(n12099), .ZN(n15443) );
  INV_X1 U11295 ( .A(n15604), .ZN(n18091) );
  AND2_X1 U11296 ( .A1(n20066), .A2(n20051), .ZN(n12795) );
  NAND2_X1 U11297 ( .A1(n12601), .A2(n12600), .ZN(n12599) );
  OR2_X1 U11298 ( .A1(n13472), .A2(n13471), .ZN(n14594) );
  INV_X1 U11299 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19616) );
  NOR2_X2 U11300 ( .A1(n14977), .A2(n14976), .ZN(n14978) );
  NAND2_X1 U11301 ( .A1(n13893), .A2(n13892), .ZN(n13901) );
  BUF_X1 U11302 ( .A(n12426), .Z(n15400) );
  NOR2_X1 U11303 ( .A1(n11531), .A2(n11530), .ZN(n18057) );
  NOR2_X1 U11304 ( .A1(n11573), .A2(n11572), .ZN(n18097) );
  NAND2_X1 U11305 ( .A1(n9970), .A2(n9848), .ZN(n17603) );
  INV_X1 U11306 ( .A(n15431), .ZN(n15429) );
  INV_X1 U11307 ( .A(n19838), .ZN(n19906) );
  OR2_X2 U11308 ( .A1(n15454), .A2(n13772), .ZN(n9783) );
  INV_X2 U11309 ( .A(n9800), .ZN(n18035) );
  OR2_X1 U11310 ( .A1(n11500), .A2(n11498), .ZN(n9841) );
  NAND2_X2 U11311 ( .A1(n17615), .A2(n15649), .ZN(n17519) );
  XNOR2_X2 U11312 ( .A(n11133), .B(n20010), .ZN(n19990) );
  AND2_X1 U11313 ( .A1(n11947), .A2(n11628), .ZN(n9784) );
  AND2_X1 U11314 ( .A1(n11947), .A2(n11628), .ZN(n9785) );
  NOR2_X2 U11315 ( .A1(n13065), .A2(n13064), .ZN(n13067) );
  NAND2_X2 U11316 ( .A1(n12634), .A2(n11127), .ZN(n11133) );
  NAND2_X2 U11317 ( .A1(n9999), .A2(n9954), .ZN(n13163) );
  NOR2_X2 U11318 ( .A1(n18921), .A2(n12962), .ZN(n18922) );
  AND2_X4 U11319 ( .A1(n12681), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9786) );
  OR2_X2 U11320 ( .A1(n14331), .A2(n11294), .ZN(n9916) );
  INV_X1 U11321 ( .A(n9801), .ZN(n9787) );
  INV_X2 U11322 ( .A(n9801), .ZN(n9788) );
  NOR2_X1 U11323 ( .A1(n16769), .A2(n11495), .ZN(n11492) );
  NOR2_X1 U11324 ( .A1(n11499), .A2(n11497), .ZN(n11566) );
  INV_X1 U11325 ( .A(n9841), .ZN(n9791) );
  NOR2_X1 U11326 ( .A1(n18708), .A2(n16402), .ZN(n9792) );
  INV_X1 U11327 ( .A(n17698), .ZN(n17713) );
  NAND2_X1 U11328 ( .A1(n15360), .A2(n15362), .ZN(n10230) );
  AND2_X1 U11329 ( .A1(n15715), .A2(n16279), .ZN(n16233) );
  INV_X1 U11330 ( .A(n13850), .ZN(n14793) );
  AND2_X1 U11331 ( .A1(n14600), .A2(n9905), .ZN(n14736) );
  NOR2_X2 U11332 ( .A1(n17409), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17408) );
  NAND2_X1 U11333 ( .A1(n17415), .A2(n10116), .ZN(n17409) );
  NAND2_X1 U11334 ( .A1(n17603), .A2(n17823), .ZN(n17514) );
  INV_X4 U11335 ( .A(n11179), .ZN(n11189) );
  AND2_X1 U11336 ( .A1(n15190), .A2(n15189), .ZN(n15192) );
  AND2_X1 U11337 ( .A1(n14667), .A2(n14666), .ZN(n14820) );
  NOR2_X1 U11338 ( .A1(n14201), .A2(n14142), .ZN(n13166) );
  NAND2_X1 U11339 ( .A1(n12583), .A2(n12582), .ZN(n12581) );
  NOR3_X1 U11340 ( .A1(n15272), .A2(n9872), .A3(n10192), .ZN(n14667) );
  NAND2_X1 U11341 ( .A1(n20323), .A2(n10081), .ZN(n10567) );
  NOR2_X1 U11342 ( .A1(n17329), .A2(n17199), .ZN(n17198) );
  OAI22_X2 U11343 ( .A1(n15743), .A2(n17278), .B1(n15742), .B2(n15741), .ZN(
        n17230) );
  OAI211_X1 U11344 ( .C1(n17648), .C2(n9951), .A(n9950), .B(n9860), .ZN(n9949)
         );
  AOI21_X2 U11345 ( .B1(n18508), .B2(n18514), .A(n18507), .ZN(n18516) );
  NAND2_X1 U11346 ( .A1(n10524), .A2(n10523), .ZN(n10532) );
  NOR2_X1 U11347 ( .A1(n17635), .A2(n10137), .ZN(n10136) );
  OAI21_X1 U11348 ( .B1(n17675), .B2(n10119), .A(n10118), .ZN(n17664) );
  CLKBUF_X2 U11349 ( .A(n17305), .Z(n9796) );
  INV_X2 U11350 ( .A(n18708), .ZN(n18062) );
  NOR2_X4 U11351 ( .A1(n11313), .A2(n11378), .ZN(n11396) );
  NAND2_X1 U11352 ( .A1(n13271), .A2(n15433), .ZN(n12948) );
  AND2_X1 U11353 ( .A1(n10434), .A2(n11286), .ZN(n10267) );
  INV_X1 U11355 ( .A(n20051), .ZN(n11286) );
  NAND2_X2 U11356 ( .A1(n20074), .A2(n10434), .ZN(n11349) );
  CLKBUF_X2 U11357 ( .A(n10415), .Z(n11078) );
  BUF_X2 U11358 ( .A(n10350), .Z(n10935) );
  CLKBUF_X2 U11359 ( .A(n12878), .Z(n17016) );
  BUF_X2 U11360 ( .A(n10494), .Z(n10930) );
  BUF_X4 U11362 ( .A(n11576), .Z(n9793) );
  INV_X1 U11363 ( .A(n11510), .ZN(n9801) );
  NAND2_X2 U11364 ( .A1(n11599), .A2(n18690), .ZN(n16769) );
  INV_X2 U11365 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11628) );
  INV_X2 U11367 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n10613) );
  AND2_X1 U11368 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U11369 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18526) );
  NAND2_X1 U11370 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13176) );
  OR2_X1 U11371 ( .A1(n11417), .A2(n15966), .ZN(n9847) );
  OAI211_X1 U11372 ( .C1(n14835), .C2(n14838), .A(n14836), .B(n14848), .ZN(
        n13513) );
  AOI21_X1 U11373 ( .B1(n14832), .B2(n19129), .A(n13648), .ZN(n13649) );
  NAND2_X1 U11374 ( .A1(n14986), .A2(n9877), .ZN(n14985) );
  NAND2_X1 U11375 ( .A1(n14294), .A2(n10257), .ZN(n9986) );
  AOI211_X1 U11376 ( .C1(n15061), .C2(n15060), .A(n15059), .B(n15058), .ZN(
        n15062) );
  NAND2_X1 U11377 ( .A1(n9968), .A2(n11189), .ZN(n14303) );
  AND2_X1 U11378 ( .A1(n9915), .A2(n10259), .ZN(n9914) );
  AOI21_X1 U11379 ( .B1(n10189), .B2(n19121), .A(n10188), .ZN(n10187) );
  NAND2_X1 U11380 ( .A1(n14331), .A2(n11188), .ZN(n15855) );
  AND2_X1 U11381 ( .A1(n9805), .A2(n9899), .ZN(n10309) );
  OAI21_X1 U11382 ( .B1(n15065), .B2(n16191), .A(n10239), .ZN(n15071) );
  XNOR2_X1 U11383 ( .A(n13897), .B(n13899), .ZN(n13893) );
  NAND2_X1 U11384 ( .A1(n14174), .A2(n10157), .ZN(n14233) );
  NAND2_X1 U11385 ( .A1(n9927), .A2(n11185), .ZN(n13165) );
  OAI211_X1 U11386 ( .C1(n14786), .C2(n9904), .A(n10291), .B(n9829), .ZN(
        n10290) );
  NAND2_X1 U11387 ( .A1(n14793), .A2(n10292), .ZN(n10291) );
  NAND2_X1 U11388 ( .A1(n9935), .A2(n13539), .ZN(n15371) );
  XNOR2_X1 U11389 ( .A(n13850), .B(n13867), .ZN(n14786) );
  AOI21_X1 U11390 ( .B1(n15067), .B2(n19126), .A(n10240), .ZN(n10239) );
  AND2_X1 U11391 ( .A1(n10271), .A2(n11134), .ZN(n9922) );
  NOR2_X1 U11392 ( .A1(n14343), .A2(n9956), .ZN(n10001) );
  OR2_X1 U11393 ( .A1(n17617), .A2(n17408), .ZN(n17398) );
  XNOR2_X1 U11394 ( .A(n13353), .B(n13323), .ZN(n13535) );
  NAND2_X1 U11395 ( .A1(n17744), .A2(n17487), .ZN(n17416) );
  NOR2_X1 U11396 ( .A1(n11174), .A2(n14375), .ZN(n14362) );
  NAND2_X1 U11397 ( .A1(n14360), .A2(n11172), .ZN(n14375) );
  NOR2_X1 U11398 ( .A1(n9839), .A2(n14074), .ZN(n14073) );
  AND2_X1 U11399 ( .A1(n10165), .A2(n10163), .ZN(n10162) );
  NAND2_X1 U11400 ( .A1(n10225), .A2(n13297), .ZN(n13329) );
  NAND2_X1 U11401 ( .A1(n11189), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14360) );
  AOI21_X1 U11402 ( .B1(n10227), .B2(n14018), .A(n10223), .ZN(n9934) );
  OR2_X2 U11403 ( .A1(n15258), .A2(n15257), .ZN(n15260) );
  AND2_X1 U11404 ( .A1(n13284), .A2(n13285), .ZN(n10036) );
  NAND2_X1 U11405 ( .A1(n10650), .A2(n10649), .ZN(n12600) );
  NOR2_X1 U11406 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17520), .ZN(
        n17538) );
  NAND2_X2 U11407 ( .A1(n14271), .A2(n11432), .ZN(n14268) );
  AND2_X1 U11408 ( .A1(n10155), .A2(n10156), .ZN(n10594) );
  INV_X2 U11409 ( .A(n19915), .ZN(n9794) );
  NOR2_X2 U11410 ( .A1(n20092), .A2(n9953), .ZN(n20610) );
  OR2_X1 U11411 ( .A1(n13244), .A2(n13255), .ZN(n19358) );
  NAND2_X1 U11412 ( .A1(n12555), .A2(n12554), .ZN(n15272) );
  INV_X1 U11413 ( .A(n11416), .ZN(n11408) );
  OR2_X1 U11414 ( .A1(n19489), .A2(n13773), .ZN(n13274) );
  NAND2_X1 U11415 ( .A1(n17616), .A2(n17617), .ZN(n17615) );
  OR2_X1 U11416 ( .A1(n13687), .A2(n13686), .ZN(n13689) );
  NAND2_X1 U11417 ( .A1(n13263), .A2(n10232), .ZN(n13311) );
  AOI221_X1 U11418 ( .B1(n9952), .B2(n17884), .C1(n17858), .C2(n17884), .A(
        n17537), .ZN(n17887) );
  NAND2_X1 U11419 ( .A1(n13263), .A2(n9940), .ZN(n19613) );
  NAND2_X1 U11420 ( .A1(n13263), .A2(n13257), .ZN(n19428) );
  OAI222_X1 U11421 ( .A1(n19759), .A2(n12430), .B1(n19756), .B2(n15410), .C1(
        n15409), .C2(n15414), .ZN(n15413) );
  AND2_X1 U11422 ( .A1(n12590), .A2(n10651), .ZN(n10155) );
  AND2_X1 U11423 ( .A1(n12243), .A2(n10195), .ZN(n12555) );
  AND2_X1 U11424 ( .A1(n9952), .A2(n15649), .ZN(n17616) );
  NAND2_X1 U11425 ( .A1(n12240), .A2(n12239), .ZN(n12243) );
  NOR2_X1 U11426 ( .A1(n16001), .A2(n16000), .ZN(n16003) );
  INV_X2 U11427 ( .A(n12320), .ZN(n9795) );
  NAND2_X1 U11428 ( .A1(n15646), .A2(n17948), .ZN(n15649) );
  INV_X1 U11429 ( .A(n12037), .ZN(n18958) );
  XNOR2_X1 U11430 ( .A(n12679), .B(n9846), .ZN(n13262) );
  NOR2_X1 U11431 ( .A1(n13424), .A2(n10076), .ZN(n13429) );
  INV_X1 U11432 ( .A(n18494), .ZN(n17914) );
  OR2_X2 U11433 ( .A1(n11245), .A2(n11244), .ZN(n15694) );
  NAND2_X2 U11434 ( .A1(n10534), .A2(n20100), .ZN(n12799) );
  NAND2_X1 U11435 ( .A1(n13406), .A2(n13407), .ZN(n13424) );
  NAND2_X1 U11436 ( .A1(n9842), .A2(n13485), .ZN(n13406) );
  NOR2_X1 U11438 ( .A1(n15431), .A2(n15430), .ZN(n19173) );
  XNOR2_X1 U11439 ( .A(n15583), .B(n9949), .ZN(n17625) );
  NAND2_X1 U11440 ( .A1(n11936), .A2(n11935), .ZN(n12433) );
  CLKBUF_X1 U11441 ( .A(n10634), .Z(n20289) );
  OR2_X1 U11442 ( .A1(n13395), .A2(n13502), .ZN(n13485) );
  NOR2_X2 U11443 ( .A1(n15590), .A2(n18517), .ZN(n18521) );
  NOR2_X2 U11444 ( .A1(n17664), .A2(n15544), .ZN(n17648) );
  NOR2_X1 U11445 ( .A1(n12757), .A2(n12756), .ZN(n16027) );
  AOI21_X1 U11446 ( .B1(n14692), .B2(n12193), .A(n12192), .ZN(n12196) );
  AOI21_X1 U11447 ( .B1(n9965), .B2(n10481), .A(n11162), .ZN(n9964) );
  NOR2_X2 U11448 ( .A1(n13325), .A2(n13324), .ZN(n13380) );
  NAND2_X1 U11449 ( .A1(n11929), .A2(n9855), .ZN(n10231) );
  XNOR2_X1 U11450 ( .A(n15530), .B(n17983), .ZN(n17675) );
  AND2_X1 U11451 ( .A1(n9966), .A2(n10632), .ZN(n9965) );
  NAND2_X2 U11452 ( .A1(n17280), .A2(n18552), .ZN(n17345) );
  XNOR2_X1 U11453 ( .A(n11314), .B(n12263), .ZN(n12814) );
  CLKBUF_X1 U11454 ( .A(n11931), .Z(n12652) );
  NOR2_X1 U11455 ( .A1(n15519), .A2(n15518), .ZN(n15530) );
  NAND3_X1 U11456 ( .A1(n10440), .A2(n10456), .A3(n10439), .ZN(n11289) );
  NAND2_X1 U11457 ( .A1(n11310), .A2(n11309), .ZN(n11314) );
  INV_X1 U11458 ( .A(n12342), .ZN(n10266) );
  INV_X1 U11459 ( .A(n11920), .ZN(n12082) );
  NAND2_X1 U11460 ( .A1(n9861), .A2(n11902), .ZN(n10287) );
  BUF_X2 U11461 ( .A(n12736), .Z(n9803) );
  AND2_X1 U11462 ( .A1(n12053), .A2(n10055), .ZN(n10233) );
  INV_X1 U11463 ( .A(n15620), .ZN(n17232) );
  AND2_X1 U11464 ( .A1(n10435), .A2(n11846), .ZN(n10448) );
  INV_X1 U11465 ( .A(n10267), .ZN(n10265) );
  NAND2_X1 U11466 ( .A1(n20079), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10554) );
  OR2_X1 U11467 ( .A1(n10438), .A2(n10437), .ZN(n15667) );
  AND3_X1 U11468 ( .A1(n10124), .A2(n15497), .A3(n15488), .ZN(n15620) );
  OR2_X2 U11469 ( .A1(n20066), .A2(n20051), .ZN(n11313) );
  BUF_X2 U11470 ( .A(n11349), .Z(n11378) );
  OR2_X1 U11471 ( .A1(n10480), .A2(n10479), .ZN(n11111) );
  NAND2_X1 U11472 ( .A1(n11686), .A2(n11685), .ZN(n12099) );
  NOR2_X2 U11473 ( .A1(n10431), .A2(n20074), .ZN(n12380) );
  INV_X2 U11474 ( .A(n10434), .ZN(n20066) );
  OR2_X1 U11475 ( .A1(n10470), .A2(n10469), .ZN(n11156) );
  NOR2_X2 U11476 ( .A1(n20045), .A2(n20044), .ZN(n20046) );
  AND4_X1 U11477 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10401) );
  AND4_X1 U11478 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10426) );
  AND4_X1 U11479 ( .A1(n10397), .A2(n10396), .A3(n10395), .A4(n10394), .ZN(
        n10398) );
  AND4_X1 U11480 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10427) );
  AND4_X1 U11481 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10428) );
  AND4_X1 U11482 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10400) );
  AND4_X1 U11483 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10399) );
  AND3_X1 U11484 ( .A1(n11689), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11687), .ZN(n10278) );
  AND2_X1 U11485 ( .A1(n11690), .A2(n11688), .ZN(n10277) );
  AND3_X1 U11486 ( .A1(n11693), .A2(n12694), .A3(n11692), .ZN(n10281) );
  AND3_X1 U11487 ( .A1(n10348), .A2(n10341), .A3(n10344), .ZN(n10262) );
  AND2_X1 U11488 ( .A1(n11694), .A2(n11691), .ZN(n10280) );
  INV_X4 U11489 ( .A(n9840), .ZN(n16971) );
  NAND2_X2 U11490 ( .A1(n18652), .A2(n18586), .ZN(n18639) );
  CLKBUF_X1 U11491 ( .A(n10912), .Z(n11022) );
  CLKBUF_X3 U11492 ( .A(n12889), .Z(n17019) );
  AND2_X2 U11493 ( .A1(n14030), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13838) );
  NAND2_X2 U11494 ( .A1(n20740), .A2(n19694), .ZN(n19743) );
  BUF_X2 U11495 ( .A(n10416), .Z(n10892) );
  INV_X2 U11496 ( .A(n16384), .ZN(U215) );
  NOR2_X4 U11497 ( .A1(n11500), .A2(n16769), .ZN(n12878) );
  NOR2_X2 U11498 ( .A1(n11499), .A2(n13176), .ZN(n17038) );
  BUF_X2 U11499 ( .A(n10559), .Z(n10464) );
  AND2_X2 U11500 ( .A1(n11627), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13768) );
  NOR2_X1 U11501 ( .A1(n18720), .A2(n18559), .ZN(n18706) );
  INV_X2 U11502 ( .A(n11633), .ZN(n11735) );
  BUF_X4 U11503 ( .A(n11085), .Z(n9811) );
  INV_X2 U11504 ( .A(n16387), .ZN(n16389) );
  INV_X2 U11505 ( .A(n15711), .ZN(n9800) );
  AND2_X2 U11506 ( .A1(n14515), .A2(n10323), .ZN(n10559) );
  NAND2_X1 U11507 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18690), .ZN(
        n11498) );
  INV_X1 U11508 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12391) );
  NOR2_X2 U11509 ( .A1(n14648), .A2(n14628), .ZN(n14614) );
  NAND2_X1 U11510 ( .A1(n10534), .A2(n10532), .ZN(n9918) );
  AND2_X1 U11511 ( .A1(n11904), .A2(n10003), .ZN(n9802) );
  AND2_X1 U11512 ( .A1(n11904), .A2(n10003), .ZN(n12424) );
  AND2_X1 U11513 ( .A1(n12038), .A2(n11963), .ZN(n11904) );
  AND4_X1 U11514 ( .A1(n13271), .A2(n12424), .A3(n10054), .A4(n9864), .ZN(
        n12736) );
  OAI222_X1 U11515 ( .A1(n9794), .A2(n14306), .B1(n14160), .B2(n19919), .C1(
        n14433), .C2(n19912), .ZN(P1_U2846) );
  AND4_X1 U11516 ( .A1(n10318), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10317), .A4(n10150), .ZN(n11085) );
  INV_X1 U11517 ( .A(n12940), .ZN(n12477) );
  OR2_X1 U11518 ( .A1(n15749), .A2(n15748), .ZN(n15751) );
  NAND2_X1 U11519 ( .A1(n15391), .A2(n13537), .ZN(n9936) );
  BUF_X1 U11520 ( .A(n12434), .Z(n13231) );
  NOR2_X2 U11521 ( .A1(n14594), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13479) );
  NAND4_X1 U11522 ( .A1(n11960), .A2(n11959), .A3(n11958), .A4(n11957), .ZN(
        n11961) );
  AND2_X2 U11523 ( .A1(n13689), .A2(n12432), .ZN(n13054) );
  INV_X1 U11524 ( .A(n14107), .ZN(n9808) );
  NAND2_X1 U11526 ( .A1(n13901), .A2(n13900), .ZN(n9805) );
  NOR2_X1 U11527 ( .A1(n14718), .A2(n10309), .ZN(n9806) );
  NOR2_X1 U11528 ( .A1(n14718), .A2(n10309), .ZN(n13952) );
  NAND2_X1 U11529 ( .A1(n9986), .A2(n9985), .ZN(n10268) );
  NAND2_X2 U11530 ( .A1(n11900), .A2(n12721), .ZN(n11937) );
  INV_X2 U11531 ( .A(n13239), .ZN(n13234) );
  XNOR2_X2 U11532 ( .A(n12489), .B(n12488), .ZN(n13239) );
  AOI211_X1 U11533 ( .C1(n17019), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16960), .B(n16959), .ZN(n16961) );
  AOI211_X1 U11534 ( .C1(n17019), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n12905), .B(n12904), .ZN(n12906) );
  NAND2_X2 U11535 ( .A1(n11901), .A2(n12948), .ZN(n11897) );
  NOR2_X2 U11536 ( .A1(n17625), .A2(n17962), .ZN(n17624) );
  OAI21_X4 U11537 ( .B1(n12799), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10516), 
        .ZN(n11109) );
  AOI211_X2 U11538 ( .C1(n15899), .C2(n14309), .A(n14308), .B(n14307), .ZN(
        n14310) );
  OAI21_X2 U11539 ( .B1(n14098), .B2(n14099), .A(n14084), .ZN(n14306) );
  OR2_X2 U11540 ( .A1(n14107), .A2(n10161), .ZN(n14084) );
  BUF_X1 U11541 ( .A(n10525), .Z(n9807) );
  AND2_X1 U11542 ( .A1(n13193), .A2(n10162), .ZN(n9809) );
  AND2_X1 U11543 ( .A1(n9808), .A2(n10162), .ZN(n14085) );
  AND2_X2 U11544 ( .A1(n14180), .A2(n10871), .ZN(n14174) );
  XNOR2_X2 U11545 ( .A(n14846), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15048) );
  OAI21_X2 U11546 ( .B1(n15020), .B2(n10207), .A(n10204), .ZN(n15349) );
  AND2_X4 U11547 ( .A1(n12381), .A2(n10256), .ZN(n10409) );
  XNOR2_X1 U11548 ( .A(n13927), .B(n9899), .ZN(n14720) );
  NOR2_X2 U11549 ( .A1(n11927), .A2(n11926), .ZN(n12023) );
  AND2_X1 U11550 ( .A1(n11947), .A2(n11948), .ZN(n13836) );
  AND2_X2 U11551 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11947) );
  AND2_X4 U11552 ( .A1(n12381), .A2(n14515), .ZN(n10494) );
  NOR2_X4 U11553 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14515) );
  AND2_X1 U11554 ( .A1(n12381), .A2(n14516), .ZN(n9812) );
  AND2_X1 U11555 ( .A1(n12381), .A2(n14516), .ZN(n9813) );
  NAND2_X2 U11556 ( .A1(n10262), .A2(n10261), .ZN(n11406) );
  AND2_X1 U11557 ( .A1(n14174), .A2(n14177), .ZN(n14175) );
  NAND2_X2 U11558 ( .A1(n18932), .A2(n12479), .ZN(n12518) );
  AOI21_X2 U11559 ( .B1(n12477), .B2(n12476), .A(n10311), .ZN(n18932) );
  AND3_X1 U11560 ( .A1(n10345), .A2(n10346), .A3(n10347), .ZN(n10260) );
  NOR2_X2 U11561 ( .A1(n13953), .A2(n13961), .ZN(n13955) );
  AND2_X1 U11562 ( .A1(n11627), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9814) );
  AND2_X2 U11563 ( .A1(n11627), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9815) );
  AND2_X4 U11564 ( .A1(n12383), .A2(n10324), .ZN(n10912) );
  OAI21_X2 U11565 ( .B1(n12641), .B2(n10770), .A(n10624), .ZN(n10625) );
  AND2_X2 U11566 ( .A1(n10625), .A2(n10641), .ZN(n10307) );
  XNOR2_X1 U11567 ( .A(n10642), .B(n12590), .ZN(n20048) );
  OAI21_X1 U11568 ( .B1(n12641), .B2(n11190), .A(n11104), .ZN(n12582) );
  OAI21_X1 U11569 ( .B1(n11109), .B2(n20066), .A(n11108), .ZN(n11115) );
  OAI222_X1 U11570 ( .A1(n9794), .A2(n14289), .B1(n13200), .B2(n19919), .C1(
        n14414), .C2(n19912), .ZN(P1_U2844) );
  NAND2_X2 U11571 ( .A1(n12580), .A2(n10641), .ZN(n12601) );
  AND2_X2 U11572 ( .A1(n13080), .A2(n13095), .ZN(n13093) );
  AND2_X2 U11573 ( .A1(n13093), .A2(n10151), .ZN(n14147) );
  NOR2_X2 U11574 ( .A1(n12779), .A2(n12934), .ZN(n12983) );
  NAND2_X2 U11575 ( .A1(n14121), .A2(n14123), .ZN(n14107) );
  NAND2_X1 U11576 ( .A1(n12082), .A2(n10285), .ZN(n10284) );
  NOR2_X1 U11577 ( .A1(n13271), .A2(n12075), .ZN(n10285) );
  AND4_X1 U11578 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11699) );
  NAND2_X1 U11579 ( .A1(n9919), .A2(n9856), .ZN(n9924) );
  NAND2_X1 U11580 ( .A1(n10272), .A2(n11151), .ZN(n9919) );
  INV_X1 U11581 ( .A(n11143), .ZN(n10272) );
  OR2_X1 U11582 ( .A1(n12212), .A2(n12211), .ZN(n13270) );
  INV_X1 U11583 ( .A(n10642), .ZN(n10156) );
  NAND2_X1 U11584 ( .A1(n10266), .A2(n10264), .ZN(n10263) );
  NAND2_X1 U11585 ( .A1(n10265), .A2(n9820), .ZN(n10264) );
  INV_X1 U11586 ( .A(n13270), .ZN(n12955) );
  AND2_X1 U11587 ( .A1(n14177), .A2(n14169), .ZN(n10159) );
  INV_X1 U11588 ( .A(n11096), .ZN(n11071) );
  INV_X1 U11589 ( .A(n10546), .ZN(n11120) );
  INV_X1 U11590 ( .A(n10632), .ZN(n9994) );
  AOI21_X1 U11591 ( .B1(n11719), .B2(n11718), .A(n11714), .ZN(n11723) );
  AND2_X1 U11592 ( .A1(n10197), .A2(n12366), .ZN(n10196) );
  INV_X1 U11593 ( .A(n13707), .ZN(n10237) );
  NOR2_X1 U11594 ( .A1(n13452), .A2(n13451), .ZN(n10063) );
  NOR2_X1 U11595 ( .A1(n11769), .A2(n11910), .ZN(n10054) );
  OR2_X1 U11596 ( .A1(n18813), .A2(n13543), .ZN(n13459) );
  NAND2_X1 U11597 ( .A1(n10038), .A2(n18895), .ZN(n13382) );
  NAND2_X1 U11598 ( .A1(n12678), .A2(n12677), .ZN(n10251) );
  NAND2_X1 U11599 ( .A1(n10249), .A2(n10248), .ZN(n10247) );
  INV_X1 U11600 ( .A(n12677), .ZN(n10248) );
  OR2_X1 U11601 ( .A1(n11499), .A2(n11495), .ZN(n15575) );
  OR2_X1 U11602 ( .A1(n16769), .A2(n11497), .ZN(n11575) );
  INV_X1 U11603 ( .A(n11492), .ZN(n16953) );
  NAND2_X1 U11604 ( .A1(n18665), .A2(n18675), .ZN(n11497) );
  OR2_X1 U11605 ( .A1(n18526), .A2(n11495), .ZN(n15485) );
  NOR2_X1 U11606 ( .A1(n15589), .A2(n16231), .ZN(n13186) );
  NAND2_X1 U11607 ( .A1(n17232), .A2(n15611), .ZN(n15532) );
  INV_X1 U11608 ( .A(n18498), .ZN(n16231) );
  OR2_X1 U11609 ( .A1(n20724), .A2(n12794), .ZN(n19857) );
  INV_X1 U11610 ( .A(n19811), .ZN(n11892) );
  AND2_X1 U11611 ( .A1(n10613), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11455) );
  NAND2_X1 U11612 ( .A1(n14382), .A2(n10001), .ZN(n9927) );
  NAND2_X1 U11613 ( .A1(n9923), .A2(n9920), .ZN(n11161) );
  OR2_X1 U11614 ( .A1(n9924), .A2(n10269), .ZN(n9923) );
  AOI21_X1 U11615 ( .B1(n9922), .B2(n19988), .A(n9921), .ZN(n9920) );
  NAND2_X1 U11616 ( .A1(n14294), .A2(n9960), .ZN(n9959) );
  NOR2_X1 U11617 ( .A1(n11189), .A2(n14401), .ZN(n9960) );
  NAND2_X1 U11618 ( .A1(n14303), .A2(n14295), .ZN(n14294) );
  INV_X1 U11619 ( .A(n9955), .ZN(n9954) );
  OAI21_X1 U11620 ( .B1(n10001), .B2(n10000), .A(n13164), .ZN(n9955) );
  NOR2_X1 U11621 ( .A1(n11212), .A2(n11199), .ZN(n11245) );
  NOR2_X1 U11622 ( .A1(n12663), .A2(n12048), .ZN(n12696) );
  NOR2_X1 U11623 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  INV_X1 U11624 ( .A(n13603), .ZN(n10299) );
  NOR2_X1 U11625 ( .A1(n14927), .A2(n10014), .ZN(n10013) );
  AND2_X1 U11626 ( .A1(n16130), .A2(n10015), .ZN(n10014) );
  INV_X1 U11627 ( .A(n14925), .ZN(n10015) );
  AOI21_X1 U11628 ( .B1(n10013), .B2(n10016), .A(n10012), .ZN(n10011) );
  INV_X1 U11629 ( .A(n16130), .ZN(n10016) );
  INV_X1 U11630 ( .A(n15243), .ZN(n10012) );
  AND2_X1 U11631 ( .A1(n12095), .A2(n12788), .ZN(n12123) );
  NAND2_X1 U11632 ( .A1(n12071), .A2(n11770), .ZN(n12701) );
  NAND2_X1 U11633 ( .A1(n11907), .A2(n12002), .ZN(n11770) );
  INV_X1 U11634 ( .A(n10610), .ZN(n10147) );
  NAND2_X1 U11635 ( .A1(n10093), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10092) );
  NAND2_X1 U11636 ( .A1(n11179), .A2(n14451), .ZN(n10093) );
  NOR2_X1 U11637 ( .A1(n10149), .A2(n10671), .ZN(n10148) );
  INV_X1 U11638 ( .A(n9892), .ZN(n10149) );
  NAND2_X1 U11639 ( .A1(n10580), .A2(n10579), .ZN(n10651) );
  NAND2_X1 U11640 ( .A1(n10438), .A2(n20074), .ZN(n10447) );
  NAND2_X1 U11641 ( .A1(n10430), .A2(n11423), .ZN(n9931) );
  NOR2_X1 U11642 ( .A1(n10521), .A2(n10081), .ZN(n10080) );
  NAND2_X1 U11643 ( .A1(n11196), .A2(n11195), .ZN(n11233) );
  OR2_X1 U11644 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20042), .ZN(
        n11232) );
  AND2_X1 U11645 ( .A1(n13384), .A2(n13379), .ZN(n10075) );
  AND2_X1 U11646 ( .A1(n10075), .A2(n10074), .ZN(n10073) );
  INV_X1 U11647 ( .A(n13048), .ZN(n10074) );
  NOR2_X1 U11648 ( .A1(n13266), .A2(n13265), .ZN(n10224) );
  NAND2_X1 U11649 ( .A1(n11589), .A2(n11593), .ZN(n9972) );
  NAND2_X1 U11650 ( .A1(n11596), .A2(n18075), .ZN(n9973) );
  INV_X1 U11651 ( .A(n11588), .ZN(n9971) );
  NOR2_X1 U11652 ( .A1(n11596), .A2(n13178), .ZN(n13177) );
  NOR4_X1 U11653 ( .A1(n11593), .A2(n13179), .A3(n11592), .A4(n18097), .ZN(
        n11595) );
  NOR2_X1 U11654 ( .A1(n15599), .A2(n11586), .ZN(n11594) );
  AND2_X1 U11655 ( .A1(n10164), .A2(n14099), .ZN(n10163) );
  INV_X1 U11656 ( .A(n14108), .ZN(n10164) );
  NOR2_X1 U11657 ( .A1(n11184), .A2(n14345), .ZN(n11185) );
  AND2_X1 U11658 ( .A1(n10771), .A2(n10154), .ZN(n10153) );
  OR2_X1 U11659 ( .A1(n13110), .A2(n13120), .ZN(n10154) );
  INV_X1 U11660 ( .A(n10770), .ZN(n10797) );
  NAND2_X1 U11661 ( .A1(n10185), .A2(n14082), .ZN(n10184) );
  AND2_X1 U11662 ( .A1(n9828), .A2(n9906), .ZN(n10177) );
  NAND2_X1 U11663 ( .A1(n9958), .A2(n9957), .ZN(n9956) );
  NOR2_X1 U11664 ( .A1(n10002), .A2(n11178), .ZN(n9957) );
  INV_X1 U11665 ( .A(n14352), .ZN(n9958) );
  NAND2_X1 U11666 ( .A1(n10672), .A2(n10671), .ZN(n11144) );
  OAI21_X1 U11667 ( .B1(n11135), .B2(n11190), .A(n11141), .ZN(n11142) );
  INV_X1 U11668 ( .A(n11313), .ZN(n11837) );
  OAI211_X1 U11669 ( .C1(n10487), .C2(n11286), .A(n10486), .B(n10485), .ZN(
        n10632) );
  NOR2_X1 U11670 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20050), .ZN(n20053) );
  NAND2_X1 U11671 ( .A1(n10436), .A2(n10448), .ZN(n9997) );
  OR2_X1 U11672 ( .A1(n11996), .A2(n11995), .ZN(n13296) );
  AND3_X1 U11673 ( .A1(n12959), .A2(n12958), .A3(n12957), .ZN(n12960) );
  NAND2_X1 U11674 ( .A1(n10069), .A2(n10068), .ZN(n13064) );
  NAND2_X1 U11675 ( .A1(n13502), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U11676 ( .A1(n12954), .A2(n11979), .ZN(n10069) );
  INV_X1 U11677 ( .A(n14552), .ZN(n12941) );
  INV_X1 U11678 ( .A(n14935), .ZN(n10062) );
  NAND2_X1 U11679 ( .A1(n10063), .A2(n9882), .ZN(n10057) );
  NAND2_X1 U11680 ( .A1(n10066), .A2(n13510), .ZN(n13453) );
  INV_X1 U11681 ( .A(n14644), .ZN(n10066) );
  CLKBUF_X1 U11682 ( .A(n13575), .Z(n13574) );
  NAND2_X1 U11683 ( .A1(n12629), .A2(n12775), .ZN(n10192) );
  INV_X1 U11684 ( .A(n12632), .ZN(n10193) );
  INV_X1 U11685 ( .A(n12512), .ZN(n10238) );
  NAND2_X1 U11686 ( .A1(n10230), .A2(n9851), .ZN(n15307) );
  AND2_X1 U11687 ( .A1(n15342), .A2(n10229), .ZN(n10228) );
  NAND2_X1 U11688 ( .A1(n10040), .A2(n9821), .ZN(n13542) );
  OR2_X1 U11689 ( .A1(n13542), .A2(n13543), .ZN(n13545) );
  INV_X1 U11690 ( .A(n13697), .ZN(n10254) );
  XNOR2_X1 U11691 ( .A(n12491), .B(n12490), .ZN(n12488) );
  OR2_X1 U11692 ( .A1(n13585), .A2(n19697), .ZN(n12446) );
  NAND2_X1 U11693 ( .A1(n10283), .A2(n10286), .ZN(n12047) );
  AND2_X1 U11694 ( .A1(n11897), .A2(n10316), .ZN(n12046) );
  NAND2_X1 U11695 ( .A1(n12054), .A2(n10055), .ZN(n12771) );
  AND2_X1 U11696 ( .A1(n12063), .A2(n12062), .ZN(n12189) );
  NAND2_X1 U11697 ( .A1(n10278), .A2(n10277), .ZN(n10282) );
  NAND2_X1 U11698 ( .A1(n10281), .A2(n10280), .ZN(n10279) );
  AND2_X1 U11699 ( .A1(n12001), .A2(n12948), .ZN(n11766) );
  INV_X1 U11700 ( .A(n15516), .ZN(n10131) );
  INV_X1 U11701 ( .A(n15511), .ZN(n10130) );
  NAND2_X1 U11702 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10134) );
  INV_X1 U11703 ( .A(n15512), .ZN(n10135) );
  AOI21_X1 U11704 ( .B1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n12878), .A(
        n10127), .ZN(n10126) );
  INV_X1 U11705 ( .A(n11496), .ZN(n17018) );
  NOR2_X1 U11706 ( .A1(n10107), .A2(n10111), .ZN(n10106) );
  INV_X1 U11707 ( .A(n10108), .ZN(n10107) );
  NOR2_X1 U11708 ( .A1(n10104), .A2(n10110), .ZN(n10103) );
  INV_X1 U11709 ( .A(n10106), .ZN(n10104) );
  NOR2_X1 U11710 ( .A1(n17473), .A2(n10096), .ZN(n10095) );
  INV_X1 U11711 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10096) );
  INV_X1 U11712 ( .A(n18075), .ZN(n11593) );
  NAND2_X1 U11713 ( .A1(n15545), .A2(n15613), .ZN(n15558) );
  XNOR2_X1 U11714 ( .A(n10128), .B(n15620), .ZN(n15517) );
  NOR2_X1 U11715 ( .A1(n18097), .A2(n18075), .ZN(n15591) );
  NOR2_X1 U11716 ( .A1(n18097), .A2(n15742), .ZN(n11597) );
  INV_X1 U11717 ( .A(n15694), .ZN(n11842) );
  AND2_X1 U11718 ( .A1(n19857), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12810) );
  AND2_X1 U11719 ( .A1(n16027), .A2(n16026), .ZN(n16029) );
  OAI21_X1 U11720 ( .B1(n14298), .B2(n12792), .A(n11034), .ZN(n14086) );
  NOR2_X1 U11721 ( .A1(n10160), .A2(n10158), .ZN(n10157) );
  INV_X1 U11722 ( .A(n9901), .ZN(n10160) );
  INV_X1 U11723 ( .A(n10159), .ZN(n10158) );
  INV_X1 U11724 ( .A(n14150), .ZN(n10805) );
  NAND2_X1 U11725 ( .A1(n13081), .A2(n10144), .ZN(n10143) );
  INV_X1 U11726 ( .A(n13074), .ZN(n10144) );
  AND2_X1 U11727 ( .A1(n14312), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10259) );
  INV_X1 U11728 ( .A(n14282), .ZN(n9969) );
  NAND2_X1 U11729 ( .A1(n13088), .A2(n11168), .ZN(n11170) );
  NAND2_X1 U11730 ( .A1(n16029), .A2(n12979), .ZN(n12989) );
  NOR2_X1 U11731 ( .A1(n10273), .A2(n10270), .ZN(n10269) );
  INV_X1 U11732 ( .A(n11151), .ZN(n10273) );
  INV_X1 U11733 ( .A(n15921), .ZN(n10270) );
  INV_X1 U11734 ( .A(n9924), .ZN(n10271) );
  NAND2_X1 U11735 ( .A1(n11142), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11143) );
  NAND2_X1 U11736 ( .A1(n19988), .A2(n11134), .ZN(n15922) );
  NAND2_X1 U11737 ( .A1(n15922), .A2(n15921), .ZN(n15920) );
  OAI211_X1 U11738 ( .C1(n9978), .C2(n12581), .A(n12635), .B(n9977), .ZN(
        n12634) );
  INV_X1 U11739 ( .A(n9978), .ZN(n9976) );
  OAI21_X1 U11740 ( .B1(n11114), .B2(n11190), .A(n11113), .ZN(n12258) );
  NOR2_X1 U11741 ( .A1(n9994), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9988) );
  AND2_X1 U11742 ( .A1(n9994), .A2(n10482), .ZN(n9992) );
  NAND2_X1 U11743 ( .A1(n9992), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U11744 ( .A1(n10481), .A2(n10632), .ZN(n9993) );
  NAND2_X1 U11745 ( .A1(n9917), .A2(n9881), .ZN(n10549) );
  NAND2_X1 U11746 ( .A1(n10552), .A2(n10551), .ZN(n20204) );
  NAND2_X1 U11747 ( .A1(n20047), .A2(n12589), .ZN(n20299) );
  INV_X1 U11749 ( .A(n20053), .ZN(n20210) );
  OR2_X1 U11750 ( .A1(n12002), .A2(n11724), .ZN(n12697) );
  NOR2_X1 U11751 ( .A1(n13445), .A2(n10072), .ZN(n10071) );
  INV_X1 U11752 ( .A(n13412), .ZN(n10077) );
  INV_X1 U11753 ( .A(n13423), .ZN(n10078) );
  NAND2_X1 U11754 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n14551), .ZN(
        n14552) );
  AND2_X1 U11755 ( .A1(n10196), .A2(n12541), .ZN(n10195) );
  OR2_X1 U11756 ( .A1(n14542), .A2(n14539), .ZN(n14541) );
  AND2_X1 U11757 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12942), .ZN(
        n14558) );
  INV_X1 U11758 ( .A(n14556), .ZN(n12942) );
  XNOR2_X1 U11759 ( .A(n13545), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15347) );
  NAND2_X1 U11760 ( .A1(n10043), .A2(n10042), .ZN(n14856) );
  NAND2_X1 U11761 ( .A1(n10049), .A2(n10051), .ZN(n10042) );
  NOR2_X1 U11762 ( .A1(n14855), .A2(n10045), .ZN(n10044) );
  NAND2_X1 U11763 ( .A1(n10053), .A2(n10052), .ZN(n14886) );
  NAND2_X1 U11764 ( .A1(n14895), .A2(n15118), .ZN(n10052) );
  NAND2_X1 U11765 ( .A1(n10048), .A2(n14893), .ZN(n10053) );
  OR2_X1 U11766 ( .A1(n14895), .A2(n15118), .ZN(n10048) );
  AND2_X1 U11767 ( .A1(n9875), .A2(n10246), .ZN(n10245) );
  INV_X1 U11768 ( .A(n14645), .ZN(n10246) );
  AOI21_X1 U11769 ( .B1(n10009), .B2(n10011), .A(n9885), .ZN(n10008) );
  AND2_X1 U11770 ( .A1(n16133), .A2(n16130), .ZN(n15242) );
  NAND2_X1 U11771 ( .A1(n15268), .A2(n14925), .ZN(n16133) );
  NOR3_X1 U11772 ( .A1(n15272), .A2(n10193), .A3(n15271), .ZN(n12776) );
  NAND2_X1 U11773 ( .A1(n10020), .A2(n15288), .ZN(n15270) );
  NAND2_X1 U11774 ( .A1(n10061), .A2(n10059), .ZN(n10020) );
  NAND2_X1 U11775 ( .A1(n15307), .A2(n13403), .ZN(n10061) );
  NAND2_X1 U11776 ( .A1(n15018), .A2(n13394), .ZN(n10209) );
  INV_X1 U11777 ( .A(n15347), .ZN(n10205) );
  OR2_X1 U11778 ( .A1(n15018), .A2(n13394), .ZN(n10208) );
  AND2_X1 U11779 ( .A1(n10230), .A2(n9887), .ZN(n15344) );
  XNOR2_X1 U11780 ( .A(n12430), .B(n12431), .ZN(n13686) );
  NAND2_X1 U11781 ( .A1(n11667), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11674) );
  NAND2_X1 U11782 ( .A1(n11672), .A2(n12694), .ZN(n11673) );
  NAND2_X1 U11783 ( .A1(n11679), .A2(n12694), .ZN(n11686) );
  NAND2_X1 U11784 ( .A1(n11684), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11685) );
  NAND2_X1 U11785 ( .A1(n13240), .A2(n13253), .ZN(n19462) );
  NOR2_X1 U11786 ( .A1(n13252), .A2(n14698), .ZN(n13253) );
  INV_X1 U11787 ( .A(n15428), .ZN(n19545) );
  INV_X1 U11788 ( .A(n19771), .ZN(n19762) );
  INV_X1 U11789 ( .A(n19361), .ZN(n19763) );
  AND2_X1 U11790 ( .A1(n12651), .A2(n12650), .ZN(n15411) );
  INV_X1 U11791 ( .A(n18085), .ZN(n17087) );
  INV_X1 U11792 ( .A(n11567), .ZN(n17015) );
  OAI21_X1 U11793 ( .B1(n13186), .B2(n12833), .A(n18706), .ZN(n15741) );
  NOR2_X1 U11794 ( .A1(n17645), .A2(n10100), .ZN(n10099) );
  AOI22_X1 U11795 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U11796 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11509) );
  AOI211_X1 U11797 ( .C1(n17016), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n11506), .B(n11505), .ZN(n11507) );
  NOR2_X1 U11798 ( .A1(n17204), .A2(n16290), .ZN(n15582) );
  OR2_X1 U11799 ( .A1(n17617), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9948) );
  OAI21_X1 U11800 ( .B1(n16289), .B2(n16290), .A(n10115), .ZN(n10114) );
  NOR2_X1 U11801 ( .A1(n18499), .A2(n17204), .ZN(n10115) );
  INV_X1 U11802 ( .A(n17894), .ZN(n17915) );
  NOR2_X1 U11803 ( .A1(n17614), .A2(n17948), .ZN(n17613) );
  INV_X1 U11804 ( .A(n10139), .ZN(n10137) );
  NAND2_X1 U11805 ( .A1(n17649), .A2(n10142), .ZN(n10139) );
  NAND2_X1 U11806 ( .A1(n10123), .A2(n10120), .ZN(n10119) );
  NAND2_X1 U11807 ( .A1(n15531), .A2(n10123), .ZN(n10118) );
  INV_X1 U11808 ( .A(n17674), .ZN(n10120) );
  OR2_X1 U11809 ( .A1(n17675), .A2(n17674), .ZN(n10122) );
  AOI21_X1 U11810 ( .B1(n12831), .B2(n12830), .A(n15601), .ZN(n18498) );
  NAND2_X1 U11811 ( .A1(n17850), .A2(n15596), .ZN(n18499) );
  NOR2_X1 U11812 ( .A1(n18722), .A2(n15589), .ZN(n18506) );
  AND2_X1 U11813 ( .A1(n12798), .A2(n12797), .ZN(n19838) );
  XNOR2_X1 U11814 ( .A(n13216), .B(n13215), .ZN(n14393) );
  NAND2_X1 U11815 ( .A1(n14271), .A2(n11444), .ZN(n14262) );
  NAND2_X1 U11816 ( .A1(n11430), .A2(n11892), .ZN(n14235) );
  OR2_X1 U11817 ( .A1(n12341), .A2(n11429), .ZN(n11430) );
  INV_X1 U11818 ( .A(n14393), .ZN(n10170) );
  XNOR2_X1 U11819 ( .A(n10084), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14400) );
  NAND2_X1 U11820 ( .A1(n10086), .A2(n10085), .ZN(n10084) );
  NAND2_X1 U11821 ( .A1(n11451), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10085) );
  NAND2_X1 U11822 ( .A1(n10268), .A2(n10087), .ZN(n10086) );
  OR2_X1 U11823 ( .A1(n20299), .A2(n20298), .ZN(n20321) );
  INV_X1 U11824 ( .A(n18952), .ZN(n18920) );
  INV_X1 U11825 ( .A(n18957), .ZN(n18939) );
  NAND2_X1 U11826 ( .A1(n10301), .A2(n12735), .ZN(n10300) );
  INV_X1 U11827 ( .A(n18973), .ZN(n10301) );
  AND2_X1 U11828 ( .A1(n18978), .A2(n18977), .ZN(n12731) );
  OR2_X1 U11829 ( .A1(n13003), .A2(n13002), .ZN(n13603) );
  AND2_X2 U11830 ( .A1(n12425), .A2(n12788), .ZN(n19000) );
  AND2_X1 U11831 ( .A1(n16186), .A2(n12034), .ZN(n16178) );
  INV_X1 U11832 ( .A(n16094), .ZN(n10189) );
  XNOR2_X1 U11833 ( .A(n14046), .B(n13627), .ZN(n19001) );
  AND2_X1 U11834 ( .A1(n14877), .A2(n10210), .ZN(n13551) );
  NOR2_X1 U11835 ( .A1(n10212), .A2(n15055), .ZN(n10210) );
  NAND2_X1 U11836 ( .A1(n10213), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10212) );
  INV_X1 U11837 ( .A(n16212), .ZN(n19129) );
  AND2_X1 U11838 ( .A1(n12123), .A2(n12119), .ZN(n19126) );
  INV_X1 U11839 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19794) );
  NOR2_X2 U11840 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19771) );
  INV_X1 U11841 ( .A(n19302), .ZN(n19279) );
  AND2_X1 U11842 ( .A1(n19367), .A2(n19545), .ZN(n19353) );
  INV_X1 U11843 ( .A(n18734), .ZN(n12788) );
  NOR2_X2 U11844 ( .A1(n16288), .A2(n17712), .ZN(n17543) );
  NAND2_X1 U11845 ( .A1(n17701), .A2(n16288), .ZN(n17606) );
  INV_X1 U11846 ( .A(n17606), .ZN(n17618) );
  XNOR2_X1 U11847 ( .A(n9946), .B(n16278), .ZN(n16261) );
  NAND2_X1 U11848 ( .A1(n9947), .A2(n16235), .ZN(n9946) );
  INV_X1 U11849 ( .A(n16233), .ZN(n9947) );
  NOR2_X2 U11850 ( .A1(n17204), .A2(n18037), .ZN(n17955) );
  NOR2_X1 U11851 ( .A1(n18022), .A2(n17914), .ZN(n18019) );
  NOR2_X1 U11852 ( .A1(n11214), .A2(n11262), .ZN(n11224) );
  NAND2_X1 U11853 ( .A1(n10226), .A2(n10055), .ZN(n10222) );
  INV_X1 U11854 ( .A(n10227), .ZN(n10220) );
  NOR2_X1 U11855 ( .A1(n13250), .A2(n13249), .ZN(n10004) );
  INV_X1 U11856 ( .A(n13267), .ZN(n10221) );
  AOI21_X1 U11857 ( .B1(n12462), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11943), .ZN(n12436) );
  NAND2_X1 U11858 ( .A1(n11942), .A2(n11941), .ZN(n11943) );
  AOI21_X1 U11859 ( .B1(n9803), .B2(P2_EBX_REG_1__SCAN_IN), .A(n10308), .ZN(
        n11941) );
  NAND2_X1 U11860 ( .A1(n9939), .A2(n9938), .ZN(n12073) );
  NAND2_X1 U11861 ( .A1(n11905), .A2(n11911), .ZN(n12078) );
  INV_X1 U11862 ( .A(n11171), .ZN(n10002) );
  OR2_X1 U11863 ( .A1(n10591), .A2(n10590), .ZN(n11146) );
  OR2_X1 U11864 ( .A1(n10500), .A2(n10499), .ZN(n11105) );
  NAND2_X1 U11865 ( .A1(n10482), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U11866 ( .A1(n9879), .A2(n20091), .ZN(n11280) );
  OR2_X1 U11867 ( .A1(n10565), .A2(n10564), .ZN(n11137) );
  NOR2_X1 U11868 ( .A1(n20051), .A2(n10081), .ZN(n10483) );
  NOR2_X1 U11869 ( .A1(n13424), .A2(n13423), .ZN(n13410) );
  AND2_X1 U11870 ( .A1(n10295), .A2(n13852), .ZN(n10292) );
  INV_X1 U11871 ( .A(n14785), .ZN(n10293) );
  OR2_X1 U11872 ( .A1(n12225), .A2(n12224), .ZN(n13046) );
  OR2_X1 U11873 ( .A1(n14893), .A2(n15118), .ZN(n10047) );
  AND2_X1 U11874 ( .A1(n10201), .A2(n14650), .ZN(n10200) );
  AOI21_X1 U11875 ( .B1(n10233), .B2(n12096), .A(n12943), .ZN(n11917) );
  INV_X1 U11876 ( .A(n11963), .ZN(n11898) );
  INV_X1 U11877 ( .A(n11653), .ZN(n11654) );
  INV_X1 U11878 ( .A(n15487), .ZN(n10127) );
  NOR2_X1 U11879 ( .A1(n11500), .A2(n18526), .ZN(n11493) );
  NAND2_X1 U11880 ( .A1(n18675), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11495) );
  NOR2_X1 U11881 ( .A1(n12828), .A2(n12827), .ZN(n11600) );
  NOR2_X1 U11882 ( .A1(n11233), .A2(n11232), .ZN(n11265) );
  NOR2_X1 U11883 ( .A1(n10765), .A2(n15827), .ZN(n10772) );
  INV_X1 U11884 ( .A(n15912), .ZN(n9921) );
  OAI211_X1 U11885 ( .C1(n10594), .C2(n10147), .A(n10146), .B(n10145), .ZN(
        n11152) );
  OR2_X1 U11886 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  AND2_X1 U11887 ( .A1(n10657), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10665) );
  NAND2_X1 U11888 ( .A1(n10664), .A2(n10672), .ZN(n11135) );
  OR2_X1 U11889 ( .A1(n10594), .A2(n9892), .ZN(n10664) );
  AND2_X1 U11890 ( .A1(n10643), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10657) );
  NOR2_X1 U11891 ( .A1(n10258), .A2(n14401), .ZN(n10257) );
  NAND2_X1 U11892 ( .A1(n11179), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10258) );
  NAND2_X1 U11893 ( .A1(n10091), .A2(n14281), .ZN(n9915) );
  NOR2_X1 U11894 ( .A1(n11389), .A2(n10186), .ZN(n10185) );
  NAND2_X1 U11895 ( .A1(n10088), .A2(n11179), .ZN(n14312) );
  AND2_X1 U11896 ( .A1(n10090), .A2(n13164), .ZN(n10089) );
  NOR2_X1 U11897 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n9925) );
  INV_X1 U11898 ( .A(n13165), .ZN(n9926) );
  INV_X1 U11899 ( .A(n11185), .ZN(n10000) );
  INV_X1 U11900 ( .A(n14184), .ZN(n10178) );
  NAND2_X1 U11901 ( .A1(n10181), .A2(n14207), .ZN(n10180) );
  INV_X1 U11902 ( .A(n13129), .ZN(n10181) );
  OR2_X1 U11903 ( .A1(n11179), .A2(n11181), .ZN(n14342) );
  INV_X1 U11904 ( .A(n11371), .ZN(n11397) );
  NAND2_X1 U11905 ( .A1(n10594), .A2(n10148), .ZN(n11164) );
  NOR2_X1 U11906 ( .A1(n20051), .A2(n20074), .ZN(n11371) );
  NAND2_X1 U11907 ( .A1(n12581), .A2(n11119), .ZN(n11126) );
  OR2_X1 U11908 ( .A1(n10578), .A2(n10577), .ZN(n11136) );
  NAND2_X1 U11909 ( .A1(n11837), .A2(n11378), .ZN(n11382) );
  NAND2_X1 U11910 ( .A1(n9983), .A2(n20019), .ZN(n9982) );
  AOI22_X1 U11911 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10344) );
  INV_X1 U11912 ( .A(n11433), .ZN(n10620) );
  AND2_X1 U11913 ( .A1(n11397), .A2(n11378), .ZN(n12262) );
  INV_X1 U11914 ( .A(n11105), .ZN(n10515) );
  OR2_X1 U11915 ( .A1(n10545), .A2(n10544), .ZN(n10546) );
  INV_X1 U11916 ( .A(n11228), .ZN(n11237) );
  AOI21_X1 U11917 ( .B1(n9807), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10526), .ZN(n10533) );
  NAND2_X1 U11918 ( .A1(n10437), .A2(n11433), .ZN(n9928) );
  AOI21_X1 U11919 ( .B1(n10431), .B2(n10381), .A(n9930), .ZN(n9929) );
  NOR2_X1 U11920 ( .A1(n9931), .A2(n10431), .ZN(n9930) );
  AND2_X1 U11921 ( .A1(n9932), .A2(n20051), .ZN(n10402) );
  INV_X1 U11922 ( .A(n11406), .ZN(n10433) );
  AOI21_X1 U11923 ( .B1(n20730), .B2(n16039), .A(n12571), .ZN(n20050) );
  INV_X1 U11924 ( .A(n10509), .ZN(n10082) );
  AND2_X1 U11925 ( .A1(n11198), .A2(n11232), .ZN(n11267) );
  OR2_X1 U11926 ( .A1(n11233), .A2(n11197), .ZN(n11198) );
  OR2_X1 U11927 ( .A1(n11228), .A2(n11190), .ZN(n11212) );
  NOR2_X1 U11928 ( .A1(n11910), .A2(n12099), .ZN(n11725) );
  NOR2_X1 U11929 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n13480), .ZN(n13484) );
  INV_X1 U11930 ( .A(n13410), .ZN(n13426) );
  AND2_X1 U11931 ( .A1(n13380), .A2(n9852), .ZN(n13396) );
  AND2_X1 U11932 ( .A1(n13502), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13048) );
  NAND2_X1 U11933 ( .A1(n13380), .A2(n10075), .ZN(n13395) );
  NAND2_X1 U11934 ( .A1(n13380), .A2(n10073), .ZN(n13389) );
  AND2_X1 U11935 ( .A1(n13380), .A2(n13379), .ZN(n13386) );
  NAND2_X1 U11936 ( .A1(n13901), .A2(n13900), .ZN(n13927) );
  NAND2_X1 U11937 ( .A1(n10290), .A2(n13899), .ZN(n13900) );
  AND2_X1 U11938 ( .A1(n14768), .A2(n14757), .ZN(n10194) );
  AND2_X1 U11939 ( .A1(n15192), .A2(n10199), .ZN(n14618) );
  AND2_X1 U11940 ( .A1(n10200), .A2(n14631), .ZN(n10199) );
  AND2_X1 U11941 ( .A1(n14618), .A2(n14619), .ZN(n14601) );
  AND2_X1 U11942 ( .A1(n10306), .A2(n10305), .ZN(n10304) );
  INV_X1 U11943 ( .A(n14724), .ZN(n10305) );
  AND2_X1 U11944 ( .A1(n14808), .A2(n15163), .ZN(n10201) );
  AND2_X1 U11945 ( .A1(n16103), .A2(n13756), .ZN(n10306) );
  NAND2_X1 U11946 ( .A1(n12734), .A2(n10297), .ZN(n14729) );
  AND2_X1 U11947 ( .A1(n10298), .A2(n10302), .ZN(n10297) );
  INV_X1 U11948 ( .A(n18970), .ZN(n10302) );
  NOR2_X1 U11949 ( .A1(n12295), .A2(n10198), .ZN(n10197) );
  INV_X1 U11950 ( .A(n12242), .ZN(n10198) );
  NOR2_X1 U11951 ( .A1(n14906), .A2(n10024), .ZN(n10023) );
  INV_X1 U11952 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10024) );
  NOR2_X1 U11953 ( .A1(n16138), .A2(n10028), .ZN(n10027) );
  NOR2_X1 U11954 ( .A1(n15026), .A2(n10031), .ZN(n10030) );
  INV_X1 U11955 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U11956 ( .A1(n13067), .A2(n12960), .ZN(n13341) );
  NAND2_X1 U11957 ( .A1(n14893), .A2(n15118), .ZN(n10050) );
  INV_X1 U11958 ( .A(n10047), .ZN(n10045) );
  OR2_X1 U11959 ( .A1(n10216), .A2(n15111), .ZN(n10215) );
  AND2_X1 U11960 ( .A1(n15192), .A2(n10200), .ZN(n14652) );
  NAND2_X1 U11961 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10216) );
  AND2_X1 U11962 ( .A1(n14820), .A2(n14818), .ZN(n15190) );
  INV_X1 U11963 ( .A(n10011), .ZN(n10010) );
  INV_X1 U11964 ( .A(n10013), .ZN(n10009) );
  NOR2_X1 U11965 ( .A1(n13402), .A2(n10060), .ZN(n10059) );
  INV_X1 U11966 ( .A(n15289), .ZN(n10060) );
  INV_X1 U11967 ( .A(n15023), .ZN(n10229) );
  INV_X1 U11968 ( .A(n13329), .ZN(n13526) );
  NAND2_X1 U11969 ( .A1(n12469), .A2(n12468), .ZN(n12490) );
  AOI21_X1 U11970 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12466), .ZN(n12491) );
  INV_X1 U11971 ( .A(n18936), .ZN(n10255) );
  NAND2_X1 U11972 ( .A1(n12467), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12440) );
  NAND2_X1 U11973 ( .A1(n12059), .A2(n12058), .ZN(n12063) );
  OR2_X1 U11974 ( .A1(n12055), .A2(n12771), .ZN(n12059) );
  NAND2_X1 U11975 ( .A1(n10003), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12060) );
  OR2_X1 U11976 ( .A1(n12215), .A2(n12214), .ZN(n12964) );
  NAND2_X1 U11977 ( .A1(n13234), .A2(n13691), .ZN(n13247) );
  NAND2_X1 U11978 ( .A1(n13234), .A2(n13262), .ZN(n13244) );
  AND2_X1 U11979 ( .A1(n13262), .A2(n13261), .ZN(n10232) );
  OR2_X1 U11980 ( .A1(n19772), .A2(n19783), .ZN(n15428) );
  INV_X1 U11981 ( .A(n12038), .ZN(n12042) );
  AND2_X1 U11982 ( .A1(n13259), .A2(n13262), .ZN(n9940) );
  INV_X1 U11983 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n20973) );
  NAND2_X1 U11984 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18665), .ZN(
        n11500) );
  NOR3_X1 U11985 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11599), .A3(
        n13176), .ZN(n11510) );
  NOR2_X1 U11986 ( .A1(n21011), .A2(n10109), .ZN(n10108) );
  AOI211_X1 U11987 ( .C1(n11592), .C2(n13181), .A(n11591), .B(n11590), .ZN(
        n15594) );
  OAI211_X1 U11988 ( .C1(n11597), .C2(n9973), .A(n9972), .B(n9971), .ZN(n11590) );
  INV_X1 U11989 ( .A(n17665), .ZN(n10123) );
  AOI22_X1 U11990 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18536), .B2(n11599), .ZN(
        n12828) );
  OR2_X1 U11991 ( .A1(n17281), .A2(n13177), .ZN(n11598) );
  AND2_X1 U11992 ( .A1(n18508), .A2(n13182), .ZN(n12832) );
  NAND3_X1 U11993 ( .A1(n11585), .A2(n11584), .A3(n11583), .ZN(n15599) );
  AOI211_X1 U11994 ( .C1(n9788), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n11582), .B(n11581), .ZN(n11583) );
  NOR3_X1 U11995 ( .A1(n13186), .A2(n13185), .A3(n15610), .ZN(n18539) );
  INV_X1 U11996 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15827) );
  INV_X1 U11997 ( .A(n12262), .ZN(n13214) );
  OR2_X1 U11998 ( .A1(n11016), .A2(n11015), .ZN(n11052) );
  INV_X1 U11999 ( .A(n14086), .ZN(n10165) );
  INV_X1 U12000 ( .A(n10163), .ZN(n10161) );
  AND2_X1 U12001 ( .A1(n10974), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10975) );
  NAND2_X1 U12002 ( .A1(n10975), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11013) );
  NOR2_X1 U12003 ( .A1(n10927), .A2(n10926), .ZN(n10928) );
  NOR2_X1 U12004 ( .A1(n10889), .A2(n15872), .ZN(n10890) );
  AND2_X1 U12005 ( .A1(n10888), .A2(n10887), .ZN(n14177) );
  AND2_X1 U12006 ( .A1(n10867), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10868) );
  NAND2_X1 U12007 ( .A1(n10868), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10889) );
  NOR2_X1 U12008 ( .A1(n21018), .A2(n10822), .ZN(n10867) );
  CLKBUF_X1 U12009 ( .A(n14134), .Z(n14191) );
  AND2_X1 U12010 ( .A1(n10806), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10821) );
  AND2_X1 U12011 ( .A1(n10787), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10806) );
  AND2_X1 U12012 ( .A1(n10772), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10787) );
  AND2_X1 U12013 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  INV_X1 U12014 ( .A(n14206), .ZN(n10152) );
  NAND2_X1 U12015 ( .A1(n10711), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10712) );
  NOR2_X1 U12016 ( .A1(n14389), .A2(n10712), .ZN(n10728) );
  NOR2_X1 U12017 ( .A1(n10697), .A2(n10696), .ZN(n10711) );
  AND4_X1 U12018 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(
        n13074) );
  NAND2_X1 U12019 ( .A1(n10673), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10697) );
  AND2_X1 U12020 ( .A1(n10665), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10673) );
  AOI21_X1 U12021 ( .B1(n11144), .B2(n10797), .A(n10680), .ZN(n12934) );
  AOI21_X1 U12022 ( .B1(n11128), .B2(n10797), .A(n10663), .ZN(n12726) );
  NOR2_X1 U12023 ( .A1(n11179), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10087) );
  INV_X1 U12024 ( .A(n9986), .ZN(n11451) );
  XNOR2_X1 U12025 ( .A(n10268), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11417) );
  NOR2_X1 U12026 ( .A1(n15751), .A2(n10183), .ZN(n14097) );
  INV_X1 U12027 ( .A(n10185), .ZN(n10183) );
  NOR2_X1 U12028 ( .A1(n15751), .A2(n11389), .ZN(n14112) );
  AND2_X1 U12029 ( .A1(n14312), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14321) );
  NAND2_X1 U12030 ( .A1(n13166), .A2(n9828), .ZN(n14187) );
  NAND2_X1 U12031 ( .A1(n13166), .A2(n11366), .ZN(n14185) );
  NAND2_X1 U12032 ( .A1(n14199), .A2(n14198), .ZN(n14201) );
  AND2_X1 U12033 ( .A1(n15882), .A2(n11177), .ZN(n14352) );
  OR2_X1 U12034 ( .A1(n15892), .A2(n14348), .ZN(n15880) );
  NOR2_X1 U12035 ( .A1(n13130), .A2(n10179), .ZN(n14199) );
  OR3_X1 U12036 ( .A1(n10180), .A2(n10182), .A3(n14151), .ZN(n10179) );
  NOR3_X1 U12037 ( .A1(n13130), .A2(n10182), .A3(n13129), .ZN(n14208) );
  NOR2_X1 U12038 ( .A1(n13130), .A2(n13129), .ZN(n13139) );
  OR2_X1 U12039 ( .A1(n13112), .A2(n13113), .ZN(n13130) );
  NAND2_X1 U12040 ( .A1(n16003), .A2(n13096), .ZN(n13112) );
  AND2_X1 U12041 ( .A1(n11169), .A2(n10313), .ZN(n10274) );
  NAND2_X1 U12042 ( .A1(n10166), .A2(n9910), .ZN(n16001) );
  INV_X1 U12043 ( .A(n12988), .ZN(n10167) );
  INV_X1 U12044 ( .A(n12989), .ZN(n10168) );
  AND2_X1 U12045 ( .A1(n10172), .A2(n11314), .ZN(n10171) );
  AND2_X1 U12046 ( .A1(n12577), .A2(n10173), .ZN(n10172) );
  INV_X1 U12047 ( .A(n12596), .ZN(n10173) );
  NAND2_X1 U12048 ( .A1(n10176), .A2(n10174), .ZN(n12597) );
  NOR2_X1 U12049 ( .A1(n11315), .A2(n10175), .ZN(n10174) );
  AND2_X1 U12050 ( .A1(n14506), .A2(n11290), .ZN(n20000) );
  AND2_X1 U12051 ( .A1(n15969), .A2(n14464), .ZN(n20001) );
  AND2_X1 U12052 ( .A1(n20001), .A2(n20024), .ZN(n13162) );
  NAND2_X1 U12053 ( .A1(n10266), .A2(n10267), .ZN(n11425) );
  NAND4_X1 U12054 ( .A1(n12795), .A2(n20083), .A3(n10620), .A4(n12380), .ZN(
        n11412) );
  NAND2_X1 U12055 ( .A1(n11278), .A2(n11892), .ZN(n11416) );
  AND3_X1 U12056 ( .A1(n12349), .A2(n12348), .A3(n12347), .ZN(n15672) );
  INV_X1 U12057 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20380) );
  OR2_X1 U12058 ( .A1(n20572), .A2(n20456), .ZN(n20458) );
  INV_X1 U12059 ( .A(n20374), .ZN(n20521) );
  NAND2_X1 U12060 ( .A1(n12590), .A2(n20047), .ZN(n20572) );
  AOI21_X1 U12061 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20489), .A(n20210), 
        .ZN(n20573) );
  INV_X1 U12062 ( .A(n9997), .ZN(n9995) );
  AND2_X1 U12063 ( .A1(n11717), .A2(n11716), .ZN(n12002) );
  OR2_X1 U12064 ( .A1(n13040), .A2(n12956), .ZN(n12001) );
  XNOR2_X1 U12065 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11999) );
  OAI21_X1 U12066 ( .B1(n13296), .B2(n12948), .A(n11998), .ZN(n12954) );
  NAND2_X1 U12067 ( .A1(n13506), .A2(n13486), .ZN(n13490) );
  NOR2_X1 U12068 ( .A1(n13490), .A2(n13491), .ZN(n13501) );
  NAND2_X1 U12069 ( .A1(n13396), .A2(n12743), .ZN(n13404) );
  NAND2_X1 U12070 ( .A1(n9862), .A2(n13067), .ZN(n13325) );
  INV_X1 U12071 ( .A(n13340), .ZN(n10067) );
  NAND2_X1 U12072 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12945) );
  AND2_X1 U12073 ( .A1(n12481), .A2(n12484), .ZN(n10288) );
  AND2_X1 U12074 ( .A1(n14600), .A2(n10194), .ZN(n14759) );
  AND2_X1 U12075 ( .A1(n14600), .A2(n14768), .ZN(n14767) );
  INV_X1 U12076 ( .A(n13857), .ZN(n10295) );
  NAND2_X1 U12077 ( .A1(n10294), .A2(n9822), .ZN(n10296) );
  INV_X1 U12078 ( .A(n14784), .ZN(n10294) );
  AND2_X1 U12079 ( .A1(n15192), .A2(n14808), .ZN(n15164) );
  NAND2_X1 U12080 ( .A1(n13754), .A2(n10306), .ZN(n16102) );
  CLKBUF_X1 U12081 ( .A(n14729), .Z(n18968) );
  NAND2_X1 U12082 ( .A1(n12243), .A2(n10196), .ZN(n15317) );
  AND2_X1 U12083 ( .A1(n12243), .A2(n10197), .ZN(n12365) );
  NAND2_X1 U12084 ( .A1(n12243), .A2(n12242), .ZN(n12294) );
  INV_X1 U12085 ( .A(n11485), .ZN(n15431) );
  XNOR2_X1 U12086 ( .A(n10035), .B(n14827), .ZN(n14825) );
  NAND2_X1 U12087 ( .A1(n14561), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10035) );
  AND2_X1 U12088 ( .A1(n14534), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14561) );
  AND2_X1 U12089 ( .A1(n14538), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14534) );
  NOR2_X1 U12090 ( .A1(n14541), .A2(n14868), .ZN(n14538) );
  AND2_X1 U12091 ( .A1(n9835), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10022) );
  NAND2_X1 U12092 ( .A1(n14558), .A2(n9835), .ZN(n14560) );
  NAND2_X1 U12093 ( .A1(n14558), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14557) );
  NAND2_X1 U12094 ( .A1(n12941), .A2(n9838), .ZN(n14556) );
  AND2_X1 U12095 ( .A1(n14978), .A2(n13757), .ZN(n14953) );
  AND2_X1 U12096 ( .A1(n12941), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14555) );
  NAND2_X1 U12097 ( .A1(n12941), .A2(n9834), .ZN(n14554) );
  AND2_X1 U12098 ( .A1(n14549), .A2(n10026), .ZN(n14551) );
  AND2_X1 U12099 ( .A1(n9836), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10026) );
  NAND2_X1 U12100 ( .A1(n14549), .A2(n9836), .ZN(n14550) );
  NAND2_X1 U12101 ( .A1(n14549), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14548) );
  NOR2_X1 U12102 ( .A1(n9817), .A2(n10236), .ZN(n10235) );
  INV_X1 U12103 ( .A(n15276), .ZN(n10236) );
  NOR2_X1 U12104 ( .A1(n16153), .A2(n14546), .ZN(n14549) );
  NOR2_X1 U12105 ( .A1(n13029), .A2(n9817), .ZN(n15275) );
  NAND2_X1 U12106 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n14547), .ZN(
        n14546) );
  AND2_X1 U12107 ( .A1(n13035), .A2(n10029), .ZN(n14547) );
  AND2_X1 U12108 ( .A1(n9827), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10029) );
  NAND2_X1 U12109 ( .A1(n13035), .A2(n9827), .ZN(n14544) );
  INV_X1 U12110 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15026) );
  NAND2_X1 U12111 ( .A1(n9845), .A2(n10253), .ZN(n10252) );
  INV_X1 U12112 ( .A(n12523), .ZN(n10253) );
  NAND2_X1 U12113 ( .A1(n13035), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13034) );
  NOR2_X1 U12114 ( .A1(n18906), .A2(n13032), .ZN(n13035) );
  NOR2_X1 U12115 ( .A1(n12945), .A2(n15036), .ZN(n13033) );
  NAND2_X1 U12116 ( .A1(n13033), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13032) );
  CLKBUF_X2 U12117 ( .A(n12197), .Z(n13624) );
  CLKBUF_X2 U12118 ( .A(n12181), .Z(n13625) );
  NOR2_X1 U12119 ( .A1(n15069), .A2(n15060), .ZN(n10213) );
  OR3_X1 U12120 ( .A1(n16045), .A2(n13543), .A3(n13643), .ZN(n14836) );
  NAND2_X1 U12121 ( .A1(n10211), .A2(n10213), .ZN(n14846) );
  INV_X1 U12122 ( .A(n15083), .ZN(n10211) );
  AND2_X1 U12123 ( .A1(n14600), .A2(n9898), .ZN(n14586) );
  OR2_X1 U12124 ( .A1(n10215), .A2(n13628), .ZN(n10214) );
  AOI21_X1 U12125 ( .B1(n14904), .B2(n14905), .A(n13475), .ZN(n14895) );
  OR2_X1 U12126 ( .A1(n14973), .A2(n10215), .ZN(n14918) );
  AOI21_X1 U12127 ( .B1(n15307), .B2(n10058), .A(n10056), .ZN(n14916) );
  AND2_X1 U12128 ( .A1(n10063), .A2(n13403), .ZN(n10058) );
  NAND2_X1 U12129 ( .A1(n10057), .A2(n9816), .ZN(n10056) );
  NAND2_X1 U12130 ( .A1(n13453), .A2(n15111), .ZN(n14933) );
  NAND2_X1 U12131 ( .A1(n14985), .A2(n10017), .ZN(n14947) );
  AND2_X1 U12132 ( .A1(n14959), .A2(n10018), .ZN(n10017) );
  OR2_X1 U12133 ( .A1(n19127), .A2(n15402), .ZN(n13645) );
  NOR2_X1 U12134 ( .A1(n14973), .A2(n15183), .ZN(n14964) );
  NOR2_X1 U12135 ( .A1(n10019), .A2(n14970), .ZN(n10018) );
  INV_X1 U12136 ( .A(n14930), .ZN(n10019) );
  NAND2_X1 U12137 ( .A1(n14985), .A2(n14930), .ZN(n14984) );
  INV_X1 U12138 ( .A(n15230), .ZN(n10191) );
  NOR3_X1 U12139 ( .A1(n15272), .A2(n10192), .A3(n10193), .ZN(n15231) );
  OR2_X1 U12140 ( .A1(n15328), .A2(n15293), .ZN(n15286) );
  NOR2_X1 U12141 ( .A1(n13029), .A2(n12512), .ZN(n15313) );
  NAND2_X1 U12142 ( .A1(n10234), .A2(n9844), .ZN(n15315) );
  NAND2_X1 U12143 ( .A1(n9936), .A2(n9937), .ZN(n9935) );
  NAND2_X1 U12144 ( .A1(n10255), .A2(n9845), .ZN(n13695) );
  NAND2_X1 U12145 ( .A1(n10255), .A2(n12499), .ZN(n18938) );
  AND2_X1 U12146 ( .A1(n13651), .A2(n13339), .ZN(n19107) );
  AND2_X1 U12147 ( .A1(n12046), .A2(n12047), .ZN(n12115) );
  OR2_X1 U12148 ( .A1(n12196), .A2(n12194), .ZN(n13060) );
  OR2_X1 U12149 ( .A1(n19772), .A2(n19780), .ZN(n19361) );
  NAND2_X1 U12150 ( .A1(n12039), .A2(n19616), .ZN(n12473) );
  NOR2_X1 U12151 ( .A1(n12027), .A2(n12026), .ZN(n12029) );
  INV_X1 U12152 ( .A(n11937), .ZN(n11938) );
  OR2_X1 U12153 ( .A1(n12430), .A2(n12431), .ZN(n12432) );
  AND3_X1 U12154 ( .A1(n12457), .A2(n12456), .A3(n12455), .ZN(n13056) );
  AND2_X1 U12155 ( .A1(n19772), .A2(n19780), .ZN(n19420) );
  CLKBUF_X1 U12156 ( .A(n12042), .Z(n12043) );
  AND2_X1 U12157 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12441), .ZN(
        n12470) );
  INV_X1 U12158 ( .A(n19173), .ZN(n19169) );
  INV_X1 U12159 ( .A(n19174), .ZN(n19171) );
  INV_X1 U12160 ( .A(n12483), .ZN(n10003) );
  NOR2_X1 U12161 ( .A1(n18521), .A2(n11598), .ZN(n18495) );
  NAND2_X1 U12162 ( .A1(n18723), .A2(n17239), .ZN(n11614) );
  INV_X1 U12163 ( .A(n11614), .ZN(n11617) );
  NOR2_X1 U12164 ( .A1(n10135), .A2(n10133), .ZN(n10132) );
  NOR3_X1 U12165 ( .A1(n15514), .A2(n10131), .A3(n10130), .ZN(n10129) );
  NOR2_X1 U12166 ( .A1(n15491), .A2(n10125), .ZN(n10124) );
  NAND2_X1 U12167 ( .A1(n18062), .A2(n18057), .ZN(n15742) );
  AOI21_X1 U12168 ( .B1(n17281), .B2(n18708), .A(n18521), .ZN(n15743) );
  NOR2_X1 U12169 ( .A1(n17277), .A2(n17238), .ZN(n17256) );
  INV_X1 U12170 ( .A(n17279), .ZN(n17281) );
  NAND2_X1 U12171 ( .A1(n10105), .A2(n10101), .ZN(n16764) );
  OR2_X1 U12172 ( .A1(n16271), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10105) );
  NOR2_X1 U12173 ( .A1(n10106), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10102) );
  NAND2_X1 U12174 ( .A1(n16271), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16242) );
  NAND2_X1 U12175 ( .A1(n17374), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17352) );
  AND2_X1 U12176 ( .A1(n17491), .A2(n9893), .ZN(n17419) );
  INV_X1 U12177 ( .A(n17438), .ZN(n10094) );
  NOR2_X1 U12178 ( .A1(n17514), .A2(n17779), .ZN(n17378) );
  NAND2_X1 U12179 ( .A1(n17491), .A2(n9830), .ZN(n17437) );
  NAND2_X1 U12180 ( .A1(n17491), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17471) );
  NOR2_X1 U12181 ( .A1(n17506), .A2(n17505), .ZN(n17491) );
  AND2_X1 U12182 ( .A1(n10098), .A2(n9831), .ZN(n17562) );
  NAND2_X1 U12183 ( .A1(n15714), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16235) );
  NAND2_X1 U12184 ( .A1(n10314), .A2(n15653), .ZN(n15654) );
  OR2_X1 U12185 ( .A1(n17399), .A2(n15647), .ZN(n10314) );
  OR2_X1 U12186 ( .A1(n17387), .A2(n17735), .ZN(n17723) );
  NAND2_X1 U12187 ( .A1(n10117), .A2(n9874), .ZN(n10116) );
  NOR2_X1 U12188 ( .A1(n17617), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17486) );
  NOR2_X1 U12189 ( .A1(n17501), .A2(n9945), .ZN(n17497) );
  OAI21_X1 U12190 ( .B1(n15651), .B2(n17848), .A(n9883), .ZN(n9945) );
  NAND2_X1 U12191 ( .A1(n17497), .A2(n17837), .ZN(n17496) );
  AOI21_X1 U12192 ( .B1(n17538), .B2(n17860), .A(n17617), .ZN(n17501) );
  INV_X1 U12193 ( .A(n15651), .ZN(n17502) );
  NOR2_X1 U12194 ( .A1(n15599), .A2(n11593), .ZN(n18508) );
  NAND2_X1 U12195 ( .A1(n15601), .A2(n15602), .ZN(n18496) );
  NAND2_X1 U12196 ( .A1(n18514), .A2(n15590), .ZN(n17876) );
  NOR2_X1 U12197 ( .A1(n11520), .A2(n11519), .ZN(n18075) );
  NOR2_X1 U12198 ( .A1(n11541), .A2(n11540), .ZN(n18080) );
  NOR2_X1 U12199 ( .A1(n11551), .A2(n11550), .ZN(n18085) );
  INV_X1 U12200 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18536) );
  INV_X1 U12201 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18360) );
  OAI21_X1 U12202 ( .B1(n17914), .B2(n16231), .A(n9858), .ZN(n18549) );
  INV_X1 U12203 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18504) );
  INV_X1 U12204 ( .A(n19897), .ZN(n15826) );
  INV_X1 U12205 ( .A(n19891), .ZN(n19878) );
  INV_X1 U12206 ( .A(n19847), .ZN(n19873) );
  AND2_X1 U12207 ( .A1(n12810), .A2(n12809), .ZN(n19901) );
  NAND2_X1 U12208 ( .A1(n11467), .A2(n11892), .ZN(n14188) );
  INV_X2 U12209 ( .A(n14188), .ZN(n19919) );
  INV_X1 U12210 ( .A(n14239), .ZN(n14264) );
  AND2_X1 U12211 ( .A1(n12728), .A2(n20043), .ZN(n14265) );
  AND2_X1 U12212 ( .A1(n12729), .A2(n14262), .ZN(n14273) );
  AND2_X1 U12213 ( .A1(n15694), .A2(n11892), .ZN(n11893) );
  INV_X2 U12214 ( .A(n19925), .ZN(n19950) );
  XNOR2_X1 U12215 ( .A(n11461), .B(n13219), .ZN(n12798) );
  AND2_X1 U12216 ( .A1(n15871), .A2(n11253), .ZN(n15899) );
  INV_X1 U12217 ( .A(n19993), .ZN(n20044) );
  OAI21_X1 U12218 ( .B1(n9984), .B2(n9961), .A(n9959), .ZN(n14275) );
  NAND2_X1 U12219 ( .A1(n14303), .A2(n14412), .ZN(n9984) );
  NAND2_X1 U12220 ( .A1(n14295), .A2(n11189), .ZN(n9961) );
  NAND2_X1 U12221 ( .A1(n11170), .A2(n11169), .ZN(n13103) );
  NAND2_X1 U12222 ( .A1(n10269), .A2(n15922), .ZN(n9962) );
  NAND2_X1 U12223 ( .A1(n15920), .A2(n11143), .ZN(n13017) );
  NOR3_X1 U12224 ( .A1(n20014), .A2(n11301), .A3(n13018), .ZN(n16014) );
  NAND2_X1 U12225 ( .A1(n9976), .A2(n9975), .ZN(n12636) );
  NAND2_X1 U12226 ( .A1(n9980), .A2(n12581), .ZN(n9975) );
  INV_X1 U12227 ( .A(n20001), .ZN(n20035) );
  INV_X1 U12228 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20489) );
  INV_X1 U12229 ( .A(n9992), .ZN(n9990) );
  OR2_X1 U12230 ( .A1(n10618), .A2(n10617), .ZN(n10619) );
  INV_X1 U12231 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20042) );
  INV_X1 U12232 ( .A(n20706), .ZN(n12571) );
  CLKBUF_X1 U12233 ( .A(n11420), .Z(n12565) );
  INV_X1 U12234 ( .A(n20157), .ZN(n20124) );
  OAI21_X1 U12235 ( .B1(n20228), .B2(n20212), .A(n20526), .ZN(n20231) );
  INV_X1 U12236 ( .A(n20288), .ZN(n20278) );
  OAI211_X1 U12237 ( .C1(n20343), .C2(n20704), .A(n20384), .B(n20328), .ZN(
        n20346) );
  INV_X1 U12238 ( .A(n20449), .ZN(n20452) );
  NOR2_X2 U12239 ( .A1(n20572), .A2(n20521), .ZN(n20621) );
  OR2_X1 U12240 ( .A1(n15691), .A2(n10081), .ZN(n19811) );
  INV_X1 U12241 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20627) );
  CLKBUF_X1 U12242 ( .A(n20667), .Z(n20739) );
  OR2_X1 U12243 ( .A1(n13444), .A2(n13467), .ZN(n14644) );
  NAND2_X1 U12244 ( .A1(n13449), .A2(n10071), .ZN(n13441) );
  NAND2_X1 U12245 ( .A1(n10034), .A2(n10033), .ZN(n18941) );
  NAND2_X1 U12246 ( .A1(n13646), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U12247 ( .A1(n14825), .A2(n12943), .ZN(n10034) );
  INV_X1 U12248 ( .A(n18941), .ZN(n18912) );
  INV_X1 U12249 ( .A(n18954), .ZN(n18907) );
  INV_X1 U12250 ( .A(n18961), .ZN(n18928) );
  CLKBUF_X1 U12251 ( .A(n12785), .Z(n18916) );
  OR2_X1 U12252 ( .A1(n12624), .A2(n12623), .ZN(n18977) );
  OR2_X1 U12253 ( .A1(n12551), .A2(n12550), .ZN(n18978) );
  INV_X1 U12254 ( .A(n14811), .ZN(n19005) );
  INV_X1 U12255 ( .A(n19791), .ZN(n19030) );
  INV_X1 U12256 ( .A(n19061), .ZN(n19038) );
  INV_X1 U12257 ( .A(n12096), .ZN(n12050) );
  AND2_X1 U12258 ( .A1(n11773), .A2(n11772), .ZN(n19089) );
  NAND2_X1 U12259 ( .A1(n14978), .A2(n9875), .ZN(n14646) );
  NAND2_X1 U12260 ( .A1(n10203), .A2(n10208), .ZN(n15348) );
  NAND2_X1 U12261 ( .A1(n15020), .A2(n10209), .ZN(n10203) );
  INV_X1 U12262 ( .A(n16178), .ZN(n19120) );
  INV_X1 U12263 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15036) );
  NAND2_X1 U12264 ( .A1(n18736), .A2(n12015), .ZN(n16186) );
  OR2_X1 U12265 ( .A1(n18736), .A2(n10055), .ZN(n16179) );
  OR2_X1 U12266 ( .A1(n18736), .A2(n14018), .ZN(n16181) );
  INV_X1 U12267 ( .A(n15400), .ZN(n14698) );
  INV_X1 U12268 ( .A(n16186), .ZN(n19104) );
  INV_X1 U12269 ( .A(n16181), .ZN(n19115) );
  XNOR2_X1 U12270 ( .A(n14847), .B(n14850), .ZN(n15051) );
  NAND2_X1 U12271 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  NOR2_X1 U12272 ( .A1(n15066), .A2(n10243), .ZN(n10242) );
  OR2_X1 U12273 ( .A1(n15070), .A2(n15069), .ZN(n10241) );
  INV_X1 U12274 ( .A(n15068), .ZN(n10243) );
  NAND2_X1 U12275 ( .A1(n10244), .A2(n9850), .ZN(n15065) );
  NAND2_X1 U12276 ( .A1(n10007), .A2(n10011), .ZN(n15007) );
  NAND2_X1 U12277 ( .A1(n15268), .A2(n10013), .ZN(n10007) );
  OR2_X1 U12278 ( .A1(n15242), .A2(n15241), .ZN(n15246) );
  NOR2_X1 U12279 ( .A1(n15272), .A2(n15271), .ZN(n12631) );
  INV_X1 U12280 ( .A(n19126), .ZN(n16209) );
  AND2_X1 U12281 ( .A1(n10061), .A2(n10064), .ZN(n15287) );
  INV_X1 U12282 ( .A(n10208), .ZN(n10207) );
  AOI21_X1 U12283 ( .B1(n10208), .B2(n10206), .A(n10205), .ZN(n10204) );
  INV_X1 U12284 ( .A(n10209), .ZN(n10206) );
  NAND2_X1 U12285 ( .A1(n10230), .A2(n13383), .ZN(n15022) );
  AND2_X1 U12286 ( .A1(n13534), .A2(n19112), .ZN(n15389) );
  INV_X1 U12287 ( .A(n16192), .ZN(n19130) );
  NAND2_X1 U12288 ( .A1(n15206), .A2(n13654), .ZN(n15402) );
  INV_X1 U12289 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19787) );
  INV_X1 U12290 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19777) );
  AND2_X1 U12291 ( .A1(n12701), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15416) );
  INV_X1 U12292 ( .A(n19780), .ZN(n19783) );
  AND4_X1 U12293 ( .A1(n19162), .A2(n19157), .A3(n12483), .A4(n12099), .ZN(
        n11707) );
  OAI21_X1 U12294 ( .B1(n19147), .B2(n19146), .A(n19145), .ZN(n19180) );
  OR2_X1 U12295 ( .A1(n19223), .A2(n19281), .ZN(n19241) );
  OAI21_X1 U12296 ( .B1(n19285), .B2(n19284), .A(n19283), .ZN(n19303) );
  OR2_X1 U12297 ( .A1(n19329), .A2(n19328), .ZN(n19354) );
  OAI21_X1 U12298 ( .B1(n19414), .B2(n19393), .A(n19624), .ZN(n19417) );
  INV_X1 U12299 ( .A(n19413), .ZN(n19415) );
  OAI21_X1 U12300 ( .B1(n19463), .B2(n19478), .A(n19624), .ZN(n19481) );
  OAI22_X1 U12301 ( .A1(n19156), .A2(n19171), .B1(n19155), .B2(n19169), .ZN(
        n19556) );
  AND2_X1 U12302 ( .A1(n19571), .A2(n19545), .ZN(n19567) );
  NAND2_X1 U12303 ( .A1(n19540), .A2(n19545), .ZN(n19596) );
  INV_X1 U12304 ( .A(n19667), .ZN(n19603) );
  OAI21_X1 U12305 ( .B1(n19584), .B2(n19583), .A(n19582), .ZN(n19609) );
  INV_X1 U12306 ( .A(n19137), .ZN(n19618) );
  INV_X1 U12307 ( .A(n19500), .ZN(n19638) );
  INV_X1 U12308 ( .A(n19507), .ZN(n19656) );
  INV_X1 U12309 ( .A(n19677), .ZN(n19663) );
  AND2_X1 U12310 ( .A1(n12470), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19669) );
  NAND2_X1 U12311 ( .A1(n19540), .A2(n19763), .ZN(n19677) );
  INV_X1 U12312 ( .A(n19666), .ZN(n19673) );
  OR2_X1 U12313 ( .A1(n12965), .A2(n19390), .ZN(n18734) );
  OR2_X1 U12314 ( .A1(n12723), .A2(n12722), .ZN(n12786) );
  OR2_X1 U12315 ( .A1(n15588), .A2(n15587), .ZN(n18722) );
  NOR2_X1 U12316 ( .A1(n18495), .A2(n17277), .ZN(n18723) );
  NAND2_X1 U12317 ( .A1(n18549), .A2(n18706), .ZN(n16402) );
  NOR2_X1 U12318 ( .A1(n16561), .A2(n16547), .ZN(n16540) );
  NOR2_X1 U12319 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16646), .ZN(n16626) );
  INV_X1 U12320 ( .A(n16768), .ZN(n16761) );
  NAND2_X1 U12321 ( .A1(n18551), .A2(n11617), .ZN(n16768) );
  INV_X1 U12322 ( .A(n16722), .ZN(n16767) );
  INV_X1 U12323 ( .A(n16745), .ZN(n16765) );
  INV_X1 U12324 ( .A(n16581), .ZN(n16777) );
  INV_X1 U12325 ( .A(n16773), .ZN(n16779) );
  INV_X2 U12326 ( .A(n17080), .ZN(n17075) );
  INV_X1 U12327 ( .A(n17093), .ZN(n17089) );
  NOR2_X1 U12328 ( .A1(n17307), .A2(n17102), .ZN(n17098) );
  NAND2_X1 U12329 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17107), .ZN(n17102) );
  INV_X1 U12330 ( .A(n17117), .ZN(n17112) );
  NAND2_X1 U12331 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17112), .ZN(n17111) );
  NOR2_X1 U12332 ( .A1(n17163), .A2(n17121), .ZN(n17118) );
  NOR2_X1 U12333 ( .A1(n20845), .A2(n17146), .ZN(n17140) );
  NOR3_X1 U12334 ( .A1(n17163), .A2(n17158), .A3(n17285), .ZN(n17150) );
  NOR2_X1 U12335 ( .A1(n20940), .A2(n17164), .ZN(n17159) );
  NAND4_X1 U12336 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n17198), .A4(n17170), .ZN(n17164) );
  INV_X1 U12337 ( .A(n18097), .ZN(n17163) );
  NOR2_X1 U12338 ( .A1(n15557), .A2(n15556), .ZN(n17211) );
  NOR2_X1 U12339 ( .A1(n15529), .A2(n15528), .ZN(n17219) );
  NAND2_X1 U12340 ( .A1(n17163), .A2(n17230), .ZN(n17225) );
  INV_X1 U12341 ( .A(n17234), .ZN(n17229) );
  INV_X1 U12342 ( .A(n17226), .ZN(n17233) );
  CLKBUF_X1 U12343 ( .A(n17266), .Z(n18703) );
  CLKBUF_X1 U12344 ( .A(n17268), .Z(n17274) );
  INV_X1 U12346 ( .A(n16764), .ZN(n16733) );
  NOR2_X1 U12347 ( .A1(n17352), .A2(n17353), .ZN(n16271) );
  NOR2_X1 U12348 ( .A1(n17392), .A2(n17393), .ZN(n17374) );
  NOR2_X1 U12349 ( .A1(n17709), .A2(n17634), .ZN(n17565) );
  INV_X1 U12350 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17533) );
  NAND2_X1 U12351 ( .A1(n17543), .A2(n17916), .ZN(n9970) );
  NAND2_X1 U12352 ( .A1(n17681), .A2(n17708), .ZN(n17634) );
  NAND2_X1 U12353 ( .A1(n10098), .A2(n10099), .ZN(n17531) );
  INV_X1 U12354 ( .A(n17543), .ZN(n17621) );
  NOR2_X1 U12355 ( .A1(n17637), .A2(n17645), .ZN(n17623) );
  INV_X1 U12356 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17645) );
  NAND2_X1 U12357 ( .A1(n17646), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17637) );
  NOR2_X1 U12358 ( .A1(n17666), .A2(n17668), .ZN(n17646) );
  INV_X1 U12359 ( .A(n18132), .ZN(n18442) );
  INV_X1 U12360 ( .A(n17712), .ZN(n17701) );
  NAND2_X1 U12361 ( .A1(n9974), .A2(n18708), .ZN(n17712) );
  INV_X1 U12362 ( .A(n16402), .ZN(n9974) );
  OAI21_X1 U12363 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18705), .A(n16402), 
        .ZN(n17708) );
  INV_X1 U12364 ( .A(n17850), .ZN(n15710) );
  INV_X1 U12365 ( .A(n10114), .ZN(n10113) );
  AND2_X1 U12366 ( .A1(n17930), .A2(n18516), .ZN(n17850) );
  INV_X1 U12367 ( .A(n18516), .ZN(n18529) );
  AOI21_X1 U12368 ( .B1(n17822), .B2(n17859), .A(n18022), .ZN(n17939) );
  INV_X1 U12369 ( .A(n17616), .ZN(n17959) );
  NAND2_X1 U12370 ( .A1(n10138), .A2(n10139), .ZN(n17636) );
  NAND2_X1 U12371 ( .A1(n17648), .A2(n10140), .ZN(n10138) );
  NAND2_X1 U12372 ( .A1(n17648), .A2(n17649), .ZN(n17647) );
  INV_X1 U12373 ( .A(n15531), .ZN(n10121) );
  INV_X1 U12374 ( .A(n10122), .ZN(n17673) );
  AND2_X1 U12375 ( .A1(n17850), .A2(n18062), .ZN(n18494) );
  INV_X1 U12376 ( .A(n18019), .ZN(n18039) );
  INV_X1 U12377 ( .A(n17876), .ZN(n18531) );
  INV_X1 U12378 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21014) );
  INV_X1 U12379 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18684) );
  CLKBUF_X1 U12380 ( .A(n18642), .Z(n18636) );
  AND2_X1 U12381 ( .A1(n11443), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20045)
         );
  OAI21_X1 U12383 ( .B1(n14400), .B2(n15966), .A(n9913), .ZN(P1_U3000) );
  AND2_X1 U12384 ( .A1(n9866), .A2(n10169), .ZN(n9913) );
  NAND2_X1 U12385 ( .A1(n10170), .A2(n20027), .ZN(n10169) );
  OR2_X1 U12386 ( .A1(n16067), .A2(n18920), .ZN(n10021) );
  NOR2_X1 U12387 ( .A1(n12732), .A2(n10300), .ZN(n13004) );
  NAND2_X1 U12388 ( .A1(n10190), .A2(n10187), .ZN(n13648) );
  NAND2_X1 U12389 ( .A1(n19001), .A2(n19126), .ZN(n10190) );
  NAND2_X1 U12390 ( .A1(n16262), .A2(n9941), .ZN(P3_U2800) );
  NAND2_X1 U12391 ( .A1(n9942), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9941) );
  NAND2_X1 U12392 ( .A1(n16263), .A2(n16265), .ZN(n9942) );
  NAND2_X1 U12393 ( .A1(n15718), .A2(n9943), .ZN(P3_U2832) );
  NAND2_X1 U12394 ( .A1(n9944), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9943) );
  NAND2_X1 U12395 ( .A1(n15719), .A2(n16276), .ZN(n9944) );
  OR2_X2 U12396 ( .A1(n16769), .A2(n13176), .ZN(n9840) );
  INV_X2 U12397 ( .A(n11979), .ZN(n13502) );
  AND2_X1 U12398 ( .A1(n14035), .A2(n12694), .ZN(n12152) );
  AND3_X1 U12399 ( .A1(n9823), .A2(n10062), .A3(n9895), .ZN(n9816) );
  INV_X4 U12400 ( .A(n13271), .ZN(n10055) );
  INV_X2 U12401 ( .A(n15647), .ZN(n17617) );
  OAI211_X1 U12402 ( .C1(n10634), .C2(n9990), .A(n9857), .B(n9987), .ZN(n11114) );
  NAND2_X1 U12403 ( .A1(n13093), .A2(n10153), .ZN(n13134) );
  NAND2_X1 U12404 ( .A1(n13093), .A2(n13110), .ZN(n13109) );
  NAND2_X1 U12405 ( .A1(n9844), .A2(n10237), .ZN(n9817) );
  OR3_X1 U12406 ( .A1(n15043), .A2(n15291), .A3(n13646), .ZN(n9818) );
  OR2_X1 U12407 ( .A1(n14858), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9819) );
  AND2_X2 U12408 ( .A1(n10324), .A2(n12381), .ZN(n10493) );
  OR2_X1 U12409 ( .A1(n20051), .A2(n11260), .ZN(n9820) );
  AND2_X1 U12410 ( .A1(n13323), .A2(n13538), .ZN(n9821) );
  NAND2_X1 U12411 ( .A1(n14793), .A2(n13852), .ZN(n9822) );
  AND4_X1 U12412 ( .A1(n13465), .A2(n14929), .A3(n14959), .A4(n14931), .ZN(
        n9823) );
  AND2_X1 U12413 ( .A1(n10004), .A2(n10226), .ZN(n9824) );
  AND2_X1 U12414 ( .A1(n11188), .A2(n9969), .ZN(n9825) );
  NAND2_X1 U12415 ( .A1(n10550), .A2(n10535), .ZN(n12324) );
  AND2_X1 U12416 ( .A1(n12518), .A2(n12481), .ZN(n9826) );
  AND2_X1 U12417 ( .A1(n10030), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9827) );
  AND2_X1 U12418 ( .A1(n11366), .A2(n10178), .ZN(n9828) );
  OR3_X1 U12419 ( .A1(n13867), .A2(n13866), .A3(n13865), .ZN(n9829) );
  AND2_X1 U12420 ( .A1(n10095), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9830) );
  AND2_X1 U12421 ( .A1(n10099), .A2(n9912), .ZN(n9831) );
  INV_X1 U12422 ( .A(n10303), .ZN(n14723) );
  NOR2_X1 U12423 ( .A1(n11179), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9832) );
  AND2_X1 U12424 ( .A1(n9832), .A2(n14412), .ZN(n9833) );
  AND2_X1 U12425 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9834) );
  AND2_X1 U12426 ( .A1(n10023), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9835) );
  AND2_X1 U12427 ( .A1(n10027), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9836) );
  AND2_X1 U12428 ( .A1(n9834), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9837) );
  NAND2_X1 U12429 ( .A1(n10168), .A2(n10167), .ZN(n13076) );
  INV_X1 U12430 ( .A(n13076), .ZN(n10166) );
  AND2_X1 U12431 ( .A1(n9837), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9838) );
  AND2_X1 U12432 ( .A1(n9786), .A2(n12694), .ZN(n11985) );
  OR3_X1 U12433 ( .A1(n15751), .A2(n10184), .A3(n13198), .ZN(n9839) );
  AND2_X2 U12434 ( .A1(n13768), .A2(n12694), .ZN(n12151) );
  OR2_X1 U12435 ( .A1(n13404), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n9842) );
  OR2_X1 U12436 ( .A1(n14973), .A2(n10216), .ZN(n14938) );
  NOR2_X1 U12437 ( .A1(n13449), .A2(n13430), .ZN(n9843) );
  AND2_X1 U12438 ( .A1(n10238), .A2(n15314), .ZN(n9844) );
  AND2_X1 U12439 ( .A1(n12499), .A2(n10254), .ZN(n9845) );
  INV_X1 U12440 ( .A(n15611), .ZN(n10128) );
  OR2_X2 U12441 ( .A1(n10380), .A2(n10379), .ZN(n10431) );
  INV_X1 U12442 ( .A(n10290), .ZN(n13897) );
  INV_X1 U12443 ( .A(n11846), .ZN(n20091) );
  OR2_X2 U12444 ( .A1(n10340), .A2(n10339), .ZN(n11846) );
  XOR2_X1 U12445 ( .A(n12677), .B(n12678), .Z(n9846) );
  INV_X1 U12446 ( .A(n11963), .ZN(n11979) );
  INV_X2 U12447 ( .A(n11910), .ZN(n19162) );
  INV_X1 U12448 ( .A(n17916), .ZN(n9952) );
  NAND2_X1 U12449 ( .A1(n14382), .A2(n11171), .ZN(n14341) );
  OR2_X1 U12450 ( .A1(n17713), .A2(n17529), .ZN(n9848) );
  NAND4_X2 U12451 ( .A1(n11907), .A2(n11727), .A3(n13271), .A4(n11919), .ZN(
        n13585) );
  NAND2_X1 U12452 ( .A1(n12041), .A2(n12040), .ZN(n12430) );
  NAND2_X1 U12453 ( .A1(n15433), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11769) );
  INV_X1 U12454 ( .A(n12105), .ZN(n19157) );
  OAI21_X1 U12455 ( .B1(n13163), .B2(n14451), .A(n11179), .ZN(n14330) );
  AND2_X1 U12456 ( .A1(n10296), .A2(n10295), .ZN(n9849) );
  NOR3_X1 U12457 ( .A1(n13424), .A2(n13423), .A3(n13412), .ZN(n13415) );
  OR2_X1 U12458 ( .A1(n13985), .A2(n13984), .ZN(n9850) );
  AND2_X1 U12459 ( .A1(n13383), .A2(n10228), .ZN(n9851) );
  AND2_X1 U12460 ( .A1(n10073), .A2(n18867), .ZN(n9852) );
  OR2_X1 U12461 ( .A1(n15751), .A2(n10184), .ZN(n9853) );
  AND2_X1 U12462 ( .A1(n11904), .A2(n12483), .ZN(n9854) );
  INV_X2 U12463 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12694) );
  INV_X1 U12464 ( .A(n14855), .ZN(n10051) );
  AND2_X1 U12465 ( .A1(n14018), .A2(n11907), .ZN(n9855) );
  INV_X1 U12466 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10317) );
  NAND2_X1 U12467 ( .A1(n13015), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9856) );
  AND2_X1 U12468 ( .A1(n9989), .A2(n9993), .ZN(n9857) );
  OR2_X1 U12469 ( .A1(n18499), .A2(n16232), .ZN(n9858) );
  NAND2_X1 U12470 ( .A1(n13322), .A2(n13321), .ZN(n13352) );
  NOR2_X1 U12471 ( .A1(n14876), .A2(n14882), .ZN(n9859) );
  AND2_X1 U12472 ( .A1(n12440), .A2(n12439), .ZN(n12678) );
  INV_X1 U12473 ( .A(n12678), .ZN(n10249) );
  INV_X1 U12474 ( .A(n10091), .ZN(n11188) );
  AOI21_X1 U12475 ( .B1(n13163), .B2(n11179), .A(n10092), .ZN(n10091) );
  NOR2_X1 U12476 ( .A1(n10554), .A2(n11165), .ZN(n11162) );
  NAND2_X1 U12477 ( .A1(n14174), .A2(n10159), .ZN(n14163) );
  NAND2_X1 U12478 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15569), .ZN(
        n9860) );
  AND2_X1 U12479 ( .A1(n9864), .A2(n9854), .ZN(n9861) );
  AND2_X1 U12480 ( .A1(n10067), .A2(n12960), .ZN(n9862) );
  INV_X1 U12481 ( .A(n10049), .ZN(n10046) );
  NAND2_X1 U12482 ( .A1(n9859), .A2(n10050), .ZN(n10049) );
  AND2_X1 U12483 ( .A1(n10039), .A2(n13542), .ZN(n9863) );
  AND2_X2 U12484 ( .A1(n15443), .A2(n19157), .ZN(n9864) );
  OR2_X1 U12485 ( .A1(n14399), .A2(n14398), .ZN(n9865) );
  NOR2_X1 U12486 ( .A1(n18506), .A2(n17876), .ZN(n17930) );
  NOR2_X1 U12487 ( .A1(n14397), .A2(n9865), .ZN(n9866) );
  AND2_X1 U12488 ( .A1(n14303), .A2(n9833), .ZN(n9867) );
  AND2_X1 U12489 ( .A1(n13378), .A2(n13377), .ZN(n13538) );
  INV_X1 U12490 ( .A(n13538), .ZN(n10037) );
  INV_X1 U12491 ( .A(n10141), .ZN(n10140) );
  NOR2_X1 U12492 ( .A1(n17649), .A2(n10142), .ZN(n10141) );
  AND2_X1 U12493 ( .A1(n10041), .A2(n10046), .ZN(n9868) );
  INV_X1 U12494 ( .A(n9981), .ZN(n9980) );
  NAND2_X1 U12495 ( .A1(n11119), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9981) );
  OR2_X1 U12496 ( .A1(n11846), .A2(n10613), .ZN(n10315) );
  INV_X1 U12497 ( .A(n11190), .ZN(n9991) );
  AND2_X1 U12498 ( .A1(n10444), .A2(n10402), .ZN(n11271) );
  AND2_X1 U12499 ( .A1(n14018), .A2(n19616), .ZN(n12197) );
  NAND2_X1 U12500 ( .A1(n18980), .A2(n12735), .ZN(n12993) );
  NAND2_X1 U12501 ( .A1(n18980), .A2(n10298), .ZN(n13722) );
  AND2_X1 U12502 ( .A1(n17491), .A2(n10095), .ZN(n9869) );
  AND2_X1 U12503 ( .A1(n13035), .A2(n10030), .ZN(n9870) );
  AND2_X1 U12504 ( .A1(n14549), .A2(n10027), .ZN(n9871) );
  AND2_X1 U12505 ( .A1(n10607), .A2(n10606), .ZN(n10671) );
  INV_X1 U12506 ( .A(n10217), .ZN(n12053) );
  OR2_X1 U12507 ( .A1(n10193), .A2(n10191), .ZN(n9872) );
  NOR2_X1 U12508 ( .A1(n12982), .A2(n13074), .ZN(n9873) );
  OR2_X1 U12509 ( .A1(n12176), .A2(n12175), .ZN(n13528) );
  OR3_X1 U12510 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17432), .ZN(n9874) );
  AND2_X1 U12511 ( .A1(n14951), .A2(n13757), .ZN(n9875) );
  AND2_X1 U12512 ( .A1(n13166), .A2(n10177), .ZN(n9876) );
  AND2_X1 U12513 ( .A1(n15192), .A2(n10201), .ZN(n14649) );
  NOR2_X1 U12514 ( .A1(n14786), .A2(n14785), .ZN(n14784) );
  AND2_X1 U12515 ( .A1(n14930), .A2(n14987), .ZN(n9877) );
  OR3_X1 U12516 ( .A1(n13130), .A2(n10180), .A3(n10182), .ZN(n9878) );
  NAND2_X1 U12517 ( .A1(n13754), .A2(n10304), .ZN(n10303) );
  AND2_X1 U12518 ( .A1(n10431), .A2(n9953), .ZN(n9879) );
  AND2_X1 U12519 ( .A1(n13528), .A2(n10222), .ZN(n9880) );
  OR2_X1 U12520 ( .A1(n11120), .A2(n10554), .ZN(n9881) );
  INV_X1 U12521 ( .A(n13402), .ZN(n10064) );
  NAND2_X1 U12522 ( .A1(n10059), .A2(n15269), .ZN(n9882) );
  NAND2_X1 U12523 ( .A1(n17617), .A2(n17848), .ZN(n9883) );
  AND2_X1 U12524 ( .A1(n13754), .A2(n13756), .ZN(n9884) );
  NAND2_X1 U12525 ( .A1(n14928), .A2(n15008), .ZN(n9885) );
  INV_X1 U12526 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10521) );
  AND3_X1 U12527 ( .A1(n9996), .A2(n11397), .A3(n11282), .ZN(n9886) );
  OR2_X1 U12528 ( .A1(n12536), .A2(n12535), .ZN(n18984) );
  AND2_X1 U12529 ( .A1(n13383), .A2(n10229), .ZN(n9887) );
  AND2_X1 U12530 ( .A1(n10148), .A2(n10147), .ZN(n9888) );
  AND2_X1 U12531 ( .A1(n10071), .A2(n10070), .ZN(n9889) );
  AND2_X1 U12532 ( .A1(n13297), .A2(n9880), .ZN(n9890) );
  AND2_X1 U12533 ( .A1(n10288), .A2(n18984), .ZN(n9891) );
  NAND2_X1 U12534 ( .A1(n10593), .A2(n10592), .ZN(n9892) );
  AND2_X1 U12535 ( .A1(n9830), .A2(n10094), .ZN(n9893) );
  NAND2_X1 U12536 ( .A1(n13270), .A2(n10055), .ZN(n10226) );
  INV_X1 U12537 ( .A(n10226), .ZN(n10223) );
  INV_X1 U12538 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18869) );
  OR2_X1 U12539 ( .A1(n13463), .A2(n15183), .ZN(n14959) );
  INV_X1 U12540 ( .A(n15430), .ZN(n19114) );
  OR2_X2 U12541 ( .A1(n12238), .A2(n12237), .ZN(n13510) );
  NOR2_X1 U12542 ( .A1(n12524), .A2(n13702), .ZN(n9894) );
  INV_X1 U12543 ( .A(n20003), .ZN(n20027) );
  INV_X1 U12544 ( .A(n11378), .ZN(n9998) );
  NAND2_X2 U12545 ( .A1(n12052), .A2(n12788), .ZN(n19056) );
  NAND2_X1 U12546 ( .A1(n18754), .A2(n13454), .ZN(n9895) );
  AND2_X1 U12547 ( .A1(n12941), .A2(n9837), .ZN(n9896) );
  AND2_X1 U12548 ( .A1(n14558), .A2(n10023), .ZN(n9897) );
  INV_X1 U12549 ( .A(n13448), .ZN(n10072) );
  AND2_X1 U12550 ( .A1(n10194), .A2(n14584), .ZN(n9898) );
  AND2_X1 U12551 ( .A1(n13924), .A2(n13947), .ZN(n9899) );
  NAND3_X1 U12552 ( .A1(n11509), .A2(n11508), .A3(n11507), .ZN(n18708) );
  AND2_X1 U12553 ( .A1(n11902), .A2(n9864), .ZN(n9900) );
  AND2_X1 U12554 ( .A1(n10925), .A2(n10924), .ZN(n9901) );
  AND2_X1 U12555 ( .A1(n10304), .A2(n14792), .ZN(n9902) );
  AND2_X1 U12556 ( .A1(n10138), .A2(n10136), .ZN(n9903) );
  NAND2_X1 U12557 ( .A1(n12518), .A2(n10288), .ZN(n10289) );
  INV_X1 U12558 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10150) );
  NAND2_X1 U12559 ( .A1(n10295), .A2(n10293), .ZN(n9904) );
  AND2_X1 U12560 ( .A1(n9898), .A2(n14570), .ZN(n9905) );
  AND2_X1 U12561 ( .A1(n14170), .A2(n14178), .ZN(n9906) );
  AND2_X1 U12562 ( .A1(n10177), .A2(n14165), .ZN(n9907) );
  INV_X1 U12563 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10081) );
  AND2_X1 U12564 ( .A1(n10176), .A2(n11314), .ZN(n9908) );
  INV_X1 U12565 ( .A(n17637), .ZN(n10098) );
  AND2_X1 U12566 ( .A1(n16271), .A2(n10108), .ZN(n9909) );
  OR2_X1 U12567 ( .A1(n11336), .A2(n11335), .ZN(n9910) );
  INV_X1 U12568 ( .A(n10381), .ZN(n9932) );
  AND2_X1 U12569 ( .A1(n10122), .A2(n10121), .ZN(n9911) );
  INV_X1 U12570 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10032) );
  INV_X1 U12571 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10070) );
  AND2_X1 U12572 ( .A1(n12018), .A2(n12943), .ZN(n18885) );
  INV_X1 U12573 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10109) );
  INV_X1 U12574 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10025) );
  INV_X1 U12575 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10110) );
  AND4_X1 U12576 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9912) );
  INV_X1 U12577 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10111) );
  INV_X1 U12578 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10100) );
  INV_X1 U12579 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10028) );
  NOR2_X1 U12580 ( .A1(n18703), .A2(n17256), .ZN(n17268) );
  OR2_X1 U12581 ( .A1(n19423), .A2(n19030), .ZN(n19421) );
  AND2_X1 U12582 ( .A1(n19423), .A2(n19030), .ZN(n19323) );
  NOR2_X1 U12583 ( .A1(n19423), .A2(n19791), .ZN(n19571) );
  AOI22_X2 U12584 ( .A1(DATAI_21_), .A2(n20046), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20090), .ZN(n20609) );
  AOI22_X2 U12585 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20090), .B1(DATAI_19_), 
        .B2(n20046), .ZN(n20597) );
  AOI22_X2 U12586 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20090), .B1(DATAI_30_), 
        .B2(n20046), .ZN(n20555) );
  NOR3_X2 U12587 ( .A1(n18410), .A2(n18536), .A3(n18291), .ZN(n18260) );
  NOR3_X2 U12588 ( .A1(n18410), .A2(n18536), .A3(n18201), .ZN(n18172) );
  NOR3_X2 U12589 ( .A1(n18410), .A2(n18536), .A3(n18386), .ZN(n18354) );
  AOI22_X2 U12590 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19173), .ZN(n19678) );
  AOI22_X2 U12591 ( .A1(DATAI_20_), .A2(n20046), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20090), .ZN(n20603) );
  NOR3_X2 U12592 ( .A1(n18410), .A2(n18362), .A3(n18386), .ZN(n18332) );
  NOR2_X2 U12593 ( .A1(n19175), .A2(n10003), .ZN(n19668) );
  NAND2_X1 U12594 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19624), .ZN(n19175) );
  NAND2_X2 U12595 ( .A1(n9916), .A2(n9914), .ZN(n14295) );
  NAND3_X1 U12596 ( .A1(n10550), .A2(n10535), .A3(n10081), .ZN(n9917) );
  NAND2_X2 U12597 ( .A1(n9918), .A2(n10530), .ZN(n10550) );
  NAND2_X2 U12598 ( .A1(n11170), .A2(n10274), .ZN(n14382) );
  NAND3_X1 U12599 ( .A1(n10402), .A2(n10444), .A3(n20066), .ZN(n11420) );
  AND3_X2 U12600 ( .A1(n10447), .A2(n9929), .A3(n9928), .ZN(n10444) );
  NAND2_X2 U12601 ( .A1(n10433), .A2(n10430), .ZN(n10381) );
  XNOR2_X2 U12602 ( .A(n13527), .B(n13329), .ZN(n15038) );
  NAND3_X1 U12603 ( .A1(n10218), .A2(n13293), .A3(n13292), .ZN(n10225) );
  NAND2_X1 U12604 ( .A1(n10202), .A2(n14018), .ZN(n9933) );
  NAND2_X1 U12605 ( .A1(n15038), .A2(n15037), .ZN(n13525) );
  NAND3_X1 U12606 ( .A1(n13534), .A2(n19112), .A3(n15386), .ZN(n15391) );
  NAND4_X1 U12607 ( .A1(n13534), .A2(n19112), .A3(n15386), .A4(n9863), .ZN(
        n9937) );
  NAND2_X1 U12608 ( .A1(n11910), .A2(n10217), .ZN(n9938) );
  AND2_X2 U12609 ( .A1(n12042), .A2(n11898), .ZN(n10217) );
  NAND2_X1 U12610 ( .A1(n12078), .A2(n19162), .ZN(n9939) );
  NAND2_X1 U12611 ( .A1(n11898), .A2(n12038), .ZN(n11911) );
  NAND2_X1 U12612 ( .A1(n12042), .A2(n11963), .ZN(n11905) );
  INV_X2 U12613 ( .A(n13262), .ZN(n13691) );
  NAND2_X2 U12614 ( .A1(n14877), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15083) );
  AND2_X2 U12615 ( .A1(n14896), .A2(n15090), .ZN(n14877) );
  NOR2_X2 U12616 ( .A1(n14973), .A2(n10214), .ZN(n14896) );
  NOR2_X2 U12617 ( .A1(n16301), .A2(n9948), .ZN(n15715) );
  INV_X1 U12618 ( .A(n9949), .ZN(n15585) );
  NAND2_X1 U12619 ( .A1(n10136), .A2(n10141), .ZN(n9950) );
  INV_X1 U12620 ( .A(n10136), .ZN(n9951) );
  NAND2_X1 U12621 ( .A1(n9953), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10770) );
  NAND4_X1 U12622 ( .A1(n11424), .A2(n20070), .A3(n20074), .A4(n9953), .ZN(
        n11840) );
  NAND2_X1 U12623 ( .A1(n12380), .A2(n9953), .ZN(n11285) );
  NAND2_X1 U12624 ( .A1(n9991), .A2(n9953), .ZN(n11288) );
  NAND2_X1 U12625 ( .A1(n11114), .A2(n9953), .ZN(n10633) );
  INV_X2 U12626 ( .A(n11423), .ZN(n9953) );
  NAND2_X1 U12627 ( .A1(n9962), .A2(n10271), .ZN(n15914) );
  NAND2_X1 U12628 ( .A1(n10634), .A2(n9965), .ZN(n9963) );
  NAND2_X1 U12629 ( .A1(n9963), .A2(n9964), .ZN(n10506) );
  NAND2_X1 U12630 ( .A1(n12582), .A2(n9967), .ZN(n9979) );
  AND2_X1 U12631 ( .A1(n12583), .A2(n20019), .ZN(n9967) );
  NAND2_X1 U12632 ( .A1(n9979), .A2(n9982), .ZN(n9978) );
  NAND2_X1 U12633 ( .A1(n9825), .A2(n14331), .ZN(n9968) );
  INV_X1 U12634 ( .A(n11119), .ZN(n9983) );
  NAND3_X1 U12635 ( .A1(n9981), .A2(n9982), .A3(n9979), .ZN(n9977) );
  NAND2_X1 U12636 ( .A1(n14295), .A2(n9867), .ZN(n9985) );
  NAND2_X1 U12637 ( .A1(n10634), .A2(n9988), .ZN(n9987) );
  NAND3_X1 U12638 ( .A1(n10436), .A2(n10448), .A3(n20079), .ZN(n11273) );
  AND2_X1 U12639 ( .A1(n9995), .A2(n11247), .ZN(n15680) );
  NAND2_X1 U12640 ( .A1(n9998), .A2(n9997), .ZN(n9996) );
  OR2_X1 U12641 ( .A1(n14382), .A2(n10000), .ZN(n9999) );
  NOR2_X2 U12642 ( .A1(n19056), .A2(n12483), .ZN(n19057) );
  NAND3_X1 U12643 ( .A1(n13268), .A2(n10221), .A3(n10004), .ZN(n10202) );
  NAND2_X1 U12644 ( .A1(n10005), .A2(n12438), .ZN(n12679) );
  NAND3_X1 U12645 ( .A1(n10005), .A2(n12438), .A3(n10251), .ZN(n10250) );
  NAND2_X1 U12646 ( .A1(n12434), .A2(n12433), .ZN(n10005) );
  OR2_X1 U12647 ( .A1(n15268), .A2(n10010), .ZN(n10006) );
  NAND2_X1 U12648 ( .A1(n10006), .A2(n10008), .ZN(n15006) );
  AND2_X1 U12649 ( .A1(n14985), .A2(n10018), .ZN(n14961) );
  NAND3_X1 U12650 ( .A1(n16066), .A2(n16065), .A3(n10021), .ZN(P2_U2826) );
  NAND2_X1 U12651 ( .A1(n14558), .A2(n10022), .ZN(n14542) );
  INV_X1 U12652 ( .A(n13353), .ZN(n10040) );
  OAI21_X1 U12653 ( .B1(n13353), .B2(n13352), .A(n10037), .ZN(n10039) );
  NAND3_X1 U12654 ( .A1(n10039), .A2(n13543), .A3(n13542), .ZN(n10038) );
  NAND2_X1 U12655 ( .A1(n14895), .A2(n10047), .ZN(n10041) );
  NAND2_X1 U12656 ( .A1(n14895), .A2(n10044), .ZN(n10043) );
  NAND2_X1 U12657 ( .A1(n12424), .A2(n19162), .ZN(n12096) );
  NAND2_X1 U12658 ( .A1(n10065), .A2(n13493), .ZN(n13495) );
  NAND2_X1 U12659 ( .A1(n9868), .A2(n9819), .ZN(n10065) );
  NAND2_X1 U12660 ( .A1(n11965), .A2(n11966), .ZN(n13065) );
  NAND2_X1 U12661 ( .A1(n13449), .A2(n13448), .ZN(n13447) );
  AND2_X2 U12662 ( .A1(n13449), .A2(n9889), .ZN(n13443) );
  NAND3_X1 U12663 ( .A1(n10078), .A2(n10077), .A3(n13416), .ZN(n10076) );
  NAND2_X1 U12664 ( .A1(n11846), .A2(n11406), .ZN(n10437) );
  NAND2_X2 U12665 ( .A1(n11846), .A2(n11423), .ZN(n11433) );
  NAND2_X1 U12666 ( .A1(n11289), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10083) );
  OAI211_X1 U12667 ( .C1(n10510), .C2(n10521), .A(n10082), .B(n10079), .ZN(
        n10511) );
  NAND2_X1 U12668 ( .A1(n11289), .A2(n10080), .ZN(n10079) );
  NAND2_X1 U12669 ( .A1(n10083), .A2(n10510), .ZN(n10525) );
  NAND2_X1 U12670 ( .A1(n13165), .A2(n10089), .ZN(n10088) );
  INV_X1 U12671 ( .A(n10092), .ZN(n10090) );
  INV_X1 U12672 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10097) );
  NAND3_X1 U12673 ( .A1(n10098), .A2(n9831), .A3(n17504), .ZN(n17506) );
  AOI21_X1 U12674 ( .B1(n16271), .B2(n10103), .A(n10102), .ZN(n10101) );
  NAND2_X1 U12675 ( .A1(n10112), .A2(n16293), .ZN(n16294) );
  NAND2_X1 U12676 ( .A1(n17346), .A2(n10113), .ZN(n10112) );
  NAND2_X1 U12677 ( .A1(n17347), .A2(n17348), .ZN(n17346) );
  NAND2_X1 U12678 ( .A1(n17365), .A2(n16301), .ZN(n17347) );
  NAND2_X1 U12679 ( .A1(n15651), .A2(n15650), .ZN(n10117) );
  NAND2_X2 U12680 ( .A1(n17496), .A2(n15647), .ZN(n17415) );
  NAND3_X1 U12681 ( .A1(n15489), .A2(n15490), .A3(n10126), .ZN(n10125) );
  NAND3_X1 U12682 ( .A1(n15513), .A2(n10132), .A3(n10129), .ZN(n15611) );
  NAND3_X1 U12683 ( .A1(n15515), .A2(n15510), .A3(n10134), .ZN(n10133) );
  INV_X1 U12684 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10142) );
  INV_X2 U12685 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18675) );
  NOR2_X2 U12686 ( .A1(n12982), .A2(n10143), .ZN(n13080) );
  NAND2_X1 U12687 ( .A1(n10594), .A2(n9888), .ZN(n10145) );
  NAND2_X1 U12688 ( .A1(n10594), .A2(n9892), .ZN(n10672) );
  AND2_X2 U12689 ( .A1(n10318), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12383) );
  AOI22_X1 U12690 ( .A1(n9810), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10319) );
  AND2_X2 U12691 ( .A1(n10323), .A2(n14516), .ZN(n10403) );
  AND2_X2 U12692 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14516) );
  NAND2_X1 U12693 ( .A1(n10156), .A2(n12590), .ZN(n10652) );
  NOR2_X1 U12694 ( .A1(n14107), .A2(n14108), .ZN(n14098) );
  NOR2_X2 U12695 ( .A1(n10150), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10256) );
  NAND2_X1 U12696 ( .A1(n12814), .A2(n11837), .ZN(n10176) );
  NAND2_X1 U12697 ( .A1(n10176), .A2(n10171), .ZN(n12757) );
  INV_X1 U12698 ( .A(n12577), .ZN(n10175) );
  NAND2_X1 U12699 ( .A1(n13166), .A2(n9907), .ZN(n15749) );
  INV_X1 U12700 ( .A(n13138), .ZN(n10182) );
  INV_X1 U12701 ( .A(n14095), .ZN(n10186) );
  NAND3_X1 U12702 ( .A1(n9818), .A2(n13647), .A3(n14826), .ZN(n10188) );
  NAND2_X1 U12704 ( .A1(n11727), .A2(n11919), .ZN(n11920) );
  NAND2_X1 U12705 ( .A1(n10217), .A2(n12105), .ZN(n10286) );
  NAND2_X1 U12706 ( .A1(n12197), .A2(n10217), .ZN(n12190) );
  NAND3_X1 U12707 ( .A1(n10219), .A2(n10225), .A3(n9890), .ZN(n13353) );
  NAND4_X1 U12708 ( .A1(n10221), .A2(n13268), .A3(n9824), .A4(n10220), .ZN(
        n10219) );
  NAND2_X1 U12709 ( .A1(n13269), .A2(n10224), .ZN(n10227) );
  NAND2_X2 U12710 ( .A1(n11930), .A2(n10231), .ZN(n12467) );
  AND3_X2 U12711 ( .A1(n11925), .A2(n11923), .A3(n11924), .ZN(n11930) );
  MUX2_X1 U12712 ( .A(n15478), .B(n10233), .S(n12096), .Z(n12097) );
  INV_X1 U12713 ( .A(n13029), .ZN(n10234) );
  NAND2_X1 U12714 ( .A1(n10234), .A2(n10235), .ZN(n15278) );
  INV_X1 U12715 ( .A(n14705), .ZN(n10244) );
  NAND2_X1 U12716 ( .A1(n14978), .A2(n10245), .ZN(n14648) );
  NAND3_X1 U12717 ( .A1(n10250), .A2(n12488), .A3(n10247), .ZN(n12494) );
  NOR2_X2 U12718 ( .A1(n18936), .A2(n10252), .ZN(n13702) );
  AND2_X2 U12720 ( .A1(n12383), .A2(n10256), .ZN(n10408) );
  AND3_X2 U12721 ( .A1(n10260), .A2(n10343), .A3(n10342), .ZN(n10261) );
  XNOR2_X2 U12722 ( .A(n11118), .B(n20036), .ZN(n12583) );
  NAND3_X1 U12723 ( .A1(n11420), .A2(n11412), .A3(n10263), .ZN(n10432) );
  NOR2_X1 U12724 ( .A1(n12342), .A2(n20051), .ZN(n11748) );
  NAND2_X1 U12725 ( .A1(n11420), .A2(n11425), .ZN(n11414) );
  INV_X1 U12726 ( .A(n11748), .ZN(n11834) );
  NAND3_X2 U12727 ( .A1(n11628), .A2(n10276), .A3(n10275), .ZN(n11633) );
  INV_X1 U12728 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10275) );
  AND2_X2 U12729 ( .A1(n10282), .A2(n10279), .ZN(n12038) );
  NAND4_X1 U12730 ( .A1(n12047), .A2(n11897), .A3(n9864), .A4(n10316), .ZN(
        n11931) );
  NAND2_X1 U12731 ( .A1(n11899), .A2(n19157), .ZN(n10283) );
  NAND4_X1 U12732 ( .A1(n11931), .A2(n11900), .A3(n10284), .A4(n10287), .ZN(
        n11903) );
  NAND2_X2 U12733 ( .A1(n11708), .A2(n12075), .ZN(n11900) );
  AND2_X2 U12734 ( .A1(n12518), .A2(n9891), .ZN(n13706) );
  INV_X1 U12735 ( .A(n10289), .ZN(n12730) );
  INV_X1 U12736 ( .A(n10296), .ZN(n13858) );
  NAND2_X1 U12738 ( .A1(n13054), .A2(n13056), .ZN(n13055) );
  NAND2_X1 U12739 ( .A1(n10307), .A2(n10640), .ZN(n12580) );
  CLKBUF_X1 U12740 ( .A(n11901), .Z(n15478) );
  NAND2_X1 U12741 ( .A1(n11660), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11661) );
  NAND2_X1 U12742 ( .A1(n14147), .A2(n10805), .ZN(n14148) );
  NAND2_X1 U12743 ( .A1(n11249), .A2(n19994), .ZN(n11258) );
  AOI211_X2 U12744 ( .C1(n15048), .C2(n19115), .A(n14843), .B(n14842), .ZN(
        n14844) );
  AOI211_X2 U12745 ( .C1(n15048), .C2(n19129), .A(n15047), .B(n15046), .ZN(
        n15049) );
  NAND2_X1 U12746 ( .A1(n13027), .A2(n13028), .ZN(n13029) );
  NAND2_X1 U12747 ( .A1(n12075), .A2(n10055), .ZN(n11901) );
  NOR2_X1 U12748 ( .A1(n11406), .A2(n10430), .ZN(n11424) );
  NAND2_X1 U12749 ( .A1(n10483), .A2(n11406), .ZN(n11228) );
  XNOR2_X1 U12750 ( .A(n13551), .B(n13646), .ZN(n14832) );
  AND2_X2 U12751 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12656) );
  XNOR2_X1 U12752 ( .A(n12940), .B(n12939), .ZN(n19423) );
  INV_X1 U12753 ( .A(n12641), .ZN(n20047) );
  AND2_X1 U12754 ( .A1(n20048), .A2(n12641), .ZN(n20425) );
  OAI21_X1 U12755 ( .B1(n13054), .B2(n13056), .A(n13055), .ZN(n19772) );
  NAND2_X1 U12756 ( .A1(n14665), .A2(n14664), .ZN(n14663) );
  AOI211_X2 U12757 ( .C1(n15899), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        n14293) );
  NAND2_X1 U12758 ( .A1(n13239), .A2(n18958), .ZN(n13251) );
  NAND2_X1 U12759 ( .A1(n11468), .A2(n19915), .ZN(n11473) );
  INV_X1 U12760 ( .A(n11468), .ZN(n14069) );
  NAND2_X1 U12761 ( .A1(n12037), .A2(n12475), .ZN(n12041) );
  NAND2_X1 U12762 ( .A1(n11734), .A2(n12694), .ZN(n11742) );
  INV_X1 U12763 ( .A(n19994), .ZN(n19817) );
  AND3_X1 U12764 ( .A1(n15694), .A2(n15680), .A3(n11248), .ZN(n19994) );
  INV_X1 U12765 ( .A(n11525), .ZN(n11567) );
  NOR2_X1 U12766 ( .A1(n11495), .A2(n11498), .ZN(n11496) );
  INV_X1 U12767 ( .A(n14147), .ZN(n14205) );
  INV_X1 U12768 ( .A(n10612), .ZN(n12792) );
  INV_X1 U12769 ( .A(n12792), .ZN(n11099) );
  AND2_X1 U12770 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10308) );
  INV_X1 U12771 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15409) );
  INV_X1 U12772 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19390) );
  AOI21_X1 U12773 ( .B1(n13263), .B2(n12475), .A(n10312), .ZN(n12938) );
  AND2_X1 U12774 ( .A1(n14396), .A2(n14395), .ZN(n10310) );
  AND2_X1 U12775 ( .A1(n12038), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10311) );
  NAND2_X1 U12776 ( .A1(n12474), .A2(n12478), .ZN(n10312) );
  OR2_X1 U12777 ( .A1(n11179), .A2(n16010), .ZN(n10313) );
  AND2_X1 U12778 ( .A1(n19919), .A2(n11846), .ZN(n19915) );
  NOR2_X1 U12779 ( .A1(n17565), .A2(n17375), .ZN(n17693) );
  INV_X1 U12780 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11452) );
  INV_X1 U12781 ( .A(n14059), .ZN(n11471) );
  INV_X1 U12782 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10318) );
  INV_X1 U12783 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21018) );
  NOR2_X1 U12784 ( .A1(n11497), .A2(n11498), .ZN(n11576) );
  INV_X1 U12785 ( .A(n11493), .ZN(n16842) );
  OR2_X1 U12786 ( .A1(n12612), .A2(n12611), .ZN(n12735) );
  INV_X1 U12787 ( .A(n14730), .ZN(n16107) );
  AND2_X1 U12788 ( .A1(n12483), .A2(n11910), .ZN(n10316) );
  INV_X1 U12789 ( .A(n10403), .ZN(n12378) );
  INV_X1 U12790 ( .A(n11207), .ZN(n11214) );
  NAND2_X1 U12791 ( .A1(n11209), .A2(n11208), .ZN(n11218) );
  OR2_X1 U12792 ( .A1(n13311), .A2(n13278), .ZN(n13279) );
  OR2_X1 U12793 ( .A1(n11218), .A2(n20066), .ZN(n11235) );
  OAI22_X1 U12794 ( .A1(n19389), .A2(n13254), .B1(n13913), .B2(n19462), .ZN(
        n13267) );
  INV_X1 U12795 ( .A(n11235), .ZN(n11236) );
  INV_X1 U12796 ( .A(n11210), .ZN(n11205) );
  NAND2_X1 U12797 ( .A1(n11713), .A2(n11712), .ZN(n11719) );
  NOR2_X1 U12798 ( .A1(n11602), .A2(n11601), .ZN(n11603) );
  OR2_X1 U12799 ( .A1(n10605), .A2(n10604), .ZN(n11154) );
  NAND2_X1 U12800 ( .A1(n20051), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10553) );
  INV_X1 U12801 ( .A(n13528), .ZN(n13298) );
  INV_X1 U12802 ( .A(n11955), .ZN(n11956) );
  INV_X1 U12803 ( .A(n13898), .ZN(n13899) );
  NOR2_X1 U12804 ( .A1(n11962), .A2(n11961), .ZN(n13294) );
  AND2_X1 U12805 ( .A1(n11723), .A2(n11722), .ZN(n13040) );
  AOI21_X1 U12806 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n21014), .A(
        n11603), .ZN(n11604) );
  NAND2_X1 U12807 ( .A1(n10525), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10443) );
  INV_X1 U12808 ( .A(n11382), .ZN(n11393) );
  NOR2_X1 U12809 ( .A1(n11052), .A2(n14288), .ZN(n11053) );
  INV_X1 U12810 ( .A(n10973), .ZN(n10974) );
  INV_X1 U12811 ( .A(n11156), .ZN(n11165) );
  NAND2_X1 U12812 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10644) );
  INV_X1 U12813 ( .A(n11111), .ZN(n10487) );
  OR2_X2 U12814 ( .A1(n10360), .A2(n10359), .ZN(n10430) );
  AOI22_X1 U12815 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11665) );
  OR2_X1 U12816 ( .A1(n13923), .A2(n13925), .ZN(n13947) );
  OR2_X1 U12817 ( .A1(n13848), .A2(n13847), .ZN(n13854) );
  AOI21_X1 U12818 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18536), .A(
        n11600), .ZN(n11602) );
  INV_X1 U12819 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n21015) );
  NAND2_X1 U12820 ( .A1(n17617), .A2(n17719), .ZN(n15653) );
  NOR2_X1 U12821 ( .A1(n17211), .A2(n15558), .ZN(n15570) );
  INV_X1 U12822 ( .A(n11267), .ZN(n11199) );
  AND2_X1 U12823 ( .A1(n11326), .A2(n11325), .ZN(n16026) );
  INV_X1 U12824 ( .A(n14181), .ZN(n10871) );
  NOR2_X1 U12825 ( .A1(n15667), .A2(n10081), .ZN(n11096) );
  AND4_X1 U12826 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10425) );
  INV_X1 U12827 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10696) );
  AND2_X1 U12828 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10611), .ZN(
        n10643) );
  AND2_X1 U12829 ( .A1(n20035), .A2(n20034), .ZN(n14487) );
  INV_X1 U12830 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20457) );
  OR2_X1 U12831 ( .A1(n12289), .A2(n12288), .ZN(n18990) );
  AND2_X1 U12832 ( .A1(n9806), .A2(n13951), .ZN(n13953) );
  INV_X1 U12833 ( .A(n12484), .ZN(n12482) );
  AND2_X1 U12834 ( .A1(n12943), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12475) );
  OR2_X1 U12835 ( .A1(n18846), .A2(n13543), .ZN(n13439) );
  INV_X1 U12836 ( .A(n13510), .ZN(n13543) );
  AND2_X1 U12837 ( .A1(n13393), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15023) );
  AND3_X1 U12838 ( .A1(n12109), .A2(n12108), .A3(n12107), .ZN(n12689) );
  AOI21_X1 U12839 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20939), .A(
        n11609), .ZN(n11612) );
  NOR2_X1 U12840 ( .A1(n13176), .A2(n18526), .ZN(n11525) );
  NOR2_X1 U12841 ( .A1(n15496), .A2(n15495), .ZN(n15497) );
  AND2_X1 U12842 ( .A1(n15612), .A2(n15617), .ZN(n15627) );
  INV_X1 U12843 ( .A(n17930), .ZN(n17847) );
  AOI21_X1 U12844 ( .B1(n11597), .B2(n12832), .A(n11598), .ZN(n18514) );
  NOR2_X1 U12845 ( .A1(n18499), .A2(n16288), .ZN(n17894) );
  INV_X1 U12846 ( .A(n18514), .ZN(n18517) );
  AND2_X1 U12847 ( .A1(n11243), .A2(n11242), .ZN(n11244) );
  INV_X1 U12848 ( .A(n13167), .ZN(n11366) );
  OR2_X1 U12849 ( .A1(n11460), .A2(n11459), .ZN(n11461) );
  NAND2_X1 U12850 ( .A1(n12810), .A2(n12804), .ZN(n19891) );
  INV_X1 U12851 ( .A(n12579), .ZN(n10640) );
  OAI21_X1 U12852 ( .B1(n14317), .B2(n12792), .A(n10995), .ZN(n14108) );
  NAND2_X1 U12853 ( .A1(n10821), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10822) );
  INV_X1 U12854 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14389) );
  INV_X1 U12855 ( .A(n13166), .ZN(n14144) );
  NOR2_X1 U12856 ( .A1(n20714), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11254) );
  INV_X1 U12857 ( .A(n19986), .ZN(n20002) );
  NAND2_X1 U12858 ( .A1(n11408), .A2(n15669), .ZN(n15969) );
  NOR2_X1 U12859 ( .A1(n20211), .A2(n20210), .ZN(n20526) );
  OR3_X1 U12860 ( .A1(n20704), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20050), 
        .ZN(n20092) );
  NAND2_X1 U12861 ( .A1(n13467), .A2(n13466), .ZN(n13472) );
  NAND2_X1 U12862 ( .A1(n12973), .A2(n12972), .ZN(n18925) );
  OR2_X1 U12863 ( .A1(n15154), .A2(n13641), .ZN(n15103) );
  AND2_X1 U12864 ( .A1(n13420), .A2(n14929), .ZN(n14997) );
  INV_X1 U12865 ( .A(n13662), .ZN(n15206) );
  NAND2_X1 U12866 ( .A1(n15416), .A2(n12943), .ZN(n11945) );
  AND2_X1 U12867 ( .A1(n19358), .A2(n19357), .ZN(n19364) );
  INV_X1 U12868 ( .A(n19420), .ZN(n19424) );
  INV_X1 U12869 ( .A(n19453), .ZN(n19491) );
  INV_X1 U12870 ( .A(n19624), .ZN(n19281) );
  OAI21_X1 U12871 ( .B1(n11610), .B2(n12829), .A(n11612), .ZN(n15601) );
  NOR2_X1 U12872 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16693), .ZN(n16668) );
  OAI21_X1 U12873 ( .B1(n18709), .B2(P3_STATEBS16_REG_SCAN_IN), .A(n11617), 
        .ZN(n16661) );
  NAND2_X1 U12874 ( .A1(n17168), .A2(n17230), .ZN(n17199) );
  NAND2_X1 U12875 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17419), .ZN(
        n17392) );
  INV_X1 U12876 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17668) );
  NAND2_X1 U12877 ( .A1(n17546), .A2(n17708), .ZN(n17457) );
  NOR2_X1 U12878 ( .A1(n15642), .A2(n17613), .ZN(n17529) );
  INV_X1 U12879 ( .A(n19857), .ZN(n15758) );
  AND2_X1 U12880 ( .A1(n12810), .A2(n12802), .ZN(n19880) );
  OR2_X1 U12881 ( .A1(n13202), .A2(n15758), .ZN(n19832) );
  AND2_X1 U12882 ( .A1(n19857), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19897) );
  NOR2_X1 U12883 ( .A1(n19919), .A2(n11469), .ZN(n11470) );
  OR2_X1 U12884 ( .A1(n14085), .A2(n13193), .ZN(n13194) );
  INV_X1 U12885 ( .A(n12394), .ZN(n19983) );
  NAND2_X1 U12886 ( .A1(n10928), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10973) );
  NAND2_X1 U12887 ( .A1(n10890), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10927) );
  NAND2_X1 U12888 ( .A1(n10728), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10765) );
  INV_X1 U12889 ( .A(n15871), .ZN(n19987) );
  AND2_X1 U12890 ( .A1(n11101), .A2(n20496), .ZN(n19993) );
  AND2_X1 U12891 ( .A1(n14354), .A2(n15881), .ZN(n15954) );
  AND2_X1 U12892 ( .A1(n11254), .A2(n10613), .ZN(n19986) );
  INV_X1 U12893 ( .A(n20024), .ZN(n14491) );
  INV_X1 U12894 ( .A(n20002), .ZN(n20033) );
  NAND2_X1 U12895 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n15694), .ZN(n20706) );
  OAI22_X1 U12896 ( .A1(n20063), .A2(n20062), .B1(n20387), .B2(n20206), .ZN(
        n20096) );
  INV_X1 U12897 ( .A(n20625), .ZN(n20094) );
  OAI22_X1 U12898 ( .A1(n20135), .A2(n20134), .B1(n20265), .B2(n20387), .ZN(
        n20159) );
  NOR2_X1 U12899 ( .A1(n20048), .A2(n20047), .ZN(n20171) );
  INV_X1 U12900 ( .A(n20213), .ZN(n20230) );
  OR2_X1 U12901 ( .A1(n20129), .A2(n20049), .ZN(n20456) );
  OR2_X1 U12902 ( .A1(n20129), .A2(n11114), .ZN(n20238) );
  INV_X1 U12903 ( .A(n20321), .ZN(n20345) );
  INV_X1 U12904 ( .A(n20423), .ZN(n20378) );
  AND2_X1 U12905 ( .A1(n20129), .A2(n11114), .ZN(n20374) );
  AND2_X1 U12906 ( .A1(n20129), .A2(n20049), .ZN(n20424) );
  INV_X1 U12907 ( .A(n20458), .ZN(n20513) );
  OAI211_X1 U12908 ( .C1(n20556), .C2(n20527), .A(n20526), .B(n20525), .ZN(
        n20559) );
  INV_X1 U12909 ( .A(n20238), .ZN(n20487) );
  OR2_X1 U12910 ( .A1(n12704), .A2(n18734), .ZN(n18730) );
  INV_X1 U12911 ( .A(n18925), .ZN(n18950) );
  AND2_X1 U12912 ( .A1(n19100), .A2(n12971), .ZN(n18952) );
  NOR2_X1 U12913 ( .A1(n14705), .A2(n14704), .ZN(n14706) );
  OR2_X1 U12914 ( .A1(n12361), .A2(n12360), .ZN(n12484) );
  INV_X1 U12915 ( .A(n18992), .ZN(n18998) );
  INV_X1 U12916 ( .A(n12776), .ZN(n12630) );
  INV_X1 U12917 ( .A(n11887), .ZN(n19100) );
  CLKBUF_X1 U12918 ( .A(n11798), .Z(n11879) );
  AND2_X1 U12919 ( .A1(n12514), .A2(n12513), .ZN(n18876) );
  INV_X1 U12920 ( .A(n16179), .ZN(n19116) );
  INV_X1 U12921 ( .A(n18905), .ZN(n19132) );
  AND2_X1 U12922 ( .A1(n12123), .A2(n12696), .ZN(n13662) );
  INV_X1 U12923 ( .A(n16191), .ZN(n19121) );
  NOR2_X1 U12924 ( .A1(n12430), .A2(n12045), .ZN(n19791) );
  NAND2_X1 U12925 ( .A1(n11945), .A2(n11944), .ZN(n19624) );
  INV_X1 U12926 ( .A(n19764), .ZN(n19756) );
  OAI21_X1 U12927 ( .B1(n19147), .B2(n19143), .A(n19142), .ZN(n19181) );
  INV_X1 U12928 ( .A(n19218), .ZN(n19240) );
  AND2_X1 U12929 ( .A1(n19367), .A2(n19453), .ZN(n19302) );
  OAI21_X1 U12930 ( .B1(n15438), .B2(n19275), .A(n15437), .ZN(n19318) );
  AND2_X1 U12931 ( .A1(n19423), .A2(n19791), .ZN(n19367) );
  INV_X1 U12932 ( .A(n19452), .ZN(n19441) );
  NOR2_X2 U12933 ( .A1(n19421), .A2(n19424), .ZN(n19480) );
  AND2_X1 U12934 ( .A1(n19772), .A2(n19783), .ZN(n19453) );
  INV_X1 U12935 ( .A(n19635), .ZN(n19588) );
  INV_X1 U12936 ( .A(n19596), .ZN(n19608) );
  OAI22_X1 U12937 ( .A1(n19172), .A2(n19171), .B1(n19170), .B2(n19169), .ZN(
        n19662) );
  INV_X1 U12938 ( .A(n19421), .ZN(n19540) );
  NAND2_X1 U12939 ( .A1(n18706), .A2(n18496), .ZN(n17277) );
  INV_X1 U12940 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n17709) );
  NOR2_X1 U12941 ( .A1(n16532), .A2(n16431), .ZN(n16507) );
  INV_X1 U12942 ( .A(n16749), .ZN(n16770) );
  NOR2_X1 U12943 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16597), .ZN(n16578) );
  NOR2_X1 U12944 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16619), .ZN(n16603) );
  NOR2_X1 U12945 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16650), .ZN(n16649) );
  NOR2_X2 U12946 ( .A1(n16667), .A2(n16661), .ZN(n16749) );
  NOR4_X1 U12947 ( .A1(n15711), .A2(n18723), .A3(n16753), .A4(n18555), .ZN(
        n16773) );
  NOR2_X1 U12948 ( .A1(n16897), .A2(n16896), .ZN(n16895) );
  NOR2_X1 U12949 ( .A1(n17302), .A2(n17111), .ZN(n17107) );
  NAND2_X1 U12950 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17159), .ZN(n17158) );
  INV_X1 U12951 ( .A(n17195), .ZN(n17189) );
  INV_X1 U12952 ( .A(n17237), .ZN(n17215) );
  INV_X1 U12953 ( .A(n18057), .ZN(n17239) );
  NOR2_X1 U12954 ( .A1(n9952), .A2(n15648), .ZN(n17856) );
  INV_X1 U12955 ( .A(n18131), .ZN(n18364) );
  INV_X1 U12956 ( .A(n17973), .ZN(n18024) );
  INV_X1 U12957 ( .A(n18022), .ZN(n18032) );
  NAND2_X1 U12958 ( .A1(n18711), .A2(n18055), .ZN(n18131) );
  INV_X1 U12959 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18720) );
  INV_X1 U12960 ( .A(n19880), .ZN(n19892) );
  OR2_X1 U12961 ( .A1(n12798), .A2(n12796), .ZN(n19847) );
  INV_X1 U12962 ( .A(n19901), .ZN(n19866) );
  INV_X2 U12963 ( .A(n14235), .ZN(n14271) );
  NAND2_X1 U12964 ( .A1(n19952), .A2(n19928), .ZN(n19925) );
  NAND2_X1 U12965 ( .A1(n11894), .A2(n11893), .ZN(n19952) );
  NOR2_X1 U12966 ( .A1(n12248), .A2(n12247), .ZN(n12320) );
  AOI21_X1 U12967 ( .B1(n13988), .B2(n19993), .A(n11463), .ZN(n11464) );
  OR2_X1 U12968 ( .A1(n19994), .A2(n11250), .ZN(n15871) );
  INV_X1 U12969 ( .A(n15899), .ZN(n19998) );
  NAND2_X1 U12970 ( .A1(n11408), .A2(n11407), .ZN(n20003) );
  AOI21_X1 U12971 ( .B1(n14491), .B2(n19999), .A(n11300), .ZN(n20014) );
  INV_X1 U12972 ( .A(n20031), .ZN(n15966) );
  INV_X1 U12973 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20375) );
  INV_X1 U12974 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12373) );
  NAND2_X1 U12975 ( .A1(n20171), .A2(n20322), .ZN(n20128) );
  NAND2_X1 U12976 ( .A1(n20171), .A2(n20487), .ZN(n20157) );
  NAND2_X1 U12977 ( .A1(n20171), .A2(n20374), .ZN(n20198) );
  OR2_X1 U12978 ( .A1(n20299), .A2(n20456), .ZN(n20259) );
  OR2_X1 U12979 ( .A1(n20299), .A2(n20238), .ZN(n20288) );
  OR2_X1 U12980 ( .A1(n20299), .A2(n20521), .ZN(n20314) );
  NAND2_X1 U12981 ( .A1(n20425), .A2(n20322), .ZN(n20373) );
  NAND2_X1 U12982 ( .A1(n20425), .A2(n20487), .ZN(n20423) );
  NAND2_X1 U12983 ( .A1(n20425), .A2(n20374), .ZN(n20449) );
  NAND2_X1 U12984 ( .A1(n20425), .A2(n20424), .ZN(n20486) );
  NAND2_X1 U12985 ( .A1(n20488), .A2(n20487), .ZN(n20562) );
  OR2_X1 U12986 ( .A1(n20572), .A2(n20298), .ZN(n20625) );
  INV_X1 U12987 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20704) );
  INV_X1 U12988 ( .A(n20703), .ZN(n20699) );
  INV_X1 U12989 ( .A(n20736), .ZN(n20667) );
  INV_X1 U12990 ( .A(n20691), .ZN(n20689) );
  INV_X1 U12991 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19683) );
  OR2_X1 U12992 ( .A1(n18949), .A2(n19616), .ZN(n18961) );
  NAND2_X1 U12993 ( .A1(n12950), .A2(n12949), .ZN(n18957) );
  AND2_X1 U12994 ( .A1(n13689), .A2(n13688), .ZN(n19780) );
  OR2_X1 U12995 ( .A1(n19056), .A2(n12053), .ZN(n19061) );
  INV_X1 U12996 ( .A(n19056), .ZN(n14810) );
  AND2_X1 U12997 ( .A1(n14811), .A2(n14049), .ZN(n19065) );
  OR2_X1 U12998 ( .A1(n19089), .A2(n19097), .ZN(n19091) );
  OR2_X1 U12999 ( .A1(n12969), .A2(n14018), .ZN(n11887) );
  INV_X1 U13000 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16138) );
  INV_X1 U13001 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16153) );
  INV_X1 U13002 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18906) );
  NAND2_X1 U13003 ( .A1(n12123), .A2(n19797), .ZN(n16192) );
  NAND2_X1 U13004 ( .A1(n19420), .A2(n19323), .ZN(n19211) );
  NAND2_X1 U13005 ( .A1(n19323), .A2(n19453), .ZN(n19263) );
  NAND2_X1 U13006 ( .A1(n19323), .A2(n19545), .ZN(n19322) );
  NAND2_X1 U13007 ( .A1(n19763), .A2(n19323), .ZN(n19380) );
  NAND2_X1 U13008 ( .A1(n19367), .A2(n19763), .ZN(n19413) );
  INV_X1 U13009 ( .A(n19480), .ZN(n19458) );
  NAND2_X1 U13010 ( .A1(n19571), .A2(n19420), .ZN(n19452) );
  NAND2_X1 U13011 ( .A1(n19571), .A2(n19453), .ZN(n19516) );
  AOI21_X1 U13012 ( .B1(n15456), .B2(n15457), .A(n15455), .ZN(n19539) );
  INV_X1 U13013 ( .A(n19626), .ZN(n19587) );
  INV_X1 U13014 ( .A(n19662), .ZN(n19606) );
  INV_X1 U13015 ( .A(n19523), .ZN(n19641) );
  NAND2_X1 U13016 ( .A1(n19571), .A2(n19763), .ZN(n19666) );
  INV_X1 U13017 ( .A(n19753), .ZN(n19679) );
  NAND2_X1 U13018 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16540), .ZN(n16532) );
  NAND2_X1 U13019 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16779), .ZN(n16745) );
  INV_X1 U13020 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16743) );
  NOR2_X1 U13021 ( .A1(n16517), .A2(n16834), .ZN(n16839) );
  AND2_X1 U13022 ( .A1(n17076), .A2(n17163), .ZN(n17080) );
  NOR2_X1 U13023 ( .A1(n15581), .A2(n15580), .ZN(n17204) );
  INV_X1 U13024 ( .A(n17225), .ZN(n17237) );
  INV_X1 U13025 ( .A(n17256), .ZN(n17276) );
  INV_X1 U13026 ( .A(n17565), .ZN(n17549) );
  INV_X1 U13027 ( .A(n17955), .ZN(n17942) );
  NAND2_X1 U13028 ( .A1(n15644), .A2(n18032), .ZN(n18037) );
  INV_X1 U13029 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18072) );
  INV_X1 U13030 ( .A(n18102), .ZN(n18446) );
  INV_X1 U13031 ( .A(n18116), .ZN(n18470) );
  INV_X1 U13032 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18711) );
  INV_X1 U13033 ( .A(n18656), .ZN(n18570) );
  INV_X1 U13034 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18584) );
  INV_X1 U13035 ( .A(n16341), .ZN(n16352) );
  NAND2_X1 U13036 ( .A1(n11473), .A2(n11472), .ZN(P1_U2842) );
  NOR2_X2 U13037 ( .A1(n10317), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10324) );
  NOR2_X4 U13038 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U13039 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10322) );
  AND2_X4 U13040 ( .A1(n12391), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12381) );
  AND2_X4 U13041 ( .A1(n14515), .A2(n12376), .ZN(n10997) );
  AOI22_X1 U13042 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13043 ( .A1(n10408), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10320) );
  NAND4_X1 U13044 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10330) );
  AOI22_X1 U13045 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10328) );
  AND2_X4 U13046 ( .A1(n12381), .A2(n14516), .ZN(n10414) );
  AOI22_X1 U13047 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9812), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13048 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10416), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10326) );
  AND2_X2 U13049 ( .A1(n12376), .A2(n14516), .ZN(n10488) );
  AOI22_X1 U13050 ( .A1(n10493), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10325) );
  NAND4_X1 U13051 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10329) );
  OR2_X2 U13052 ( .A1(n10330), .A2(n10329), .ZN(n11423) );
  AOI22_X1 U13053 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13054 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13055 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10416), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13056 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10331) );
  NAND4_X1 U13057 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10340) );
  AOI22_X1 U13058 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10408), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13059 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13060 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13061 ( .A1(n10493), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10335) );
  NAND4_X1 U13062 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10339) );
  AOI22_X1 U13063 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13064 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10416), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13065 ( .A1(n9810), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13066 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13067 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10408), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13068 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13069 ( .A1(n10493), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13070 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10494), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10354) );
  AOI22_X1 U13071 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10353) );
  AOI22_X1 U13072 ( .A1(n10493), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13073 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10351) );
  NAND4_X1 U13074 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10360) );
  AOI22_X1 U13075 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9813), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13076 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10416), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13077 ( .A1(n10408), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13078 ( .A1(n9810), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10355) );
  NAND4_X1 U13079 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10359) );
  AOI22_X1 U13080 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13081 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10416), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13082 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13083 ( .A1(n10493), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10361) );
  NAND4_X1 U13084 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10370) );
  AOI22_X1 U13085 ( .A1(n10408), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10494), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13086 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U13087 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13088 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10365) );
  NAND4_X1 U13089 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10369) );
  AOI22_X1 U13090 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13091 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10349), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U13092 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10416), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13093 ( .A1(n9810), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10371) );
  NAND4_X1 U13094 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10380) );
  AOI22_X1 U13095 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10408), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13096 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13097 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13098 ( .A1(n10493), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10488), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U13099 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10379) );
  NAND2_X1 U13100 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10385) );
  NAND2_X1 U13101 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10384) );
  NAND2_X1 U13102 ( .A1(n10408), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10383) );
  NAND2_X1 U13103 ( .A1(n10559), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U13104 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10389) );
  NAND2_X1 U13105 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10388) );
  NAND2_X1 U13106 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10387) );
  NAND2_X1 U13107 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10386) );
  NAND2_X1 U13108 ( .A1(n10493), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10393) );
  NAND2_X1 U13109 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10392) );
  NAND2_X1 U13110 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10391) );
  NAND2_X1 U13111 ( .A1(n10488), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10390) );
  NAND2_X1 U13112 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10397) );
  NAND2_X1 U13113 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10396) );
  NAND2_X1 U13114 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10395) );
  NAND2_X1 U13115 ( .A1(n10403), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10394) );
  AND4_X4 U13116 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n20051) );
  NAND2_X1 U13117 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10407) );
  NAND2_X1 U13118 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10406) );
  NAND2_X1 U13119 ( .A1(n10349), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10405) );
  NAND2_X1 U13120 ( .A1(n10403), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13121 ( .A1(n10408), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10413) );
  NAND2_X1 U13122 ( .A1(n10493), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10412) );
  NAND2_X1 U13123 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10411) );
  NAND2_X1 U13124 ( .A1(n10559), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10410) );
  NAND2_X1 U13125 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10420) );
  NAND2_X1 U13126 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10419) );
  NAND2_X1 U13127 ( .A1(n10350), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10418) );
  NAND2_X1 U13128 ( .A1(n10416), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10417) );
  NAND2_X1 U13129 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10424) );
  NAND2_X1 U13130 ( .A1(n10913), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U13131 ( .A1(n10488), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10422) );
  NAND2_X1 U13132 ( .A1(n10997), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10421) );
  NAND4_X4 U13133 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        n10434) );
  INV_X1 U13134 ( .A(n11840), .ZN(n10429) );
  NAND2_X2 U13135 ( .A1(n10429), .A2(n11846), .ZN(n12342) );
  NAND2_X1 U13136 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20637) );
  OAI21_X1 U13137 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20637), .ZN(n11260) );
  NAND2_X1 U13138 ( .A1(n10432), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10510) );
  OR2_X2 U13139 ( .A1(n20051), .A2(n10434), .ZN(n20729) );
  OR2_X1 U13141 ( .A1(n10381), .A2(n11349), .ZN(n12326) );
  NAND2_X1 U13142 ( .A1(n20051), .A2(n10434), .ZN(n12800) );
  OAI211_X1 U13143 ( .C1(n20729), .C2(n20079), .A(n12326), .B(n12800), .ZN(
        n10453) );
  NOR2_X1 U13144 ( .A1(n10453), .A2(n12380), .ZN(n10440) );
  OR2_X1 U13145 ( .A1(n10381), .A2(n11423), .ZN(n10436) );
  NAND2_X1 U13146 ( .A1(n20083), .A2(n11423), .ZN(n10435) );
  NAND2_X1 U13147 ( .A1(n11273), .A2(n15667), .ZN(n10456) );
  MUX2_X1 U13148 ( .A(n20070), .B(n10444), .S(n20051), .Z(n10439) );
  NAND2_X1 U13149 ( .A1(n20627), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15691) );
  NAND2_X1 U13150 ( .A1(n20627), .A2(n20704), .ZN(n20714) );
  MUX2_X1 U13151 ( .A(n15691), .B(n11254), .S(n20489), .Z(n10441) );
  INV_X1 U13152 ( .A(n10441), .ZN(n10442) );
  NAND2_X2 U13153 ( .A1(n10443), .A2(n10442), .ZN(n10513) );
  INV_X1 U13154 ( .A(n10444), .ZN(n10446) );
  NOR2_X1 U13155 ( .A1(n20070), .A2(n20051), .ZN(n10445) );
  AOI21_X1 U13156 ( .B1(n10446), .B2(n12795), .A(n10445), .ZN(n11284) );
  INV_X1 U13157 ( .A(n12795), .ZN(n11428) );
  AND2_X1 U13158 ( .A1(n11428), .A2(n11349), .ZN(n11754) );
  NAND2_X1 U13159 ( .A1(n11754), .A2(n10447), .ZN(n10452) );
  NOR2_X1 U13160 ( .A1(n20714), .A2(n10081), .ZN(n10451) );
  INV_X1 U13161 ( .A(n10448), .ZN(n10449) );
  NAND2_X1 U13162 ( .A1(n11889), .A2(n10449), .ZN(n10450) );
  NAND4_X1 U13163 ( .A1(n10452), .A2(n10451), .A3(n11285), .A4(n10450), .ZN(
        n10454) );
  NOR2_X1 U13164 ( .A1(n10454), .A2(n10453), .ZN(n10455) );
  OAI211_X1 U13165 ( .C1(n10456), .C2(n20066), .A(n11284), .B(n10455), .ZN(
        n10512) );
  INV_X1 U13166 ( .A(n10512), .ZN(n10457) );
  XNOR2_X2 U13167 ( .A(n10513), .B(n10457), .ZN(n10634) );
  AOI22_X1 U13168 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10409), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13169 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9811), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13170 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U13171 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10460) );
  NAND4_X1 U13172 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10470) );
  AOI22_X1 U13173 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13174 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10416), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13175 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13176 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10465) );
  NAND4_X1 U13177 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .ZN(
        n10469) );
  NOR2_X1 U13178 ( .A1(n10554), .A2(n11156), .ZN(n10502) );
  AOI22_X1 U13179 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13180 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13181 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10350), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13182 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10471) );
  NAND4_X1 U13183 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10480) );
  AOI22_X1 U13184 ( .A1(n10415), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U13185 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U13186 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U13187 ( .A1(n10892), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10475) );
  NAND4_X1 U13188 ( .A1(n10478), .A2(n10477), .A3(n10476), .A4(n10475), .ZN(
        n10479) );
  MUX2_X1 U13189 ( .A(n10502), .B(n11162), .S(n10487), .Z(n10481) );
  INV_X1 U13190 ( .A(n10481), .ZN(n10482) );
  INV_X1 U13191 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10484) );
  OR2_X1 U13192 ( .A1(n11228), .A2(n10484), .ZN(n10486) );
  AOI21_X1 U13193 ( .B1(n20079), .B2(n11156), .A(n10081), .ZN(n10485) );
  AOI22_X1 U13194 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13195 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9811), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13196 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13197 ( .A1(n10459), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10489) );
  NAND4_X1 U13198 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10500) );
  AOI22_X1 U13199 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13200 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13201 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13202 ( .A1(n10409), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10495) );
  NAND4_X1 U13203 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10499) );
  INV_X1 U13204 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10501) );
  OR2_X1 U13205 ( .A1(n11228), .A2(n10501), .ZN(n10504) );
  INV_X1 U13206 ( .A(n10502), .ZN(n10503) );
  OAI211_X1 U13207 ( .C1(n10515), .C2(n10553), .A(n10504), .B(n10503), .ZN(
        n10505) );
  NAND2_X1 U13208 ( .A1(n10506), .A2(n10505), .ZN(n10507) );
  NAND2_X2 U13209 ( .A1(n10517), .A2(n10507), .ZN(n10626) );
  INV_X1 U13210 ( .A(n10626), .ZN(n10520) );
  INV_X1 U13211 ( .A(n11254), .ZN(n10508) );
  NAND2_X1 U13212 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10528) );
  OAI21_X1 U13213 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10528), .ZN(n20381) );
  NAND2_X1 U13214 ( .A1(n15691), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10522) );
  OAI21_X1 U13215 ( .B1(n10508), .B2(n20381), .A(n10522), .ZN(n10509) );
  XNOR2_X2 U13216 ( .A(n10511), .B(n10524), .ZN(n20165) );
  NAND2_X1 U13217 ( .A1(n10513), .A2(n10512), .ZN(n10514) );
  OR2_X2 U13218 ( .A1(n20165), .A2(n10514), .ZN(n10534) );
  NAND2_X1 U13219 ( .A1(n20165), .A2(n10514), .ZN(n20100) );
  OR2_X1 U13220 ( .A1(n10554), .A2(n10515), .ZN(n10516) );
  INV_X1 U13221 ( .A(n11109), .ZN(n10519) );
  INV_X1 U13222 ( .A(n10517), .ZN(n10518) );
  AOI21_X2 U13223 ( .B1(n10520), .B2(n10519), .A(n10518), .ZN(n10617) );
  NAND2_X1 U13224 ( .A1(n10522), .A2(n10521), .ZN(n10523) );
  AND2_X1 U13225 ( .A1(n15691), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10526) );
  INV_X1 U13226 ( .A(n10528), .ZN(n10527) );
  NAND2_X1 U13227 ( .A1(n10527), .A2(n20375), .ZN(n20163) );
  NAND2_X1 U13228 ( .A1(n10528), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10529) );
  NAND2_X1 U13229 ( .A1(n20163), .A2(n10529), .ZN(n20060) );
  NAND2_X1 U13230 ( .A1(n11254), .A2(n20060), .ZN(n10531) );
  NAND2_X1 U13231 ( .A1(n10533), .A2(n10531), .ZN(n10530) );
  NAND4_X1 U13232 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n10535) );
  AOI22_X1 U13233 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13234 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13235 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13236 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10536) );
  NAND4_X1 U13237 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10545) );
  AOI22_X1 U13238 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13239 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13240 ( .A1(n10494), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13241 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10540) );
  NAND4_X1 U13242 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10544) );
  INV_X1 U13243 ( .A(n10553), .ZN(n10547) );
  AOI22_X1 U13244 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10547), .B2(n10546), .ZN(n10548) );
  XNOR2_X2 U13245 ( .A(n10549), .B(n10548), .ZN(n10618) );
  NAND2_X2 U13246 ( .A1(n10617), .A2(n10618), .ZN(n10642) );
  NAND2_X1 U13247 ( .A1(n9807), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10552) );
  NOR3_X1 U13248 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20375), .A3(
        n20457), .ZN(n20297) );
  NAND2_X1 U13249 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20297), .ZN(
        n20292) );
  NAND3_X1 U13250 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20570) );
  NOR2_X1 U13251 ( .A1(n20489), .A2(n20570), .ZN(n20616) );
  AOI21_X1 U13252 ( .B1(n20380), .B2(n20292), .A(n20616), .ZN(n20324) );
  AOI22_X1 U13253 ( .A1(n11254), .A2(n20324), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15691), .ZN(n10551) );
  XNOR2_X2 U13254 ( .A(n10550), .B(n20204), .ZN(n20323) );
  AOI22_X1 U13255 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13256 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13257 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13258 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10555) );
  NAND4_X1 U13259 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10565) );
  AOI22_X1 U13260 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13261 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13262 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13263 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10560) );
  NAND4_X1 U13264 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(
        n10564) );
  AOI22_X1 U13265 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11207), .B2(n11137), .ZN(n10566) );
  INV_X1 U13266 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10568) );
  OR2_X1 U13267 ( .A1(n11228), .A2(n10568), .ZN(n10580) );
  AOI22_X1 U13268 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13269 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11078), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13270 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10414), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13271 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10569) );
  NAND4_X1 U13272 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10578) );
  AOI22_X1 U13273 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n9799), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13274 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U13275 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13276 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10573) );
  NAND4_X1 U13277 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n10577) );
  NAND2_X1 U13278 ( .A1(n11207), .A2(n11136), .ZN(n10579) );
  INV_X1 U13279 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10581) );
  OR2_X1 U13280 ( .A1(n11228), .A2(n10581), .ZN(n10593) );
  AOI22_X1 U13281 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13282 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13283 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U13284 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10582) );
  NAND4_X1 U13285 ( .A1(n10585), .A2(n10584), .A3(n10583), .A4(n10582), .ZN(
        n10591) );
  AOI22_X1 U13286 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13287 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13288 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13289 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10586) );
  NAND4_X1 U13290 ( .A1(n10589), .A2(n10588), .A3(n10587), .A4(n10586), .ZN(
        n10590) );
  NAND2_X1 U13291 ( .A1(n11207), .A2(n11146), .ZN(n10592) );
  INV_X1 U13292 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10595) );
  OR2_X1 U13293 ( .A1(n11228), .A2(n10595), .ZN(n10607) );
  AOI22_X1 U13294 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13295 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13296 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13297 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10596) );
  NAND4_X1 U13298 ( .A1(n10599), .A2(n10598), .A3(n10597), .A4(n10596), .ZN(
        n10605) );
  AOI22_X1 U13299 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13300 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13301 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13302 ( .A1(n10459), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10600) );
  NAND4_X1 U13303 ( .A1(n10603), .A2(n10602), .A3(n10601), .A4(n10600), .ZN(
        n10604) );
  NAND2_X1 U13304 ( .A1(n11207), .A2(n11154), .ZN(n10606) );
  INV_X1 U13305 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13306 ( .A1(n11207), .A2(n11156), .ZN(n10608) );
  OAI21_X1 U13307 ( .B1(n11228), .B2(n10609), .A(n10608), .ZN(n10610) );
  INV_X1 U13308 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10615) );
  INV_X1 U13309 ( .A(n10644), .ZN(n10611) );
  OAI21_X1 U13310 ( .B1(n10673), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n10697), .ZN(n19859) );
  NOR2_X1 U13311 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13312 ( .A1(n19859), .A2(n11099), .B1(n11455), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10614) );
  OAI21_X1 U13313 ( .B1(n10315), .B2(n10615), .A(n10614), .ZN(n10616) );
  AOI21_X1 U13314 ( .B1(n11152), .B2(n10797), .A(n10616), .ZN(n12984) );
  INV_X1 U13315 ( .A(n12984), .ZN(n10681) );
  NAND2_X2 U13316 ( .A1(n10619), .A2(n10642), .ZN(n12641) );
  NAND2_X1 U13317 ( .A1(n10620), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10655) );
  XNOR2_X1 U13318 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12928) );
  AOI21_X1 U13319 ( .B1(n10612), .B2(n12928), .A(n11455), .ZN(n10622) );
  NAND2_X1 U13320 ( .A1(n10957), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10621) );
  OAI211_X1 U13321 ( .C1(n10655), .C2(n10318), .A(n10622), .B(n10621), .ZN(
        n10623) );
  INV_X1 U13322 ( .A(n10623), .ZN(n10624) );
  NAND2_X1 U13323 ( .A1(n11455), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10641) );
  XNOR2_X2 U13324 ( .A(n10626), .B(n11109), .ZN(n20129) );
  NAND2_X1 U13325 ( .A1(n20129), .A2(n10797), .ZN(n10631) );
  AOI22_X1 U13326 ( .A1(n10957), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n10613), .ZN(n10629) );
  INV_X1 U13327 ( .A(n10655), .ZN(n10627) );
  NAND2_X1 U13328 ( .A1(n10627), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10628) );
  AND2_X1 U13329 ( .A1(n10629), .A2(n10628), .ZN(n10630) );
  NAND2_X1 U13330 ( .A1(n10631), .A2(n10630), .ZN(n12273) );
  NAND2_X1 U13331 ( .A1(n10633), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12252) );
  INV_X2 U13332 ( .A(n10315), .ZN(n10957) );
  NAND2_X1 U13333 ( .A1(n10957), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10636) );
  NAND2_X1 U13334 ( .A1(n10613), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10635) );
  OAI211_X1 U13335 ( .C1(n10655), .C2(n10150), .A(n10636), .B(n10635), .ZN(
        n10637) );
  AOI21_X1 U13336 ( .B1(n20289), .B2(n10797), .A(n10637), .ZN(n10638) );
  OR2_X1 U13337 ( .A1(n12252), .A2(n10638), .ZN(n12253) );
  INV_X1 U13338 ( .A(n10638), .ZN(n12254) );
  OR2_X1 U13339 ( .A1(n12254), .A2(n12792), .ZN(n10639) );
  NAND2_X1 U13340 ( .A1(n12253), .A2(n10639), .ZN(n12272) );
  NAND2_X1 U13341 ( .A1(n12273), .A2(n12272), .ZN(n12579) );
  NAND2_X1 U13342 ( .A1(n20048), .A2(n10797), .ZN(n10650) );
  INV_X1 U13343 ( .A(n10643), .ZN(n10659) );
  INV_X1 U13344 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20866) );
  NAND2_X1 U13345 ( .A1(n20866), .A2(n10644), .ZN(n10645) );
  NAND2_X1 U13346 ( .A1(n10659), .A2(n10645), .ZN(n12917) );
  AOI22_X1 U13347 ( .A1(n12917), .A2(n11099), .B1(n11455), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U13348 ( .A1(n10957), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n10646) );
  OAI211_X1 U13349 ( .C1(n10655), .C2(n12391), .A(n10647), .B(n10646), .ZN(
        n10648) );
  INV_X1 U13350 ( .A(n10648), .ZN(n10649) );
  XNOR2_X1 U13351 ( .A(n10652), .B(n10651), .ZN(n11128) );
  NAND2_X1 U13352 ( .A1(n10613), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10654) );
  NAND2_X1 U13353 ( .A1(n10957), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n10653) );
  OAI211_X1 U13354 ( .C1(n10655), .C2(n12373), .A(n10654), .B(n10653), .ZN(
        n10656) );
  NAND2_X1 U13355 ( .A1(n10656), .A2(n12792), .ZN(n10662) );
  INV_X1 U13356 ( .A(n10657), .ZN(n10667) );
  INV_X1 U13357 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U13358 ( .A1(n10659), .A2(n10658), .ZN(n10660) );
  NAND2_X1 U13359 ( .A1(n10667), .A2(n10660), .ZN(n19997) );
  NAND2_X1 U13360 ( .A1(n19997), .A2(n11099), .ZN(n10661) );
  NAND2_X1 U13361 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  NOR2_X2 U13362 ( .A1(n12599), .A2(n12726), .ZN(n12781) );
  INV_X1 U13363 ( .A(n10665), .ZN(n10675) );
  INV_X1 U13364 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U13365 ( .A1(n10667), .A2(n10666), .ZN(n10668) );
  NAND2_X1 U13366 ( .A1(n10675), .A2(n10668), .ZN(n19889) );
  AOI22_X1 U13367 ( .A1(n19889), .A2(n11099), .B1(n11455), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U13368 ( .A1(n10957), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n10669) );
  OAI211_X1 U13369 ( .C1(n11135), .C2(n10770), .A(n10670), .B(n10669), .ZN(
        n12780) );
  NAND2_X1 U13370 ( .A1(n12781), .A2(n12780), .ZN(n12779) );
  INV_X1 U13371 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10679) );
  INV_X1 U13372 ( .A(n10673), .ZN(n10677) );
  INV_X1 U13373 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U13374 ( .A1(n10675), .A2(n10674), .ZN(n10676) );
  NAND2_X1 U13375 ( .A1(n10677), .A2(n10676), .ZN(n19876) );
  AOI22_X1 U13376 ( .A1(n19876), .A2(n11099), .B1(n11455), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10678) );
  OAI21_X1 U13377 ( .B1(n10315), .B2(n10679), .A(n10678), .ZN(n10680) );
  NAND2_X1 U13378 ( .A1(n10681), .A2(n12983), .ZN(n12982) );
  AOI22_X1 U13379 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13380 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13381 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13382 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10682) );
  NAND4_X1 U13383 ( .A1(n10685), .A2(n10684), .A3(n10683), .A4(n10682), .ZN(
        n10691) );
  AOI22_X1 U13384 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13385 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13386 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13387 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10686) );
  NAND4_X1 U13388 ( .A1(n10689), .A2(n10688), .A3(n10687), .A4(n10686), .ZN(
        n10690) );
  OAI21_X1 U13389 ( .B1(n10691), .B2(n10690), .A(n10797), .ZN(n10695) );
  NAND2_X1 U13390 ( .A1(n10957), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10694) );
  XNOR2_X1 U13391 ( .A(n10697), .B(n10696), .ZN(n19846) );
  NAND2_X1 U13392 ( .A1(n19846), .A2(n11099), .ZN(n10693) );
  NAND2_X1 U13393 ( .A1(n11455), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10692) );
  XOR2_X1 U13394 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10711), .Z(n19837) );
  AOI22_X1 U13395 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13396 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13397 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13398 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10698) );
  NAND4_X1 U13399 ( .A1(n10701), .A2(n10700), .A3(n10699), .A4(n10698), .ZN(
        n10707) );
  AOI22_X1 U13400 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13401 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13402 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U13403 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10702) );
  NAND4_X1 U13404 ( .A1(n10705), .A2(n10704), .A3(n10703), .A4(n10702), .ZN(
        n10706) );
  OR2_X1 U13405 ( .A1(n10707), .A2(n10706), .ZN(n10708) );
  AOI22_X1 U13406 ( .A1(n10797), .A2(n10708), .B1(n11455), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10710) );
  NAND2_X1 U13407 ( .A1(n10957), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10709) );
  OAI211_X1 U13408 ( .C1(n19837), .C2(n12792), .A(n10710), .B(n10709), .ZN(
        n13081) );
  AOI21_X1 U13409 ( .B1(n10712), .B2(n14389), .A(n10728), .ZN(n15847) );
  OR2_X1 U13410 ( .A1(n15847), .A2(n12792), .ZN(n10727) );
  AOI22_X1 U13411 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13412 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13413 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13414 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10713) );
  NAND4_X1 U13415 ( .A1(n10716), .A2(n10715), .A3(n10714), .A4(n10713), .ZN(
        n10722) );
  AOI22_X1 U13416 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13417 ( .A1(n9813), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13418 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13419 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10717) );
  NAND4_X1 U13420 ( .A1(n10720), .A2(n10719), .A3(n10718), .A4(n10717), .ZN(
        n10721) );
  OAI21_X1 U13421 ( .B1(n10722), .B2(n10721), .A(n10797), .ZN(n10725) );
  NAND2_X1 U13422 ( .A1(n10957), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10724) );
  NAND2_X1 U13423 ( .A1(n11455), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10723) );
  AND3_X1 U13424 ( .A1(n10725), .A2(n10724), .A3(n10723), .ZN(n10726) );
  NAND2_X1 U13425 ( .A1(n10727), .A2(n10726), .ZN(n13095) );
  INV_X1 U13426 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13117) );
  OR2_X1 U13427 ( .A1(n10315), .A2(n13117), .ZN(n10730) );
  OAI21_X1 U13428 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10728), .A(
        n10765), .ZN(n15910) );
  AOI22_X1 U13429 ( .A1(n11099), .A2(n15910), .B1(n11455), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10729) );
  NAND2_X1 U13430 ( .A1(n10730), .A2(n10729), .ZN(n13110) );
  AOI22_X1 U13431 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13432 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13433 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13434 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10731) );
  NAND4_X1 U13435 ( .A1(n10734), .A2(n10733), .A3(n10732), .A4(n10731), .ZN(
        n10740) );
  AOI22_X1 U13436 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U13437 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U13438 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13439 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10735) );
  NAND4_X1 U13440 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n10739) );
  OR2_X1 U13441 ( .A1(n10740), .A2(n10739), .ZN(n10741) );
  AND2_X1 U13442 ( .A1(n10797), .A2(n10741), .ZN(n13120) );
  XOR2_X1 U13443 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10772), .Z(
        n13144) );
  AOI22_X1 U13444 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10788), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13445 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13446 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13447 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10742) );
  NAND4_X1 U13448 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10751) );
  AOI22_X1 U13449 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9811), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13450 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13451 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13452 ( .A1(n10459), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10746) );
  NAND4_X1 U13453 ( .A1(n10749), .A2(n10748), .A3(n10747), .A4(n10746), .ZN(
        n10750) );
  OR2_X1 U13454 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  AOI22_X1 U13455 ( .A1(n10797), .A2(n10752), .B1(n11455), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10754) );
  NAND2_X1 U13456 ( .A1(n10957), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n10753) );
  OAI211_X1 U13457 ( .C1(n13144), .C2(n12792), .A(n10754), .B(n10753), .ZN(
        n13133) );
  AOI22_X1 U13458 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13459 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13460 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11022), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13461 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10755) );
  NAND4_X1 U13462 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10764) );
  AOI22_X1 U13463 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9799), .B1(
        n11078), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U13464 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10935), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13465 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13466 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10759) );
  NAND4_X1 U13467 ( .A1(n10762), .A2(n10761), .A3(n10760), .A4(n10759), .ZN(
        n10763) );
  NOR2_X1 U13468 ( .A1(n10764), .A2(n10763), .ZN(n10769) );
  XNOR2_X1 U13469 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10765), .ZN(
        n15898) );
  INV_X1 U13470 ( .A(n15898), .ZN(n10766) );
  AOI22_X1 U13471 ( .A1(n11455), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11099), .B2(n10766), .ZN(n10768) );
  NAND2_X1 U13472 ( .A1(n10957), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n10767) );
  OAI211_X1 U13473 ( .C1(n10770), .C2(n10769), .A(n10768), .B(n10767), .ZN(
        n13123) );
  AND2_X1 U13474 ( .A1(n13133), .A2(n13123), .ZN(n10771) );
  XNOR2_X1 U13475 ( .A(n10787), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15817) );
  AOI22_X1 U13476 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13477 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9811), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13478 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13479 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10773) );
  NAND4_X1 U13480 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        n10782) );
  AOI22_X1 U13481 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13482 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U13483 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13484 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10777) );
  NAND4_X1 U13485 ( .A1(n10780), .A2(n10779), .A3(n10778), .A4(n10777), .ZN(
        n10781) );
  OAI21_X1 U13486 ( .B1(n10782), .B2(n10781), .A(n10797), .ZN(n10785) );
  NAND2_X1 U13487 ( .A1(n10957), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10784) );
  NAND2_X1 U13488 ( .A1(n11455), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10783) );
  NAND3_X1 U13489 ( .A1(n10785), .A2(n10784), .A3(n10783), .ZN(n10786) );
  AOI21_X1 U13490 ( .B1(n15817), .B2(n11099), .A(n10786), .ZN(n14206) );
  XOR2_X1 U13491 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n10806), .Z(
        n15893) );
  INV_X1 U13492 ( .A(n15893), .ZN(n10804) );
  AOI22_X1 U13493 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13494 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13495 ( .A1(n9813), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U13496 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10789) );
  NAND4_X1 U13497 ( .A1(n10792), .A2(n10791), .A3(n10790), .A4(n10789), .ZN(
        n10799) );
  AOI22_X1 U13498 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13499 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13500 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10794) );
  AOI22_X1 U13501 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10793) );
  NAND4_X1 U13502 ( .A1(n10796), .A2(n10795), .A3(n10794), .A4(n10793), .ZN(
        n10798) );
  OAI21_X1 U13503 ( .B1(n10799), .B2(n10798), .A(n10797), .ZN(n10802) );
  NAND2_X1 U13504 ( .A1(n10957), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10801) );
  NAND2_X1 U13505 ( .A1(n11455), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10800) );
  NAND3_X1 U13506 ( .A1(n10802), .A2(n10801), .A3(n10800), .ZN(n10803) );
  AOI21_X1 U13507 ( .B1(n10804), .B2(n11099), .A(n10803), .ZN(n14150) );
  INV_X1 U13508 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14356) );
  XNOR2_X1 U13509 ( .A(n10821), .B(n14356), .ZN(n15809) );
  INV_X1 U13510 ( .A(n15809), .ZN(n10820) );
  AOI22_X1 U13511 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13512 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13513 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13514 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10807) );
  NAND4_X1 U13515 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10816) );
  AOI22_X1 U13516 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13517 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13518 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U13519 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10811) );
  NAND4_X1 U13520 ( .A1(n10814), .A2(n10813), .A3(n10812), .A4(n10811), .ZN(
        n10815) );
  OAI21_X1 U13521 ( .B1(n10816), .B2(n10815), .A(n11096), .ZN(n10818) );
  AOI22_X1 U13522 ( .A1(n10957), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10613), .ZN(n10817) );
  AOI21_X1 U13523 ( .B1(n10818), .B2(n10817), .A(n10612), .ZN(n10819) );
  AOI21_X1 U13524 ( .B1(n10820), .B2(n11099), .A(n10819), .ZN(n14196) );
  NOR2_X2 U13525 ( .A1(n14148), .A2(n14196), .ZN(n14133) );
  AOI21_X1 U13526 ( .B1(n21018), .B2(n10822), .A(n10867), .ZN(n15887) );
  OR2_X1 U13527 ( .A1(n15887), .A2(n12792), .ZN(n10837) );
  AOI22_X1 U13528 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10826) );
  AOI22_X1 U13529 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9812), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13530 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13531 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10823) );
  NAND4_X1 U13532 ( .A1(n10826), .A2(n10825), .A3(n10824), .A4(n10823), .ZN(
        n10832) );
  AOI22_X1 U13533 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13534 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13535 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11079), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13536 ( .A1(n10459), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10827) );
  NAND4_X1 U13537 ( .A1(n10830), .A2(n10829), .A3(n10828), .A4(n10827), .ZN(
        n10831) );
  OR2_X1 U13538 ( .A1(n10832), .A2(n10831), .ZN(n10835) );
  INV_X1 U13539 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14258) );
  INV_X1 U13540 ( .A(n11455), .ZN(n10833) );
  OAI22_X1 U13541 ( .A1(n10315), .A2(n14258), .B1(n10833), .B2(n21018), .ZN(
        n10834) );
  AOI21_X1 U13542 ( .B1(n11096), .B2(n10835), .A(n10834), .ZN(n10836) );
  NAND2_X1 U13543 ( .A1(n10837), .A2(n10836), .ZN(n14135) );
  NAND2_X1 U13544 ( .A1(n14133), .A2(n14135), .ZN(n14134) );
  INV_X1 U13545 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14336) );
  XNOR2_X1 U13546 ( .A(n10867), .B(n14336), .ZN(n15798) );
  NAND2_X1 U13547 ( .A1(n15798), .A2(n11099), .ZN(n10852) );
  AOI22_X1 U13548 ( .A1(n9813), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13549 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13550 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13551 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10838) );
  NAND4_X1 U13552 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n10847) );
  AOI22_X1 U13553 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13554 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13555 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11079), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13556 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10842) );
  NAND4_X1 U13557 ( .A1(n10845), .A2(n10844), .A3(n10843), .A4(n10842), .ZN(
        n10846) );
  NOR2_X1 U13558 ( .A1(n10847), .A2(n10846), .ZN(n10850) );
  AOI21_X1 U13559 ( .B1(n14336), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10848) );
  AOI21_X1 U13560 ( .B1(n10957), .B2(P1_EAX_REG_18__SCAN_IN), .A(n10848), .ZN(
        n10849) );
  OAI21_X1 U13561 ( .B1(n11071), .B2(n10850), .A(n10849), .ZN(n10851) );
  NAND2_X1 U13562 ( .A1(n10852), .A2(n10851), .ZN(n14190) );
  NOR2_X2 U13563 ( .A1(n14134), .A2(n14190), .ZN(n14180) );
  AOI22_X1 U13564 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13565 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11078), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13566 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13567 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10853) );
  NAND4_X1 U13568 ( .A1(n10856), .A2(n10855), .A3(n10854), .A4(n10853), .ZN(
        n10862) );
  AOI22_X1 U13569 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U13570 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13571 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13572 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10857) );
  NAND4_X1 U13573 ( .A1(n10860), .A2(n10859), .A3(n10858), .A4(n10857), .ZN(
        n10861) );
  NOR2_X1 U13574 ( .A1(n10862), .A2(n10861), .ZN(n10866) );
  NAND2_X1 U13575 ( .A1(n10613), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10863) );
  NAND2_X1 U13576 ( .A1(n12792), .A2(n10863), .ZN(n10864) );
  AOI21_X1 U13577 ( .B1(n10957), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10864), .ZN(
        n10865) );
  OAI21_X1 U13578 ( .B1(n11071), .B2(n10866), .A(n10865), .ZN(n10870) );
  OAI21_X1 U13579 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n10868), .A(
        n10889), .ZN(n15879) );
  OR2_X1 U13580 ( .A1(n12792), .A2(n15879), .ZN(n10869) );
  NAND2_X1 U13581 ( .A1(n10870), .A2(n10869), .ZN(n14181) );
  AOI22_X1 U13582 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13583 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11022), .B1(
        n11078), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U13584 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13585 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10872) );
  NAND4_X1 U13586 ( .A1(n10875), .A2(n10874), .A3(n10873), .A4(n10872), .ZN(
        n10881) );
  AOI22_X1 U13587 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n9799), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13588 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11076), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13589 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13590 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10876) );
  NAND4_X1 U13591 ( .A1(n10879), .A2(n10878), .A3(n10877), .A4(n10876), .ZN(
        n10880) );
  NOR2_X1 U13592 ( .A1(n10881), .A2(n10880), .ZN(n10884) );
  INV_X1 U13593 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15872) );
  AOI21_X1 U13594 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15872), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10882) );
  AOI21_X1 U13595 ( .B1(n10957), .B2(P1_EAX_REG_20__SCAN_IN), .A(n10882), .ZN(
        n10883) );
  OAI21_X1 U13596 ( .B1(n11071), .B2(n10884), .A(n10883), .ZN(n10888) );
  INV_X1 U13597 ( .A(n10889), .ZN(n10885) );
  XNOR2_X1 U13598 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n10885), .ZN(
        n15865) );
  INV_X1 U13599 ( .A(n15865), .ZN(n10886) );
  NAND2_X1 U13600 ( .A1(n10886), .A2(n11099), .ZN(n10887) );
  OR2_X1 U13601 ( .A1(n10890), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10891) );
  NAND2_X1 U13602 ( .A1(n10891), .A2(n10927), .ZN(n15864) );
  INV_X1 U13603 ( .A(n15864), .ZN(n10907) );
  AOI22_X1 U13604 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13605 ( .A1(n11022), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10895) );
  AOI22_X1 U13606 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11079), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13607 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10893) );
  NAND4_X1 U13608 ( .A1(n10896), .A2(n10895), .A3(n10894), .A4(n10893), .ZN(
        n10902) );
  AOI22_X1 U13609 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13610 ( .A1(n9813), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13611 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13612 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10897) );
  NAND4_X1 U13613 ( .A1(n10900), .A2(n10899), .A3(n10898), .A4(n10897), .ZN(
        n10901) );
  OR2_X1 U13614 ( .A1(n10902), .A2(n10901), .ZN(n10905) );
  INV_X1 U13615 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U13616 ( .A1(n10613), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10903) );
  OAI211_X1 U13617 ( .C1(n10315), .C2(n14245), .A(n12792), .B(n10903), .ZN(
        n10904) );
  AOI21_X1 U13618 ( .B1(n11096), .B2(n10905), .A(n10904), .ZN(n10906) );
  AOI21_X1 U13619 ( .B1(n10907), .B2(n11099), .A(n10906), .ZN(n14169) );
  AOI22_X1 U13620 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13621 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13622 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13623 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10908) );
  NAND4_X1 U13624 ( .A1(n10911), .A2(n10910), .A3(n10909), .A4(n10908), .ZN(
        n10919) );
  AOI22_X1 U13625 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13626 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13627 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U13628 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10914) );
  NAND4_X1 U13629 ( .A1(n10917), .A2(n10916), .A3(n10915), .A4(n10914), .ZN(
        n10918) );
  NOR2_X1 U13630 ( .A1(n10919), .A2(n10918), .ZN(n10923) );
  NAND2_X1 U13631 ( .A1(n10613), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10920) );
  NAND2_X1 U13632 ( .A1(n12792), .A2(n10920), .ZN(n10921) );
  AOI21_X1 U13633 ( .B1(n10957), .B2(P1_EAX_REG_22__SCAN_IN), .A(n10921), .ZN(
        n10922) );
  OAI21_X1 U13634 ( .B1(n11071), .B2(n10923), .A(n10922), .ZN(n10925) );
  XNOR2_X1 U13635 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n10927), .ZN(
        n15766) );
  NAND2_X1 U13636 ( .A1(n15766), .A2(n11099), .ZN(n10924) );
  INV_X1 U13637 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10926) );
  OR2_X1 U13638 ( .A1(n10928), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10929) );
  NAND2_X1 U13639 ( .A1(n10973), .A2(n10929), .ZN(n15859) );
  AOI22_X1 U13640 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13641 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13642 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13643 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10931) );
  NAND4_X1 U13644 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10941) );
  AOI22_X1 U13645 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13646 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10414), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13647 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13648 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10936) );
  NAND4_X1 U13649 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10940) );
  NOR2_X1 U13650 ( .A1(n10941), .A2(n10940), .ZN(n10969) );
  AOI22_X1 U13651 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13652 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13653 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13654 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10942) );
  NAND4_X1 U13655 ( .A1(n10945), .A2(n10944), .A3(n10943), .A4(n10942), .ZN(
        n10951) );
  AOI22_X1 U13656 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9813), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U13657 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13658 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13659 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10946) );
  NAND4_X1 U13660 ( .A1(n10949), .A2(n10948), .A3(n10947), .A4(n10946), .ZN(
        n10950) );
  NOR2_X1 U13661 ( .A1(n10951), .A2(n10950), .ZN(n10968) );
  XNOR2_X1 U13662 ( .A(n10969), .B(n10968), .ZN(n10954) );
  INV_X1 U13663 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15746) );
  AOI21_X1 U13664 ( .B1(n15746), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10952) );
  AOI21_X1 U13665 ( .B1(n10957), .B2(P1_EAX_REG_23__SCAN_IN), .A(n10952), .ZN(
        n10953) );
  OAI21_X1 U13666 ( .B1(n11071), .B2(n10954), .A(n10953), .ZN(n10955) );
  OAI21_X1 U13667 ( .B1(n15859), .B2(n12792), .A(n10955), .ZN(n14232) );
  NOR2_X2 U13668 ( .A1(n14233), .A2(n14232), .ZN(n14121) );
  XNOR2_X1 U13669 ( .A(n10973), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14328) );
  INV_X1 U13670 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14324) );
  NOR2_X1 U13671 ( .A1(n14324), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10956) );
  AOI211_X1 U13672 ( .C1(n10957), .C2(P1_EAX_REG_24__SCAN_IN), .A(n10612), .B(
        n10956), .ZN(n10972) );
  AOI22_X1 U13673 ( .A1(n10414), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13674 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13675 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13676 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10958) );
  NAND4_X1 U13677 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10967) );
  AOI22_X1 U13678 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U13679 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U13680 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U13681 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10962) );
  NAND4_X1 U13682 ( .A1(n10965), .A2(n10964), .A3(n10963), .A4(n10962), .ZN(
        n10966) );
  OR2_X1 U13683 ( .A1(n10967), .A2(n10966), .ZN(n10990) );
  NOR2_X1 U13684 ( .A1(n10969), .A2(n10968), .ZN(n10991) );
  XOR2_X1 U13685 ( .A(n10990), .B(n10991), .Z(n10970) );
  NAND2_X1 U13686 ( .A1(n10970), .A2(n11096), .ZN(n10971) );
  AOI22_X1 U13687 ( .A1(n14328), .A2(n11099), .B1(n10972), .B2(n10971), .ZN(
        n14123) );
  INV_X1 U13688 ( .A(n10975), .ZN(n10977) );
  INV_X1 U13689 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U13690 ( .A1(n10977), .A2(n10976), .ZN(n10978) );
  NAND2_X1 U13691 ( .A1(n11013), .A2(n10978), .ZN(n14317) );
  AOI22_X1 U13692 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U13693 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U13694 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10979), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U13695 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10980) );
  NAND4_X1 U13696 ( .A1(n10983), .A2(n10982), .A3(n10981), .A4(n10980), .ZN(
        n10989) );
  AOI22_X1 U13697 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U13698 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11078), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U13699 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U13700 ( .A1(n9813), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10984) );
  NAND4_X1 U13701 ( .A1(n10987), .A2(n10986), .A3(n10985), .A4(n10984), .ZN(
        n10988) );
  NOR2_X1 U13702 ( .A1(n10989), .A2(n10988), .ZN(n11009) );
  NAND2_X1 U13703 ( .A1(n10991), .A2(n10990), .ZN(n11008) );
  XNOR2_X1 U13704 ( .A(n11009), .B(n11008), .ZN(n10994) );
  AOI21_X1 U13705 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n10613), .A(
        n10612), .ZN(n10993) );
  NAND2_X1 U13706 ( .A1(n10957), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n10992) );
  OAI211_X1 U13707 ( .C1(n10994), .C2(n11071), .A(n10993), .B(n10992), .ZN(
        n10995) );
  XNOR2_X1 U13708 ( .A(n11013), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14309) );
  INV_X1 U13709 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14305) );
  NOR2_X1 U13710 ( .A1(n14305), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10996) );
  AOI211_X1 U13711 ( .C1(n10957), .C2(P1_EAX_REG_26__SCAN_IN), .A(n11099), .B(
        n10996), .ZN(n11012) );
  AOI22_X1 U13712 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U13713 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U13714 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10997), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U13715 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10998) );
  NAND4_X1 U13716 ( .A1(n11001), .A2(n11000), .A3(n10999), .A4(n10998), .ZN(
        n11007) );
  AOI22_X1 U13717 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U13718 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U13719 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U13720 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11002) );
  NAND4_X1 U13721 ( .A1(n11005), .A2(n11004), .A3(n11003), .A4(n11002), .ZN(
        n11006) );
  OR2_X1 U13722 ( .A1(n11007), .A2(n11006), .ZN(n11029) );
  NOR2_X1 U13723 ( .A1(n11009), .A2(n11008), .ZN(n11030) );
  XOR2_X1 U13724 ( .A(n11029), .B(n11030), .Z(n11010) );
  NAND2_X1 U13725 ( .A1(n11010), .A2(n11096), .ZN(n11011) );
  AOI22_X1 U13726 ( .A1(n14309), .A2(n11099), .B1(n11012), .B2(n11011), .ZN(
        n14099) );
  INV_X1 U13727 ( .A(n11013), .ZN(n11014) );
  NAND2_X1 U13728 ( .A1(n11014), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11016) );
  INV_X1 U13729 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11015) );
  NAND2_X1 U13730 ( .A1(n11016), .A2(n11015), .ZN(n11017) );
  NAND2_X1 U13731 ( .A1(n11052), .A2(n11017), .ZN(n14298) );
  AOI22_X1 U13732 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10788), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U13733 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n9799), .B1(
        n11078), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U13734 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10935), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U13735 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10403), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11018) );
  NAND4_X1 U13736 ( .A1(n11021), .A2(n11020), .A3(n11019), .A4(n11018), .ZN(
        n11028) );
  AOI22_X1 U13737 ( .A1(n11076), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10930), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U13738 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11022), .B1(
        n9813), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11025) );
  AOI22_X1 U13739 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11024) );
  AOI22_X1 U13740 ( .A1(n11079), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11023) );
  NAND4_X1 U13741 ( .A1(n11026), .A2(n11025), .A3(n11024), .A4(n11023), .ZN(
        n11027) );
  NOR2_X1 U13742 ( .A1(n11028), .A2(n11027), .ZN(n11048) );
  NAND2_X1 U13743 ( .A1(n11030), .A2(n11029), .ZN(n11047) );
  XNOR2_X1 U13744 ( .A(n11048), .B(n11047), .ZN(n11033) );
  AOI21_X1 U13745 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n10613), .A(
        n10612), .ZN(n11032) );
  NAND2_X1 U13746 ( .A1(n10957), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n11031) );
  OAI211_X1 U13747 ( .C1(n11033), .C2(n11071), .A(n11032), .B(n11031), .ZN(
        n11034) );
  INV_X1 U13748 ( .A(n11052), .ZN(n11035) );
  XOR2_X1 U13749 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n11035), .Z(
        n14292) );
  INV_X1 U13750 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14288) );
  NOR2_X1 U13751 ( .A1(n14288), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11036) );
  AOI211_X1 U13752 ( .C1(n10957), .C2(P1_EAX_REG_28__SCAN_IN), .A(n10612), .B(
        n11036), .ZN(n11051) );
  AOI22_X1 U13753 ( .A1(n9812), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11040) );
  AOI22_X1 U13754 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U13755 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U13756 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11037) );
  NAND4_X1 U13757 ( .A1(n11040), .A2(n11039), .A3(n11038), .A4(n11037), .ZN(
        n11046) );
  AOI22_X1 U13758 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U13759 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10464), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U13760 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11079), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U13761 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11041) );
  NAND4_X1 U13762 ( .A1(n11044), .A2(n11043), .A3(n11042), .A4(n11041), .ZN(
        n11045) );
  OR2_X1 U13763 ( .A1(n11046), .A2(n11045), .ZN(n11057) );
  NOR2_X1 U13764 ( .A1(n11048), .A2(n11047), .ZN(n11058) );
  XOR2_X1 U13765 ( .A(n11057), .B(n11058), .Z(n11049) );
  NAND2_X1 U13766 ( .A1(n11049), .A2(n11096), .ZN(n11050) );
  AOI22_X1 U13767 ( .A1(n14292), .A2(n11099), .B1(n11051), .B2(n11050), .ZN(
        n13193) );
  NAND2_X1 U13768 ( .A1(n9809), .A2(n9808), .ZN(n14071) );
  NAND2_X1 U13769 ( .A1(n11053), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11460) );
  INV_X1 U13770 ( .A(n11053), .ZN(n11055) );
  INV_X1 U13771 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11054) );
  NAND2_X1 U13772 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  NAND2_X1 U13773 ( .A1(n11460), .A2(n11056), .ZN(n14277) );
  NAND2_X1 U13774 ( .A1(n11058), .A2(n11057), .ZN(n11074) );
  AOI22_X1 U13775 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U13776 ( .A1(n9813), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U13777 ( .A1(n9799), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U13778 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11059) );
  NAND4_X1 U13779 ( .A1(n11062), .A2(n11061), .A3(n11060), .A4(n11059), .ZN(
        n11068) );
  AOI22_X1 U13780 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11078), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U13781 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U13782 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11079), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U13783 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11063) );
  NAND4_X1 U13784 ( .A1(n11066), .A2(n11065), .A3(n11064), .A4(n11063), .ZN(
        n11067) );
  NOR2_X1 U13785 ( .A1(n11068), .A2(n11067), .ZN(n11075) );
  XNOR2_X1 U13786 ( .A(n11074), .B(n11075), .ZN(n11072) );
  INV_X1 U13787 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20207) );
  OAI21_X1 U13788 ( .B1(n20207), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n10613), .ZN(n11070) );
  NAND2_X1 U13789 ( .A1(n10957), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11069) );
  OAI211_X1 U13790 ( .C1(n11072), .C2(n11071), .A(n11070), .B(n11069), .ZN(
        n11073) );
  OAI21_X1 U13791 ( .B1(n14277), .B2(n12792), .A(n11073), .ZN(n14072) );
  NOR2_X2 U13792 ( .A1(n14071), .A2(n14072), .ZN(n11454) );
  XNOR2_X1 U13794 ( .A(n11460), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14060) );
  NOR2_X1 U13795 ( .A1(n11075), .A2(n11074), .ZN(n11093) );
  AOI22_X1 U13796 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U13797 ( .A1(n11078), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9799), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U13798 ( .A1(n10912), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10892), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U13799 ( .A1(n10458), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11079), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11080) );
  NAND4_X1 U13800 ( .A1(n11083), .A2(n11082), .A3(n11081), .A4(n11080), .ZN(
        n11091) );
  AOI22_X1 U13801 ( .A1(n9813), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U13802 ( .A1(n10788), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10559), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U13803 ( .A1(n10930), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10459), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U13804 ( .A1(n9811), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11084), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11086) );
  NAND4_X1 U13805 ( .A1(n11089), .A2(n11088), .A3(n11087), .A4(n11086), .ZN(
        n11090) );
  NOR2_X1 U13806 ( .A1(n11091), .A2(n11090), .ZN(n11092) );
  XNOR2_X1 U13807 ( .A(n11093), .B(n11092), .ZN(n11097) );
  INV_X1 U13808 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n11446) );
  NOR2_X1 U13809 ( .A1(n20207), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11094) );
  OAI22_X1 U13810 ( .A1(n10315), .A2(n11446), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11094), .ZN(n11095) );
  AOI21_X1 U13811 ( .B1(n11097), .B2(n11096), .A(n11095), .ZN(n11098) );
  AOI21_X1 U13812 ( .B1(n14060), .B2(n11099), .A(n11098), .ZN(n11453) );
  INV_X1 U13813 ( .A(n11453), .ZN(n11100) );
  XNOR2_X2 U13814 ( .A(n14070), .B(n11100), .ZN(n11468) );
  NAND3_X1 U13815 ( .A1(n10081), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16037) );
  INV_X1 U13816 ( .A(n16037), .ZN(n11101) );
  NOR2_X2 U13817 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20496) );
  NAND2_X1 U13818 ( .A1(n11468), .A2(n19993), .ZN(n11259) );
  NAND2_X1 U13819 ( .A1(n12325), .A2(n10434), .ZN(n11190) );
  NAND2_X1 U13820 ( .A1(n11105), .A2(n11111), .ZN(n11121) );
  XNOR2_X1 U13821 ( .A(n11121), .B(n11120), .ZN(n11103) );
  NAND2_X1 U13822 ( .A1(n20051), .A2(n20074), .ZN(n11110) );
  INV_X1 U13823 ( .A(n11110), .ZN(n11102) );
  AOI21_X1 U13824 ( .B1(n11103), .B2(n11889), .A(n11102), .ZN(n11104) );
  OAI21_X1 U13825 ( .B1(n11111), .B2(n11105), .A(n11121), .ZN(n11106) );
  OAI211_X1 U13826 ( .C1(n11106), .C2(n20729), .A(n20070), .B(n12325), .ZN(
        n11107) );
  INV_X1 U13827 ( .A(n11107), .ZN(n11108) );
  OAI21_X1 U13828 ( .B1(n20729), .B2(n11111), .A(n11110), .ZN(n11112) );
  INV_X1 U13829 ( .A(n11112), .ZN(n11113) );
  NAND2_X1 U13830 ( .A1(n12258), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12257) );
  XNOR2_X1 U13831 ( .A(n11115), .B(n12257), .ZN(n12275) );
  NAND2_X1 U13832 ( .A1(n12275), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12276) );
  INV_X1 U13833 ( .A(n11115), .ZN(n11116) );
  OR2_X1 U13834 ( .A1(n12257), .A2(n11116), .ZN(n11117) );
  NAND2_X2 U13835 ( .A1(n12276), .A2(n11117), .ZN(n11118) );
  INV_X1 U13836 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20036) );
  NAND2_X1 U13837 ( .A1(n11118), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11119) );
  INV_X1 U13838 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20019) );
  NAND2_X1 U13839 ( .A1(n20048), .A2(n9991), .ZN(n11125) );
  NAND2_X1 U13840 ( .A1(n11121), .A2(n11120), .ZN(n11139) );
  INV_X1 U13841 ( .A(n11137), .ZN(n11122) );
  XNOR2_X1 U13842 ( .A(n11139), .B(n11122), .ZN(n11123) );
  NAND2_X1 U13843 ( .A1(n11123), .A2(n11889), .ZN(n11124) );
  NAND2_X1 U13844 ( .A1(n11125), .A2(n11124), .ZN(n12635) );
  NAND2_X1 U13845 ( .A1(n11126), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11127) );
  INV_X1 U13846 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20010) );
  NAND2_X1 U13847 ( .A1(n11128), .A2(n9991), .ZN(n11132) );
  NAND2_X1 U13848 ( .A1(n11139), .A2(n11137), .ZN(n11129) );
  XNOR2_X1 U13849 ( .A(n11129), .B(n11136), .ZN(n11130) );
  NAND2_X1 U13850 ( .A1(n11130), .A2(n11889), .ZN(n11131) );
  NAND2_X1 U13851 ( .A1(n11132), .A2(n11131), .ZN(n19989) );
  NAND2_X1 U13852 ( .A1(n19990), .A2(n19989), .ZN(n19988) );
  NAND2_X1 U13853 ( .A1(n11133), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11134) );
  AND2_X1 U13854 ( .A1(n11137), .A2(n11136), .ZN(n11138) );
  NAND2_X1 U13855 ( .A1(n11139), .A2(n11138), .ZN(n11145) );
  XNOR2_X1 U13856 ( .A(n11145), .B(n11146), .ZN(n11140) );
  NAND2_X1 U13857 ( .A1(n11140), .A2(n11889), .ZN(n11141) );
  INV_X1 U13858 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13018) );
  XNOR2_X1 U13859 ( .A(n11142), .B(n13018), .ZN(n15921) );
  NAND3_X1 U13860 ( .A1(n11164), .A2(n9991), .A3(n11144), .ZN(n11150) );
  INV_X1 U13861 ( .A(n11145), .ZN(n11147) );
  NAND2_X1 U13862 ( .A1(n11147), .A2(n11146), .ZN(n11153) );
  XNOR2_X1 U13863 ( .A(n11153), .B(n11154), .ZN(n11148) );
  NAND2_X1 U13864 ( .A1(n11148), .A2(n11889), .ZN(n11149) );
  NAND2_X1 U13865 ( .A1(n11150), .A2(n11149), .ZN(n13015) );
  OR2_X1 U13866 ( .A1(n13015), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11151) );
  NAND2_X1 U13867 ( .A1(n11152), .A2(n9991), .ZN(n11159) );
  INV_X1 U13868 ( .A(n11153), .ZN(n11155) );
  NAND2_X1 U13869 ( .A1(n11155), .A2(n11154), .ZN(n11166) );
  XNOR2_X1 U13870 ( .A(n11166), .B(n11156), .ZN(n11157) );
  NAND2_X1 U13871 ( .A1(n11157), .A2(n11889), .ZN(n11158) );
  NAND2_X1 U13872 ( .A1(n11159), .A2(n11158), .ZN(n11160) );
  OR2_X1 U13873 ( .A1(n11160), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15912) );
  NAND2_X1 U13874 ( .A1(n11160), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15911) );
  NAND2_X1 U13875 ( .A1(n11161), .A2(n15911), .ZN(n13088) );
  AND2_X1 U13876 ( .A1(n11162), .A2(n9991), .ZN(n11163) );
  NAND2_X4 U13877 ( .A1(n11164), .A2(n11163), .ZN(n11179) );
  OR3_X1 U13878 ( .A1(n11166), .A2(n11165), .A3(n20729), .ZN(n11167) );
  NAND2_X1 U13879 ( .A1(n11179), .A2(n11167), .ZN(n13086) );
  OR2_X1 U13880 ( .A1(n13086), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11168) );
  NAND2_X1 U13881 ( .A1(n13086), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11169) );
  INV_X1 U13882 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16010) );
  NAND2_X1 U13883 ( .A1(n11179), .A2(n16010), .ZN(n11171) );
  INV_X1 U13884 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15980) );
  NAND2_X1 U13885 ( .A1(n11179), .A2(n15980), .ZN(n11172) );
  INV_X1 U13886 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U13887 ( .A1(n11179), .A2(n11180), .ZN(n14374) );
  NAND2_X1 U13888 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11173) );
  NAND2_X1 U13889 ( .A1(n11179), .A2(n11173), .ZN(n14372) );
  NAND2_X1 U13890 ( .A1(n14374), .A2(n14372), .ZN(n11174) );
  INV_X1 U13891 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20982) );
  NAND2_X1 U13892 ( .A1(n11179), .A2(n20982), .ZN(n11175) );
  NAND2_X1 U13893 ( .A1(n14362), .A2(n11175), .ZN(n14343) );
  NAND2_X1 U13894 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11176) );
  AND2_X1 U13895 ( .A1(n11179), .A2(n11176), .ZN(n11178) );
  OR2_X1 U13896 ( .A1(n11179), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15882) );
  NAND2_X1 U13897 ( .A1(n11179), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11177) );
  INV_X1 U13898 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15961) );
  NAND2_X1 U13899 ( .A1(n15957), .A2(n15961), .ZN(n14349) );
  OAI21_X1 U13900 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14349), .A(
        n11189), .ZN(n11182) );
  NOR2_X1 U13901 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14370) );
  AND2_X1 U13902 ( .A1(n14370), .A2(n11180), .ZN(n11181) );
  NAND2_X1 U13903 ( .A1(n11182), .A2(n14342), .ZN(n11184) );
  OR2_X1 U13904 ( .A1(n11179), .A2(n20982), .ZN(n11183) );
  NAND2_X1 U13905 ( .A1(n14360), .A2(n11183), .ZN(n14345) );
  XNOR2_X1 U13906 ( .A(n11179), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13164) );
  NAND3_X1 U13907 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14451) );
  INV_X1 U13908 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11186) );
  INV_X1 U13909 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15730) );
  NAND2_X1 U13910 ( .A1(n11186), .A2(n15730), .ZN(n11187) );
  NAND3_X1 U13911 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14281) );
  INV_X1 U13912 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21047) );
  INV_X1 U13913 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14457) );
  INV_X1 U13914 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n20954) );
  NAND3_X1 U13915 ( .A1(n21047), .A2(n14457), .A3(n20954), .ZN(n14282) );
  AND2_X1 U13916 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14411) );
  NOR2_X1 U13917 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14412) );
  INV_X1 U13918 ( .A(n11417), .ZN(n11249) );
  XNOR2_X1 U13919 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U13920 ( .A1(n20489), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11210) );
  NAND2_X1 U13921 ( .A1(n11206), .A2(n11205), .ZN(n11192) );
  NAND2_X1 U13922 ( .A1(n20457), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11191) );
  NAND2_X1 U13923 ( .A1(n11192), .A2(n11191), .ZN(n11203) );
  XNOR2_X1 U13924 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U13925 ( .A1(n11203), .A2(n11202), .ZN(n11194) );
  NAND2_X1 U13926 ( .A1(n20375), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11193) );
  NAND2_X1 U13927 ( .A1(n11194), .A2(n11193), .ZN(n11201) );
  XNOR2_X1 U13928 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11200) );
  NAND2_X1 U13929 ( .A1(n11201), .A2(n11200), .ZN(n11196) );
  NAND2_X1 U13930 ( .A1(n20380), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11195) );
  NOR2_X1 U13931 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12373), .ZN(
        n11197) );
  NAND2_X1 U13932 ( .A1(n11267), .A2(n11207), .ZN(n11243) );
  INV_X1 U13933 ( .A(n11212), .ZN(n11231) );
  XNOR2_X1 U13934 ( .A(n11201), .B(n11200), .ZN(n11264) );
  XNOR2_X1 U13935 ( .A(n11203), .B(n11202), .ZN(n11262) );
  INV_X1 U13936 ( .A(n11224), .ZN(n11227) );
  OAI21_X1 U13937 ( .B1(n20051), .B2(n12325), .A(n20066), .ZN(n11226) );
  INV_X1 U13938 ( .A(n11262), .ZN(n11204) );
  OAI21_X1 U13939 ( .B1(n11204), .B2(n11228), .A(n11226), .ZN(n11223) );
  XNOR2_X1 U13940 ( .A(n11206), .B(n11205), .ZN(n11263) );
  NAND2_X1 U13941 ( .A1(n11207), .A2(n10434), .ZN(n11209) );
  NAND2_X1 U13942 ( .A1(n20083), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11208) );
  NOR2_X1 U13943 ( .A1(n11263), .A2(n11218), .ZN(n11217) );
  OAI21_X1 U13944 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20489), .A(
        n11210), .ZN(n11213) );
  INV_X1 U13945 ( .A(n11213), .ZN(n11211) );
  OAI211_X1 U13946 ( .C1(n20051), .C2(n10381), .A(n11226), .B(n11211), .ZN(
        n11216) );
  OAI21_X1 U13947 ( .B1(n11214), .B2(n11213), .A(n11212), .ZN(n11215) );
  NAND2_X1 U13948 ( .A1(n11216), .A2(n11215), .ZN(n11219) );
  NAND2_X1 U13949 ( .A1(n11217), .A2(n11219), .ZN(n11222) );
  INV_X1 U13950 ( .A(n11218), .ZN(n11220) );
  OAI211_X1 U13951 ( .C1(n11220), .C2(n11219), .A(n11263), .B(n11235), .ZN(
        n11221) );
  OAI211_X1 U13952 ( .C1(n11224), .C2(n11223), .A(n11222), .B(n11221), .ZN(
        n11225) );
  OAI21_X1 U13953 ( .B1(n11227), .B2(n11226), .A(n11225), .ZN(n11230) );
  NAND2_X1 U13954 ( .A1(n11228), .A2(n11264), .ZN(n11229) );
  AOI22_X1 U13955 ( .A1(n11231), .A2(n11264), .B1(n11230), .B2(n11229), .ZN(
        n11240) );
  INV_X1 U13956 ( .A(n11265), .ZN(n11234) );
  NOR2_X1 U13957 ( .A1(n11237), .A2(n11234), .ZN(n11239) );
  NAND3_X1 U13958 ( .A1(n11237), .A2(n11236), .A3(n11265), .ZN(n11238) );
  OAI21_X1 U13959 ( .B1(n11240), .B2(n11239), .A(n11238), .ZN(n11241) );
  AOI21_X1 U13960 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n10081), .A(
        n11241), .ZN(n11242) );
  NAND2_X1 U13961 ( .A1(n20070), .A2(n20074), .ZN(n11246) );
  AOI21_X1 U13962 ( .B1(n15667), .B2(n20051), .A(n11246), .ZN(n11247) );
  NOR2_X1 U13963 ( .A1(n10381), .A2(n19811), .ZN(n11248) );
  INV_X1 U13964 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11459) );
  OR2_X1 U13965 ( .A1(n11254), .A2(n20496), .ZN(n20725) );
  AND2_X1 U13966 ( .A1(n20725), .A2(n10081), .ZN(n11250) );
  NAND2_X1 U13967 ( .A1(n10081), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11252) );
  NAND2_X1 U13968 ( .A1(n20207), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11251) );
  AND2_X1 U13969 ( .A1(n11252), .A2(n11251), .ZN(n12256) );
  INV_X1 U13970 ( .A(n12256), .ZN(n11253) );
  NAND2_X1 U13971 ( .A1(n14060), .A2(n15899), .ZN(n11255) );
  NAND2_X1 U13972 ( .A1(n20033), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n11409) );
  OAI211_X1 U13973 ( .C1(n11459), .C2(n15871), .A(n11255), .B(n11409), .ZN(
        n11256) );
  INV_X1 U13974 ( .A(n11256), .ZN(n11257) );
  NAND3_X1 U13975 ( .A1(n11259), .A2(n11258), .A3(n11257), .ZN(P1_U2969) );
  OR2_X1 U13976 ( .A1(n11260), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n12344) );
  INV_X1 U13977 ( .A(n12344), .ZN(n15720) );
  NAND2_X1 U13978 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20726) );
  OAI21_X1 U13979 ( .B1(n10434), .B2(n15720), .A(n20726), .ZN(n12803) );
  OAI211_X1 U13980 ( .C1(n12342), .C2(n12803), .A(n11286), .B(n11433), .ZN(
        n11261) );
  NAND2_X1 U13981 ( .A1(n15694), .A2(n11261), .ZN(n11270) );
  NOR4_X1 U13982 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n11266) );
  NOR2_X1 U13983 ( .A1(n11267), .A2(n11266), .ZN(n11833) );
  NAND2_X1 U13984 ( .A1(n11833), .A2(n20726), .ZN(n11422) );
  AND2_X1 U13985 ( .A1(n10434), .A2(n12344), .ZN(n11268) );
  OR2_X1 U13986 ( .A1(n11422), .A2(n11268), .ZN(n11269) );
  MUX2_X1 U13987 ( .A(n11270), .B(n11269), .S(n10431), .Z(n11277) );
  INV_X1 U13988 ( .A(n11271), .ZN(n11835) );
  AND2_X1 U13989 ( .A1(n11288), .A2(n11286), .ZN(n11272) );
  NAND2_X1 U13990 ( .A1(n11273), .A2(n11272), .ZN(n11283) );
  NAND2_X1 U13991 ( .A1(n11283), .A2(n15680), .ZN(n11274) );
  NAND2_X1 U13992 ( .A1(n11835), .A2(n11274), .ZN(n12339) );
  INV_X1 U13993 ( .A(n11288), .ZN(n11275) );
  NAND2_X1 U13994 ( .A1(n11842), .A2(n11275), .ZN(n11276) );
  NAND3_X1 U13995 ( .A1(n11277), .A2(n12339), .A3(n11276), .ZN(n11278) );
  AND2_X1 U13996 ( .A1(n11271), .A2(n10434), .ZN(n15669) );
  INV_X1 U13997 ( .A(n12380), .ZN(n12330) );
  NAND2_X1 U13998 ( .A1(n10381), .A2(n20051), .ZN(n11279) );
  NAND3_X1 U13999 ( .A1(n12330), .A2(n11280), .A3(n11279), .ZN(n11281) );
  NAND2_X1 U14000 ( .A1(n11281), .A2(n10434), .ZN(n11282) );
  AND3_X1 U14001 ( .A1(n11284), .A2(n9886), .A3(n11283), .ZN(n12328) );
  OAI211_X1 U14002 ( .C1(n12326), .C2(n11286), .A(n12328), .B(n11285), .ZN(
        n11287) );
  NAND2_X1 U14003 ( .A1(n11408), .A2(n11287), .ZN(n14464) );
  NOR2_X1 U14004 ( .A1(n11289), .A2(n11288), .ZN(n12334) );
  NAND2_X1 U14005 ( .A1(n11408), .A2(n12334), .ZN(n20024) );
  NAND2_X1 U14006 ( .A1(n20002), .A2(n11416), .ZN(n14506) );
  INV_X1 U14007 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20023) );
  INV_X1 U14008 ( .A(n14464), .ZN(n14479) );
  NAND2_X1 U14009 ( .A1(n20023), .A2(n14479), .ZN(n11290) );
  NAND2_X1 U14010 ( .A1(n13162), .A2(n20000), .ZN(n16012) );
  INV_X1 U14011 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15874) );
  NOR2_X1 U14012 ( .A1(n15730), .A2(n15874), .ZN(n14469) );
  INV_X1 U14013 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11362) );
  NAND4_X1 U14014 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13171) );
  NOR2_X1 U14015 ( .A1(n11362), .A2(n13171), .ZN(n14453) );
  AND3_X1 U14016 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15993) );
  AND3_X1 U14017 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15993), .ZN(n14488) );
  NAND2_X1 U14018 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14488), .ZN(
        n14490) );
  INV_X1 U14019 ( .A(n14490), .ZN(n14493) );
  AND2_X1 U14020 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14493), .ZN(
        n14477) );
  NAND2_X1 U14021 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11301) );
  AOI21_X1 U14022 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11299) );
  NOR3_X1 U14023 ( .A1(n11301), .A2(n13018), .A3(n11299), .ZN(n13019) );
  AND2_X1 U14024 ( .A1(n14477), .A2(n13019), .ZN(n14466) );
  NAND3_X1 U14025 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14453), .A3(
        n14466), .ZN(n14467) );
  INV_X1 U14026 ( .A(n11301), .ZN(n20005) );
  NAND3_X1 U14027 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20005), .ZN(n13020) );
  NOR2_X1 U14028 ( .A1(n13018), .A2(n13020), .ZN(n15990) );
  NAND2_X1 U14029 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14477), .ZN(
        n14455) );
  INV_X1 U14030 ( .A(n14455), .ZN(n13159) );
  AND2_X1 U14031 ( .A1(n15990), .A2(n13159), .ZN(n15970) );
  NAND2_X1 U14032 ( .A1(n15970), .A2(n14453), .ZN(n14468) );
  INV_X1 U14033 ( .A(n14468), .ZN(n15938) );
  OAI21_X1 U14034 ( .B1(n20001), .B2(n15938), .A(n20000), .ZN(n11291) );
  AOI21_X1 U14035 ( .B1(n14491), .B2(n14467), .A(n11291), .ZN(n15729) );
  INV_X1 U14036 ( .A(n16012), .ZN(n14422) );
  AOI21_X1 U14037 ( .B1(n14469), .B2(n15729), .A(n14422), .ZN(n15703) );
  NAND2_X1 U14038 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14474) );
  OR2_X1 U14039 ( .A1(n15703), .A2(n14474), .ZN(n11292) );
  NAND2_X1 U14040 ( .A1(n16012), .A2(n11292), .ZN(n15932) );
  NAND2_X1 U14041 ( .A1(n14491), .A2(n21047), .ZN(n11293) );
  NAND2_X1 U14042 ( .A1(n15932), .A2(n11293), .ZN(n14456) );
  INV_X1 U14043 ( .A(n14281), .ZN(n11294) );
  NOR2_X1 U14044 ( .A1(n13162), .A2(n11294), .ZN(n11295) );
  NOR2_X1 U14045 ( .A1(n14456), .A2(n11295), .ZN(n14439) );
  NAND2_X1 U14046 ( .A1(n14439), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14436) );
  INV_X1 U14047 ( .A(n14411), .ZN(n14401) );
  OR2_X1 U14048 ( .A1(n14436), .A2(n14401), .ZN(n11296) );
  NAND2_X1 U14049 ( .A1(n11296), .A2(n16012), .ZN(n14405) );
  OAI21_X1 U14050 ( .B1(n13162), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11297) );
  INV_X1 U14051 ( .A(n11297), .ZN(n11298) );
  NAND2_X1 U14052 ( .A1(n14405), .A2(n11298), .ZN(n14394) );
  INV_X1 U14053 ( .A(n14394), .ZN(n11419) );
  INV_X1 U14054 ( .A(n11299), .ZN(n19999) );
  NAND2_X1 U14055 ( .A1(n15969), .A2(n20023), .ZN(n20034) );
  NAND3_X1 U14056 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14487), .ZN(n13021) );
  INV_X1 U14057 ( .A(n13021), .ZN(n11300) );
  NAND2_X1 U14058 ( .A1(n13159), .A2(n16014), .ZN(n15942) );
  NAND3_X1 U14059 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11302) );
  NOR2_X1 U14060 ( .A1(n14451), .A2(n11302), .ZN(n11303) );
  NAND2_X1 U14061 ( .A1(n14453), .A2(n11303), .ZN(n11304) );
  NOR2_X1 U14062 ( .A1(n15942), .A2(n11304), .ZN(n14444) );
  AND2_X1 U14063 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U14064 ( .A1(n14444), .A2(n11305), .ZN(n14410) );
  NAND2_X1 U14065 ( .A1(n14411), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11306) );
  OR2_X1 U14066 ( .A1(n14410), .A2(n11306), .ZN(n14396) );
  INV_X1 U14067 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14395) );
  MUX2_X1 U14068 ( .A(n11396), .B(n11371), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n11307) );
  INV_X1 U14069 ( .A(n11307), .ZN(n11310) );
  NAND2_X1 U14070 ( .A1(n11371), .A2(n11313), .ZN(n11346) );
  NAND3_X1 U14071 ( .A1(n11313), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n11378), .ZN(n11308) );
  AND2_X1 U14072 ( .A1(n11346), .A2(n11308), .ZN(n11309) );
  NAND2_X1 U14073 ( .A1(n11397), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11312) );
  INV_X1 U14074 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12558) );
  NAND2_X1 U14075 ( .A1(n11378), .A2(n12558), .ZN(n11311) );
  NAND2_X1 U14076 ( .A1(n11312), .A2(n11311), .ZN(n12263) );
  INV_X1 U14077 ( .A(n11314), .ZN(n11315) );
  MUX2_X1 U14078 ( .A(n11396), .B(n11371), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11316) );
  INV_X1 U14079 ( .A(n11316), .ZN(n11319) );
  NAND2_X1 U14080 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11313), .ZN(
        n11317) );
  AND2_X1 U14081 ( .A1(n11346), .A2(n11317), .ZN(n11318) );
  NAND2_X1 U14082 ( .A1(n11319), .A2(n11318), .ZN(n12577) );
  MUX2_X1 U14083 ( .A(n11382), .B(n11378), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11321) );
  NAND2_X1 U14084 ( .A1(n12262), .A2(n20019), .ZN(n11320) );
  NAND2_X1 U14085 ( .A1(n11321), .A2(n11320), .ZN(n12596) );
  MUX2_X1 U14086 ( .A(n11396), .B(n11371), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11323) );
  OAI21_X1 U14087 ( .B1(n11837), .B2(n20010), .A(n11346), .ZN(n11322) );
  NOR2_X1 U14088 ( .A1(n11323), .A2(n11322), .ZN(n12756) );
  INV_X1 U14089 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19918) );
  NAND2_X1 U14090 ( .A1(n11393), .A2(n19918), .ZN(n11326) );
  NAND2_X1 U14091 ( .A1(n11378), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11324) );
  OAI211_X1 U14092 ( .C1(n11313), .C2(P1_EBX_REG_5__SCAN_IN), .A(n11397), .B(
        n11324), .ZN(n11325) );
  MUX2_X1 U14093 ( .A(n11396), .B(n11371), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11327) );
  INV_X1 U14094 ( .A(n11327), .ZN(n11330) );
  NAND2_X1 U14095 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11313), .ZN(
        n11328) );
  AND2_X1 U14096 ( .A1(n11346), .A2(n11328), .ZN(n11329) );
  NAND2_X1 U14097 ( .A1(n11330), .A2(n11329), .ZN(n12979) );
  INV_X1 U14098 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19864) );
  NAND2_X1 U14099 ( .A1(n11393), .A2(n19864), .ZN(n11333) );
  NAND2_X1 U14100 ( .A1(n11378), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11331) );
  OAI211_X1 U14101 ( .C1(n11313), .C2(P1_EBX_REG_7__SCAN_IN), .A(n11397), .B(
        n11331), .ZN(n11332) );
  NAND2_X1 U14102 ( .A1(n11333), .A2(n11332), .ZN(n12988) );
  MUX2_X1 U14103 ( .A(n11396), .B(n11371), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11336) );
  NAND2_X1 U14104 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n11313), .ZN(
        n11334) );
  NAND2_X1 U14105 ( .A1(n11346), .A2(n11334), .ZN(n11335) );
  INV_X1 U14106 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19911) );
  NAND2_X1 U14107 ( .A1(n11393), .A2(n19911), .ZN(n11339) );
  NAND2_X1 U14108 ( .A1(n11378), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11337) );
  OAI211_X1 U14109 ( .C1(n11313), .C2(P1_EBX_REG_9__SCAN_IN), .A(n11397), .B(
        n11337), .ZN(n11338) );
  NAND2_X1 U14110 ( .A1(n11339), .A2(n11338), .ZN(n16000) );
  INV_X1 U14111 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15841) );
  NAND2_X1 U14112 ( .A1(n11396), .A2(n15841), .ZN(n11342) );
  INV_X1 U14113 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14385) );
  NAND2_X1 U14114 ( .A1(n11397), .A2(n14385), .ZN(n11340) );
  OAI211_X1 U14115 ( .C1(n11313), .C2(P1_EBX_REG_10__SCAN_IN), .A(n11340), .B(
        n11349), .ZN(n11341) );
  NAND2_X1 U14116 ( .A1(n11342), .A2(n11341), .ZN(n13096) );
  MUX2_X1 U14117 ( .A(n11382), .B(n11378), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11344) );
  INV_X1 U14118 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U14119 ( .A1(n15988), .A2(n12262), .ZN(n11343) );
  NAND2_X1 U14120 ( .A1(n11344), .A2(n11343), .ZN(n13113) );
  MUX2_X1 U14121 ( .A(n11396), .B(n11371), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11348) );
  NAND2_X1 U14122 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n11313), .ZN(
        n11345) );
  NAND2_X1 U14123 ( .A1(n11346), .A2(n11345), .ZN(n11347) );
  NOR2_X1 U14124 ( .A1(n11348), .A2(n11347), .ZN(n13129) );
  MUX2_X1 U14125 ( .A(n11393), .B(n9998), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11351) );
  NOR2_X1 U14126 ( .A1(n13214), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11350) );
  NOR2_X1 U14127 ( .A1(n11351), .A2(n11350), .ZN(n13138) );
  INV_X1 U14128 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15815) );
  NAND2_X1 U14129 ( .A1(n11396), .A2(n15815), .ZN(n11354) );
  NAND2_X1 U14130 ( .A1(n11397), .A2(n20982), .ZN(n11352) );
  OAI211_X1 U14131 ( .C1(n11313), .C2(P1_EBX_REG_14__SCAN_IN), .A(n11352), .B(
        n11378), .ZN(n11353) );
  NAND2_X1 U14132 ( .A1(n11354), .A2(n11353), .ZN(n14207) );
  MUX2_X1 U14133 ( .A(n11382), .B(n11378), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11356) );
  NAND2_X1 U14134 ( .A1(n12262), .A2(n15961), .ZN(n11355) );
  NAND2_X1 U14135 ( .A1(n11356), .A2(n11355), .ZN(n14151) );
  INV_X1 U14136 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15812) );
  NAND2_X1 U14137 ( .A1(n11396), .A2(n15812), .ZN(n11359) );
  NAND2_X1 U14138 ( .A1(n11397), .A2(n15957), .ZN(n11357) );
  OAI211_X1 U14139 ( .C1(n11313), .C2(P1_EBX_REG_16__SCAN_IN), .A(n11357), .B(
        n11378), .ZN(n11358) );
  NAND2_X1 U14140 ( .A1(n11359), .A2(n11358), .ZN(n14198) );
  MUX2_X1 U14141 ( .A(n11382), .B(n11378), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11361) );
  INV_X1 U14142 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15943) );
  NAND2_X1 U14143 ( .A1(n12262), .A2(n15943), .ZN(n11360) );
  NAND2_X1 U14144 ( .A1(n11361), .A2(n11360), .ZN(n14142) );
  INV_X1 U14145 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15794) );
  NAND2_X1 U14146 ( .A1(n11396), .A2(n15794), .ZN(n11365) );
  NAND2_X1 U14147 ( .A1(n11397), .A2(n11362), .ZN(n11363) );
  OAI211_X1 U14148 ( .C1(n11313), .C2(P1_EBX_REG_18__SCAN_IN), .A(n11363), .B(
        n11349), .ZN(n11364) );
  AND2_X1 U14149 ( .A1(n11365), .A2(n11364), .ZN(n13167) );
  MUX2_X1 U14150 ( .A(n11382), .B(n11378), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11368) );
  NAND2_X1 U14151 ( .A1(n12262), .A2(n15874), .ZN(n11367) );
  NAND2_X1 U14152 ( .A1(n11368), .A2(n11367), .ZN(n14184) );
  MUX2_X1 U14153 ( .A(n11382), .B(n11349), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11370) );
  NAND2_X1 U14154 ( .A1(n12262), .A2(n11186), .ZN(n11369) );
  AND2_X1 U14155 ( .A1(n11370), .A2(n11369), .ZN(n14170) );
  MUX2_X1 U14156 ( .A(n11396), .B(n11371), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n11372) );
  INV_X1 U14157 ( .A(n11372), .ZN(n11374) );
  NAND2_X1 U14158 ( .A1(n11313), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11373) );
  NAND2_X1 U14159 ( .A1(n11374), .A2(n11373), .ZN(n14178) );
  INV_X1 U14160 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15769) );
  NAND2_X1 U14161 ( .A1(n11396), .A2(n15769), .ZN(n11377) );
  INV_X1 U14162 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14447) );
  NAND2_X1 U14163 ( .A1(n11397), .A2(n14447), .ZN(n11375) );
  OAI211_X1 U14164 ( .C1(n11313), .C2(P1_EBX_REG_22__SCAN_IN), .A(n11375), .B(
        n11378), .ZN(n11376) );
  NAND2_X1 U14165 ( .A1(n11377), .A2(n11376), .ZN(n14165) );
  INV_X1 U14166 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15852) );
  NAND2_X1 U14167 ( .A1(n11393), .A2(n15852), .ZN(n11381) );
  NAND2_X1 U14168 ( .A1(n11378), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11379) );
  OAI211_X1 U14169 ( .C1(n11313), .C2(P1_EBX_REG_23__SCAN_IN), .A(n11397), .B(
        n11379), .ZN(n11380) );
  NAND2_X1 U14170 ( .A1(n11381), .A2(n11380), .ZN(n15748) );
  MUX2_X1 U14171 ( .A(n11382), .B(n11378), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11384) );
  NAND2_X1 U14172 ( .A1(n12262), .A2(n20954), .ZN(n11383) );
  NAND2_X1 U14173 ( .A1(n11384), .A2(n11383), .ZN(n14109) );
  INV_X1 U14174 ( .A(n14109), .ZN(n11388) );
  INV_X1 U14175 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14126) );
  NAND2_X1 U14176 ( .A1(n11396), .A2(n14126), .ZN(n11387) );
  NAND2_X1 U14177 ( .A1(n11397), .A2(n14457), .ZN(n11385) );
  OAI211_X1 U14178 ( .C1(n11313), .C2(P1_EBX_REG_24__SCAN_IN), .A(n11385), .B(
        n11378), .ZN(n11386) );
  NAND2_X1 U14179 ( .A1(n11387), .A2(n11386), .ZN(n14124) );
  NAND2_X1 U14180 ( .A1(n11388), .A2(n14124), .ZN(n11389) );
  INV_X1 U14181 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14160) );
  NAND2_X1 U14182 ( .A1(n11396), .A2(n14160), .ZN(n11392) );
  INV_X1 U14183 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14430) );
  NAND2_X1 U14184 ( .A1(n11397), .A2(n14430), .ZN(n11390) );
  OAI211_X1 U14185 ( .C1(n11313), .C2(P1_EBX_REG_26__SCAN_IN), .A(n11390), .B(
        n11378), .ZN(n11391) );
  NAND2_X1 U14186 ( .A1(n11392), .A2(n11391), .ZN(n14095) );
  MUX2_X1 U14187 ( .A(n11393), .B(n9998), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11395) );
  NOR2_X1 U14188 ( .A1(n13214), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11394) );
  NOR2_X1 U14189 ( .A1(n11395), .A2(n11394), .ZN(n14082) );
  INV_X1 U14190 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n13200) );
  NAND2_X1 U14191 ( .A1(n11396), .A2(n13200), .ZN(n11400) );
  INV_X1 U14192 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14286) );
  NAND2_X1 U14193 ( .A1(n11397), .A2(n14286), .ZN(n11398) );
  OAI211_X1 U14194 ( .C1(n11313), .C2(P1_EBX_REG_28__SCAN_IN), .A(n11398), .B(
        n11378), .ZN(n11399) );
  AND2_X1 U14195 ( .A1(n11400), .A2(n11399), .ZN(n13198) );
  INV_X1 U14196 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n11401) );
  NAND2_X1 U14197 ( .A1(n11837), .A2(n11401), .ZN(n11402) );
  OAI21_X1 U14198 ( .B1(n13214), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11402), .ZN(n11403) );
  MUX2_X1 U14199 ( .A(n11403), .B(n11402), .S(n9998), .Z(n14074) );
  OAI22_X1 U14200 ( .A1(n14073), .A2(n11378), .B1(n11403), .B2(n9839), .ZN(
        n11405) );
  AOI22_X1 U14201 ( .A1(n13214), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n11313), .ZN(n13213) );
  INV_X1 U14202 ( .A(n13213), .ZN(n11404) );
  XNOR2_X1 U14203 ( .A(n11405), .B(n11404), .ZN(n14059) );
  OAI22_X1 U14204 ( .A1(n12342), .A2(n20729), .B1(n11412), .B2(n11406), .ZN(
        n11407) );
  OAI21_X1 U14205 ( .B1(n14059), .B2(n20003), .A(n11409), .ZN(n11410) );
  INV_X1 U14206 ( .A(n11410), .ZN(n11418) );
  NAND2_X1 U14207 ( .A1(n11428), .A2(n10381), .ZN(n11411) );
  NAND2_X1 U14208 ( .A1(n15680), .A2(n11411), .ZN(n11839) );
  OAI21_X1 U14209 ( .B1(n20079), .B2(n11412), .A(n11839), .ZN(n11413) );
  NOR2_X1 U14210 ( .A1(n11414), .A2(n11413), .ZN(n11415) );
  NOR2_X2 U14211 ( .A1(n11416), .A2(n11415), .ZN(n20031) );
  OAI211_X1 U14212 ( .C1(n11419), .C2(n10310), .A(n11418), .B(n9847), .ZN(
        P1_U3001) );
  AND2_X1 U14213 ( .A1(n15680), .A2(n12795), .ZN(n12333) );
  NAND2_X1 U14214 ( .A1(n12333), .A2(n15694), .ZN(n11421) );
  OAI21_X1 U14215 ( .B1(n12565), .B2(n11422), .A(n11421), .ZN(n12341) );
  NAND4_X1 U14216 ( .A1(n12380), .A2(n11424), .A3(n20091), .A4(n11423), .ZN(
        n11465) );
  INV_X1 U14217 ( .A(n11425), .ZN(n11426) );
  NAND3_X1 U14218 ( .A1(n11426), .A2(n20726), .A3(n15694), .ZN(n11427) );
  OAI21_X1 U14219 ( .B1(n11465), .B2(n11428), .A(n11427), .ZN(n11429) );
  AND2_X1 U14220 ( .A1(n20083), .A2(n11846), .ZN(n11444) );
  INV_X1 U14221 ( .A(n11444), .ZN(n11431) );
  AND2_X1 U14222 ( .A1(n11431), .A2(n11433), .ZN(n11432) );
  NOR2_X1 U14223 ( .A1(n14235), .A2(n11433), .ZN(n12728) );
  NOR4_X1 U14224 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n11437) );
  NOR4_X1 U14225 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n11436) );
  NOR4_X1 U14226 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n11435) );
  NOR4_X1 U14227 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n11434) );
  AND4_X1 U14228 ( .A1(n11437), .A2(n11436), .A3(n11435), .A4(n11434), .ZN(
        n11442) );
  NOR4_X1 U14229 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n11440) );
  NOR4_X1 U14230 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_24__SCAN_IN), .A3(P1_ADDRESS_REG_23__SCAN_IN), .A4(
        P1_ADDRESS_REG_22__SCAN_IN), .ZN(n11439) );
  NOR4_X1 U14231 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(
        P1_ADDRESS_REG_3__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n11438) );
  INV_X1 U14232 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20648) );
  AND4_X1 U14233 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n20648), .ZN(
        n11441) );
  NAND2_X1 U14234 ( .A1(n11442), .A2(n11441), .ZN(n11443) );
  NAND2_X1 U14235 ( .A1(n12728), .A2(n20045), .ZN(n14239) );
  INV_X1 U14236 ( .A(DATAI_14_), .ZN(n11445) );
  INV_X1 U14237 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n11860) );
  MUX2_X1 U14238 ( .A(n11445), .B(n11860), .S(n20045), .Z(n19967) );
  OAI22_X1 U14239 ( .A1(n14262), .A2(n19967), .B1(n14271), .B2(n11446), .ZN(
        n11447) );
  AOI21_X1 U14240 ( .B1(n14264), .B2(BUF1_REG_30__SCAN_IN), .A(n11447), .ZN(
        n11449) );
  INV_X1 U14241 ( .A(n20045), .ZN(n20043) );
  NAND2_X1 U14242 ( .A1(n14265), .A2(DATAI_30_), .ZN(n11448) );
  AND2_X1 U14243 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  OAI21_X1 U14244 ( .B1(n14069), .B2(n14268), .A(n11450), .ZN(P1_U2874) );
  NAND2_X1 U14245 ( .A1(n11454), .A2(n11453), .ZN(n11458) );
  AOI22_X1 U14246 ( .A1(n10957), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11455), .ZN(n11456) );
  INV_X1 U14247 ( .A(n11456), .ZN(n11457) );
  XNOR2_X2 U14248 ( .A(n11458), .B(n11457), .ZN(n13988) );
  INV_X1 U14249 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13219) );
  INV_X1 U14250 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20694) );
  NOR2_X1 U14251 ( .A1(n20002), .A2(n20694), .ZN(n14398) );
  AOI21_X1 U14252 ( .B1(n19987), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14398), .ZN(n11462) );
  OAI21_X1 U14253 ( .B1(n12798), .B2(n19998), .A(n11462), .ZN(n11463) );
  OAI21_X1 U14254 ( .B1(n14400), .B2(n19817), .A(n11464), .ZN(P1_U2968) );
  NAND2_X1 U14255 ( .A1(n12334), .A2(n11842), .ZN(n12349) );
  OR2_X1 U14256 ( .A1(n11313), .A2(n11465), .ZN(n11466) );
  NAND2_X1 U14257 ( .A1(n12349), .A2(n11466), .ZN(n11467) );
  NAND2_X2 U14258 ( .A1(n19919), .A2(n20091), .ZN(n19912) );
  INV_X1 U14259 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n11469) );
  AOI21_X1 U14260 ( .B1(n11471), .B2(n19908), .A(n11470), .ZN(n11472) );
  INV_X1 U14261 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20737) );
  NOR3_X1 U14262 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20737), .ZN(n11475) );
  NOR4_X1 U14263 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n11474) );
  NAND4_X1 U14264 ( .A1(n20045), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n11475), .A4(
        n11474), .ZN(U214) );
  NOR4_X1 U14265 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n11479) );
  NOR4_X1 U14266 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n11478) );
  NOR4_X1 U14267 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11477) );
  NOR4_X1 U14268 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n11476) );
  NAND4_X1 U14269 ( .A1(n11479), .A2(n11478), .A3(n11477), .A4(n11476), .ZN(
        n11484) );
  NOR4_X1 U14270 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n11482) );
  NOR4_X1 U14271 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n11481) );
  NOR4_X1 U14272 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n11480) );
  INV_X1 U14273 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19699) );
  NAND4_X1 U14274 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n19699), .ZN(
        n11483) );
  OAI21_X1 U14275 ( .B1(n11484), .B2(n11483), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n11485) );
  NOR2_X1 U14276 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n11487) );
  NOR4_X1 U14277 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14278 ( .A1(P2_W_R_N_REG_SCAN_IN), .A2(P2_M_IO_N_REG_SCAN_IN), 
        .A3(n11487), .A4(n11486), .ZN(n11488) );
  NOR2_X1 U14279 ( .A1(n15429), .A2(n11488), .ZN(n16307) );
  NAND2_X1 U14280 ( .A1(n16307), .A2(U214), .ZN(U212) );
  NOR2_X1 U14281 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n11488), .ZN(n16378)
         );
  INV_X1 U14282 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U14283 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17473) );
  INV_X1 U14284 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21011) );
  NAND2_X1 U14285 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17666) );
  NAND2_X1 U14286 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17534) );
  NOR2_X1 U14287 ( .A1(n17534), .A2(n17533), .ZN(n17504) );
  NAND2_X1 U14288 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17505) );
  NOR2_X1 U14289 ( .A1(n21011), .A2(n17471), .ZN(n17470) );
  INV_X1 U14290 ( .A(n17470), .ZN(n16568) );
  NOR2_X1 U14291 ( .A1(n17473), .A2(n16568), .ZN(n17434) );
  INV_X1 U14292 ( .A(n17434), .ZN(n16544) );
  NOR2_X1 U14293 ( .A1(n10097), .A2(n16544), .ZN(n11490) );
  NAND2_X1 U14294 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11490), .ZN(
        n11489) );
  NOR2_X1 U14295 ( .A1(n11616), .A2(n11489), .ZN(n17389) );
  AOI21_X1 U14296 ( .B1(n11616), .B2(n11489), .A(n17389), .ZN(n17436) );
  OAI21_X1 U14297 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11490), .A(
        n11489), .ZN(n17444) );
  INV_X1 U14298 ( .A(n17444), .ZN(n16525) );
  AOI21_X1 U14299 ( .B1(n10097), .B2(n16544), .A(n11490), .ZN(n17461) );
  NOR2_X1 U14300 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21011), .ZN(
        n16754) );
  NAND2_X1 U14301 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17438) );
  NAND2_X1 U14302 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17393) );
  NAND2_X1 U14303 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17353) );
  AOI21_X1 U14304 ( .B1(n9869), .B2(n16754), .A(n16764), .ZN(n16538) );
  NOR2_X1 U14305 ( .A1(n17461), .A2(n16538), .ZN(n16537) );
  NOR2_X1 U14306 ( .A1(n16537), .A2(n16764), .ZN(n16524) );
  NOR2_X1 U14307 ( .A1(n16525), .A2(n16524), .ZN(n16523) );
  NOR2_X1 U14308 ( .A1(n16523), .A2(n16764), .ZN(n11491) );
  NOR2_X1 U14309 ( .A1(n17436), .A2(n11491), .ZN(n16426) );
  NOR3_X1 U14310 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18569) );
  AND2_X1 U14311 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18569), .ZN(n16753) );
  INV_X1 U14312 ( .A(n16753), .ZN(n18565) );
  AOI211_X1 U14313 ( .C1(n17436), .C2(n11491), .A(n16426), .B(n18565), .ZN(
        n11625) );
  NOR3_X1 U14314 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16747) );
  NAND2_X1 U14315 ( .A1(n16747), .A2(n16743), .ZN(n16740) );
  NOR2_X1 U14316 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16740), .ZN(n16724) );
  INV_X1 U14317 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17060) );
  NAND2_X1 U14318 ( .A1(n16724), .A2(n17060), .ZN(n16714) );
  NOR2_X1 U14319 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16714), .ZN(n16696) );
  INV_X1 U14320 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16969) );
  NAND2_X1 U14321 ( .A1(n16696), .A2(n16969), .ZN(n16693) );
  INV_X1 U14322 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16995) );
  NAND2_X1 U14323 ( .A1(n16668), .A2(n16995), .ZN(n16650) );
  INV_X1 U14324 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16997) );
  NAND2_X1 U14325 ( .A1(n16649), .A2(n16997), .ZN(n16646) );
  INV_X1 U14326 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16620) );
  NAND2_X1 U14327 ( .A1(n16626), .A2(n16620), .ZN(n16619) );
  INV_X1 U14328 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16598) );
  NAND2_X1 U14329 ( .A1(n16603), .A2(n16598), .ZN(n16597) );
  INV_X1 U14330 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16577) );
  NAND2_X1 U14331 ( .A1(n16578), .A2(n16577), .ZN(n16574) );
  NOR2_X1 U14332 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16574), .ZN(n16559) );
  INV_X1 U14333 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16556) );
  NAND2_X1 U14334 ( .A1(n16559), .A2(n16556), .ZN(n16553) );
  NOR2_X1 U14335 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16553), .ZN(n16534) );
  INV_X1 U14336 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16526) );
  NAND2_X1 U14337 ( .A1(n16534), .A2(n16526), .ZN(n16529) );
  NOR2_X1 U14338 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16529), .ZN(n16518) );
  INV_X2 U14339 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18690) );
  INV_X2 U14340 ( .A(n16953), .ZN(n17035) );
  INV_X2 U14341 ( .A(n15485), .ZN(n17003) );
  AOI22_X1 U14342 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11494) );
  OAI21_X1 U14343 ( .B1(n9840), .B2(n21015), .A(n11494), .ZN(n11506) );
  INV_X4 U14344 ( .A(n16899), .ZN(n16924) );
  AOI22_X1 U14345 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11504) );
  NOR2_X2 U14346 ( .A1(n18526), .A2(n11497), .ZN(n12889) );
  AOI22_X1 U14347 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11503) );
  INV_X2 U14348 ( .A(n17018), .ZN(n17039) );
  AOI22_X1 U14349 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11502) );
  NOR2_X2 U14350 ( .A1(n11500), .A2(n11499), .ZN(n15492) );
  AOI22_X1 U14351 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11501) );
  NAND4_X1 U14352 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11505) );
  NAND2_X1 U14353 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18708), .ZN(n16667) );
  NAND2_X1 U14354 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18702) );
  INV_X1 U14355 ( .A(n18702), .ZN(n18709) );
  AOI22_X1 U14356 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U14357 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14358 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14359 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11511) );
  NAND4_X1 U14360 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(
        n11520) );
  AOI22_X1 U14361 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14362 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14363 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11516) );
  INV_X2 U14364 ( .A(n15575), .ZN(n17004) );
  AOI22_X1 U14365 ( .A1(n17004), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11515) );
  NAND4_X1 U14366 ( .A1(n11518), .A2(n11517), .A3(n11516), .A4(n11515), .ZN(
        n11519) );
  AOI22_X1 U14367 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14368 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14369 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14370 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11521) );
  NAND4_X1 U14371 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11531) );
  AOI22_X1 U14372 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14373 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14374 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11527) );
  INV_X2 U14375 ( .A(n11567), .ZN(n17046) );
  AOI22_X1 U14376 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11526) );
  NAND4_X1 U14377 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11530) );
  AOI22_X1 U14378 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14379 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14380 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11533) );
  INV_X2 U14381 ( .A(n15575), .ZN(n15551) );
  AOI22_X1 U14382 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11532) );
  NAND4_X1 U14383 ( .A1(n11535), .A2(n11534), .A3(n11533), .A4(n11532), .ZN(
        n11541) );
  AOI22_X1 U14384 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14385 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14386 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14387 ( .A1(n9790), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11536) );
  NAND4_X1 U14388 ( .A1(n11539), .A2(n11538), .A3(n11537), .A4(n11536), .ZN(
        n11540) );
  NAND2_X1 U14389 ( .A1(n18057), .A2(n18080), .ZN(n13179) );
  AOI22_X1 U14390 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14391 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14392 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14393 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11542) );
  NAND4_X1 U14394 ( .A1(n11545), .A2(n11544), .A3(n11543), .A4(n11542), .ZN(
        n11551) );
  AOI22_X1 U14395 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14396 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14397 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14398 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11546) );
  NAND4_X1 U14399 ( .A1(n11549), .A2(n11548), .A3(n11547), .A4(n11546), .ZN(
        n11550) );
  AOI22_X1 U14400 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14401 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14402 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11552) );
  OAI21_X1 U14403 ( .B1(n17018), .B2(n20973), .A(n11552), .ZN(n11558) );
  AOI22_X1 U14404 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14405 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14406 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14407 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9787), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11553) );
  NAND4_X1 U14408 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n11557) );
  AOI211_X1 U14409 ( .C1(n17003), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n11558), .B(n11557), .ZN(n11559) );
  NAND3_X1 U14410 ( .A1(n11561), .A2(n11560), .A3(n11559), .ZN(n15604) );
  NAND2_X1 U14411 ( .A1(n17087), .A2(n15604), .ZN(n11592) );
  AOI22_X1 U14412 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14413 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11564) );
  INV_X2 U14414 ( .A(n11575), .ZN(n17020) );
  AOI22_X1 U14415 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14416 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11562) );
  NAND4_X1 U14417 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11573) );
  AOI22_X1 U14418 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14419 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14420 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14421 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11568) );
  NAND4_X1 U14422 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11572) );
  NAND2_X1 U14423 ( .A1(n18080), .A2(n18091), .ZN(n11586) );
  AOI22_X1 U14424 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14425 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16924), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14426 ( .A1(n17004), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11574) );
  OAI21_X1 U14427 ( .B1(n11575), .B2(n18072), .A(n11574), .ZN(n11582) );
  AOI22_X1 U14428 ( .A1(n9790), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14429 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14430 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14431 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11577) );
  NAND4_X1 U14432 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11581) );
  INV_X1 U14433 ( .A(n15599), .ZN(n18069) );
  NAND2_X1 U14434 ( .A1(n18057), .A2(n18708), .ZN(n11596) );
  OAI211_X1 U14435 ( .C1(n18085), .C2(n11586), .A(n18069), .B(n11596), .ZN(
        n13181) );
  NOR2_X1 U14436 ( .A1(n18085), .A2(n15599), .ZN(n12826) );
  INV_X1 U14437 ( .A(n12826), .ZN(n15595) );
  NOR2_X1 U14438 ( .A1(n15595), .A2(n18091), .ZN(n15598) );
  OAI21_X1 U14439 ( .B1(n11594), .B2(n15598), .A(n18057), .ZN(n11587) );
  INV_X1 U14440 ( .A(n11587), .ZN(n11591) );
  NOR2_X1 U14441 ( .A1(n15604), .A2(n18085), .ZN(n18530) );
  NOR2_X1 U14442 ( .A1(n18708), .A2(n18057), .ZN(n15587) );
  OAI21_X1 U14443 ( .B1(n18097), .B2(n18530), .A(n15587), .ZN(n13183) );
  OAI21_X1 U14444 ( .B1(n12826), .B2(n11594), .A(n13183), .ZN(n11589) );
  AOI21_X1 U14445 ( .B1(n17163), .B2(n11592), .A(n18080), .ZN(n11588) );
  INV_X1 U14446 ( .A(n11596), .ZN(n15588) );
  NAND2_X1 U14447 ( .A1(n11595), .A2(n15594), .ZN(n15590) );
  NOR2_X1 U14448 ( .A1(n17087), .A2(n18091), .ZN(n13182) );
  NAND4_X1 U14449 ( .A1(n15591), .A2(n18085), .A3(n11594), .A4(n17239), .ZN(
        n17279) );
  NAND2_X1 U14450 ( .A1(n15599), .A2(n11595), .ZN(n13178) );
  NAND2_X1 U14451 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17709), .ZN(n18559) );
  NAND2_X1 U14452 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18360), .ZN(
        n12827) );
  OAI22_X1 U14453 ( .A1(n18675), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21014), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11601) );
  XNOR2_X1 U14454 ( .A(n11602), .B(n11601), .ZN(n11610) );
  AOI22_X1 U14455 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18504), .B1(
        n11604), .B2(n18665), .ZN(n11606) );
  INV_X1 U14456 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18543) );
  NOR2_X1 U14457 ( .A1(n11604), .A2(n18665), .ZN(n11607) );
  NAND2_X1 U14458 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18504), .ZN(
        n11605) );
  OAI22_X1 U14459 ( .A1(n11606), .A2(n18543), .B1(n11607), .B2(n11605), .ZN(
        n12829) );
  INV_X1 U14460 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20939) );
  OAI21_X1 U14461 ( .B1(n18543), .B2(n11607), .A(n11606), .ZN(n11608) );
  INV_X1 U14462 ( .A(n11608), .ZN(n11609) );
  INV_X1 U14463 ( .A(n12827), .ZN(n11613) );
  NAND2_X1 U14464 ( .A1(n11613), .A2(n12828), .ZN(n11611) );
  OAI211_X1 U14465 ( .C1(n11613), .C2(n12828), .A(n11612), .B(n11611), .ZN(
        n15602) );
  AOI211_X1 U14466 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16529), .A(n16518), .B(
        n16770), .ZN(n11624) );
  NAND2_X1 U14467 ( .A1(n17709), .A2(n18684), .ZN(n18670) );
  NOR3_X1 U14468 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18670), .ZN(n15711) );
  NAND2_X1 U14469 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18720), .ZN(n18560) );
  NOR2_X1 U14470 ( .A1(n18559), .A2(n18560), .ZN(n18555) );
  NAND2_X1 U14471 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18584), .ZN(n18718) );
  INV_X2 U14472 ( .A(n18718), .ZN(n18652) );
  NAND2_X1 U14473 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18652), .ZN(n18642) );
  NOR2_X1 U14474 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n16396) );
  INV_X1 U14475 ( .A(n16396), .ZN(n18571) );
  NAND3_X1 U14476 ( .A1(n18584), .A2(n18636), .A3(n18571), .ZN(n18577) );
  AOI211_X1 U14477 ( .C1(n18577), .C2(n18062), .A(n18709), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18551) );
  AOI211_X4 U14478 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18708), .A(n18551), .B(
        n11614), .ZN(n16722) );
  INV_X1 U14479 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n11615) );
  OAI22_X1 U14480 ( .A1(n11616), .A2(n16745), .B1(n16767), .B2(n11615), .ZN(
        n11623) );
  INV_X1 U14481 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18612) );
  INV_X1 U14482 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18609) );
  INV_X1 U14483 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18606) );
  NAND3_X1 U14484 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n16707) );
  NAND2_X1 U14485 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n16652) );
  INV_X1 U14486 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18601) );
  NAND2_X1 U14487 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16688) );
  NOR2_X1 U14488 ( .A1(n18601), .A2(n16688), .ZN(n16653) );
  NAND3_X1 U14489 ( .A1(n16653), .A2(P3_REIP_REG_10__SCAN_IN), .A3(
        P3_REIP_REG_9__SCAN_IN), .ZN(n16635) );
  NOR4_X1 U14490 ( .A1(n18606), .A2(n16707), .A3(n16652), .A4(n16635), .ZN(
        n16625) );
  NAND2_X1 U14491 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16625), .ZN(n16604) );
  NOR3_X1 U14492 ( .A1(n18612), .A2(n18609), .A3(n16604), .ZN(n11618) );
  NAND2_X1 U14493 ( .A1(n16761), .A2(n11618), .ZN(n16566) );
  INV_X1 U14494 ( .A(n16566), .ZN(n16596) );
  NAND4_X1 U14495 ( .A1(n16596), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16561) );
  NAND2_X1 U14496 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16547) );
  INV_X1 U14497 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18626) );
  NOR2_X1 U14498 ( .A1(n16532), .A2(n18626), .ZN(n11621) );
  NAND3_X1 U14499 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n11619) );
  NAND2_X1 U14500 ( .A1(n11618), .A2(n16779), .ZN(n16580) );
  NOR2_X1 U14501 ( .A1(n11619), .A2(n16580), .ZN(n16548) );
  NAND4_X1 U14502 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_20__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n16548), .ZN(n16536) );
  NOR2_X1 U14503 ( .A1(n16761), .A2(n16773), .ZN(n16581) );
  OAI21_X1 U14504 ( .B1(n18626), .B2(n16536), .A(n16777), .ZN(n16533) );
  INV_X1 U14505 ( .A(n16533), .ZN(n11620) );
  MUX2_X1 U14506 ( .A(n11621), .B(n11620), .S(P3_REIP_REG_22__SCAN_IN), .Z(
        n11622) );
  OR4_X1 U14507 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        P3_U2649) );
  AND2_X4 U14508 ( .A1(n12656), .A2(n10276), .ZN(n14034) );
  AOI22_X1 U14509 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11632) );
  INV_X1 U14510 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11626) );
  AND2_X2 U14511 ( .A1(n11626), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11627) );
  AND3_X4 U14512 ( .A1(n11628), .A2(n10276), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U14513 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11631) );
  AND2_X4 U14514 ( .A1(n11627), .A2(n11628), .ZN(n13767) );
  AND2_X4 U14515 ( .A1(n12681), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11955) );
  AOI22_X1 U14516 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11630) );
  AND2_X4 U14517 ( .A1(n12656), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14036) );
  AOI22_X1 U14518 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9785), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11629) );
  NAND4_X1 U14519 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11639) );
  INV_X2 U14520 ( .A(n11633), .ZN(n14035) );
  AOI22_X1 U14521 ( .A1(n14035), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14522 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14523 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14524 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11634) );
  NAND4_X1 U14525 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11638) );
  MUX2_X2 U14526 ( .A(n11639), .B(n11638), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15433) );
  INV_X2 U14527 ( .A(n15433), .ZN(n12075) );
  AOI22_X1 U14528 ( .A1(n14035), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14529 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14530 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14531 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9785), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11640) );
  NAND4_X1 U14532 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n11649) );
  AOI22_X1 U14533 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14534 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14535 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14536 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9784), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11644) );
  NAND4_X1 U14537 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11648) );
  MUX2_X2 U14538 ( .A(n11649), .B(n11648), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11910) );
  AOI22_X1 U14539 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14540 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14541 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9784), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11650) );
  NAND3_X1 U14542 ( .A1(n11652), .A2(n11651), .A3(n11650), .ZN(n11655) );
  AOI22_X1 U14543 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11653) );
  OAI21_X2 U14544 ( .B1(n11655), .B2(n11654), .A(n12694), .ZN(n11662) );
  AOI22_X1 U14545 ( .A1(n14035), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14546 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14547 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14548 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11656) );
  NAND4_X1 U14549 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11660) );
  NAND2_X2 U14550 ( .A1(n11662), .A2(n11661), .ZN(n12105) );
  AOI22_X1 U14551 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14552 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14553 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11663) );
  NAND4_X1 U14554 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n11667) );
  AOI22_X1 U14555 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13767), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14556 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14557 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14036), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14558 ( .A1(n11955), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11668) );
  NAND4_X1 U14559 ( .A1(n11671), .A2(n11670), .A3(n11669), .A4(n11668), .ZN(
        n11672) );
  NAND2_X4 U14560 ( .A1(n11674), .A2(n11673), .ZN(n12483) );
  AOI22_X1 U14561 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14562 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14563 ( .A1(n14035), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14564 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11675) );
  NAND4_X1 U14565 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11679) );
  AOI22_X1 U14566 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14567 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14568 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9785), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14569 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11680) );
  NAND4_X1 U14570 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n11684) );
  AOI22_X1 U14571 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14572 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14573 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14574 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9784), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14575 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14576 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14577 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9785), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14578 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14579 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14580 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14581 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14582 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9785), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11695) );
  NAND2_X1 U14583 ( .A1(n11699), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11706) );
  AOI22_X1 U14584 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14585 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9786), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U14586 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14587 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11700) );
  NAND2_X1 U14588 ( .A1(n11704), .A2(n12694), .ZN(n11705) );
  NAND2_X2 U14589 ( .A1(n11706), .A2(n11705), .ZN(n11963) );
  INV_X1 U14590 ( .A(n11911), .ZN(n11918) );
  INV_X1 U14591 ( .A(n15479), .ZN(n11708) );
  NAND2_X1 U14592 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19794), .ZN(
        n11755) );
  INV_X1 U14593 ( .A(n11755), .ZN(n11709) );
  NAND2_X1 U14594 ( .A1(n11999), .A2(n11709), .ZN(n11711) );
  NAND2_X1 U14595 ( .A1(n19787), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11710) );
  NAND2_X1 U14596 ( .A1(n11711), .A2(n11710), .ZN(n11721) );
  XNOR2_X1 U14597 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11720) );
  NAND2_X1 U14598 ( .A1(n11721), .A2(n11720), .ZN(n11713) );
  NAND2_X1 U14599 ( .A1(n19777), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11712) );
  XNOR2_X1 U14600 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11718) );
  NOR2_X1 U14601 ( .A1(n12694), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11714) );
  INV_X1 U14602 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15740) );
  NAND2_X1 U14603 ( .A1(n15740), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11715) );
  NAND2_X1 U14604 ( .A1(n11723), .A2(n11715), .ZN(n11717) );
  INV_X1 U14605 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15482) );
  NAND2_X1 U14606 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15482), .ZN(
        n11716) );
  XNOR2_X1 U14607 ( .A(n11999), .B(n11755), .ZN(n11756) );
  XNOR2_X1 U14608 ( .A(n11719), .B(n11718), .ZN(n12956) );
  XNOR2_X1 U14609 ( .A(n11721), .B(n11720), .ZN(n11997) );
  NOR2_X1 U14610 ( .A1(n15740), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11722) );
  NOR3_X1 U14611 ( .A1(n12956), .A2(n11997), .A3(n13040), .ZN(n12007) );
  AND2_X1 U14612 ( .A1(n11756), .A2(n12007), .ZN(n11724) );
  NAND2_X1 U14613 ( .A1(n15409), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12965) );
  OR2_X1 U14614 ( .A1(n12697), .A2(n18734), .ZN(n11728) );
  OR2_X1 U14615 ( .A1(n11900), .A2(n11728), .ZN(n14703) );
  INV_X1 U14616 ( .A(n14703), .ZN(n18964) );
  INV_X1 U14617 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n19808) );
  AND2_X2 U14618 ( .A1(n12483), .A2(n12105), .ZN(n11726) );
  AND2_X2 U14619 ( .A1(n11726), .A2(n11725), .ZN(n11919) );
  INV_X1 U14620 ( .A(n11905), .ZN(n11727) );
  OR2_X1 U14621 ( .A1(n12721), .A2(n11728), .ZN(n12969) );
  NOR2_X1 U14622 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19764) );
  NOR2_X1 U14623 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19756), .ZN(n12018) );
  INV_X1 U14624 ( .A(n12018), .ZN(n11729) );
  AND2_X1 U14625 ( .A1(n12969), .A2(n11729), .ZN(n11744) );
  OAI21_X1 U14626 ( .B1(n18964), .B2(n19808), .A(n11744), .ZN(P2_U2814) );
  INV_X1 U14627 ( .A(n12697), .ZN(n12083) );
  NAND2_X1 U14628 ( .A1(n11937), .A2(n12083), .ZN(n12704) );
  AOI22_X1 U14629 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11733) );
  AOI22_X1 U14630 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14631 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14632 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11730) );
  NAND4_X1 U14633 ( .A1(n11733), .A2(n11732), .A3(n11731), .A4(n11730), .ZN(
        n11734) );
  AOI22_X1 U14634 ( .A1(n11735), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14635 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14636 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11950), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14637 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9784), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11736) );
  NAND4_X1 U14638 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n11740) );
  NAND2_X1 U14639 ( .A1(n11740), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11741) );
  INV_X1 U14640 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n11743) );
  NAND3_X1 U14641 ( .A1(n11744), .A2(n14703), .A3(n11743), .ZN(n11745) );
  OAI21_X1 U14642 ( .B1(n18730), .B2(n11897), .A(n11745), .ZN(n11746) );
  INV_X1 U14643 ( .A(n11746), .ZN(P2_U3612) );
  AND2_X1 U14644 ( .A1(n11833), .A2(n11892), .ZN(n11747) );
  NAND2_X1 U14645 ( .A1(n11271), .A2(n11747), .ZN(n11750) );
  INV_X1 U14646 ( .A(n11750), .ZN(n11749) );
  INV_X1 U14647 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20738) );
  NAND3_X1 U14648 ( .A1(n15694), .A2(n11892), .A3(n11748), .ZN(n12248) );
  NAND2_X1 U14649 ( .A1(n20496), .A2(n20627), .ZN(n19814) );
  OAI211_X1 U14650 ( .C1(n11749), .C2(n20738), .A(n12248), .B(n19814), .ZN(
        P1_U2801) );
  NAND2_X1 U14651 ( .A1(n12248), .A2(n11750), .ZN(n20724) );
  INV_X1 U14652 ( .A(n20724), .ZN(n11753) );
  INV_X1 U14653 ( .A(n19814), .ZN(n11751) );
  OAI21_X1 U14654 ( .B1(n11751), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n11753), 
        .ZN(n11752) );
  OAI21_X1 U14655 ( .B1(n11754), .B2(n11753), .A(n11752), .ZN(P1_U3487) );
  INV_X1 U14656 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n11878) );
  OAI21_X1 U14657 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19794), .A(
        n11755), .ZN(n11757) );
  INV_X1 U14658 ( .A(n11757), .ZN(n12008) );
  OAI211_X1 U14659 ( .C1(n14018), .C2(n12008), .A(n12075), .B(n11756), .ZN(
        n11760) );
  INV_X1 U14660 ( .A(n11999), .ZN(n11758) );
  INV_X1 U14661 ( .A(n12948), .ZN(n11764) );
  OAI21_X1 U14662 ( .B1(n11758), .B2(n11757), .A(n11764), .ZN(n11759) );
  OAI211_X1 U14663 ( .C1(n15478), .C2(n11997), .A(n11760), .B(n11759), .ZN(
        n11763) );
  NAND2_X1 U14664 ( .A1(n11769), .A2(n14018), .ZN(n11761) );
  MUX2_X1 U14665 ( .A(n12948), .B(n11761), .S(n11997), .Z(n11762) );
  AOI21_X1 U14666 ( .B1(n11763), .B2(n11762), .A(n12956), .ZN(n11767) );
  AOI21_X1 U14667 ( .B1(n11764), .B2(n13040), .A(n12002), .ZN(n11765) );
  OAI21_X1 U14668 ( .B1(n11767), .B2(n11766), .A(n11765), .ZN(n11768) );
  MUX2_X1 U14669 ( .A(n11768), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n12943), .Z(n12071) );
  NAND2_X1 U14670 ( .A1(n12701), .A2(n14018), .ZN(n12647) );
  OR2_X1 U14671 ( .A1(n11900), .A2(n18734), .ZN(n11771) );
  OAI21_X1 U14672 ( .B1(n12647), .B2(n11771), .A(n11887), .ZN(n11773) );
  NOR2_X1 U14673 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20741) );
  INV_X1 U14674 ( .A(n20741), .ZN(n19690) );
  NAND2_X1 U14675 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19683), .ZN(n19806) );
  INV_X2 U14676 ( .A(n19806), .ZN(n20740) );
  NAND2_X2 U14677 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20740), .ZN(n19741) );
  NAND3_X1 U14678 ( .A1(n19683), .A2(n19690), .A3(n19741), .ZN(n19681) );
  INV_X1 U14679 ( .A(n19681), .ZN(n11772) );
  NAND2_X1 U14680 ( .A1(n19089), .A2(n11907), .ZN(n11795) );
  NAND2_X1 U14681 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n16225) );
  NOR2_X1 U14682 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16225), .ZN(n19088) );
  CLKBUF_X1 U14683 ( .A(n19088), .Z(n19097) );
  INV_X2 U14684 ( .A(n19091), .ZN(n19094) );
  AOI22_X1 U14685 ( .A1(n19088), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11774) );
  OAI21_X1 U14686 ( .B1(n11878), .B2(n11795), .A(n11774), .ZN(P2_U2925) );
  INV_X1 U14687 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14795) );
  AOI22_X1 U14688 ( .A1(n19088), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n11775) );
  OAI21_X1 U14689 ( .B1(n14795), .B2(n11795), .A(n11775), .ZN(P2_U2929) );
  INV_X1 U14690 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14773) );
  AOI22_X1 U14691 ( .A1(n19088), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n11776) );
  OAI21_X1 U14692 ( .B1(n14773), .B2(n11795), .A(n11776), .ZN(P2_U2926) );
  INV_X1 U14693 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14694 ( .A1(n19088), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11777) );
  OAI21_X1 U14695 ( .B1(n11778), .B2(n11795), .A(n11777), .ZN(P2_U2928) );
  INV_X1 U14696 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U14697 ( .A1(n19088), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n11779) );
  OAI21_X1 U14698 ( .B1(n14809), .B2(n11795), .A(n11779), .ZN(P2_U2932) );
  INV_X1 U14699 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14700 ( .A1(n19088), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n11780) );
  OAI21_X1 U14701 ( .B1(n11781), .B2(n11795), .A(n11780), .ZN(P2_U2931) );
  INV_X1 U14702 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14703 ( .A1(n19088), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11782) );
  OAI21_X1 U14704 ( .B1(n11871), .B2(n11795), .A(n11782), .ZN(P2_U2927) );
  INV_X1 U14705 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14706 ( .A1(n19088), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n11783) );
  OAI21_X1 U14707 ( .B1(n11784), .B2(n11795), .A(n11783), .ZN(P2_U2930) );
  INV_X1 U14708 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14709 ( .A1(n19097), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11785) );
  OAI21_X1 U14710 ( .B1(n11852), .B2(n11795), .A(n11785), .ZN(P2_U2923) );
  INV_X1 U14711 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14712 ( .A1(n19097), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11786) );
  OAI21_X1 U14713 ( .B1(n11787), .B2(n11795), .A(n11786), .ZN(P2_U2924) );
  INV_X1 U14714 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14715 ( .A1(n19097), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11788) );
  OAI21_X1 U14716 ( .B1(n11864), .B2(n11795), .A(n11788), .ZN(P2_U2921) );
  INV_X1 U14717 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14718 ( .A1(n19097), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11789) );
  OAI21_X1 U14719 ( .B1(n11790), .B2(n11795), .A(n11789), .ZN(P2_U2922) );
  INV_X1 U14720 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14721 ( .A1(n19097), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n11791) );
  OAI21_X1 U14722 ( .B1(n11792), .B2(n11795), .A(n11791), .ZN(P2_U2934) );
  INV_X1 U14723 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14724 ( .A1(n19097), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n11793) );
  OAI21_X1 U14725 ( .B1(n11880), .B2(n11795), .A(n11793), .ZN(P2_U2935) );
  INV_X1 U14726 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14727 ( .A1(n19097), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n11794) );
  OAI21_X1 U14728 ( .B1(n11796), .B2(n11795), .A(n11794), .ZN(P2_U2933) );
  NAND2_X1 U14729 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n15735) );
  INV_X1 U14730 ( .A(n12969), .ZN(n11797) );
  OAI21_X1 U14731 ( .B1(n10055), .B2(n15735), .A(n11797), .ZN(n11853) );
  AOI22_X1 U14732 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11800) );
  INV_X1 U14733 ( .A(n15735), .ZN(n19680) );
  NOR3_X1 U14734 ( .A1(n12969), .A2(n10055), .A3(n19680), .ZN(n11798) );
  AOI22_X1 U14735 ( .A1(n15431), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15429), .ZN(n19176) );
  INV_X1 U14736 ( .A(n19176), .ZN(n11799) );
  NAND2_X1 U14737 ( .A1(n11879), .A2(n11799), .ZN(n11805) );
  NAND2_X1 U14738 ( .A1(n11800), .A2(n11805), .ZN(P2_U2958) );
  AOI22_X1 U14739 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14740 ( .A1(n15431), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15429), .ZN(n15460) );
  INV_X1 U14741 ( .A(n15460), .ZN(n14787) );
  NAND2_X1 U14742 ( .A1(n11879), .A2(n14787), .ZN(n11814) );
  NAND2_X1 U14743 ( .A1(n11801), .A2(n11814), .ZN(P2_U2974) );
  INV_X1 U14744 ( .A(n11853), .ZN(n11885) );
  INV_X1 U14745 ( .A(n11885), .ZN(n19101) );
  AOI22_X1 U14746 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14747 ( .A1(n15431), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15429), .ZN(n19158) );
  INV_X1 U14748 ( .A(n19158), .ZN(n11802) );
  NAND2_X1 U14749 ( .A1(n11879), .A2(n11802), .ZN(n11808) );
  NAND2_X1 U14750 ( .A1(n11803), .A2(n11808), .ZN(P2_U2955) );
  AOI22_X1 U14751 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U14752 ( .A1(n15431), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15429), .ZN(n19150) );
  INV_X1 U14753 ( .A(n19150), .ZN(n14817) );
  NAND2_X1 U14754 ( .A1(n11879), .A2(n14817), .ZN(n11812) );
  NAND2_X1 U14755 ( .A1(n11804), .A2(n11812), .ZN(P2_U2968) );
  AOI22_X1 U14756 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n11806) );
  NAND2_X1 U14757 ( .A1(n11806), .A2(n11805), .ZN(P2_U2973) );
  AOI22_X1 U14758 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14759 ( .A1(n15431), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15429), .ZN(n19166) );
  INV_X1 U14760 ( .A(n19166), .ZN(n14802) );
  NAND2_X1 U14761 ( .A1(n11879), .A2(n14802), .ZN(n11810) );
  NAND2_X1 U14762 ( .A1(n11807), .A2(n11810), .ZN(P2_U2957) );
  AOI22_X1 U14763 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n11809) );
  NAND2_X1 U14764 ( .A1(n11809), .A2(n11808), .ZN(P2_U2970) );
  AOI22_X1 U14765 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U14766 ( .A1(n11811), .A2(n11810), .ZN(P2_U2972) );
  AOI22_X1 U14767 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n11813) );
  NAND2_X1 U14768 ( .A1(n11813), .A2(n11812), .ZN(P2_U2953) );
  AOI22_X1 U14769 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11815) );
  NAND2_X1 U14770 ( .A1(n11815), .A2(n11814), .ZN(P2_U2959) );
  AOI22_X1 U14771 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n11819) );
  INV_X1 U14772 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n11816) );
  OR2_X1 U14773 ( .A1(n15429), .A2(n11816), .ZN(n11818) );
  NAND2_X1 U14774 ( .A1(n15429), .A2(BUF2_REG_9__SCAN_IN), .ZN(n11817) );
  NAND2_X1 U14775 ( .A1(n11818), .A2(n11817), .ZN(n14776) );
  NAND2_X1 U14776 ( .A1(n11879), .A2(n14776), .ZN(n11827) );
  NAND2_X1 U14777 ( .A1(n11819), .A2(n11827), .ZN(P2_U2961) );
  AOI22_X1 U14778 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11822) );
  INV_X1 U14779 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n12403) );
  OR2_X1 U14780 ( .A1(n15429), .A2(n12403), .ZN(n11821) );
  NAND2_X1 U14781 ( .A1(n15429), .A2(BUF2_REG_13__SCAN_IN), .ZN(n11820) );
  NAND2_X1 U14782 ( .A1(n11821), .A2(n11820), .ZN(n14738) );
  NAND2_X1 U14783 ( .A1(n11879), .A2(n14738), .ZN(n11831) );
  NAND2_X1 U14784 ( .A1(n11822), .A2(n11831), .ZN(P2_U2980) );
  AOI22_X1 U14785 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11826) );
  INV_X1 U14786 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n11823) );
  OR2_X1 U14787 ( .A1(n15429), .A2(n11823), .ZN(n11825) );
  NAND2_X1 U14788 ( .A1(n15429), .A2(BUF2_REG_11__SCAN_IN), .ZN(n11824) );
  NAND2_X1 U14789 ( .A1(n11825), .A2(n11824), .ZN(n14750) );
  NAND2_X1 U14790 ( .A1(n11879), .A2(n14750), .ZN(n11829) );
  NAND2_X1 U14791 ( .A1(n11826), .A2(n11829), .ZN(P2_U2978) );
  AOI22_X1 U14792 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11828) );
  NAND2_X1 U14793 ( .A1(n11828), .A2(n11827), .ZN(P2_U2976) );
  AOI22_X1 U14794 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11830) );
  NAND2_X1 U14795 ( .A1(n11830), .A2(n11829), .ZN(P2_U2963) );
  AOI22_X1 U14796 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11832) );
  NAND2_X1 U14797 ( .A1(n11832), .A2(n11831), .ZN(P2_U2965) );
  INV_X1 U14798 ( .A(n11833), .ZN(n11841) );
  OAI21_X1 U14799 ( .B1(n11835), .B2(n11841), .A(n11834), .ZN(n11836) );
  OAI21_X1 U14800 ( .B1(n12795), .B2(n15694), .A(n11836), .ZN(n19812) );
  NOR3_X1 U14801 ( .A1(n11837), .A2(n12795), .A3(n15720), .ZN(n11838) );
  INV_X1 U14802 ( .A(n20726), .ZN(n20635) );
  NOR2_X1 U14803 ( .A1(n11838), .A2(n20635), .ZN(n20728) );
  NOR2_X1 U14804 ( .A1(n19812), .A2(n20728), .ZN(n15681) );
  NOR2_X1 U14805 ( .A1(n15681), .A2(n19811), .ZN(n19819) );
  INV_X1 U14806 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n11850) );
  NAND2_X1 U14807 ( .A1(n12334), .A2(n15694), .ZN(n11845) );
  OAI21_X1 U14808 ( .B1(n20051), .B2(n11840), .A(n11839), .ZN(n11843) );
  AOI22_X1 U14809 ( .A1(n11843), .A2(n11842), .B1(n11271), .B2(n11841), .ZN(
        n11844) );
  NAND2_X1 U14810 ( .A1(n11845), .A2(n11844), .ZN(n11847) );
  NAND2_X1 U14811 ( .A1(n11847), .A2(n11846), .ZN(n15683) );
  INV_X1 U14812 ( .A(n15683), .ZN(n11848) );
  NAND2_X1 U14813 ( .A1(n19819), .A2(n11848), .ZN(n11849) );
  OAI21_X1 U14814 ( .B1(n19819), .B2(n11850), .A(n11849), .ZN(P1_U3484) );
  MUX2_X1 U14815 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n15429), .Z(n19016) );
  NAND2_X1 U14816 ( .A1(n11879), .A2(n19016), .ZN(n19102) );
  NAND2_X1 U14817 ( .A1(n19101), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n11851) );
  OAI211_X1 U14818 ( .C1(n11852), .C2(n11887), .A(n19102), .B(n11851), .ZN(
        P2_U2964) );
  AOI22_X1 U14819 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n11853), .B1(n19100), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n11854) );
  INV_X1 U14820 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16347) );
  INV_X1 U14821 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18068) );
  AOI22_X1 U14822 ( .A1(n15431), .A2(n16347), .B1(n18068), .B2(n15429), .ZN(
        n16115) );
  NAND2_X1 U14823 ( .A1(n11879), .A2(n16115), .ZN(n11855) );
  NAND2_X1 U14824 ( .A1(n11854), .A2(n11855), .ZN(P2_U2969) );
  AOI22_X1 U14825 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11856) );
  NAND2_X1 U14826 ( .A1(n11856), .A2(n11855), .ZN(P2_U2954) );
  AOI22_X1 U14827 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11857) );
  INV_X1 U14828 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16344) );
  INV_X1 U14829 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U14830 ( .A1(n15431), .A2(n16344), .B1(n18079), .B2(n15429), .ZN(
        n19028) );
  NAND2_X1 U14831 ( .A1(n11879), .A2(n19028), .ZN(n11858) );
  NAND2_X1 U14832 ( .A1(n11857), .A2(n11858), .ZN(P2_U2956) );
  AOI22_X1 U14833 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11859) );
  NAND2_X1 U14834 ( .A1(n11859), .A2(n11858), .ZN(P2_U2971) );
  OR2_X1 U14835 ( .A1(n15429), .A2(n11860), .ZN(n11862) );
  NAND2_X1 U14836 ( .A1(n15429), .A2(BUF2_REG_14__SCAN_IN), .ZN(n11861) );
  NAND2_X1 U14837 ( .A1(n11862), .A2(n11861), .ZN(n14048) );
  NAND2_X1 U14838 ( .A1(n11879), .A2(n14048), .ZN(n11873) );
  NAND2_X1 U14839 ( .A1(n19101), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n11863) );
  OAI211_X1 U14840 ( .C1(n11864), .C2(n11887), .A(n11873), .B(n11863), .ZN(
        P2_U2966) );
  INV_X1 U14841 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19076) );
  INV_X1 U14842 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n21043) );
  OR2_X1 U14843 ( .A1(n15429), .A2(n21043), .ZN(n11866) );
  NAND2_X1 U14844 ( .A1(n15429), .A2(BUF2_REG_10__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U14845 ( .A1(n11866), .A2(n11865), .ZN(n19019) );
  NAND2_X1 U14846 ( .A1(n11879), .A2(n19019), .ZN(n11877) );
  NAND2_X1 U14847 ( .A1(n19101), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n11867) );
  OAI211_X1 U14848 ( .C1(n19076), .C2(n11887), .A(n11877), .B(n11867), .ZN(
        P2_U2977) );
  INV_X1 U14849 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16338) );
  OR2_X1 U14850 ( .A1(n15429), .A2(n16338), .ZN(n11869) );
  NAND2_X1 U14851 ( .A1(n15429), .A2(BUF2_REG_8__SCAN_IN), .ZN(n11868) );
  NAND2_X1 U14852 ( .A1(n11869), .A2(n11868), .ZN(n14780) );
  NAND2_X1 U14853 ( .A1(n11879), .A2(n14780), .ZN(n11875) );
  NAND2_X1 U14854 ( .A1(n19101), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n11870) );
  OAI211_X1 U14855 ( .C1(n11871), .C2(n11887), .A(n11875), .B(n11870), .ZN(
        P2_U2960) );
  INV_X1 U14856 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19069) );
  NAND2_X1 U14857 ( .A1(n19101), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n11872) );
  OAI211_X1 U14858 ( .C1(n19069), .C2(n11887), .A(n11873), .B(n11872), .ZN(
        P2_U2981) );
  INV_X1 U14859 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19079) );
  NAND2_X1 U14860 ( .A1(n19101), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n11874) );
  OAI211_X1 U14861 ( .C1(n19079), .C2(n11887), .A(n11875), .B(n11874), .ZN(
        P2_U2975) );
  NAND2_X1 U14862 ( .A1(n19101), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n11876) );
  OAI211_X1 U14863 ( .C1(n11878), .C2(n11887), .A(n11877), .B(n11876), .ZN(
        P2_U2962) );
  INV_X1 U14864 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16353) );
  INV_X1 U14865 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18054) );
  AOI22_X1 U14866 ( .A1(n15431), .A2(n16353), .B1(n18054), .B2(n15429), .ZN(
        n19004) );
  INV_X1 U14867 ( .A(n19004), .ZN(n15439) );
  INV_X1 U14868 ( .A(n11879), .ZN(n11884) );
  INV_X1 U14869 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n11881) );
  OAI222_X1 U14870 ( .A1(n15439), .A2(n11884), .B1(n11881), .B2(n11885), .C1(
        n11887), .C2(n11880), .ZN(P2_U2952) );
  INV_X1 U14871 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n11883) );
  INV_X1 U14872 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U14873 ( .A1(n15431), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15429), .ZN(n19015) );
  OAI222_X1 U14874 ( .A1(n11887), .A2(n11883), .B1(n11882), .B2(n11885), .C1(
        n11884), .C2(n19015), .ZN(P2_U2982) );
  INV_X1 U14875 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11888) );
  INV_X1 U14876 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n11886) );
  OAI222_X1 U14877 ( .A1(n11888), .A2(n11887), .B1(n11886), .B2(n11885), .C1(
        n11884), .C2(n15439), .ZN(P2_U2967) );
  NAND2_X1 U14878 ( .A1(n15669), .A2(n15720), .ZN(n12343) );
  NAND2_X1 U14879 ( .A1(n11889), .A2(n15720), .ZN(n11890) );
  NOR2_X1 U14880 ( .A1(n12342), .A2(n11890), .ZN(n15693) );
  INV_X1 U14881 ( .A(n15693), .ZN(n11891) );
  NAND2_X1 U14882 ( .A1(n12343), .A2(n11891), .ZN(n11894) );
  OR2_X1 U14883 ( .A1(n19952), .A2(n20051), .ZN(n19920) );
  INV_X1 U14884 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n20828) );
  INV_X1 U14885 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n20948) );
  NAND2_X1 U14886 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16039) );
  OR2_X1 U14887 ( .A1(n16039), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19928) );
  INV_X1 U14888 ( .A(P1_UWORD_REG_4__SCAN_IN), .ZN(n20989) );
  OAI22_X1 U14889 ( .A1(n20948), .A2(n19925), .B1(n20989), .B2(n19928), .ZN(
        n11895) );
  INV_X1 U14890 ( .A(n11895), .ZN(n11896) );
  OAI21_X1 U14891 ( .B1(n19920), .B2(n20828), .A(n11896), .ZN(P1_U2916) );
  NOR2_X1 U14892 ( .A1(n11905), .A2(n15433), .ZN(n11899) );
  INV_X1 U14893 ( .A(n11901), .ZN(n11902) );
  AND2_X2 U14894 ( .A1(n11903), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U14895 ( .A1(n12073), .A2(n12483), .ZN(n12103) );
  AND2_X2 U14896 ( .A1(n11917), .A2(n11929), .ZN(n11906) );
  AOI21_X2 U14897 ( .B1(n12462), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11906), .ZN(n12030) );
  INV_X4 U14898 ( .A(n12736), .ZN(n13598) );
  INV_X1 U14899 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11909) );
  INV_X1 U14900 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n11908) );
  OAI22_X1 U14901 ( .A1(n13598), .A2(n11909), .B1(n13585), .B2(n11908), .ZN(
        n11927) );
  NAND2_X1 U14902 ( .A1(n12053), .A2(n12105), .ZN(n11914) );
  MUX2_X1 U14903 ( .A(n12038), .B(n12483), .S(n11910), .Z(n11913) );
  AND2_X1 U14904 ( .A1(n11911), .A2(n15443), .ZN(n11912) );
  NAND3_X1 U14905 ( .A1(n11914), .A2(n11913), .A3(n11912), .ZN(n11915) );
  NAND3_X1 U14906 ( .A1(n11915), .A2(n12075), .A3(n15479), .ZN(n12102) );
  INV_X1 U14907 ( .A(n12102), .ZN(n11916) );
  NAND2_X1 U14908 ( .A1(n11916), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11925) );
  NAND2_X1 U14909 ( .A1(n11917), .A2(n12075), .ZN(n11924) );
  NAND2_X1 U14910 ( .A1(n11919), .A2(n11918), .ZN(n12005) );
  NAND3_X1 U14911 ( .A1(n12005), .A2(n15443), .A3(n13271), .ZN(n11921) );
  NAND2_X1 U14912 ( .A1(n11921), .A2(n11920), .ZN(n12116) );
  INV_X1 U14913 ( .A(n12116), .ZN(n11922) );
  NAND2_X1 U14914 ( .A1(n11922), .A2(n11907), .ZN(n11923) );
  INV_X1 U14915 ( .A(n11930), .ZN(n11926) );
  OAI21_X1 U14916 ( .B1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n15409), .A(
        n12965), .ZN(n11928) );
  NAND3_X1 U14917 ( .A1(n12030), .A2(n12023), .A3(n11928), .ZN(n11936) );
  NAND2_X1 U14918 ( .A1(n12467), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11934) );
  INV_X1 U14919 ( .A(n12652), .ZN(n11932) );
  NAND2_X1 U14920 ( .A1(n11932), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12028) );
  NOR2_X1 U14921 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12718) );
  NAND2_X1 U14922 ( .A1(n12718), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11933) );
  NAND4_X1 U14923 ( .A1(n11934), .A2(n13598), .A3(n12028), .A4(n11933), .ZN(
        n11935) );
  NAND2_X1 U14924 ( .A1(n12467), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11940) );
  NAND2_X2 U14925 ( .A1(n11938), .A2(n10287), .ZN(n12668) );
  AOI22_X1 U14926 ( .A1(n12668), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n12718), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U14927 ( .A1(n11940), .A2(n11939), .ZN(n12435) );
  NAND2_X1 U14928 ( .A1(n13595), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11942) );
  INV_X1 U14929 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14697) );
  XNOR2_X1 U14930 ( .A(n12435), .B(n12436), .ZN(n12434) );
  XNOR2_X1 U14931 ( .A(n12433), .B(n13231), .ZN(n12426) );
  AOI21_X1 U14932 ( .B1(n15409), .B2(n19390), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n14526) );
  NAND2_X1 U14933 ( .A1(n14526), .A2(n16225), .ZN(n11944) );
  INV_X1 U14934 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12944) );
  AND2_X1 U14935 ( .A1(n11946), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12205) );
  AND2_X1 U14936 ( .A1(n14034), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12206) );
  AOI22_X1 U14937 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12205), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11954) );
  AND2_X1 U14938 ( .A1(n11946), .A2(n12694), .ZN(n12170) );
  AND2_X1 U14939 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U14940 ( .A1(n12170), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n13836), .ZN(n11953) );
  BUF_X1 U14941 ( .A(n13767), .Z(n11949) );
  AND2_X2 U14942 ( .A1(n11949), .A2(n12694), .ZN(n12279) );
  AND2_X2 U14943 ( .A1(n11949), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12200) );
  AOI22_X1 U14944 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12279), .B1(
        n12200), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11952) );
  AND2_X2 U14945 ( .A1(n14030), .A2(n12694), .ZN(n13791) );
  AOI22_X1 U14946 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11951) );
  NAND4_X1 U14947 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11962) );
  AND2_X1 U14948 ( .A1(n14034), .A2(n12694), .ZN(n11986) );
  AOI22_X1 U14949 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11960) );
  AND2_X1 U14950 ( .A1(n13768), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12165) );
  AOI22_X1 U14951 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n12165), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U14952 ( .A1(n13837), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11958) );
  AND2_X2 U14953 ( .A1(n14036), .A2(n12694), .ZN(n12654) );
  AOI22_X1 U14954 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11957) );
  MUX2_X1 U14955 ( .A(n13294), .B(P2_EBX_REG_1__SCAN_IN), .S(n13502), .Z(
        n11964) );
  INV_X1 U14956 ( .A(n11964), .ZN(n11965) );
  NAND2_X1 U14957 ( .A1(n13502), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11966) );
  INV_X1 U14958 ( .A(n11966), .ZN(n11980) );
  NAND2_X1 U14959 ( .A1(n11980), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11967) );
  AND2_X1 U14960 ( .A1(n13065), .A2(n11967), .ZN(n14693) );
  AOI22_X1 U14961 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U14962 ( .A1(n13837), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U14963 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U14964 ( .A1(n12279), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13836), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11968) );
  NAND4_X1 U14965 ( .A1(n11971), .A2(n11970), .A3(n11969), .A4(n11968), .ZN(
        n11977) );
  AOI22_X1 U14966 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11985), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U14967 ( .A1(n12152), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U14968 ( .A1(n12205), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U14969 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11972) );
  NAND4_X1 U14970 ( .A1(n11975), .A2(n11974), .A3(n11973), .A4(n11972), .ZN(
        n11976) );
  NOR2_X1 U14971 ( .A1(n11977), .A2(n11976), .ZN(n12055) );
  NOR2_X1 U14972 ( .A1(n12948), .A2(n13502), .ZN(n13041) );
  INV_X1 U14973 ( .A(n13041), .ZN(n11978) );
  OR2_X1 U14974 ( .A1(n12055), .A2(n11978), .ZN(n11982) );
  AND2_X1 U14975 ( .A1(n11979), .A2(n12948), .ZN(n13039) );
  AOI21_X1 U14976 ( .B1(n13039), .B2(n12008), .A(n11980), .ZN(n11981) );
  NAND2_X1 U14977 ( .A1(n11982), .A2(n11981), .ZN(n18953) );
  NAND2_X1 U14978 ( .A1(n18953), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13333) );
  XOR2_X1 U14979 ( .A(n14693), .B(n13333), .Z(n11983) );
  NOR2_X1 U14980 ( .A1(n12944), .A2(n11983), .ZN(n13334) );
  AOI21_X1 U14981 ( .B1(n12944), .B2(n11983), .A(n13334), .ZN(n15398) );
  AOI22_X1 U14982 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11985), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U14983 ( .A1(n13837), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U14984 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11986), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U14985 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12205), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11987) );
  NAND4_X1 U14986 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11996) );
  AOI22_X1 U14987 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12151), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U14988 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12279), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U14989 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n13836), .ZN(n11992) );
  AOI22_X1 U14990 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13791), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11991) );
  NAND4_X1 U14991 ( .A1(n11994), .A2(n11993), .A3(n11992), .A4(n11991), .ZN(
        n11995) );
  NAND2_X1 U14992 ( .A1(n12948), .A2(n11997), .ZN(n11998) );
  NAND2_X1 U14993 ( .A1(n12008), .A2(n11999), .ZN(n12000) );
  NAND2_X1 U14994 ( .A1(n12954), .A2(n12000), .ZN(n12004) );
  INV_X1 U14995 ( .A(n12001), .ZN(n12003) );
  AOI21_X1 U14996 ( .B1(n12004), .B2(n12003), .A(n12002), .ZN(n19801) );
  AND2_X1 U14997 ( .A1(n10055), .A2(n15433), .ZN(n12079) );
  INV_X1 U14998 ( .A(n12079), .ZN(n12006) );
  NOR2_X1 U14999 ( .A1(n12005), .A2(n12006), .ZN(n19796) );
  NAND2_X1 U15000 ( .A1(n19801), .A2(n19796), .ZN(n12012) );
  INV_X1 U15001 ( .A(n12005), .ZN(n12709) );
  AOI21_X1 U15002 ( .B1(n12008), .B2(n12007), .A(n12697), .ZN(n12009) );
  INV_X1 U15003 ( .A(n12009), .ZN(n12010) );
  INV_X1 U15004 ( .A(n12165), .ZN(n13794) );
  AOI21_X1 U15005 ( .B1(n11947), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15477) );
  AOI21_X1 U15006 ( .B1(n13794), .B2(n15477), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n16226) );
  MUX2_X1 U15007 ( .A(n12010), .B(n16226), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n15738) );
  INV_X1 U15008 ( .A(n15738), .ZN(n19798) );
  NAND3_X1 U15009 ( .A1(n12709), .A2(n19798), .A3(n14018), .ZN(n12011) );
  NAND2_X1 U15010 ( .A1(n12012), .A2(n12011), .ZN(n12090) );
  AND2_X1 U15011 ( .A1(n15433), .A2(n12788), .ZN(n12013) );
  NAND2_X1 U15012 ( .A1(n12090), .A2(n12013), .ZN(n18736) );
  XOR2_X1 U15013 ( .A(n12055), .B(n13294), .Z(n13515) );
  OR2_X1 U15014 ( .A1(n12055), .A2(n14018), .ZN(n13295) );
  NAND2_X1 U15015 ( .A1(n13295), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13514) );
  XNOR2_X1 U15016 ( .A(n13515), .B(n13514), .ZN(n12014) );
  NAND2_X1 U15017 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12014), .ZN(
        n13517) );
  OAI21_X1 U15018 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12014), .A(
        n13517), .ZN(n15395) );
  OR2_X1 U15019 ( .A1(n19771), .A2(n19764), .ZN(n19790) );
  NAND2_X1 U15020 ( .A1(n19790), .A2(n12943), .ZN(n12015) );
  INV_X1 U15021 ( .A(n12475), .ZN(n12017) );
  NAND2_X1 U15022 ( .A1(n19574), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U15023 ( .A1(n12017), .A2(n12016), .ZN(n12034) );
  MUX2_X1 U15024 ( .A(n19120), .B(n16186), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n12020) );
  INV_X2 U15025 ( .A(n18885), .ZN(n18905) );
  INV_X1 U15026 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19696) );
  AND2_X1 U15027 ( .A1(n19132), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15397) );
  INV_X1 U15028 ( .A(n15397), .ZN(n12019) );
  OAI211_X1 U15029 ( .C1(n15395), .C2(n16181), .A(n12020), .B(n12019), .ZN(
        n12021) );
  AOI21_X1 U15030 ( .B1(n15398), .B2(n19116), .A(n12021), .ZN(n12022) );
  OAI21_X1 U15031 ( .B1(n14698), .B2(n15430), .A(n12022), .ZN(P2_U3013) );
  INV_X1 U15032 ( .A(n12023), .ZN(n12027) );
  INV_X1 U15033 ( .A(n12718), .ZN(n12025) );
  NAND2_X1 U15034 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12024) );
  NAND3_X1 U15035 ( .A1(n13598), .A2(n12025), .A3(n12024), .ZN(n12026) );
  NAND3_X1 U15036 ( .A1(n12030), .A2(n12029), .A3(n12028), .ZN(n12031) );
  AND2_X2 U15037 ( .A1(n12433), .A2(n12031), .ZN(n12037) );
  OAI21_X1 U15038 ( .B1(n13295), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13514), .ZN(n12124) );
  INV_X1 U15039 ( .A(n12124), .ZN(n12033) );
  OAI21_X1 U15040 ( .B1(n18953), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13333), .ZN(n12114) );
  NAND2_X1 U15041 ( .A1(n18885), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12121) );
  OAI21_X1 U15042 ( .B1(n16179), .B2(n12114), .A(n12121), .ZN(n12032) );
  AOI21_X1 U15043 ( .B1(n19115), .B2(n12033), .A(n12032), .ZN(n12036) );
  OAI21_X1 U15044 ( .B1(n19104), .B2(n12034), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12035) );
  OAI211_X1 U15045 ( .C1(n18958), .C2(n15430), .A(n12036), .B(n12035), .ZN(
        P2_U3014) );
  NAND2_X1 U15046 ( .A1(n12038), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15047 ( .A1(n12473), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19771), .B2(n19794), .ZN(n12040) );
  NAND2_X1 U15048 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12044) );
  AND4_X1 U15049 ( .A1(n12043), .A2(n12044), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19616), .ZN(n12045) );
  NAND2_X1 U15050 ( .A1(n12047), .A2(n12046), .ZN(n12663) );
  NAND3_X1 U15051 ( .A1(n11979), .A2(n10055), .A3(n15443), .ZN(n12048) );
  NAND2_X1 U15052 ( .A1(n11897), .A2(n15735), .ZN(n12702) );
  NOR2_X1 U15053 ( .A1(n12704), .A2(n12702), .ZN(n12049) );
  AOI21_X1 U15054 ( .B1(n12701), .B2(n12696), .A(n12049), .ZN(n12646) );
  NAND2_X1 U15055 ( .A1(n12050), .A2(n9900), .ZN(n12051) );
  NAND2_X1 U15056 ( .A1(n12646), .A2(n12051), .ZN(n12052) );
  AOI21_X1 U15057 ( .B1(n19030), .B2(n19038), .A(n19057), .ZN(n12070) );
  NOR2_X1 U15058 ( .A1(n11963), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12054) );
  AND2_X1 U15059 ( .A1(n12483), .A2(n19616), .ZN(n12184) );
  INV_X1 U15060 ( .A(n12184), .ZN(n12056) );
  OAI21_X1 U15061 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19616), .A(
        n12056), .ZN(n12057) );
  AND2_X1 U15062 ( .A1(n12057), .A2(n12190), .ZN(n12058) );
  NAND3_X1 U15063 ( .A1(n12184), .A2(n10055), .A3(n11963), .ZN(n12150) );
  AOI21_X1 U15064 ( .B1(n14018), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12061) );
  OAI211_X1 U15065 ( .C1(n12150), .C2(n11908), .A(n12061), .B(n12060), .ZN(
        n12062) );
  NOR2_X1 U15066 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  NOR2_X1 U15067 ( .A1(n12189), .A2(n12064), .ZN(n18951) );
  INV_X1 U15068 ( .A(n18951), .ZN(n19029) );
  NOR3_X1 U15069 ( .A1(n19030), .A2(n18951), .A3(n19061), .ZN(n12065) );
  AOI21_X1 U15070 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19056), .A(n12065), .ZN(
        n12069) );
  NAND2_X1 U15071 ( .A1(n13502), .A2(n12483), .ZN(n12066) );
  OR2_X1 U15072 ( .A1(n19056), .A2(n12066), .ZN(n14811) );
  NAND2_X1 U15073 ( .A1(n12038), .A2(n12483), .ZN(n12067) );
  OR2_X1 U15074 ( .A1(n19056), .A2(n12067), .ZN(n14049) );
  INV_X1 U15075 ( .A(n19065), .ZN(n19020) );
  NAND2_X1 U15076 ( .A1(n19020), .A2(n19004), .ZN(n12068) );
  OAI211_X1 U15077 ( .C1(n12070), .C2(n19029), .A(n12069), .B(n12068), .ZN(
        P2_U2919) );
  INV_X1 U15078 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15408) );
  NOR2_X1 U15079 ( .A1(n19681), .A2(n19680), .ZN(n12716) );
  NAND2_X1 U15080 ( .A1(n12099), .A2(n12716), .ZN(n12094) );
  AOI21_X1 U15081 ( .B1(n12071), .B2(n12075), .A(n19162), .ZN(n12072) );
  NAND2_X1 U15082 ( .A1(n12647), .A2(n12072), .ZN(n12093) );
  NAND2_X1 U15083 ( .A1(n12073), .A2(n15443), .ZN(n12074) );
  NAND2_X1 U15084 ( .A1(n12074), .A2(n11900), .ZN(n12086) );
  OAI21_X1 U15085 ( .B1(n19162), .B2(n14018), .A(n12075), .ZN(n12076) );
  NAND2_X1 U15086 ( .A1(n12076), .A2(n12483), .ZN(n12077) );
  AOI21_X1 U15087 ( .B1(n12077), .B2(n15443), .A(n9864), .ZN(n12081) );
  NAND2_X1 U15088 ( .A1(n12078), .A2(n12483), .ZN(n12080) );
  NAND2_X1 U15089 ( .A1(n12080), .A2(n12079), .ZN(n12104) );
  AND2_X1 U15090 ( .A1(n12081), .A2(n12104), .ZN(n12085) );
  NAND3_X1 U15091 ( .A1(n12082), .A2(n12083), .A3(n12716), .ZN(n12084) );
  AND3_X1 U15092 ( .A1(n12086), .A2(n12085), .A3(n12084), .ZN(n12644) );
  MUX2_X1 U15093 ( .A(n12082), .B(n12099), .S(n10055), .Z(n12088) );
  NOR2_X1 U15094 ( .A1(n12697), .A2(n19680), .ZN(n12087) );
  NAND2_X1 U15095 ( .A1(n12088), .A2(n12087), .ZN(n12089) );
  NAND2_X1 U15096 ( .A1(n12644), .A2(n12089), .ZN(n12091) );
  NOR2_X1 U15097 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  OAI211_X1 U15098 ( .C1(n12647), .C2(n12094), .A(n12093), .B(n12092), .ZN(
        n12095) );
  NAND2_X1 U15099 ( .A1(n12097), .A2(n11897), .ZN(n12098) );
  NAND2_X1 U15100 ( .A1(n12098), .A2(n9864), .ZN(n12109) );
  INV_X1 U15101 ( .A(n11897), .ZN(n12100) );
  AOI22_X1 U15102 ( .A1(n12100), .A2(n11910), .B1(n15433), .B2(n12099), .ZN(
        n12101) );
  AND2_X1 U15103 ( .A1(n12102), .A2(n12101), .ZN(n12108) );
  NAND2_X1 U15104 ( .A1(n12103), .A2(n14018), .ZN(n12664) );
  NAND2_X1 U15105 ( .A1(n12664), .A2(n12104), .ZN(n12106) );
  NAND2_X1 U15106 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  INV_X1 U15107 ( .A(n9802), .ZN(n12110) );
  NAND2_X1 U15108 ( .A1(n12689), .A2(n12110), .ZN(n12111) );
  NAND2_X1 U15109 ( .A1(n12123), .A2(n12111), .ZN(n13654) );
  NAND2_X1 U15110 ( .A1(n12668), .A2(n10055), .ZN(n12112) );
  NAND2_X1 U15111 ( .A1(n12112), .A2(n12652), .ZN(n12113) );
  NAND2_X1 U15112 ( .A1(n12123), .A2(n12113), .ZN(n16191) );
  NOR2_X1 U15113 ( .A1(n12005), .A2(n12948), .ZN(n19797) );
  INV_X1 U15114 ( .A(n12114), .ZN(n12120) );
  AND2_X1 U15115 ( .A1(n12116), .A2(n12115), .ZN(n12698) );
  INV_X1 U15116 ( .A(n12698), .ZN(n12118) );
  NAND2_X1 U15117 ( .A1(n11937), .A2(n14018), .ZN(n12117) );
  NAND2_X1 U15118 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  AOI22_X1 U15119 ( .A1(n19130), .A2(n12120), .B1(n19126), .B2(n18951), .ZN(
        n12122) );
  OAI211_X1 U15120 ( .C1(n16191), .C2(n18958), .A(n12122), .B(n12121), .ZN(
        n12126) );
  NOR2_X1 U15121 ( .A1(n12123), .A2(n18885), .ZN(n15399) );
  INV_X1 U15122 ( .A(n15399), .ZN(n13657) );
  NAND2_X1 U15123 ( .A1(n12123), .A2(n19796), .ZN(n16212) );
  OAI22_X1 U15124 ( .A1(n13657), .A2(n15408), .B1(n16212), .B2(n12124), .ZN(
        n12125) );
  AOI211_X1 U15125 ( .C1(n15408), .C2(n15402), .A(n12126), .B(n12125), .ZN(
        n12127) );
  INV_X1 U15126 ( .A(n12127), .ZN(P2_U3046) );
  INV_X1 U15127 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12129) );
  INV_X2 U15128 ( .A(n19928), .ZN(n20727) );
  AOI22_X1 U15129 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12128) );
  OAI21_X1 U15130 ( .B1(n12129), .B2(n19920), .A(n12128), .ZN(P1_U2912) );
  INV_X1 U15131 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15132 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12130) );
  OAI21_X1 U15133 ( .B1(n12131), .B2(n19920), .A(n12130), .ZN(P1_U2913) );
  INV_X1 U15134 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n20884) );
  AOI22_X1 U15135 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12132) );
  OAI21_X1 U15136 ( .B1(n20884), .B2(n19920), .A(n12132), .ZN(P1_U2914) );
  INV_X1 U15137 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15138 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12133) );
  OAI21_X1 U15139 ( .B1(n12134), .B2(n19920), .A(n12133), .ZN(P1_U2911) );
  INV_X1 U15140 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15141 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12135) );
  OAI21_X1 U15142 ( .B1(n12136), .B2(n19920), .A(n12135), .ZN(P1_U2917) );
  INV_X1 U15143 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15144 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12137) );
  OAI21_X1 U15145 ( .B1(n12138), .B2(n19920), .A(n12137), .ZN(P1_U2920) );
  INV_X1 U15146 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14212) );
  AOI22_X1 U15147 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12139) );
  OAI21_X1 U15148 ( .B1(n14212), .B2(n19920), .A(n12139), .ZN(P1_U2907) );
  INV_X1 U15149 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15150 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12140) );
  OAI21_X1 U15151 ( .B1(n12141), .B2(n19920), .A(n12140), .ZN(P1_U2908) );
  AOI22_X1 U15152 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12142) );
  OAI21_X1 U15153 ( .B1(n14258), .B2(n19920), .A(n12142), .ZN(P1_U2919) );
  INV_X1 U15154 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15155 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12143) );
  OAI21_X1 U15156 ( .B1(n12144), .B2(n19920), .A(n12143), .ZN(P1_U2910) );
  INV_X1 U15157 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15158 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n12145) );
  OAI21_X1 U15159 ( .B1(n12146), .B2(n19920), .A(n12145), .ZN(P1_U2918) );
  INV_X1 U15160 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15161 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12147) );
  OAI21_X1 U15162 ( .B1(n12148), .B2(n19920), .A(n12147), .ZN(P1_U2909) );
  AOI22_X1 U15163 ( .A1(n20727), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n19950), .ZN(n12149) );
  OAI21_X1 U15164 ( .B1(n19920), .B2(n14245), .A(n12149), .ZN(P1_U2915) );
  INV_X1 U15165 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15380) );
  NOR2_X1 U15166 ( .A1(n12483), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15167 ( .A1(n13625), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13624), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15168 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12151), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15169 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13836), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15170 ( .A1(n12279), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15171 ( .A1(n12152), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U15172 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12162) );
  AOI22_X1 U15173 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11985), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15174 ( .A1(n13837), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15175 ( .A1(n11986), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15176 ( .A1(n12170), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12157) );
  NAND4_X1 U15177 ( .A1(n12160), .A2(n12159), .A3(n12158), .A4(n12157), .ZN(
        n12161) );
  NOR2_X1 U15178 ( .A1(n12162), .A2(n12161), .ZN(n13320) );
  OR2_X1 U15179 ( .A1(n12771), .A2(n13320), .ZN(n12163) );
  OAI211_X1 U15180 ( .C1(n13621), .C2(n15380), .A(n12164), .B(n12163), .ZN(
        n15377) );
  INV_X1 U15181 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15182 ( .A1(n13625), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13624), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15183 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12200), .B1(
        n12151), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15184 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n13836), .ZN(n12168) );
  AOI22_X1 U15185 ( .A1(n12279), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15186 ( .A1(n12152), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U15187 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12176) );
  AOI22_X1 U15188 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11985), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15189 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15190 ( .A1(n12206), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15191 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12170), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12171) );
  NAND4_X1 U15192 ( .A1(n12174), .A2(n12173), .A3(n12172), .A4(n12171), .ZN(
        n12175) );
  OR2_X1 U15193 ( .A1(n12771), .A2(n13298), .ZN(n12177) );
  OAI211_X1 U15194 ( .C1(n13621), .C2(n12179), .A(n12178), .B(n12177), .ZN(
        n12180) );
  INV_X1 U15195 ( .A(n12180), .ZN(n18921) );
  AOI22_X1 U15196 ( .A1(n12181), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12197), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12182) );
  OAI21_X1 U15197 ( .B1(n13621), .B2(n19696), .A(n12182), .ZN(n12188) );
  INV_X1 U15198 ( .A(n12188), .ZN(n12183) );
  XNOR2_X1 U15199 ( .A(n12189), .B(n12183), .ZN(n14688) );
  OR2_X1 U15200 ( .A1(n13294), .A2(n12771), .ZN(n12186) );
  AOI22_X1 U15201 ( .A1(n12053), .A2(n12184), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12185) );
  NAND2_X1 U15202 ( .A1(n12186), .A2(n12185), .ZN(n14689) );
  INV_X1 U15203 ( .A(n14689), .ZN(n12187) );
  NAND2_X1 U15204 ( .A1(n14688), .A2(n12187), .ZN(n14692) );
  OR2_X1 U15205 ( .A1(n12189), .A2(n12188), .ZN(n12193) );
  INV_X1 U15206 ( .A(n13296), .ZN(n13520) );
  OR2_X1 U15207 ( .A1(n12771), .A2(n13520), .ZN(n12191) );
  OAI211_X1 U15208 ( .C1(n19616), .C2(n19777), .A(n12191), .B(n12190), .ZN(
        n12192) );
  AND3_X1 U15209 ( .A1(n14692), .A2(n12193), .A3(n12192), .ZN(n12194) );
  INV_X1 U15210 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19697) );
  AOI22_X1 U15211 ( .A1(n13625), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13624), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12195) );
  OAI21_X1 U15212 ( .B1(n13621), .B2(n19697), .A(n12195), .ZN(n13059) );
  NOR2_X1 U15213 ( .A1(n13060), .A2(n13059), .ZN(n13061) );
  NOR2_X1 U15214 ( .A1(n12196), .A2(n13061), .ZN(n12963) );
  INV_X1 U15215 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15216 ( .A1(n13624), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12198) );
  OAI21_X1 U15217 ( .B1(n13621), .B2(n12199), .A(n12198), .ZN(n12215) );
  AOI22_X1 U15218 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12151), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15219 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12279), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15220 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n13836), .ZN(n12202) );
  AOI22_X1 U15221 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13791), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12201) );
  NAND4_X1 U15222 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12212) );
  AOI22_X1 U15223 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11985), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15224 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15225 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12170), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15226 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n12205), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12207) );
  NAND4_X1 U15227 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(
        n12211) );
  NAND2_X1 U15228 ( .A1(n13625), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12213) );
  OAI21_X1 U15229 ( .B1(n12771), .B2(n12955), .A(n12213), .ZN(n12214) );
  NAND2_X1 U15230 ( .A1(n12963), .A2(n12964), .ZN(n12962) );
  NAND2_X1 U15231 ( .A1(n15377), .A2(n18922), .ZN(n12227) );
  AOI22_X1 U15232 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15233 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n13836), .ZN(n12218) );
  AOI22_X1 U15234 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15235 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12216) );
  NAND4_X1 U15236 ( .A1(n12219), .A2(n12218), .A3(n12217), .A4(n12216), .ZN(
        n12225) );
  AOI22_X1 U15237 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15238 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15239 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11986), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15240 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12654), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12220) );
  NAND4_X1 U15241 ( .A1(n12223), .A2(n12222), .A3(n12221), .A4(n12220), .ZN(
        n12224) );
  INV_X1 U15242 ( .A(n13046), .ZN(n13376) );
  OR2_X1 U15243 ( .A1(n12771), .A2(n13376), .ZN(n12226) );
  NAND2_X1 U15244 ( .A1(n12227), .A2(n12226), .ZN(n12246) );
  INV_X1 U15245 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19702) );
  AOI22_X1 U15246 ( .A1(n13625), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13624), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12228) );
  OAI21_X1 U15247 ( .B1(n13621), .B2(n19702), .A(n12228), .ZN(n12245) );
  NAND2_X1 U15248 ( .A1(n12246), .A2(n12245), .ZN(n12240) );
  AOI22_X1 U15249 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15250 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n13836), .ZN(n12231) );
  AOI22_X1 U15251 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15252 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12229) );
  NAND4_X1 U15253 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12238) );
  AOI22_X1 U15254 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15255 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15256 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11986), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15257 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12206), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12233) );
  NAND4_X1 U15258 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n12237) );
  OR2_X1 U15259 ( .A1(n12771), .A2(n13543), .ZN(n12239) );
  INV_X1 U15260 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19703) );
  AOI22_X1 U15261 ( .A1(n13625), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13624), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12241) );
  OAI21_X1 U15262 ( .B1(n13621), .B2(n19703), .A(n12241), .ZN(n12242) );
  OR2_X1 U15263 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  NAND2_X1 U15264 ( .A1(n12244), .A2(n12294), .ZN(n18888) );
  OR2_X1 U15265 ( .A1(n19038), .A2(n19057), .ZN(n19025) );
  INV_X1 U15266 ( .A(n19025), .ZN(n19023) );
  INV_X1 U15267 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19081) );
  OAI222_X1 U15268 ( .A1(n18888), .A2(n19023), .B1(n15460), .B2(n19065), .C1(
        n19081), .C2(n14810), .ZN(P2_U2912) );
  XNOR2_X1 U15269 ( .A(n12246), .B(n12245), .ZN(n18904) );
  INV_X1 U15270 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19083) );
  OAI222_X1 U15271 ( .A1(n18904), .A2(n19023), .B1(n14810), .B2(n19083), .C1(
        n19065), .C2(n19176), .ZN(P2_U2913) );
  AND2_X1 U15272 ( .A1(n20729), .A2(n20635), .ZN(n12247) );
  OR2_X1 U15273 ( .A1(n9795), .A2(n10434), .ZN(n12394) );
  INV_X1 U15274 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19926) );
  NOR2_X2 U15275 ( .A1(n9795), .A2(n20066), .ZN(n19969) );
  INV_X1 U15276 ( .A(n19969), .ZN(n12251) );
  INV_X1 U15277 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12249) );
  NOR2_X1 U15278 ( .A1(n20043), .A2(n12249), .ZN(n12250) );
  AOI21_X1 U15279 ( .B1(DATAI_15_), .B2(n20043), .A(n12250), .ZN(n14269) );
  INV_X1 U15280 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19927) );
  OAI222_X1 U15281 ( .A1(n12394), .A2(n19926), .B1(n12251), .B2(n14269), .C1(
        n12320), .C2(n19927), .ZN(P1_U2967) );
  INV_X1 U15282 ( .A(n12252), .ZN(n12255) );
  OAI21_X1 U15283 ( .B1(n12255), .B2(n12254), .A(n12253), .ZN(n12825) );
  NAND2_X1 U15284 ( .A1(n12256), .A2(n15871), .ZN(n12260) );
  AND2_X1 U15285 ( .A1(n20033), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n12265) );
  OAI21_X1 U15286 ( .B1(n12258), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12257), .ZN(n12271) );
  NOR2_X1 U15287 ( .A1(n12271), .A2(n19817), .ZN(n12259) );
  AOI211_X1 U15288 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n12260), .A(
        n12265), .B(n12259), .ZN(n12261) );
  OAI21_X1 U15289 ( .B1(n20044), .B2(n12825), .A(n12261), .ZN(P1_U2999) );
  AOI21_X1 U15290 ( .B1(n15969), .B2(n14506), .A(n20023), .ZN(n12268) );
  NAND2_X1 U15291 ( .A1(n12262), .A2(n20023), .ZN(n12264) );
  AND2_X1 U15292 ( .A1(n12264), .A2(n12263), .ZN(n12820) );
  INV_X1 U15293 ( .A(n12820), .ZN(n12559) );
  INV_X1 U15294 ( .A(n12265), .ZN(n12266) );
  OAI21_X1 U15295 ( .B1(n20003), .B2(n12559), .A(n12266), .ZN(n12267) );
  NOR2_X1 U15296 ( .A1(n12268), .A2(n12267), .ZN(n12270) );
  NAND2_X1 U15297 ( .A1(n14464), .A2(n20024), .ZN(n12269) );
  NAND2_X1 U15298 ( .A1(n12269), .A2(n20023), .ZN(n14507) );
  OAI211_X1 U15299 ( .C1(n12271), .C2(n15966), .A(n12270), .B(n14507), .ZN(
        P1_U3031) );
  OAI21_X1 U15300 ( .B1(n12273), .B2(n12272), .A(n12579), .ZN(n12819) );
  INV_X1 U15301 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12817) );
  NAND2_X1 U15302 ( .A1(n20033), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14505) );
  OAI21_X1 U15303 ( .B1(n15871), .B2(n12817), .A(n14505), .ZN(n12274) );
  AOI21_X1 U15304 ( .B1(n15899), .B2(n12817), .A(n12274), .ZN(n12278) );
  OR2_X1 U15305 ( .A1(n12275), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14503) );
  NAND3_X1 U15306 ( .A1(n14503), .A2(n12276), .A3(n19994), .ZN(n12277) );
  OAI211_X1 U15307 ( .C1(n12819), .C2(n20044), .A(n12278), .B(n12277), .ZN(
        P1_U2998) );
  INV_X1 U15308 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15309 ( .A1(n13625), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13624), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15310 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12279), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15311 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13836), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15312 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15313 ( .A1(n12152), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12280) );
  NAND4_X1 U15314 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12289) );
  AOI22_X1 U15315 ( .A1(n13837), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11985), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15316 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15317 ( .A1(n12170), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15318 ( .A1(n12206), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12284) );
  NAND4_X1 U15319 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12288) );
  INV_X1 U15320 ( .A(n18990), .ZN(n12290) );
  OR2_X1 U15321 ( .A1(n12771), .A2(n12290), .ZN(n12291) );
  OAI211_X1 U15322 ( .C1(n13621), .C2(n12293), .A(n12292), .B(n12291), .ZN(
        n12298) );
  INV_X1 U15323 ( .A(n12294), .ZN(n12297) );
  INV_X1 U15324 ( .A(n12298), .ZN(n12295) );
  INV_X1 U15325 ( .A(n12365), .ZN(n12296) );
  OAI21_X1 U15326 ( .B1(n12298), .B2(n12297), .A(n12296), .ZN(n15351) );
  INV_X1 U15327 ( .A(n14780), .ZN(n12299) );
  OAI222_X1 U15328 ( .A1(n15351), .A2(n19023), .B1(n12299), .B2(n19065), .C1(
        n19079), .C2(n14810), .ZN(P2_U2911) );
  INV_X1 U15329 ( .A(n12394), .ZN(n19959) );
  AOI22_X1 U15330 ( .A1(n19959), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n9795), .ZN(n12303) );
  NAND2_X1 U15331 ( .A1(n20043), .A2(DATAI_5_), .ZN(n12301) );
  NAND2_X1 U15332 ( .A1(n20045), .A2(BUF1_REG_5__SCAN_IN), .ZN(n12300) );
  AND2_X1 U15333 ( .A1(n12301), .A2(n12300), .ZN(n20084) );
  INV_X1 U15334 ( .A(n20084), .ZN(n12302) );
  NAND2_X1 U15335 ( .A1(n19969), .A2(n12302), .ZN(n12401) );
  NAND2_X1 U15336 ( .A1(n12303), .A2(n12401), .ZN(P1_U2957) );
  AOI22_X1 U15337 ( .A1(n19959), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n9795), .ZN(n12307) );
  NAND2_X1 U15338 ( .A1(n20043), .A2(DATAI_2_), .ZN(n12305) );
  NAND2_X1 U15339 ( .A1(n20045), .A2(BUF1_REG_2__SCAN_IN), .ZN(n12304) );
  AND2_X1 U15340 ( .A1(n12305), .A2(n12304), .ZN(n20071) );
  INV_X1 U15341 ( .A(n20071), .ZN(n12306) );
  NAND2_X1 U15342 ( .A1(n19969), .A2(n12306), .ZN(n12411) );
  NAND2_X1 U15343 ( .A1(n12307), .A2(n12411), .ZN(P1_U2954) );
  AOI22_X1 U15344 ( .A1(n19959), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n9795), .ZN(n12311) );
  NAND2_X1 U15345 ( .A1(n20043), .A2(DATAI_3_), .ZN(n12309) );
  NAND2_X1 U15346 ( .A1(n20045), .A2(BUF1_REG_3__SCAN_IN), .ZN(n12308) );
  AND2_X1 U15347 ( .A1(n12309), .A2(n12308), .ZN(n20076) );
  INV_X1 U15348 ( .A(n20076), .ZN(n12310) );
  NAND2_X1 U15349 ( .A1(n19969), .A2(n12310), .ZN(n12419) );
  NAND2_X1 U15350 ( .A1(n12311), .A2(n12419), .ZN(P1_U2955) );
  AOI22_X1 U15351 ( .A1(n19959), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n9795), .ZN(n12315) );
  NAND2_X1 U15352 ( .A1(n20043), .A2(DATAI_4_), .ZN(n12313) );
  NAND2_X1 U15353 ( .A1(n20045), .A2(BUF1_REG_4__SCAN_IN), .ZN(n12312) );
  AND2_X1 U15354 ( .A1(n12313), .A2(n12312), .ZN(n20080) );
  INV_X1 U15355 ( .A(n20080), .ZN(n12314) );
  NAND2_X1 U15356 ( .A1(n19969), .A2(n12314), .ZN(n12395) );
  NAND2_X1 U15357 ( .A1(n12315), .A2(n12395), .ZN(P1_U2956) );
  AOI22_X1 U15358 ( .A1(n19959), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n9795), .ZN(n12319) );
  NAND2_X1 U15359 ( .A1(n20043), .A2(DATAI_6_), .ZN(n12317) );
  NAND2_X1 U15360 ( .A1(n20045), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12316) );
  AND2_X1 U15361 ( .A1(n12317), .A2(n12316), .ZN(n20087) );
  INV_X1 U15362 ( .A(n20087), .ZN(n12318) );
  NAND2_X1 U15363 ( .A1(n19969), .A2(n12318), .ZN(n12407) );
  NAND2_X1 U15364 ( .A1(n12319), .A2(n12407), .ZN(P1_U2958) );
  AOI22_X1 U15365 ( .A1(n19959), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n9795), .ZN(n12323) );
  NAND2_X1 U15366 ( .A1(n20043), .A2(DATAI_7_), .ZN(n12322) );
  NAND2_X1 U15367 ( .A1(n20045), .A2(BUF1_REG_7__SCAN_IN), .ZN(n12321) );
  AND2_X1 U15368 ( .A1(n12322), .A2(n12321), .ZN(n20095) );
  INV_X1 U15369 ( .A(n20095), .ZN(n14236) );
  NAND2_X1 U15370 ( .A1(n19969), .A2(n14236), .ZN(n12409) );
  NAND2_X1 U15371 ( .A1(n12323), .A2(n12409), .ZN(P1_U2959) );
  AND2_X1 U15372 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  AND2_X1 U15373 ( .A1(n12565), .A2(n12327), .ZN(n12329) );
  NAND2_X1 U15374 ( .A1(n12329), .A2(n12328), .ZN(n14521) );
  INV_X1 U15375 ( .A(n14521), .ZN(n15668) );
  XNOR2_X1 U15376 ( .A(n10521), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12332) );
  XNOR2_X1 U15377 ( .A(n14516), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12337) );
  NOR3_X1 U15378 ( .A1(n14521), .A2(n12330), .A3(n12337), .ZN(n12331) );
  AOI21_X1 U15379 ( .B1(n15669), .B2(n12332), .A(n12331), .ZN(n12336) );
  OR2_X1 U15380 ( .A1(n12334), .A2(n12333), .ZN(n12374) );
  NAND2_X1 U15381 ( .A1(n12374), .A2(n12337), .ZN(n12335) );
  OAI211_X1 U15382 ( .C1(n12324), .C2(n15668), .A(n12336), .B(n12335), .ZN(
        n12560) );
  INV_X1 U15383 ( .A(n20714), .ZN(n12390) );
  INV_X1 U15384 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20022) );
  AOI22_X1 U15385 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20022), .B2(n11452), .ZN(
        n14523) );
  NOR2_X1 U15386 ( .A1(n20627), .A2(n20023), .ZN(n20708) );
  INV_X1 U15387 ( .A(n12337), .ZN(n12338) );
  AOI222_X1 U15388 ( .A1(n12560), .A2(n12390), .B1(n14523), .B2(n20708), .C1(
        n12571), .C2(n12338), .ZN(n12351) );
  OAI21_X1 U15389 ( .B1(n12800), .B2(n10431), .A(n12339), .ZN(n12340) );
  NOR2_X1 U15390 ( .A1(n12341), .A2(n12340), .ZN(n12348) );
  NAND2_X1 U15391 ( .A1(n12343), .A2(n12342), .ZN(n12346) );
  AOI21_X1 U15392 ( .B1(n11313), .B2(n12344), .A(n20635), .ZN(n12345) );
  NAND3_X1 U15393 ( .A1(n12346), .A2(n12345), .A3(n15694), .ZN(n12347) );
  INV_X1 U15394 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19818) );
  NOR2_X1 U15395 ( .A1(n10081), .A2(n16039), .ZN(n12570) );
  INV_X1 U15396 ( .A(n12570), .ZN(n16043) );
  OAI22_X1 U15397 ( .A1(n15672), .A2(n19811), .B1(n19818), .B2(n16043), .ZN(
        n12371) );
  AOI21_X1 U15398 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n10081), .A(n12371), 
        .ZN(n20711) );
  NAND2_X1 U15399 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20711), .ZN(
        n12350) );
  OAI21_X1 U15400 ( .B1(n12351), .B2(n20711), .A(n12350), .ZN(P1_U3472) );
  INV_X1 U15401 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15402 ( .A1(n13625), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13624), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15403 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13836), .ZN(n12355) );
  AOI22_X1 U15404 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15405 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15406 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12352) );
  NAND4_X1 U15407 ( .A1(n12355), .A2(n12354), .A3(n12353), .A4(n12352), .ZN(
        n12361) );
  AOI22_X1 U15408 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15409 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15410 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12205), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15411 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12206), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12356) );
  NAND4_X1 U15412 ( .A1(n12359), .A2(n12358), .A3(n12357), .A4(n12356), .ZN(
        n12360) );
  OR2_X1 U15413 ( .A1(n12771), .A2(n12482), .ZN(n12362) );
  OAI211_X1 U15414 ( .C1(n13621), .C2(n12364), .A(n12363), .B(n12362), .ZN(
        n12366) );
  OAI21_X1 U15415 ( .B1(n12366), .B2(n12365), .A(n15317), .ZN(n18880) );
  INV_X1 U15416 ( .A(n14776), .ZN(n12367) );
  INV_X1 U15417 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20882) );
  OAI222_X1 U15418 ( .A1(n18880), .A2(n19023), .B1(n12367), .B2(n19065), .C1(
        n20882), .C2(n14810), .ZN(P2_U2910) );
  INV_X1 U15419 ( .A(n20711), .ZN(n20709) );
  INV_X1 U15420 ( .A(n12565), .ZN(n12370) );
  INV_X1 U15421 ( .A(n20204), .ZN(n20461) );
  OR2_X1 U15422 ( .A1(n10550), .A2(n20461), .ZN(n12368) );
  XNOR2_X1 U15423 ( .A(n12368), .B(n12373), .ZN(n19894) );
  INV_X1 U15424 ( .A(n19894), .ZN(n12369) );
  NAND4_X1 U15425 ( .A1(n12371), .A2(n12390), .A3(n12370), .A4(n12369), .ZN(
        n12372) );
  OAI21_X1 U15426 ( .B1(n12373), .B2(n20709), .A(n12372), .ZN(P1_U3468) );
  NAND2_X1 U15427 ( .A1(n20323), .A2(n14521), .ZN(n12388) );
  MUX2_X1 U15428 ( .A(n12383), .B(n12391), .S(n14516), .Z(n12375) );
  OAI21_X1 U15429 ( .B1(n12381), .B2(n12375), .A(n12374), .ZN(n12386) );
  NOR2_X1 U15430 ( .A1(n14516), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12377) );
  NOR2_X1 U15431 ( .A1(n12377), .A2(n12376), .ZN(n12379) );
  AND2_X1 U15432 ( .A1(n12379), .A2(n12378), .ZN(n12389) );
  NAND3_X1 U15433 ( .A1(n15668), .A2(n12380), .A3(n12389), .ZN(n12385) );
  MUX2_X1 U15434 ( .A(n12381), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n10521), .Z(n12382) );
  OAI21_X1 U15435 ( .B1(n12383), .B2(n12382), .A(n15669), .ZN(n12384) );
  AND3_X1 U15436 ( .A1(n12386), .A2(n12385), .A3(n12384), .ZN(n12387) );
  NAND2_X1 U15437 ( .A1(n12388), .A2(n12387), .ZN(n12561) );
  AOI22_X1 U15438 ( .A1(n12561), .A2(n12390), .B1(n12389), .B2(n12571), .ZN(
        n12392) );
  MUX2_X1 U15439 ( .A(n12392), .B(n12391), .S(n20711), .Z(n12393) );
  INV_X1 U15440 ( .A(n12393), .ZN(P1_U3469) );
  AOI22_X1 U15441 ( .A1(n19983), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n9795), .ZN(n12396) );
  NAND2_X1 U15442 ( .A1(n12396), .A2(n12395), .ZN(P1_U2941) );
  AOI22_X1 U15443 ( .A1(n19983), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n9795), .ZN(n12400) );
  NAND2_X1 U15444 ( .A1(n20043), .A2(DATAI_1_), .ZN(n12398) );
  NAND2_X1 U15445 ( .A1(n20045), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12397) );
  AND2_X1 U15446 ( .A1(n12398), .A2(n12397), .ZN(n20067) );
  INV_X1 U15447 ( .A(n20067), .ZN(n12399) );
  NAND2_X1 U15448 ( .A1(n19969), .A2(n12399), .ZN(n12421) );
  NAND2_X1 U15449 ( .A1(n12400), .A2(n12421), .ZN(P1_U2938) );
  AOI22_X1 U15450 ( .A1(n19983), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n9795), .ZN(n12402) );
  NAND2_X1 U15451 ( .A1(n12402), .A2(n12401), .ZN(P1_U2942) );
  AOI22_X1 U15452 ( .A1(n19983), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n9795), .ZN(n12406) );
  INV_X1 U15453 ( .A(DATAI_13_), .ZN(n12404) );
  MUX2_X1 U15454 ( .A(n12404), .B(n12403), .S(n20045), .Z(n14213) );
  INV_X1 U15455 ( .A(n14213), .ZN(n12405) );
  NAND2_X1 U15456 ( .A1(n19969), .A2(n12405), .ZN(n19981) );
  NAND2_X1 U15457 ( .A1(n12406), .A2(n19981), .ZN(P1_U2950) );
  AOI22_X1 U15458 ( .A1(n19983), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n9795), .ZN(n12408) );
  NAND2_X1 U15459 ( .A1(n12408), .A2(n12407), .ZN(P1_U2943) );
  AOI22_X1 U15460 ( .A1(n19983), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n9795), .ZN(n12410) );
  NAND2_X1 U15461 ( .A1(n12410), .A2(n12409), .ZN(P1_U2944) );
  AOI22_X1 U15462 ( .A1(n19983), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n9795), .ZN(n12412) );
  NAND2_X1 U15463 ( .A1(n12412), .A2(n12411), .ZN(P1_U2939) );
  AOI22_X1 U15464 ( .A1(n19983), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n9795), .ZN(n12416) );
  NAND2_X1 U15465 ( .A1(n20043), .A2(DATAI_0_), .ZN(n12414) );
  NAND2_X1 U15466 ( .A1(n20045), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12413) );
  AND2_X1 U15467 ( .A1(n12414), .A2(n12413), .ZN(n20058) );
  INV_X1 U15468 ( .A(n20058), .ZN(n12415) );
  NAND2_X1 U15469 ( .A1(n19969), .A2(n12415), .ZN(n12417) );
  NAND2_X1 U15470 ( .A1(n12416), .A2(n12417), .ZN(P1_U2937) );
  AOI22_X1 U15471 ( .A1(n19983), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n9795), .ZN(n12418) );
  NAND2_X1 U15472 ( .A1(n12418), .A2(n12417), .ZN(P1_U2952) );
  AOI22_X1 U15473 ( .A1(n19983), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n9795), .ZN(n12420) );
  NAND2_X1 U15474 ( .A1(n12420), .A2(n12419), .ZN(P1_U2940) );
  AOI22_X1 U15475 ( .A1(n19983), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n9795), .ZN(n12422) );
  NAND2_X1 U15476 ( .A1(n12422), .A2(n12421), .ZN(P1_U2953) );
  INV_X1 U15477 ( .A(n12701), .ZN(n12423) );
  NAND2_X1 U15478 ( .A1(n12423), .A2(n12698), .ZN(n12645) );
  NAND2_X1 U15479 ( .A1(n12689), .A2(n9802), .ZN(n12653) );
  NAND2_X1 U15480 ( .A1(n12645), .A2(n12653), .ZN(n12425) );
  INV_X1 U15481 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n18867) );
  NAND2_X1 U15482 ( .A1(n12426), .A2(n12475), .ZN(n12428) );
  XNOR2_X1 U15483 ( .A(n19794), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15450) );
  AND2_X1 U15484 ( .A1(n15450), .A2(n19771), .ZN(n19214) );
  AOI21_X1 U15485 ( .B1(n12473), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19214), .ZN(n12427) );
  NAND2_X1 U15486 ( .A1(n12428), .A2(n12427), .ZN(n13687) );
  NAND3_X1 U15487 ( .A1(n12043), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14018), 
        .ZN(n13922) );
  INV_X1 U15488 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12429) );
  NOR2_X1 U15489 ( .A1(n13922), .A2(n12429), .ZN(n12431) );
  INV_X1 U15490 ( .A(n12435), .ZN(n12437) );
  NAND2_X1 U15491 ( .A1(n12437), .A2(n12436), .ZN(n12438) );
  AOI21_X1 U15492 ( .B1(n12943), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12439) );
  NAND2_X1 U15493 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19572) );
  INV_X1 U15494 ( .A(n19572), .ZN(n12441) );
  INV_X1 U15495 ( .A(n12470), .ZN(n12443) );
  NAND2_X1 U15496 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19485) );
  NAND2_X1 U15497 ( .A1(n19485), .A2(n19777), .ZN(n12442) );
  NAND2_X1 U15498 ( .A1(n12443), .A2(n12442), .ZN(n15451) );
  NOR2_X1 U15499 ( .A1(n19762), .A2(n15451), .ZN(n12444) );
  AOI21_X1 U15500 ( .B1(n12473), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12444), .ZN(n12453) );
  INV_X1 U15501 ( .A(n13922), .ZN(n13948) );
  NAND2_X1 U15502 ( .A1(n13948), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12458) );
  AND2_X1 U15503 ( .A1(n12453), .A2(n12458), .ZN(n12449) );
  NAND2_X1 U15504 ( .A1(n10249), .A2(n12449), .ZN(n12451) );
  OR2_X1 U15505 ( .A1(n12679), .A2(n12451), .ZN(n12457) );
  INV_X1 U15506 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n12447) );
  NAND2_X1 U15507 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12445) );
  OAI211_X1 U15508 ( .C1(n13598), .C2(n12447), .A(n12446), .B(n12445), .ZN(
        n12448) );
  INV_X1 U15510 ( .A(n12449), .ZN(n12450) );
  OAI22_X1 U15511 ( .A1(n12451), .A2(n12677), .B1(n10249), .B2(n12450), .ZN(
        n12452) );
  NAND2_X1 U15512 ( .A1(n12679), .A2(n12452), .ZN(n12456) );
  INV_X1 U15513 ( .A(n12453), .ZN(n12459) );
  OAI21_X1 U15514 ( .B1(n12459), .B2(n12475), .A(n12458), .ZN(n12454) );
  OAI21_X1 U15515 ( .B1(n12458), .B2(n12459), .A(n12454), .ZN(n12455) );
  INV_X1 U15516 ( .A(n12458), .ZN(n12460) );
  NAND2_X1 U15517 ( .A1(n12460), .A2(n12459), .ZN(n12461) );
  AND2_X2 U15518 ( .A1(n13055), .A2(n12461), .ZN(n12940) );
  INV_X1 U15519 ( .A(n12462), .ZN(n13575) );
  INV_X4 U15520 ( .A(n13575), .ZN(n13600) );
  INV_X1 U15521 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12465) );
  INV_X4 U15522 ( .A(n13585), .ZN(n13595) );
  NAND2_X1 U15523 ( .A1(n13595), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12464) );
  NAND2_X1 U15524 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12463) );
  OAI211_X1 U15525 ( .C1(n13598), .C2(n12465), .A(n12464), .B(n12463), .ZN(
        n12466) );
  NAND2_X1 U15526 ( .A1(n12467), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12469) );
  NAND2_X1 U15527 ( .A1(n12718), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12468) );
  INV_X1 U15528 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13248) );
  NOR2_X1 U15529 ( .A1(n13922), .A2(n13248), .ZN(n12935) );
  INV_X1 U15530 ( .A(n12935), .ZN(n12474) );
  OAI21_X1 U15531 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12470), .A(
        n19771), .ZN(n12471) );
  NOR2_X1 U15532 ( .A1(n12471), .A2(n19669), .ZN(n12472) );
  AOI21_X1 U15533 ( .B1(n12473), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12472), .ZN(n12478) );
  INV_X1 U15534 ( .A(n12938), .ZN(n12476) );
  INV_X1 U15535 ( .A(n12478), .ZN(n12936) );
  NAND2_X1 U15536 ( .A1(n12936), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12479) );
  AND2_X1 U15537 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12519) );
  NAND4_X1 U15538 ( .A1(n18990), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .A4(n12519), .ZN(n12480) );
  NOR2_X1 U15539 ( .A1(n13922), .A2(n12480), .ZN(n12481) );
  NAND2_X1 U15540 ( .A1(n19000), .A2(n12483), .ZN(n18992) );
  OAI211_X1 U15541 ( .C1(n9826), .C2(n12484), .A(n10289), .B(n18998), .ZN(
        n12516) );
  NAND2_X1 U15542 ( .A1(n13595), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12486) );
  NAND2_X1 U15543 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12485) );
  OAI211_X1 U15544 ( .C1(n13598), .C2(n18867), .A(n12486), .B(n12485), .ZN(
        n12487) );
  AOI21_X1 U15545 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12487), .ZN(n12512) );
  INV_X1 U15546 ( .A(n12490), .ZN(n12492) );
  NAND2_X1 U15547 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  NAND2_X1 U15548 ( .A1(n12494), .A2(n12493), .ZN(n18936) );
  INV_X1 U15549 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12497) );
  NAND2_X1 U15550 ( .A1(n13595), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12496) );
  NAND2_X1 U15551 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12495) );
  OAI211_X1 U15552 ( .C1(n13598), .C2(n12497), .A(n12496), .B(n12495), .ZN(
        n12498) );
  AOI21_X1 U15553 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12498), .ZN(n18935) );
  INV_X1 U15554 ( .A(n18935), .ZN(n12499) );
  INV_X1 U15555 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U15556 ( .A1(n13595), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12501) );
  NAND2_X1 U15557 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12500) );
  OAI211_X1 U15558 ( .C1(n13598), .C2(n12502), .A(n12501), .B(n12500), .ZN(
        n12503) );
  AOI21_X1 U15559 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12503), .ZN(n13697) );
  INV_X1 U15560 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18894) );
  NAND2_X1 U15561 ( .A1(n13595), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12505) );
  NAND2_X1 U15562 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12504) );
  OAI211_X1 U15563 ( .C1(n13598), .C2(n18894), .A(n12505), .B(n12504), .ZN(
        n12506) );
  AOI21_X1 U15564 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n12506), .ZN(n12523) );
  INV_X1 U15565 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13047) );
  NAND2_X1 U15566 ( .A1(n13600), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12508) );
  AOI22_X1 U15567 ( .A1(n13595), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12507) );
  OAI211_X1 U15568 ( .C1(n13047), .C2(n13598), .A(n12508), .B(n12507), .ZN(
        n13701) );
  INV_X1 U15569 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12511) );
  NAND2_X1 U15570 ( .A1(n13600), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12510) );
  AOI22_X1 U15571 ( .A1(n13595), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12509) );
  OAI211_X1 U15572 ( .C1(n12511), .C2(n13598), .A(n12510), .B(n12509), .ZN(
        n13028) );
  NAND2_X1 U15573 ( .A1(n12512), .A2(n13029), .ZN(n12514) );
  INV_X1 U15574 ( .A(n15313), .ZN(n12513) );
  NAND2_X1 U15575 ( .A1(n18876), .A2(n19000), .ZN(n12515) );
  OAI211_X1 U15576 ( .C1(n19000), .C2(n18867), .A(n12516), .B(n12515), .ZN(
        P2_U2878) );
  INV_X1 U15577 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12517) );
  NOR2_X1 U15578 ( .A1(n13922), .A2(n12517), .ZN(n18930) );
  NAND2_X1 U15579 ( .A1(n12518), .A2(n18930), .ZN(n18934) );
  INV_X1 U15580 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13306) );
  NOR2_X1 U15581 ( .A1(n18934), .A2(n13306), .ZN(n12522) );
  INV_X1 U15582 ( .A(n12519), .ZN(n12520) );
  NOR2_X1 U15583 ( .A1(n18934), .A2(n12520), .ZN(n18991) );
  INV_X1 U15584 ( .A(n18991), .ZN(n12521) );
  OAI211_X1 U15585 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n12522), .A(
        n12521), .B(n18998), .ZN(n12526) );
  AND2_X1 U15586 ( .A1(n13695), .A2(n12523), .ZN(n12524) );
  NAND2_X1 U15587 ( .A1(n9894), .A2(n19000), .ZN(n12525) );
  OAI211_X1 U15588 ( .C1(n19000), .C2(n18894), .A(n12526), .B(n12525), .ZN(
        P2_U2881) );
  INV_X1 U15589 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19074) );
  INV_X1 U15590 ( .A(n14750), .ZN(n12556) );
  INV_X1 U15591 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U15592 ( .A1(n13625), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U15593 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12165), .B1(
        n12200), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15594 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12151), .B1(
        n12279), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15595 ( .A1(n13838), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n13836), .ZN(n12528) );
  AOI22_X1 U15596 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12527) );
  NAND4_X1 U15597 ( .A1(n12530), .A2(n12529), .A3(n12528), .A4(n12527), .ZN(
        n12536) );
  AOI22_X1 U15598 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11985), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U15599 ( .A1(n13837), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U15600 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n12206), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15601 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12205), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12531) );
  NAND4_X1 U15602 ( .A1(n12534), .A2(n12533), .A3(n12532), .A4(n12531), .ZN(
        n12535) );
  INV_X1 U15603 ( .A(n18984), .ZN(n12537) );
  OR2_X1 U15604 ( .A1(n12771), .A2(n12537), .ZN(n12538) );
  OAI211_X1 U15605 ( .C1(n12150), .C2(n12540), .A(n12539), .B(n12538), .ZN(
        n12541) );
  INV_X1 U15606 ( .A(n12541), .ZN(n15318) );
  AOI22_X1 U15607 ( .A1(n13625), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12553) );
  INV_X1 U15608 ( .A(n12771), .ZN(n13604) );
  AOI22_X1 U15609 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n13836), .ZN(n12545) );
  AOI22_X1 U15610 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15611 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15612 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12542) );
  NAND4_X1 U15613 ( .A1(n12545), .A2(n12544), .A3(n12543), .A4(n12542), .ZN(
        n12551) );
  AOI22_X1 U15614 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15615 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15616 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12205), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15617 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n12206), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12546) );
  NAND4_X1 U15618 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12550) );
  AOI22_X1 U15619 ( .A1(n13604), .A2(n18978), .B1(n13626), .B2(
        P2_REIP_REG_11__SCAN_IN), .ZN(n12552) );
  NAND2_X1 U15620 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  OAI21_X1 U15621 ( .B1(n12555), .B2(n12554), .A(n15272), .ZN(n15298) );
  OAI222_X1 U15622 ( .A1(n14810), .A2(n19074), .B1(n12556), .B2(n19065), .C1(
        n15298), .C2(n19023), .ZN(P2_U2908) );
  XNOR2_X1 U15623 ( .A(n12814), .B(n11313), .ZN(n14504) );
  INV_X1 U15624 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12557) );
  OAI222_X1 U15625 ( .A1(n14504), .A2(n19912), .B1(n19919), .B2(n12557), .C1(
        n12819), .C2(n9794), .ZN(P1_U2871) );
  OAI222_X1 U15626 ( .A1(n12559), .A2(n19912), .B1(n12558), .B2(n19919), .C1(
        n12825), .C2(n9794), .ZN(P1_U2872) );
  NOR2_X1 U15627 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20627), .ZN(n12566) );
  MUX2_X1 U15628 ( .A(n12560), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15672), .Z(n15677) );
  AOI22_X1 U15629 ( .A1(n12566), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15677), .B2(n20627), .ZN(n12563) );
  INV_X1 U15630 ( .A(n15672), .ZN(n12564) );
  MUX2_X1 U15631 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n12561), .S(
        n12564), .Z(n15666) );
  AOI22_X1 U15632 ( .A1(n12566), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20627), .B2(n15666), .ZN(n12562) );
  NOR2_X1 U15633 ( .A1(n12563), .A2(n12562), .ZN(n15687) );
  INV_X1 U15634 ( .A(n15687), .ZN(n12569) );
  OAI21_X1 U15635 ( .B1(n19894), .B2(n12565), .A(n12564), .ZN(n12568) );
  AOI21_X1 U15636 ( .B1(n15672), .B2(n12373), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n12567) );
  AOI22_X1 U15637 ( .A1(n12568), .A2(n12567), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n12566), .ZN(n15685) );
  OAI21_X1 U15638 ( .B1(n12569), .B2(n14515), .A(n15685), .ZN(n12573) );
  OAI21_X1 U15639 ( .B1(n12573), .B2(P1_FLUSH_REG_SCAN_IN), .A(n12570), .ZN(
        n12572) );
  NAND2_X1 U15640 ( .A1(n10613), .A2(n20627), .ZN(n20730) );
  NAND2_X1 U15641 ( .A1(n12572), .A2(n20210), .ZN(n20041) );
  NOR2_X1 U15642 ( .A1(n12573), .A2(n16039), .ZN(n15697) );
  INV_X1 U15643 ( .A(n20496), .ZN(n20565) );
  INV_X1 U15644 ( .A(n20289), .ZN(n20166) );
  NAND2_X1 U15645 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20704), .ZN(n12588) );
  INV_X1 U15646 ( .A(n12588), .ZN(n12574) );
  OAI22_X1 U15647 ( .A1(n11114), .A2(n20565), .B1(n20166), .B2(n12574), .ZN(
        n12575) );
  OAI21_X1 U15648 ( .B1(n15697), .B2(n12575), .A(n20041), .ZN(n12576) );
  OAI21_X1 U15649 ( .B1(n20041), .B2(n20489), .A(n12576), .ZN(P1_U3478) );
  OR2_X1 U15650 ( .A1(n9908), .A2(n12577), .ZN(n12578) );
  NAND2_X1 U15651 ( .A1(n12597), .A2(n12578), .ZN(n20021) );
  INV_X1 U15652 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n20814) );
  OAI21_X1 U15653 ( .B1(n10307), .B2(n10640), .A(n12580), .ZN(n12933) );
  OAI222_X1 U15654 ( .A1(n20021), .A2(n19912), .B1(n19919), .B2(n20814), .C1(
        n12933), .C2(n9794), .ZN(P1_U2870) );
  OAI21_X1 U15655 ( .B1(n12583), .B2(n12582), .A(n12581), .ZN(n20029) );
  INV_X1 U15656 ( .A(n12933), .ZN(n12586) );
  AOI22_X1 U15657 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20033), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n12584) );
  OAI21_X1 U15658 ( .B1(n19998), .B2(n12928), .A(n12584), .ZN(n12585) );
  AOI21_X1 U15659 ( .B1(n12586), .B2(n19993), .A(n12585), .ZN(n12587) );
  OAI21_X1 U15660 ( .B1(n19817), .B2(n20029), .A(n12587), .ZN(P1_U2997) );
  INV_X1 U15661 ( .A(n20323), .ZN(n12595) );
  NAND2_X1 U15662 ( .A1(n20041), .A2(n12588), .ZN(n13230) );
  NAND2_X1 U15663 ( .A1(n20129), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20295) );
  INV_X1 U15664 ( .A(n12590), .ZN(n12589) );
  OR2_X1 U15665 ( .A1(n20129), .A2(n20207), .ZN(n20351) );
  OR2_X1 U15666 ( .A1(n20572), .A2(n20351), .ZN(n20493) );
  NAND2_X1 U15667 ( .A1(n20048), .A2(n20207), .ZN(n12591) );
  OAI211_X1 U15668 ( .C1(n20295), .C2(n20299), .A(n20493), .B(n12591), .ZN(
        n12592) );
  NAND2_X1 U15669 ( .A1(n20041), .A2(n20496), .ZN(n12643) );
  INV_X1 U15670 ( .A(n12643), .ZN(n13226) );
  OAI21_X1 U15671 ( .B1(n20425), .B2(n12592), .A(n13226), .ZN(n12594) );
  INV_X1 U15672 ( .A(n20041), .ZN(n13227) );
  NAND2_X1 U15673 ( .A1(n13227), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12593) );
  OAI211_X1 U15674 ( .C1(n12595), .C2(n13230), .A(n12594), .B(n12593), .ZN(
        P1_U3475) );
  NAND2_X1 U15675 ( .A1(n12597), .A2(n12596), .ZN(n12598) );
  NAND2_X1 U15676 ( .A1(n12757), .A2(n12598), .ZN(n20011) );
  INV_X1 U15677 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12602) );
  OAI21_X1 U15678 ( .B1(n12601), .B2(n12600), .A(n12599), .ZN(n12921) );
  OAI222_X1 U15679 ( .A1(n20011), .A2(n19912), .B1(n12602), .B2(n19919), .C1(
        n12921), .C2(n9794), .ZN(P1_U2869) );
  INV_X1 U15680 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n18834) );
  AOI22_X1 U15681 ( .A1(n13625), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15682 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13836), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15683 ( .A1(n12279), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15684 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15685 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12603) );
  NAND4_X1 U15686 ( .A1(n12606), .A2(n12605), .A3(n12604), .A4(n12603), .ZN(
        n12612) );
  AOI22_X1 U15687 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15688 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15689 ( .A1(n12205), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U15690 ( .A1(n12206), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12607) );
  NAND4_X1 U15691 ( .A1(n12610), .A2(n12609), .A3(n12608), .A4(n12607), .ZN(
        n12611) );
  INV_X1 U15692 ( .A(n12735), .ZN(n12733) );
  OR2_X1 U15693 ( .A1(n12771), .A2(n12733), .ZN(n12613) );
  OAI211_X1 U15694 ( .C1(n12150), .C2(n18834), .A(n12614), .B(n12613), .ZN(
        n12632) );
  INV_X1 U15695 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U15696 ( .A1(n13625), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U15697 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12165), .B1(
        n12279), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15698 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n13836), .ZN(n12617) );
  AOI22_X1 U15699 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15700 ( .A1(n12152), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12615) );
  NAND4_X1 U15701 ( .A1(n12618), .A2(n12617), .A3(n12616), .A4(n12615), .ZN(
        n12624) );
  AOI22_X1 U15702 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11985), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15703 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15704 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12205), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15705 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12654), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12619) );
  NAND4_X1 U15706 ( .A1(n12622), .A2(n12621), .A3(n12620), .A4(n12619), .ZN(
        n12623) );
  INV_X1 U15707 ( .A(n18977), .ZN(n12625) );
  OR2_X1 U15708 ( .A1(n12771), .A2(n12625), .ZN(n12626) );
  OAI211_X1 U15709 ( .C1(n12150), .C2(n12628), .A(n12627), .B(n12626), .ZN(
        n12629) );
  INV_X1 U15710 ( .A(n12629), .ZN(n15271) );
  OAI21_X1 U15711 ( .B1(n12632), .B2(n12631), .A(n12630), .ZN(n18845) );
  INV_X1 U15712 ( .A(n14738), .ZN(n12633) );
  INV_X1 U15713 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19071) );
  OAI222_X1 U15714 ( .A1(n18845), .A2(n19023), .B1(n12633), .B2(n19065), .C1(
        n19071), .C2(n14810), .ZN(P2_U2906) );
  OAI21_X1 U15715 ( .B1(n12636), .B2(n12635), .A(n12634), .ZN(n12637) );
  INV_X1 U15716 ( .A(n12637), .ZN(n20016) );
  NAND2_X1 U15717 ( .A1(n20016), .A2(n19994), .ZN(n12640) );
  AND2_X1 U15718 ( .A1(n20033), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20012) );
  NOR2_X1 U15719 ( .A1(n19998), .A2(n12917), .ZN(n12638) );
  AOI211_X1 U15720 ( .C1(n19987), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20012), .B(n12638), .ZN(n12639) );
  OAI211_X1 U15721 ( .C1(n20044), .C2(n12921), .A(n12640), .B(n12639), .ZN(
        P1_U2996) );
  XNOR2_X1 U15722 ( .A(n12641), .B(n20295), .ZN(n12642) );
  OAI222_X1 U15723 ( .A1(n13230), .A2(n12324), .B1(n20041), .B2(n20375), .C1(
        n12643), .C2(n12642), .ZN(P1_U3476) );
  AND3_X1 U15724 ( .A1(n12646), .A2(n12645), .A3(n12644), .ZN(n12651) );
  INV_X1 U15725 ( .A(n12647), .ZN(n12649) );
  INV_X1 U15726 ( .A(n11900), .ZN(n12648) );
  NAND3_X1 U15727 ( .A1(n12649), .A2(n12648), .A3(n12716), .ZN(n12650) );
  NAND2_X1 U15728 ( .A1(n12653), .A2(n12652), .ZN(n12686) );
  INV_X1 U15729 ( .A(n12654), .ZN(n12655) );
  OAI21_X1 U15730 ( .B1(n14036), .B2(n12694), .A(n12655), .ZN(n12661) );
  NOR2_X1 U15731 ( .A1(n12698), .A2(n12696), .ZN(n12683) );
  NOR2_X1 U15732 ( .A1(n12656), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12680) );
  XNOR2_X1 U15733 ( .A(n12680), .B(n12694), .ZN(n12658) );
  INV_X1 U15734 ( .A(n12668), .ZN(n12682) );
  XNOR2_X1 U15735 ( .A(n11947), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12657) );
  OAI22_X1 U15736 ( .A1(n12683), .A2(n12658), .B1(n12682), .B2(n12657), .ZN(
        n12660) );
  NOR2_X1 U15737 ( .A1(n13234), .A2(n12689), .ZN(n12659) );
  AOI211_X1 U15738 ( .C1(n12686), .C2(n12661), .A(n12660), .B(n12659), .ZN(
        n15421) );
  INV_X1 U15739 ( .A(n12689), .ZN(n12671) );
  NAND2_X1 U15740 ( .A1(n15400), .A2(n12671), .ZN(n12667) );
  NOR2_X1 U15741 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12662) );
  NOR2_X1 U15742 ( .A1(n12656), .A2(n12662), .ZN(n12665) );
  NAND2_X1 U15743 ( .A1(n12664), .A2(n12663), .ZN(n12669) );
  AOI22_X1 U15744 ( .A1(n12665), .A2(n12669), .B1(n12668), .B2(n10275), .ZN(
        n12666) );
  NAND2_X1 U15745 ( .A1(n12667), .A2(n12666), .ZN(n15418) );
  MUX2_X1 U15746 ( .A(n12669), .B(n12668), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n12670) );
  AOI21_X1 U15747 ( .B1(n12037), .B2(n12671), .A(n12670), .ZN(n15410) );
  NAND2_X1 U15748 ( .A1(n15410), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12672) );
  NOR2_X1 U15749 ( .A1(n15418), .A2(n12672), .ZN(n12676) );
  AND2_X1 U15750 ( .A1(n15418), .A2(n12672), .ZN(n12674) );
  INV_X1 U15751 ( .A(n15411), .ZN(n12673) );
  OAI21_X1 U15752 ( .B1(n12674), .B2(n19787), .A(n12673), .ZN(n12675) );
  AOI211_X1 U15753 ( .C1(n15421), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n12676), .B(n12675), .ZN(n12693) );
  NOR2_X1 U15754 ( .A1(n12680), .A2(n14036), .ZN(n12687) );
  NOR3_X1 U15755 ( .A1(n12682), .A2(n12681), .A3(n11947), .ZN(n12685) );
  NOR2_X1 U15756 ( .A1(n12683), .A2(n12687), .ZN(n12684) );
  AOI211_X1 U15757 ( .C1(n12687), .C2(n12686), .A(n12685), .B(n12684), .ZN(
        n12688) );
  OAI21_X1 U15758 ( .B1(n13691), .B2(n12689), .A(n12688), .ZN(n19754) );
  NAND2_X1 U15759 ( .A1(n15411), .A2(n10276), .ZN(n12690) );
  OAI21_X1 U15760 ( .B1(n19754), .B2(n15411), .A(n12690), .ZN(n12712) );
  NOR2_X1 U15761 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19213) );
  INV_X1 U15762 ( .A(n19213), .ZN(n19244) );
  NOR2_X1 U15763 ( .A1(n12712), .A2(n19244), .ZN(n12692) );
  INV_X1 U15764 ( .A(n12712), .ZN(n12691) );
  OAI22_X1 U15765 ( .A1(n12693), .A2(n12692), .B1(n12691), .B2(n19777), .ZN(
        n12695) );
  MUX2_X1 U15766 ( .A(n15421), .B(n12694), .S(n15411), .Z(n12713) );
  AOI221_X1 U15767 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12695), 
        .C1(n12713), .C2(n12695), .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12715) );
  INV_X1 U15768 ( .A(n12696), .ZN(n12700) );
  AOI22_X1 U15769 ( .A1(n12701), .A2(n12698), .B1(n11937), .B2(n12697), .ZN(
        n12699) );
  OAI21_X1 U15770 ( .B1(n12701), .B2(n12700), .A(n12699), .ZN(n19802) );
  INV_X1 U15771 ( .A(n19802), .ZN(n12711) );
  NOR3_X1 U15772 ( .A1(n15479), .A2(n15477), .A3(n15478), .ZN(n12708) );
  INV_X1 U15773 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12706) );
  INV_X1 U15774 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n12705) );
  INV_X1 U15775 ( .A(n12702), .ZN(n12703) );
  OR3_X1 U15776 ( .A1(n12704), .A2(n12703), .A3(n12716), .ZN(n18733) );
  AOI21_X1 U15777 ( .B1(n12706), .B2(n12705), .A(n18733), .ZN(n12707) );
  AOI211_X1 U15778 ( .C1(n12709), .C2(n15433), .A(n12708), .B(n12707), .ZN(
        n12710) );
  OAI211_X1 U15779 ( .C1(n12713), .C2(n12712), .A(n12711), .B(n12710), .ZN(
        n12714) );
  AOI211_X1 U15780 ( .C1(n15411), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n12715), .B(n12714), .ZN(n16230) );
  AOI21_X1 U15781 ( .B1(n16230), .B2(n15409), .A(n12943), .ZN(n12723) );
  INV_X1 U15782 ( .A(n12716), .ZN(n12717) );
  NOR2_X1 U15783 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12717), .ZN(n12971) );
  NAND2_X1 U15784 ( .A1(n10055), .A2(n12971), .ZN(n12720) );
  OR2_X1 U15785 ( .A1(n12718), .A2(n19390), .ZN(n14529) );
  INV_X1 U15786 ( .A(n14529), .ZN(n12719) );
  OAI21_X1 U15787 ( .B1(n12721), .B2(n12720), .A(n12719), .ZN(n12722) );
  INV_X1 U15788 ( .A(n12786), .ZN(n16227) );
  OAI21_X1 U15789 ( .B1(n16227), .B2(n12943), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12725) );
  NOR2_X1 U15790 ( .A1(n12943), .A2(n16225), .ZN(n15739) );
  INV_X1 U15791 ( .A(n15739), .ZN(n12724) );
  NAND2_X1 U15792 ( .A1(n12725), .A2(n12724), .ZN(P2_U3593) );
  INV_X1 U15793 ( .A(n12726), .ZN(n12727) );
  XNOR2_X1 U15794 ( .A(n12727), .B(n12599), .ZN(n19992) );
  INV_X1 U15795 ( .A(n19992), .ZN(n12760) );
  INV_X1 U15796 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19943) );
  INV_X1 U15797 ( .A(n12728), .ZN(n12729) );
  OAI222_X1 U15798 ( .A1(n14268), .A2(n12760), .B1(n14271), .B2(n19943), .C1(
        n14273), .C2(n20080), .ZN(P1_U2900) );
  INV_X1 U15799 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U15800 ( .A1(n13706), .A2(n12731), .ZN(n12732) );
  INV_X1 U15801 ( .A(n12732), .ZN(n18980) );
  INV_X1 U15802 ( .A(n12732), .ZN(n12734) );
  OAI211_X1 U15803 ( .C1(n18980), .C2(n12735), .A(n18998), .B(n12993), .ZN(
        n12754) );
  NAND2_X1 U15804 ( .A1(n13600), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12740) );
  AOI22_X1 U15805 ( .A1(n13595), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12738) );
  NAND2_X1 U15806 ( .A1(n9803), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12737) );
  AND2_X1 U15807 ( .A1(n12738), .A2(n12737), .ZN(n12739) );
  NAND2_X1 U15808 ( .A1(n12740), .A2(n12739), .ZN(n15276) );
  INV_X1 U15809 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U15810 ( .A1(n13600), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12742) );
  AOI22_X1 U15811 ( .A1(n13595), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12741) );
  OAI211_X1 U15812 ( .C1(n13598), .C2(n12743), .A(n12742), .B(n12741), .ZN(
        n15314) );
  INV_X1 U15813 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15814 ( .A1(n13595), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U15815 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12744) );
  OAI211_X1 U15816 ( .C1(n13598), .C2(n12746), .A(n12745), .B(n12744), .ZN(
        n12747) );
  AOI21_X1 U15817 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12747), .ZN(n13707) );
  NAND2_X1 U15818 ( .A1(n13595), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U15819 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12748) );
  OAI211_X1 U15820 ( .C1(n13598), .C2(n12755), .A(n12749), .B(n12748), .ZN(
        n12750) );
  AOI21_X1 U15821 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12750), .ZN(n12751) );
  OR2_X2 U15822 ( .A1(n15278), .A2(n12751), .ZN(n15258) );
  NAND2_X1 U15823 ( .A1(n15278), .A2(n12751), .ZN(n12752) );
  AND2_X1 U15824 ( .A1(n15258), .A2(n12752), .ZN(n18842) );
  NAND2_X1 U15825 ( .A1(n18842), .A2(n19000), .ZN(n12753) );
  OAI211_X1 U15826 ( .C1(n19000), .C2(n12755), .A(n12754), .B(n12753), .ZN(
        P2_U2874) );
  AND2_X1 U15827 ( .A1(n12757), .A2(n12756), .ZN(n12758) );
  OR2_X1 U15828 ( .A1(n12758), .A2(n16027), .ZN(n20004) );
  INV_X1 U15829 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n12759) );
  OAI222_X1 U15830 ( .A1(n20004), .A2(n19912), .B1(n9794), .B2(n12760), .C1(
        n12759), .C2(n19919), .ZN(P1_U2868) );
  INV_X1 U15831 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15832 ( .A1(n13625), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15833 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12151), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15834 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12279), .B1(
        n12200), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15835 ( .A1(n13838), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n13836), .ZN(n12762) );
  AOI22_X1 U15836 ( .A1(n12152), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12761) );
  NAND4_X1 U15837 ( .A1(n12764), .A2(n12763), .A3(n12762), .A4(n12761), .ZN(
        n12770) );
  AOI22_X1 U15838 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11985), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U15839 ( .A1(n13837), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U15840 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11986), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U15841 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12170), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12765) );
  NAND4_X1 U15842 ( .A1(n12768), .A2(n12767), .A3(n12766), .A4(n12765), .ZN(
        n12769) );
  NOR2_X1 U15843 ( .A1(n12770), .A2(n12769), .ZN(n18973) );
  OR2_X1 U15844 ( .A1(n12771), .A2(n18973), .ZN(n12772) );
  OAI211_X1 U15845 ( .C1(n12150), .C2(n12774), .A(n12773), .B(n12772), .ZN(
        n12775) );
  NOR2_X1 U15846 ( .A1(n12775), .A2(n12776), .ZN(n12777) );
  NOR2_X1 U15847 ( .A1(n12777), .A2(n15231), .ZN(n15261) );
  INV_X1 U15848 ( .A(n15261), .ZN(n18827) );
  INV_X1 U15849 ( .A(n14048), .ZN(n12778) );
  OAI222_X1 U15850 ( .A1(n18827), .A2(n19023), .B1(n12778), .B2(n19065), .C1(
        n19069), .C2(n14810), .ZN(P2_U2905) );
  INV_X1 U15851 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19949) );
  OAI222_X1 U15852 ( .A1(n14268), .A2(n12819), .B1(n20067), .B2(n14273), .C1(
        n14271), .C2(n19949), .ZN(P1_U2903) );
  INV_X1 U15853 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19945) );
  OAI222_X1 U15854 ( .A1(n14268), .A2(n12921), .B1(n20076), .B2(n14273), .C1(
        n14271), .C2(n19945), .ZN(P1_U2901) );
  INV_X1 U15855 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19953) );
  OAI222_X1 U15856 ( .A1(n14268), .A2(n12825), .B1(n20058), .B2(n14273), .C1(
        n14271), .C2(n19953), .ZN(P1_U2904) );
  INV_X1 U15857 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19947) );
  OAI222_X1 U15858 ( .A1(n14268), .A2(n12933), .B1(n20071), .B2(n14273), .C1(
        n14271), .C2(n19947), .ZN(P1_U2902) );
  OR2_X1 U15859 ( .A1(n12781), .A2(n12780), .ZN(n12782) );
  AND2_X1 U15860 ( .A1(n12779), .A2(n12782), .ZN(n19916) );
  INV_X1 U15861 ( .A(n19916), .ZN(n12783) );
  INV_X1 U15862 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19941) );
  OAI222_X1 U15863 ( .A1(n14268), .A2(n12783), .B1(n20084), .B2(n14273), .C1(
        n14271), .C2(n19941), .ZN(P1_U2899) );
  NOR2_X1 U15864 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12943), .ZN(n12784) );
  NOR2_X1 U15865 ( .A1(n12786), .A2(n15735), .ZN(n16219) );
  AOI21_X1 U15866 ( .B1(n19680), .B2(n12784), .A(n16219), .ZN(n12790) );
  NOR4_X1 U15867 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n15409), .ZN(n12785) );
  INV_X1 U15868 ( .A(n18916), .ZN(n18967) );
  NOR2_X1 U15869 ( .A1(n12943), .A2(n19756), .ZN(n18729) );
  AND2_X1 U15870 ( .A1(n15735), .A2(n18729), .ZN(n12787) );
  OAI21_X1 U15871 ( .B1(n12788), .B2(n12787), .A(n12786), .ZN(n12789) );
  OAI211_X1 U15872 ( .C1(n12790), .C2(n15409), .A(n18967), .B(n12789), .ZN(
        P2_U3177) );
  NAND2_X1 U15873 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n10081), .ZN(n12793) );
  NOR2_X1 U15874 ( .A1(n20704), .A2(n20730), .ZN(n15696) );
  NAND2_X1 U15875 ( .A1(n15696), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12791) );
  OAI211_X1 U15876 ( .C1(n12793), .C2(n12792), .A(n20002), .B(n12791), .ZN(
        n12794) );
  NAND2_X1 U15877 ( .A1(n19857), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12796) );
  AOI21_X1 U15878 ( .B1(n12795), .B2(n12810), .A(n19873), .ZN(n19884) );
  INV_X1 U15879 ( .A(n12796), .ZN(n12797) );
  INV_X1 U15880 ( .A(n12800), .ZN(n12801) );
  NAND2_X1 U15881 ( .A1(n12810), .A2(n12801), .ZN(n19893) );
  INV_X1 U15882 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14157) );
  NOR2_X1 U15883 ( .A1(n11313), .A2(n14157), .ZN(n12805) );
  NAND2_X1 U15884 ( .A1(n20726), .A2(n20207), .ZN(n15689) );
  AND2_X1 U15885 ( .A1(n12805), .A2(n15689), .ZN(n12802) );
  OR2_X1 U15886 ( .A1(n12803), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12806) );
  NOR2_X1 U15887 ( .A1(n12806), .A2(n20051), .ZN(n12804) );
  NOR2_X1 U15888 ( .A1(n19891), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n12813) );
  OR2_X1 U15889 ( .A1(n12805), .A2(n20051), .ZN(n12808) );
  INV_X1 U15890 ( .A(n12806), .ZN(n12807) );
  NOR2_X1 U15891 ( .A1(n12808), .A2(n12807), .ZN(n12809) );
  AOI22_X1 U15892 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n19901), .B1(n15758), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n12811) );
  OAI21_X1 U15893 ( .B1(n15826), .B2(n12817), .A(n12811), .ZN(n12812) );
  AOI211_X1 U15894 ( .C1(n19880), .C2(n12814), .A(n12813), .B(n12812), .ZN(
        n12815) );
  OAI21_X1 U15895 ( .B1(n12799), .B2(n19893), .A(n12815), .ZN(n12816) );
  AOI21_X1 U15896 ( .B1(n19838), .B2(n12817), .A(n12816), .ZN(n12818) );
  OAI21_X1 U15897 ( .B1(n19884), .B2(n12819), .A(n12818), .ZN(P1_U2839) );
  INV_X1 U15898 ( .A(n19893), .ZN(n12931) );
  NAND2_X1 U15899 ( .A1(n19891), .A2(n19857), .ZN(n19885) );
  INV_X1 U15900 ( .A(n19885), .ZN(n14137) );
  INV_X1 U15901 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20721) );
  AOI22_X1 U15902 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(n19901), .B1(n19880), .B2(
        n12820), .ZN(n12821) );
  OAI21_X1 U15903 ( .B1(n14137), .B2(n20721), .A(n12821), .ZN(n12822) );
  AOI21_X1 U15904 ( .B1(n20289), .B2(n12931), .A(n12822), .ZN(n12824) );
  OAI21_X1 U15905 ( .B1(n19838), .B2(n19897), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12823) );
  OAI211_X1 U15906 ( .C1(n19884), .C2(n12825), .A(n12824), .B(n12823), .ZN(
        P1_U2840) );
  AND2_X1 U15907 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n13152) );
  NOR2_X1 U15908 ( .A1(n18080), .A2(n15604), .ZN(n18509) );
  NAND3_X1 U15909 ( .A1(n15591), .A2(n12826), .A3(n18509), .ZN(n15589) );
  OAI21_X1 U15910 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18360), .A(
        n12827), .ZN(n15600) );
  NOR2_X1 U15911 ( .A1(n15600), .A2(n12828), .ZN(n12831) );
  INV_X1 U15912 ( .A(n12829), .ZN(n12830) );
  AND3_X1 U15913 ( .A1(n18097), .A2(n18080), .A3(n12832), .ZN(n12833) );
  NOR3_X1 U15914 ( .A1(n18062), .A2(n18057), .A3(n15741), .ZN(n17076) );
  NAND2_X1 U15915 ( .A1(n18097), .A2(n17076), .ZN(n17082) );
  INV_X1 U15916 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16496) );
  INV_X1 U15917 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16517) );
  INV_X1 U15918 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16897) );
  INV_X1 U15919 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17068) );
  NAND2_X1 U15920 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17071) );
  NOR3_X1 U15921 ( .A1(n16743), .A2(n17068), .A3(n17071), .ZN(n17065) );
  NAND2_X1 U15922 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17065), .ZN(n17057) );
  INV_X1 U15923 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17012) );
  NAND2_X1 U15924 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17054) );
  NAND2_X1 U15925 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .ZN(n16970) );
  NOR4_X1 U15926 ( .A1(n16997), .A2(n17012), .A3(n17054), .A4(n16970), .ZN(
        n12834) );
  NAND3_X1 U15927 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n12834), .ZN(n15474) );
  NAND4_X1 U15928 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(P3_EBX_REG_13__SCAN_IN), .ZN(n12835)
         );
  NOR3_X1 U15929 ( .A1(n17057), .A2(n15474), .A3(n12835), .ZN(n16921) );
  NAND3_X1 U15930 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17076), .A3(n16921), 
        .ZN(n16896) );
  NAND2_X1 U15931 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16895), .ZN(n16893) );
  NOR2_X1 U15932 ( .A1(n17163), .A2(n16893), .ZN(n16880) );
  NAND2_X1 U15933 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16880), .ZN(n16868) );
  NOR2_X1 U15934 ( .A1(n16526), .A2(n16868), .ZN(n16840) );
  NAND2_X1 U15935 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16840), .ZN(n16834) );
  NAND2_X1 U15936 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16839), .ZN(n16824) );
  NOR2_X1 U15937 ( .A1(n16496), .A2(n16824), .ZN(n16828) );
  NAND2_X1 U15938 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16828), .ZN(n16818) );
  NAND2_X1 U15939 ( .A1(n17075), .A2(n16818), .ZN(n12836) );
  OAI21_X1 U15940 ( .B1(n13152), .B2(n17082), .A(n12836), .ZN(n16813) );
  AOI22_X1 U15941 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U15942 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U15943 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U15944 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12837) );
  NAND4_X1 U15945 ( .A1(n12840), .A2(n12839), .A3(n12838), .A4(n12837), .ZN(
        n12846) );
  AOI22_X1 U15946 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12844) );
  AOI22_X1 U15947 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U15948 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15949 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12841) );
  NAND4_X1 U15950 ( .A1(n12844), .A2(n12843), .A3(n12842), .A4(n12841), .ZN(
        n12845) );
  NOR2_X1 U15951 ( .A1(n12846), .A2(n12845), .ZN(n12909) );
  AOI22_X1 U15952 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U15953 ( .A1(n9790), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U15954 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12848) );
  AOI22_X1 U15955 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12847) );
  NAND4_X1 U15956 ( .A1(n12850), .A2(n12849), .A3(n12848), .A4(n12847), .ZN(
        n12856) );
  AOI22_X1 U15957 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U15958 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U15959 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15960 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12851) );
  NAND4_X1 U15961 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12855) );
  NOR2_X1 U15962 ( .A1(n12856), .A2(n12855), .ZN(n16820) );
  AOI22_X1 U15963 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12860) );
  AOI22_X1 U15964 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12859) );
  AOI22_X1 U15965 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U15966 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12857) );
  NAND4_X1 U15967 ( .A1(n12860), .A2(n12859), .A3(n12858), .A4(n12857), .ZN(
        n12866) );
  AOI22_X1 U15968 ( .A1(n17004), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U15969 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U15970 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U15971 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12861) );
  NAND4_X1 U15972 ( .A1(n12864), .A2(n12863), .A3(n12862), .A4(n12861), .ZN(
        n12865) );
  NOR2_X1 U15973 ( .A1(n12866), .A2(n12865), .ZN(n16830) );
  AOI22_X1 U15974 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U15975 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12875) );
  INV_X1 U15976 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18061) );
  AOI22_X1 U15977 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12867) );
  OAI21_X1 U15978 ( .B1(n9840), .B2(n18061), .A(n12867), .ZN(n12873) );
  AOI22_X1 U15979 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U15980 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U15981 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U15982 ( .A1(n9790), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12868) );
  NAND4_X1 U15983 ( .A1(n12871), .A2(n12870), .A3(n12869), .A4(n12868), .ZN(
        n12872) );
  AOI211_X1 U15984 ( .C1(n17036), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n12873), .B(n12872), .ZN(n12874) );
  NAND3_X1 U15985 ( .A1(n12876), .A2(n12875), .A3(n12874), .ZN(n16836) );
  AOI22_X1 U15986 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U15987 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12886) );
  INV_X1 U15988 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n21017) );
  AOI22_X1 U15989 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12877) );
  OAI21_X1 U15990 ( .B1(n16899), .B2(n21017), .A(n12877), .ZN(n12884) );
  AOI22_X1 U15991 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12882) );
  AOI22_X1 U15992 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12881) );
  AOI22_X1 U15993 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U15994 ( .A1(n17004), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12879) );
  NAND4_X1 U15995 ( .A1(n12882), .A2(n12881), .A3(n12880), .A4(n12879), .ZN(
        n12883) );
  AOI211_X1 U15996 ( .C1(n9790), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n12884), .B(n12883), .ZN(n12885) );
  NAND3_X1 U15997 ( .A1(n12887), .A2(n12886), .A3(n12885), .ZN(n16837) );
  NAND2_X1 U15998 ( .A1(n16836), .A2(n16837), .ZN(n16835) );
  NOR2_X1 U15999 ( .A1(n16830), .A2(n16835), .ZN(n16829) );
  AOI22_X1 U16000 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n17015), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16001 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n15486), .B1(
        P3_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n17004), .ZN(n12897) );
  AOI22_X1 U16002 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n17021), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12888) );
  OAI21_X1 U16003 ( .B1(n9840), .B2(n18072), .A(n12888), .ZN(n12895) );
  AOI22_X1 U16004 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__2__SCAN_IN), .B2(n15546), .ZN(n12893) );
  AOI22_X1 U16005 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U16006 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__2__SCAN_IN), .B2(n17036), .ZN(n12891) );
  AOI22_X1 U16007 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n17003), .B1(
        P3_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n9787), .ZN(n12890) );
  NAND4_X1 U16008 ( .A1(n12893), .A2(n12892), .A3(n12891), .A4(n12890), .ZN(
        n12894) );
  AOI211_X1 U16009 ( .C1(n17035), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n12895), .B(n12894), .ZN(n12896) );
  NAND3_X1 U16010 ( .A1(n12898), .A2(n12897), .A3(n12896), .ZN(n16826) );
  NAND2_X1 U16011 ( .A1(n16829), .A2(n16826), .ZN(n16825) );
  NOR2_X1 U16012 ( .A1(n16820), .A2(n16825), .ZN(n16819) );
  AOI22_X1 U16013 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U16014 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12907) );
  INV_X1 U16015 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18083) );
  AOI22_X1 U16016 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12899) );
  OAI21_X1 U16017 ( .B1(n9840), .B2(n18083), .A(n12899), .ZN(n12905) );
  AOI22_X1 U16018 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U16019 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U16020 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U16021 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12900) );
  NAND4_X1 U16022 ( .A1(n12903), .A2(n12902), .A3(n12901), .A4(n12900), .ZN(
        n12904) );
  NAND3_X1 U16023 ( .A1(n12908), .A2(n12907), .A3(n12906), .ZN(n16816) );
  NAND2_X1 U16024 ( .A1(n16819), .A2(n16816), .ZN(n16815) );
  NOR2_X1 U16025 ( .A1(n12909), .A2(n16815), .ZN(n16809) );
  AOI21_X1 U16026 ( .B1(n12909), .B2(n16815), .A(n16809), .ZN(n17097) );
  AOI22_X1 U16027 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16813), .B1(n17097), 
        .B2(n17080), .ZN(n12912) );
  INV_X1 U16028 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n12910) );
  INV_X1 U16029 ( .A(n16818), .ZN(n16823) );
  NAND3_X1 U16030 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n12910), .A3(n16823), 
        .ZN(n12911) );
  NAND2_X1 U16031 ( .A1(n12912), .A2(n12911), .ZN(P3_U2675) );
  INV_X1 U16032 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20649) );
  NAND4_X1 U16033 ( .A1(n19878), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .A4(n20649), .ZN(n12913) );
  OAI21_X1 U16034 ( .B1(n15826), .B2(n20866), .A(n12913), .ZN(n12915) );
  NAND2_X1 U16035 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n12923) );
  AOI21_X1 U16036 ( .B1(n19878), .B2(n12923), .A(n15758), .ZN(n12927) );
  NOR2_X1 U16037 ( .A1(n12927), .A2(n20649), .ZN(n12914) );
  AOI211_X1 U16038 ( .C1(n19901), .C2(P1_EBX_REG_3__SCAN_IN), .A(n12915), .B(
        n12914), .ZN(n12916) );
  OAI21_X1 U16039 ( .B1(n19892), .B2(n20011), .A(n12916), .ZN(n12919) );
  NOR2_X1 U16040 ( .A1(n19906), .A2(n12917), .ZN(n12918) );
  AOI211_X1 U16041 ( .C1(n12931), .C2(n20323), .A(n12919), .B(n12918), .ZN(
        n12920) );
  OAI21_X1 U16042 ( .B1(n19884), .B2(n12921), .A(n12920), .ZN(P1_U2837) );
  INV_X1 U16043 ( .A(n12324), .ZN(n20055) );
  INV_X1 U16044 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n12926) );
  INV_X1 U16045 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20991) );
  OAI22_X1 U16046 ( .A1(n20991), .A2(n15826), .B1(n19892), .B2(n20021), .ZN(
        n12922) );
  AOI21_X1 U16047 ( .B1(n19901), .B2(P1_EBX_REG_2__SCAN_IN), .A(n12922), .ZN(
        n12925) );
  NAND3_X1 U16048 ( .A1(n19878), .A2(n12923), .A3(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n12924) );
  OAI211_X1 U16049 ( .C1(n12927), .C2(n12926), .A(n12925), .B(n12924), .ZN(
        n12930) );
  NOR2_X1 U16050 ( .A1(n19906), .A2(n12928), .ZN(n12929) );
  AOI211_X1 U16051 ( .C1(n12931), .C2(n20055), .A(n12930), .B(n12929), .ZN(
        n12932) );
  OAI21_X1 U16052 ( .B1(n19884), .B2(n12933), .A(n12932), .ZN(P1_U2838) );
  XOR2_X1 U16053 ( .A(n12779), .B(n12934), .Z(n19874) );
  INV_X1 U16054 ( .A(n19874), .ZN(n12981) );
  OAI222_X1 U16055 ( .A1(n14268), .A2(n12981), .B1(n14271), .B2(n10679), .C1(
        n14273), .C2(n20087), .ZN(P1_U2898) );
  NAND2_X1 U16056 ( .A1(n12936), .A2(n12935), .ZN(n12937) );
  NAND2_X1 U16057 ( .A1(n12937), .A2(n12476), .ZN(n12939) );
  AOI21_X1 U16058 ( .B1(n15036), .B2(n12945), .A(n13033), .ZN(n15034) );
  INV_X1 U16059 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13646) );
  INV_X1 U16060 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18812) );
  INV_X1 U16061 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14965) );
  INV_X1 U16062 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14906) );
  INV_X1 U16063 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14887) );
  INV_X1 U16064 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14539) );
  INV_X1 U16065 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14868) );
  INV_X1 U16066 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14827) );
  INV_X1 U16067 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18959) );
  INV_X1 U16068 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16069 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15408), .B1(n18959), 
        .B2(n12943), .ZN(n15407) );
  AOI22_X1 U16070 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12944), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12943), .ZN(n14687) );
  NOR2_X1 U16071 ( .A1(n15407), .A2(n14687), .ZN(n14686) );
  OAI21_X1 U16072 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12945), .ZN(n13673) );
  NAND2_X1 U16073 ( .A1(n14686), .A2(n13673), .ZN(n13031) );
  NAND2_X1 U16074 ( .A1(n18912), .A2(n13031), .ZN(n12946) );
  XNOR2_X1 U16075 ( .A(n15034), .B(n12946), .ZN(n12947) );
  NAND2_X1 U16076 ( .A1(n12947), .A2(n18916), .ZN(n12978) );
  OR2_X1 U16077 ( .A1(n18730), .A2(n12948), .ZN(n12953) );
  INV_X1 U16078 ( .A(n12953), .ZN(n12950) );
  INV_X1 U16079 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19574) );
  NAND2_X1 U16080 ( .A1(n19574), .A2(n15735), .ZN(n12951) );
  INV_X1 U16081 ( .A(n12951), .ZN(n12949) );
  NAND2_X1 U16082 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12951), .ZN(n12952) );
  NOR2_X2 U16083 ( .A1(n12953), .A2(n12952), .ZN(n18954) );
  NAND2_X1 U16084 ( .A1(n13041), .A2(n12955), .ZN(n12959) );
  NAND2_X1 U16085 ( .A1(n13039), .A2(n12956), .ZN(n12958) );
  NAND2_X1 U16086 ( .A1(n13502), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n12957) );
  OR2_X1 U16087 ( .A1(n13067), .A2(n12960), .ZN(n12961) );
  NAND2_X1 U16088 ( .A1(n13341), .A2(n12961), .ZN(n13330) );
  OAI21_X1 U16089 ( .B1(n12964), .B2(n12963), .A(n12962), .ZN(n19033) );
  INV_X1 U16090 ( .A(n19033), .ZN(n19767) );
  NAND2_X1 U16091 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19390), .ZN(n19184) );
  NOR2_X1 U16092 ( .A1(n12965), .A2(n19184), .ZN(n16224) );
  OR2_X1 U16093 ( .A1(n19132), .A2(n18916), .ZN(n12966) );
  NOR2_X1 U16094 ( .A1(n16224), .A2(n12966), .ZN(n12967) );
  AND2_X2 U16095 ( .A1(n18730), .A2(n12967), .ZN(n18949) );
  AOI22_X1 U16096 ( .A1(n18952), .A2(n19767), .B1(n18928), .B2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12975) );
  INV_X1 U16097 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16093) );
  OAI21_X1 U16098 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19680), .A(n16093), 
        .ZN(n12968) );
  NOR2_X1 U16099 ( .A1(n12969), .A2(n12968), .ZN(n12970) );
  OR2_X1 U16100 ( .A1(n19100), .A2(n12970), .ZN(n12973) );
  INV_X1 U16101 ( .A(n12971), .ZN(n12972) );
  AOI22_X1 U16102 ( .A1(n18950), .A2(P2_EBX_REG_3__SCAN_IN), .B1(n18949), .B2(
        P2_REIP_REG_3__SCAN_IN), .ZN(n12974) );
  OAI211_X1 U16103 ( .C1(n18907), .C2(n13330), .A(n12975), .B(n12974), .ZN(
        n12976) );
  AOI21_X1 U16104 ( .B1(n13263), .B2(n18939), .A(n12976), .ZN(n12977) );
  OAI211_X1 U16105 ( .C1(n19423), .C2(n14703), .A(n12978), .B(n12977), .ZN(
        P2_U2852) );
  OR2_X1 U16106 ( .A1(n16029), .A2(n12979), .ZN(n12980) );
  NAND2_X1 U16107 ( .A1(n12989), .A2(n12980), .ZN(n19865) );
  INV_X1 U16108 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19867) );
  OAI222_X1 U16109 ( .A1(n19865), .A2(n19912), .B1(n19919), .B2(n19867), .C1(
        n9794), .C2(n12981), .ZN(P1_U2866) );
  INV_X1 U16110 ( .A(n12983), .ZN(n12985) );
  NAND2_X1 U16111 ( .A1(n12985), .A2(n12984), .ZN(n12986) );
  AND2_X1 U16112 ( .A1(n12982), .A2(n12986), .ZN(n19861) );
  INV_X1 U16113 ( .A(n19861), .ZN(n12987) );
  OAI222_X1 U16114 ( .A1(n12987), .A2(n14268), .B1(n14271), .B2(n10615), .C1(
        n20095), .C2(n14273), .ZN(P1_U2897) );
  NAND2_X1 U16115 ( .A1(n12989), .A2(n12988), .ZN(n12990) );
  NAND2_X1 U16116 ( .A1(n13076), .A2(n12990), .ZN(n19855) );
  OAI22_X1 U16117 ( .A1(n19855), .A2(n19912), .B1(n19864), .B2(n19919), .ZN(
        n12991) );
  AOI21_X1 U16118 ( .B1(n19861), .B2(n19915), .A(n12991), .ZN(n12992) );
  INV_X1 U16119 ( .A(n12992), .ZN(P1_U2865) );
  INV_X1 U16120 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n18811) );
  AOI22_X1 U16121 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n13836), .ZN(n12997) );
  AOI22_X1 U16122 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U16123 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U16124 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12994) );
  NAND4_X1 U16125 ( .A1(n12997), .A2(n12996), .A3(n12995), .A4(n12994), .ZN(
        n13003) );
  AOI22_X1 U16126 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U16127 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U16128 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11986), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U16129 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12206), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12998) );
  NAND4_X1 U16130 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13002) );
  OAI211_X1 U16131 ( .C1(n13004), .C2(n13603), .A(n13722), .B(n18998), .ZN(
        n13014) );
  INV_X1 U16132 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n18824) );
  NAND2_X1 U16133 ( .A1(n13595), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n13006) );
  NAND2_X1 U16134 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13005) );
  OAI211_X1 U16135 ( .C1(n13598), .C2(n18824), .A(n13006), .B(n13005), .ZN(
        n13007) );
  AOI21_X1 U16136 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n13007), .ZN(n15257) );
  NAND2_X1 U16137 ( .A1(n13595), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n13009) );
  NAND2_X1 U16138 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n13008) );
  OAI211_X1 U16139 ( .C1(n13598), .C2(n18811), .A(n13009), .B(n13008), .ZN(
        n13010) );
  AOI21_X1 U16140 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n13010), .ZN(n13011) );
  NOR2_X4 U16141 ( .A1(n15260), .A2(n13011), .ZN(n14665) );
  AND2_X1 U16142 ( .A1(n15260), .A2(n13011), .ZN(n13012) );
  NOR2_X1 U16143 ( .A1(n14665), .A2(n13012), .ZN(n18817) );
  NAND2_X1 U16144 ( .A1(n18817), .A2(n19000), .ZN(n13013) );
  OAI211_X1 U16145 ( .C1(n19000), .C2(n18811), .A(n13014), .B(n13013), .ZN(
        P2_U2872) );
  XNOR2_X1 U16146 ( .A(n13015), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13016) );
  XNOR2_X1 U16147 ( .A(n13017), .B(n13016), .ZN(n15917) );
  INV_X1 U16148 ( .A(n15917), .ZN(n13026) );
  NAND2_X1 U16149 ( .A1(n20005), .A2(n13018), .ZN(n16035) );
  OAI21_X1 U16150 ( .B1(n13019), .B2(n20024), .A(n20000), .ZN(n15992) );
  AOI21_X1 U16151 ( .B1(n20035), .B2(n13020), .A(n15992), .ZN(n16030) );
  OAI211_X1 U16152 ( .C1(n13021), .C2(n16035), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16030), .ZN(n16011) );
  OAI21_X1 U16153 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16014), .A(
        n16011), .ZN(n13025) );
  INV_X1 U16154 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n13022) );
  OAI22_X1 U16155 ( .A1(n19865), .A2(n20003), .B1(n20002), .B2(n13022), .ZN(
        n13023) );
  INV_X1 U16156 ( .A(n13023), .ZN(n13024) );
  OAI211_X1 U16157 ( .C1(n13026), .C2(n15966), .A(n13025), .B(n13024), .ZN(
        P1_U3025) );
  OR2_X1 U16158 ( .A1(n13027), .A2(n13028), .ZN(n13030) );
  NAND2_X1 U16159 ( .A1(n13030), .A2(n13029), .ZN(n18997) );
  AOI21_X1 U16160 ( .B1(n15026), .B2(n13034), .A(n9870), .ZN(n18882) );
  AOI21_X1 U16161 ( .B1(n18906), .B2(n13032), .A(n13035), .ZN(n18914) );
  NOR2_X1 U16162 ( .A1(n15034), .A2(n13031), .ZN(n18940) );
  OAI21_X1 U16163 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13033), .A(
        n13032), .ZN(n19119) );
  NAND2_X1 U16164 ( .A1(n18940), .A2(n19119), .ZN(n18911) );
  NOR2_X1 U16165 ( .A1(n18914), .A2(n18911), .ZN(n18898) );
  OAI21_X1 U16166 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13035), .A(
        n13034), .ZN(n18899) );
  NAND2_X1 U16167 ( .A1(n18898), .A2(n18899), .ZN(n18881) );
  NOR2_X1 U16168 ( .A1(n18882), .A2(n18881), .ZN(n14545) );
  NOR2_X1 U16169 ( .A1(n18941), .A2(n14545), .ZN(n13036) );
  OAI21_X1 U16170 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n9870), .A(
        n14544), .ZN(n16170) );
  XNOR2_X1 U16171 ( .A(n13036), .B(n16170), .ZN(n13037) );
  NAND2_X1 U16172 ( .A1(n13037), .A2(n18916), .ZN(n13053) );
  AOI22_X1 U16173 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18928), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18949), .ZN(n13038) );
  OAI211_X1 U16174 ( .C1(n18920), .C2(n15351), .A(n13038), .B(n18905), .ZN(
        n13051) );
  INV_X1 U16175 ( .A(n13039), .ZN(n13045) );
  INV_X1 U16176 ( .A(n13040), .ZN(n13044) );
  NAND2_X1 U16177 ( .A1(n13041), .A2(n13298), .ZN(n13043) );
  NAND2_X1 U16178 ( .A1(n13502), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13042) );
  OAI211_X1 U16179 ( .C1(n13045), .C2(n13044), .A(n13043), .B(n13042), .ZN(
        n13340) );
  MUX2_X1 U16180 ( .A(n13320), .B(P2_EBX_REG_5__SCAN_IN), .S(n13502), .Z(
        n13324) );
  MUX2_X1 U16181 ( .A(n13046), .B(n18894), .S(n13502), .Z(n13379) );
  MUX2_X1 U16182 ( .A(n13510), .B(n13047), .S(n13502), .Z(n13384) );
  NAND2_X1 U16183 ( .A1(n13395), .A2(n13048), .ZN(n13049) );
  NAND2_X1 U16184 ( .A1(n13389), .A2(n13049), .ZN(n13387) );
  NOR2_X1 U16185 ( .A1(n13387), .A2(n18907), .ZN(n13050) );
  AOI211_X1 U16186 ( .C1(n18950), .C2(P2_EBX_REG_8__SCAN_IN), .A(n13051), .B(
        n13050), .ZN(n13052) );
  OAI211_X1 U16187 ( .C1(n18957), .C2(n18997), .A(n13053), .B(n13052), .ZN(
        P2_U2847) );
  NOR2_X1 U16188 ( .A1(n18941), .A2(n14686), .ZN(n13057) );
  XNOR2_X1 U16189 ( .A(n13057), .B(n13673), .ZN(n13058) );
  NAND2_X1 U16190 ( .A1(n13058), .A2(n18916), .ZN(n13073) );
  NAND2_X1 U16191 ( .A1(n13060), .A2(n13059), .ZN(n13063) );
  INV_X1 U16192 ( .A(n13061), .ZN(n13062) );
  NAND2_X1 U16193 ( .A1(n13063), .A2(n13062), .ZN(n19775) );
  AND2_X1 U16194 ( .A1(n13065), .A2(n13064), .ZN(n13066) );
  NOR2_X1 U16195 ( .A1(n13067), .A2(n13066), .ZN(n13336) );
  NAND2_X1 U16196 ( .A1(n13336), .A2(n18954), .ZN(n13069) );
  AOI22_X1 U16197 ( .A1(n18949), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18928), .ZN(n13068) );
  OAI211_X1 U16198 ( .C1(n12447), .C2(n18925), .A(n13069), .B(n13068), .ZN(
        n13071) );
  NOR2_X1 U16199 ( .A1(n13691), .A2(n18957), .ZN(n13070) );
  AOI211_X1 U16200 ( .C1(n18952), .C2(n19775), .A(n13071), .B(n13070), .ZN(
        n13072) );
  OAI211_X1 U16201 ( .C1(n14703), .C2(n19772), .A(n13073), .B(n13072), .ZN(
        P2_U2853) );
  AND2_X1 U16202 ( .A1(n12982), .A2(n13074), .ZN(n13075) );
  OR2_X1 U16203 ( .A1(n13075), .A2(n9873), .ZN(n19848) );
  INV_X1 U16204 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13077) );
  OAI21_X1 U16205 ( .B1(n10166), .B2(n9910), .A(n16001), .ZN(n19844) );
  OAI222_X1 U16206 ( .A1(n19848), .A2(n9794), .B1(n19919), .B2(n13077), .C1(
        n19844), .C2(n19912), .ZN(P1_U2864) );
  INV_X1 U16207 ( .A(DATAI_8_), .ZN(n13078) );
  MUX2_X1 U16208 ( .A(n13078), .B(n16338), .S(n20045), .Z(n19954) );
  INV_X1 U16209 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13079) );
  OAI222_X1 U16210 ( .A1(n14268), .A2(n19848), .B1(n19954), .B2(n14273), .C1(
        n13079), .C2(n14271), .ZN(P1_U2896) );
  NOR2_X1 U16211 ( .A1(n9873), .A2(n13081), .ZN(n13082) );
  OR2_X1 U16212 ( .A1(n13080), .A2(n13082), .ZN(n19836) );
  INV_X1 U16213 ( .A(n14273), .ZN(n13127) );
  INV_X1 U16214 ( .A(DATAI_9_), .ZN(n13084) );
  NAND2_X1 U16215 ( .A1(n20045), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13083) );
  OAI21_X1 U16216 ( .B1(n20045), .B2(n13084), .A(n13083), .ZN(n19957) );
  AOI22_X1 U16217 ( .A1(n13127), .A2(n19957), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14235), .ZN(n13085) );
  OAI21_X1 U16218 ( .B1(n19836), .B2(n14268), .A(n13085), .ZN(P1_U2895) );
  XOR2_X1 U16219 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13086), .Z(
        n13087) );
  XNOR2_X1 U16220 ( .A(n13088), .B(n13087), .ZN(n16013) );
  INV_X1 U16221 ( .A(n19848), .ZN(n13091) );
  AOI22_X1 U16222 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20033), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13089) );
  OAI21_X1 U16223 ( .B1(n19998), .B2(n19846), .A(n13089), .ZN(n13090) );
  AOI21_X1 U16224 ( .B1(n13091), .B2(n19993), .A(n13090), .ZN(n13092) );
  OAI21_X1 U16225 ( .B1(n16013), .B2(n19817), .A(n13092), .ZN(P1_U2991) );
  INV_X1 U16226 ( .A(n13093), .ZN(n13094) );
  OAI21_X1 U16227 ( .B1(n13080), .B2(n13095), .A(n13094), .ZN(n15845) );
  OR2_X1 U16228 ( .A1(n16003), .A2(n13096), .ZN(n13097) );
  NAND2_X1 U16229 ( .A1(n13112), .A2(n13097), .ZN(n15994) );
  OAI22_X1 U16230 ( .A1(n15994), .A2(n19912), .B1(n15841), .B2(n19919), .ZN(
        n13098) );
  INV_X1 U16231 ( .A(n13098), .ZN(n13099) );
  OAI21_X1 U16232 ( .B1(n15845), .B2(n9794), .A(n13099), .ZN(P1_U2862) );
  INV_X1 U16233 ( .A(DATAI_10_), .ZN(n13100) );
  MUX2_X1 U16234 ( .A(n13100), .B(n21043), .S(n20045), .Z(n19960) );
  INV_X1 U16235 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13101) );
  OAI222_X1 U16236 ( .A1(n14268), .A2(n15845), .B1(n19960), .B2(n14273), .C1(
        n13101), .C2(n14271), .ZN(P1_U2894) );
  XNOR2_X1 U16237 ( .A(n11179), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13102) );
  XNOR2_X1 U16238 ( .A(n13103), .B(n13102), .ZN(n15999) );
  INV_X1 U16239 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13105) );
  INV_X1 U16240 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n13104) );
  OAI22_X1 U16241 ( .A1(n15871), .A2(n13105), .B1(n20002), .B2(n13104), .ZN(
        n13107) );
  NOR2_X1 U16242 ( .A1(n19836), .A2(n20044), .ZN(n13106) );
  AOI211_X1 U16243 ( .C1(n15899), .C2(n19837), .A(n13107), .B(n13106), .ZN(
        n13108) );
  OAI21_X1 U16244 ( .B1(n15999), .B2(n19817), .A(n13108), .ZN(P1_U2990) );
  OAI21_X1 U16245 ( .B1(n13093), .B2(n13110), .A(n13109), .ZN(n13122) );
  XNOR2_X1 U16246 ( .A(n13122), .B(n13120), .ZN(n15907) );
  INV_X1 U16247 ( .A(n15907), .ZN(n13119) );
  INV_X1 U16248 ( .A(n13130), .ZN(n13111) );
  AOI21_X1 U16249 ( .B1(n13113), .B2(n13112), .A(n13111), .ZN(n15982) );
  INV_X1 U16250 ( .A(n19912), .ZN(n19908) );
  AOI22_X1 U16251 ( .A1(n15982), .A2(n19908), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14188), .ZN(n13114) );
  OAI21_X1 U16252 ( .B1(n13119), .B2(n9794), .A(n13114), .ZN(P1_U2861) );
  INV_X1 U16253 ( .A(DATAI_11_), .ZN(n13116) );
  NAND2_X1 U16254 ( .A1(n20045), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13115) );
  OAI21_X1 U16255 ( .B1(n20045), .B2(n13116), .A(n13115), .ZN(n19963) );
  INV_X1 U16256 ( .A(n19963), .ZN(n13118) );
  OAI222_X1 U16257 ( .A1(n13119), .A2(n14268), .B1(n13118), .B2(n14273), .C1(
        n13117), .C2(n14271), .ZN(P1_U2893) );
  INV_X1 U16258 ( .A(n13120), .ZN(n13121) );
  OAI21_X1 U16259 ( .B1(n13122), .B2(n13121), .A(n13109), .ZN(n13124) );
  NAND2_X1 U16260 ( .A1(n13124), .A2(n13123), .ZN(n13137) );
  OAI21_X1 U16261 ( .B1(n13124), .B2(n13123), .A(n13137), .ZN(n15829) );
  INV_X1 U16262 ( .A(DATAI_12_), .ZN(n13126) );
  NAND2_X1 U16263 ( .A1(n20045), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13125) );
  OAI21_X1 U16264 ( .B1(n20045), .B2(n13126), .A(n13125), .ZN(n19965) );
  AOI22_X1 U16265 ( .A1(n13127), .A2(n19965), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14235), .ZN(n13128) );
  OAI21_X1 U16266 ( .B1(n15829), .B2(n14268), .A(n13128), .ZN(P1_U2892) );
  INV_X1 U16267 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n13132) );
  AND2_X1 U16268 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  OR2_X1 U16269 ( .A1(n13131), .A2(n13139), .ZN(n15825) );
  OAI222_X1 U16270 ( .A1(n15829), .A2(n9794), .B1(n13132), .B2(n19919), .C1(
        n19912), .C2(n15825), .ZN(P1_U2860) );
  INV_X1 U16271 ( .A(n13133), .ZN(n13136) );
  INV_X1 U16272 ( .A(n13134), .ZN(n13135) );
  AOI21_X1 U16273 ( .B1(n13137), .B2(n13136), .A(n13135), .ZN(n14380) );
  INV_X1 U16274 ( .A(n14380), .ZN(n13143) );
  INV_X1 U16275 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n13141) );
  NOR2_X1 U16276 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  OR2_X1 U16277 ( .A1(n14208), .A2(n13140), .ZN(n13145) );
  OAI222_X1 U16278 ( .A1(n9794), .A2(n13143), .B1(n13141), .B2(n19919), .C1(
        n13145), .C2(n19912), .ZN(P1_U2859) );
  INV_X1 U16279 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n13142) );
  OAI222_X1 U16280 ( .A1(n14268), .A2(n13143), .B1(n14213), .B2(n14273), .C1(
        n13142), .C2(n14271), .ZN(P1_U2891) );
  NAND4_X1 U16281 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(P1_REIP_REG_10__SCAN_IN), .A4(P1_REIP_REG_9__SCAN_IN), .ZN(n13201)
         );
  INV_X1 U16282 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20654) );
  INV_X1 U16283 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20647) );
  NAND3_X1 U16284 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19890) );
  NOR2_X1 U16285 ( .A1(n20647), .A2(n19890), .ZN(n19877) );
  NAND3_X1 U16286 ( .A1(n19877), .A2(P1_REIP_REG_6__SCAN_IN), .A3(
        P1_REIP_REG_5__SCAN_IN), .ZN(n19854) );
  NOR2_X1 U16287 ( .A1(n20654), .A2(n19854), .ZN(n19841) );
  NAND2_X1 U16288 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19841), .ZN(n13202) );
  NOR2_X1 U16289 ( .A1(n19891), .A2(n13202), .ZN(n15840) );
  INV_X1 U16290 ( .A(n15840), .ZN(n19834) );
  NOR3_X1 U16291 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n13201), .A3(n19834), 
        .ZN(n13150) );
  INV_X1 U16292 ( .A(n13144), .ZN(n14378) );
  INV_X1 U16293 ( .A(n13145), .ZN(n15976) );
  NOR2_X2 U16294 ( .A1(n15758), .A2(n19814), .ZN(n19895) );
  INV_X1 U16295 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20662) );
  OAI21_X1 U16296 ( .B1(n13201), .B2(n19832), .A(n19885), .ZN(n15832) );
  AOI22_X1 U16297 ( .A1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19897), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(n19901), .ZN(n13146) );
  OAI21_X1 U16298 ( .B1(n20662), .B2(n15832), .A(n13146), .ZN(n13147) );
  AOI211_X1 U16299 ( .C1(n19880), .C2(n15976), .A(n19895), .B(n13147), .ZN(
        n13148) );
  OAI21_X1 U16300 ( .B1(n14378), .B2(n19906), .A(n13148), .ZN(n13149) );
  AOI211_X1 U16301 ( .C1(n14380), .C2(n19873), .A(n13150), .B(n13149), .ZN(
        n13151) );
  INV_X1 U16302 ( .A(n13151), .ZN(P1_U2827) );
  INV_X1 U16303 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n13155) );
  NAND3_X1 U16304 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n13152), .ZN(n16810) );
  INV_X1 U16305 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n13153) );
  NOR2_X1 U16306 ( .A1(n13153), .A2(n16893), .ZN(n16855) );
  NAND4_X1 U16307 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n16855), .ZN(n13154) );
  NOR4_X1 U16308 ( .A1(n13155), .A2(n16517), .A3(n16810), .A4(n13154), .ZN(
        n16804) );
  NAND2_X1 U16309 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16804), .ZN(n13156) );
  NOR2_X1 U16310 ( .A1(n17163), .A2(n13156), .ZN(n13158) );
  NAND2_X1 U16311 ( .A1(n17075), .A2(n13156), .ZN(n16805) );
  INV_X1 U16312 ( .A(n16805), .ZN(n13157) );
  MUX2_X1 U16313 ( .A(n13158), .B(n13157), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  NAND2_X1 U16314 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15950) );
  NOR2_X1 U16315 ( .A1(n15943), .A2(n15950), .ZN(n13161) );
  INV_X1 U16316 ( .A(n13162), .ZN(n14511) );
  AOI221_X1 U16317 ( .B1(n13159), .B2(n20001), .C1(n20024), .C2(n20001), .A(
        n15970), .ZN(n13160) );
  AOI211_X1 U16318 ( .C1(n20982), .C2(n14511), .A(n13160), .B(n15992), .ZN(
        n15960) );
  OAI21_X1 U16319 ( .B1(n13162), .B2(n13161), .A(n15960), .ZN(n15945) );
  INV_X1 U16320 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20671) );
  NOR2_X1 U16321 ( .A1(n20002), .A2(n20671), .ZN(n13170) );
  OAI21_X1 U16322 ( .B1(n13165), .B2(n13164), .A(n13163), .ZN(n14340) );
  NAND2_X1 U16323 ( .A1(n14144), .A2(n13167), .ZN(n13168) );
  NAND2_X1 U16324 ( .A1(n14185), .A2(n13168), .ZN(n15802) );
  OAI22_X1 U16325 ( .A1(n14340), .A2(n15966), .B1(n20003), .B2(n15802), .ZN(
        n13169) );
  AOI211_X1 U16326 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15945), .A(
        n13170), .B(n13169), .ZN(n13175) );
  INV_X1 U16327 ( .A(n13171), .ZN(n13173) );
  INV_X1 U16328 ( .A(n15942), .ZN(n13172) );
  NAND3_X1 U16329 ( .A1(n13173), .A2(n11362), .A3(n13172), .ZN(n13174) );
  NAND2_X1 U16330 ( .A1(n13175), .A2(n13174), .ZN(P1_U3013) );
  OAI21_X1 U16331 ( .B1(n13176), .B2(n11599), .A(n18504), .ZN(n13189) );
  NAND2_X1 U16332 ( .A1(n18521), .A2(n13189), .ZN(n18503) );
  NOR2_X1 U16333 ( .A1(n18670), .A2(n18503), .ZN(n13188) );
  NOR2_X1 U16334 ( .A1(n18708), .A2(n17279), .ZN(n18552) );
  INV_X1 U16335 ( .A(n18577), .ZN(n18707) );
  OAI21_X1 U16336 ( .B1(n13177), .B2(n18552), .A(n18707), .ZN(n17238) );
  INV_X1 U16337 ( .A(n18496), .ZN(n16401) );
  AOI211_X1 U16338 ( .C1(n15743), .C2(n17238), .A(n16401), .B(n18709), .ZN(
        n13185) );
  INV_X1 U16339 ( .A(n13178), .ZN(n16392) );
  OAI211_X1 U16340 ( .C1(n18080), .C2(n18530), .A(n15591), .B(n13179), .ZN(
        n13180) );
  NOR3_X1 U16341 ( .A1(n13182), .A2(n13181), .A3(n13180), .ZN(n13184) );
  OAI21_X1 U16342 ( .B1(n16392), .B2(n13184), .A(n13183), .ZN(n15610) );
  INV_X1 U16343 ( .A(n18539), .ZN(n18528) );
  NOR2_X1 U16344 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18684), .ZN(n18056) );
  INV_X1 U16345 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16403) );
  NAND3_X1 U16346 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18658)
         );
  NOR2_X1 U16347 ( .A1(n16403), .A2(n18658), .ZN(n13187) );
  AOI211_X2 U16348 ( .C1(n18706), .C2(n18528), .A(n18056), .B(n13187), .ZN(
        n18689) );
  MUX2_X1 U16349 ( .A(n13188), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18689), .Z(P3_U3284) );
  NOR2_X1 U16350 ( .A1(n16924), .A2(n13189), .ZN(n18041) );
  NOR2_X1 U16351 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18684), .ZN(
        n18686) );
  INV_X1 U16352 ( .A(n18686), .ZN(n13190) );
  OAI221_X1 U16353 ( .B1(n18720), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n17709), .A(n13190), .ZN(n18055) );
  OAI221_X1 U16354 ( .B1(n18658), .B2(n18041), .C1(n18658), .C2(n16403), .A(
        n18131), .ZN(n18053) );
  INV_X1 U16355 ( .A(n18053), .ZN(n18044) );
  NAND2_X1 U16356 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17681) );
  INV_X1 U16357 ( .A(n17681), .ZN(n17667) );
  OAI21_X1 U16358 ( .B1(n17709), .B2(n18720), .A(n18684), .ZN(n18705) );
  NOR2_X1 U16359 ( .A1(n17667), .A2(n18705), .ZN(n18046) );
  AOI21_X1 U16360 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18046), .ZN(n18048) );
  NOR2_X1 U16361 ( .A1(n18044), .A2(n18048), .ZN(n13192) );
  INV_X1 U16362 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16397) );
  NAND2_X1 U16363 ( .A1(n18684), .A2(n18720), .ZN(n16394) );
  NOR2_X1 U16364 ( .A1(n16397), .A2(n16394), .ZN(n18315) );
  NAND2_X1 U16365 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18360), .ZN(n18104) );
  NAND2_X1 U16366 ( .A1(n18104), .A2(n18053), .ZN(n18045) );
  OR2_X1 U16367 ( .A1(n18315), .A2(n18045), .ZN(n13191) );
  MUX2_X1 U16368 ( .A(n13192), .B(n13191), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NAND2_X1 U16369 ( .A1(n13194), .A2(n14071), .ZN(n14289) );
  INV_X1 U16370 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n14746) );
  INV_X1 U16371 ( .A(n14262), .ZN(n14237) );
  AOI22_X1 U16372 ( .A1(n14237), .A2(n19965), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n14235), .ZN(n13195) );
  OAI21_X1 U16373 ( .B1(n14746), .B2(n14239), .A(n13195), .ZN(n13196) );
  AOI21_X1 U16374 ( .B1(n14265), .B2(DATAI_28_), .A(n13196), .ZN(n13197) );
  OAI21_X1 U16375 ( .B1(n14289), .B2(n14268), .A(n13197), .ZN(P1_U2876) );
  NAND2_X1 U16376 ( .A1(n9853), .A2(n13198), .ZN(n13199) );
  NAND2_X1 U16377 ( .A1(n9839), .A2(n13199), .ZN(n14414) );
  INV_X1 U16378 ( .A(n14414), .ZN(n13211) );
  INV_X1 U16379 ( .A(n14292), .ZN(n13209) );
  INV_X1 U16380 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20681) );
  INV_X1 U16381 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20672) );
  NOR2_X1 U16382 ( .A1(n20662), .A2(n13201), .ZN(n15813) );
  NAND2_X1 U16383 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15813), .ZN(n14136) );
  NOR2_X1 U16384 ( .A1(n13202), .A2(n14136), .ZN(n14139) );
  NAND4_X1 U16385 ( .A1(n14139), .A2(P1_REIP_REG_17__SCAN_IN), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n15788) );
  NOR3_X1 U16386 ( .A1(n20672), .A2(n20671), .A3(n15788), .ZN(n15757) );
  INV_X1 U16387 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20677) );
  NAND2_X1 U16388 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15761) );
  NOR2_X1 U16389 ( .A1(n20677), .A2(n15761), .ZN(n15745) );
  NAND3_X1 U16390 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n15757), .A3(n15745), 
        .ZN(n14125) );
  NOR2_X1 U16391 ( .A1(n20681), .A2(n14125), .ZN(n13205) );
  AND2_X1 U16392 ( .A1(n19878), .A2(n13205), .ZN(n14116) );
  NAND2_X1 U16393 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14116), .ZN(n14102) );
  NAND2_X1 U16394 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n13203) );
  NOR2_X1 U16395 ( .A1(n14102), .A2(n13203), .ZN(n13220) );
  AND2_X1 U16396 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n13204) );
  AND3_X1 U16397 ( .A1(n19857), .A2(n13205), .A3(n13204), .ZN(n14087) );
  NAND3_X1 U16398 ( .A1(n14087), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U16399 ( .A1(n19885), .A2(n13206), .ZN(n13218) );
  INV_X1 U16400 ( .A(n13218), .ZN(n14076) );
  OAI21_X1 U16401 ( .B1(n13220), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14076), 
        .ZN(n13208) );
  AOI22_X1 U16402 ( .A1(n19901), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19897), .ZN(n13207) );
  OAI211_X1 U16403 ( .C1(n19906), .C2(n13209), .A(n13208), .B(n13207), .ZN(
        n13210) );
  AOI21_X1 U16404 ( .B1(n13211), .B2(n19880), .A(n13210), .ZN(n13212) );
  OAI21_X1 U16405 ( .B1(n14289), .B2(n19847), .A(n13212), .ZN(P1_U2812) );
  MUX2_X1 U16406 ( .A(n11378), .B(n13213), .S(n14073), .Z(n13216) );
  AOI22_X1 U16407 ( .A1(n13214), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11313), .ZN(n13215) );
  NAND2_X1 U16408 ( .A1(n13988), .A2(n19873), .ZN(n13225) );
  NAND2_X1 U16409 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n13221) );
  NAND2_X1 U16410 ( .A1(n19885), .A2(n13221), .ZN(n13217) );
  NAND2_X1 U16411 ( .A1(n13218), .A2(n13217), .ZN(n14062) );
  OAI22_X1 U16412 ( .A1(n19866), .A2(n14157), .B1(n13219), .B2(n15826), .ZN(
        n13223) );
  NAND2_X1 U16413 ( .A1(n13220), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14075) );
  NOR3_X1 U16414 ( .A1(n14075), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n13221), 
        .ZN(n13222) );
  AOI211_X1 U16415 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14062), .A(n13223), 
        .B(n13222), .ZN(n13224) );
  OAI211_X1 U16416 ( .C1(n14393), .C2(n19892), .A(n13225), .B(n13224), .ZN(
        P1_U2809) );
  OAI211_X1 U16417 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20129), .A(n13226), 
        .B(n20295), .ZN(n13229) );
  NAND2_X1 U16418 ( .A1(n13227), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13228) );
  OAI211_X1 U16419 ( .C1(n13230), .C2(n12799), .A(n13229), .B(n13228), .ZN(
        P1_U3477) );
  INV_X1 U16420 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13902) );
  NAND2_X1 U16421 ( .A1(n13231), .A2(n12037), .ZN(n13255) );
  INV_X1 U16422 ( .A(n13231), .ZN(n13232) );
  NAND2_X1 U16423 ( .A1(n13232), .A2(n12037), .ZN(n13256) );
  INV_X1 U16424 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13233) );
  OAI22_X1 U16425 ( .A1(n13902), .A2(n19358), .B1(n15435), .B2(n13233), .ZN(
        n13238) );
  INV_X1 U16426 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U16427 ( .A1(n15400), .A2(n18958), .ZN(n13245) );
  OR2_X2 U16428 ( .A1(n13247), .A2(n13256), .ZN(n19185) );
  INV_X1 U16429 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13235) );
  OAI22_X1 U16430 ( .A1(n13236), .A2(n19327), .B1(n19185), .B2(n13235), .ZN(
        n13237) );
  NOR2_X1 U16431 ( .A1(n13238), .A2(n13237), .ZN(n13269) );
  INV_X1 U16432 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13912) );
  INV_X1 U16433 ( .A(n13251), .ZN(n13240) );
  INV_X1 U16434 ( .A(n13691), .ZN(n13252) );
  NAND2_X1 U16435 ( .A1(n13240), .A2(n13252), .ZN(n13241) );
  OR2_X2 U16436 ( .A1(n13241), .A2(n15400), .ZN(n15454) );
  OR2_X2 U16437 ( .A1(n13241), .A2(n14698), .ZN(n19578) );
  INV_X1 U16438 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13242) );
  OAI22_X1 U16439 ( .A1(n13912), .A2(n15454), .B1(n19578), .B2(n13242), .ZN(
        n13243) );
  INV_X1 U16440 ( .A(n13243), .ZN(n13268) );
  INV_X1 U16441 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13903) );
  OR2_X1 U16442 ( .A1(n15400), .A2(n12037), .ZN(n13246) );
  OR2_X2 U16444 ( .A1(n13247), .A2(n13255), .ZN(n19246) );
  INV_X1 U16445 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13905) );
  OAI22_X1 U16446 ( .A1(n13903), .A2(n13305), .B1(n19246), .B2(n13905), .ZN(
        n13250) );
  INV_X1 U16447 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13904) );
  OR2_X2 U16448 ( .A1(n13247), .A2(n13246), .ZN(n13363) );
  OAI22_X1 U16449 ( .A1(n13904), .A2(n19212), .B1(n13363), .B2(n13248), .ZN(
        n13249) );
  INV_X1 U16450 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13254) );
  INV_X1 U16451 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13913) );
  INV_X1 U16452 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13911) );
  INV_X1 U16453 ( .A(n13255), .ZN(n13259) );
  INV_X1 U16454 ( .A(n13256), .ZN(n13261) );
  AND2_X1 U16455 ( .A1(n13691), .A2(n13261), .ZN(n13257) );
  INV_X1 U16456 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13258) );
  OAI22_X1 U16457 ( .A1(n13911), .A2(n19613), .B1(n19428), .B2(n13258), .ZN(
        n13266) );
  INV_X1 U16458 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13914) );
  AND2_X1 U16459 ( .A1(n13691), .A2(n13259), .ZN(n13260) );
  NAND2_X2 U16460 ( .A1(n13263), .A2(n13260), .ZN(n19489) );
  INV_X1 U16461 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13264) );
  OAI22_X1 U16462 ( .A1(n13914), .A2(n19489), .B1(n13311), .B2(n13264), .ZN(
        n13265) );
  INV_X1 U16463 ( .A(n19578), .ZN(n19581) );
  INV_X1 U16464 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13763) );
  INV_X1 U16465 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13272) );
  OAI21_X1 U16466 ( .B1(n19613), .B2(n13272), .A(n13271), .ZN(n13273) );
  INV_X1 U16467 ( .A(n13273), .ZN(n13275) );
  INV_X1 U16468 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13773) );
  OAI211_X1 U16469 ( .C1(n19212), .C2(n13763), .A(n13275), .B(n13274), .ZN(
        n13276) );
  AOI21_X1 U16470 ( .B1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n19581), .A(
        n13276), .ZN(n13293) );
  INV_X1 U16471 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13761) );
  INV_X1 U16472 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n21044) );
  OAI22_X1 U16473 ( .A1(n13761), .A2(n19358), .B1(n19462), .B2(n21044), .ZN(
        n13283) );
  INV_X1 U16474 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13281) );
  INV_X1 U16475 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13277) );
  OR2_X1 U16476 ( .A1(n19428), .A2(n13277), .ZN(n13280) );
  INV_X1 U16477 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13278) );
  OAI211_X1 U16478 ( .C1(n19389), .C2(n13281), .A(n13280), .B(n13279), .ZN(
        n13282) );
  NOR2_X1 U16479 ( .A1(n13283), .A2(n13282), .ZN(n13292) );
  INV_X1 U16480 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13772) );
  INV_X1 U16481 ( .A(n19246), .ZN(n19249) );
  NAND2_X1 U16482 ( .A1(n19249), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13285) );
  NAND2_X1 U16484 ( .A1(n19144), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13284) );
  INV_X1 U16485 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13287) );
  INV_X1 U16486 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13286) );
  OAI22_X1 U16487 ( .A1(n13287), .A2(n19327), .B1(n15435), .B2(n13286), .ZN(
        n13290) );
  INV_X1 U16488 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13762) );
  INV_X1 U16489 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13288) );
  OAI22_X1 U16490 ( .A1(n13762), .A2(n13305), .B1(n19185), .B2(n13288), .ZN(
        n13289) );
  NOR2_X1 U16491 ( .A1(n13290), .A2(n13289), .ZN(n13291) );
  NOR2_X1 U16492 ( .A1(n13295), .A2(n13294), .ZN(n13519) );
  OR2_X1 U16493 ( .A1(n13519), .A2(n13296), .ZN(n13297) );
  INV_X1 U16494 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13963) );
  INV_X1 U16495 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13792) );
  OAI22_X1 U16496 ( .A1(n13963), .A2(n19358), .B1(n15435), .B2(n13792), .ZN(
        n13302) );
  INV_X1 U16497 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13300) );
  INV_X1 U16498 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13299) );
  OAI22_X1 U16499 ( .A1(n13300), .A2(n19327), .B1(n19185), .B2(n13299), .ZN(
        n13301) );
  NOR2_X1 U16500 ( .A1(n13302), .A2(n13301), .ZN(n13319) );
  INV_X1 U16501 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13973) );
  INV_X1 U16502 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13303) );
  OAI22_X1 U16503 ( .A1(n13973), .A2(n15454), .B1(n19578), .B2(n13303), .ZN(
        n13304) );
  INV_X1 U16504 ( .A(n13304), .ZN(n13318) );
  INV_X1 U16505 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13964) );
  INV_X1 U16506 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13966) );
  OAI22_X1 U16507 ( .A1(n13964), .A2(n13305), .B1(n19246), .B2(n13966), .ZN(
        n13308) );
  INV_X1 U16508 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13965) );
  OAI22_X1 U16509 ( .A1(n13965), .A2(n19212), .B1(n13363), .B2(n13306), .ZN(
        n13307) );
  NOR2_X1 U16510 ( .A1(n13308), .A2(n13307), .ZN(n13317) );
  INV_X1 U16511 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13974) );
  INV_X1 U16512 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13309) );
  OAI22_X1 U16513 ( .A1(n13974), .A2(n19462), .B1(n19389), .B2(n13309), .ZN(
        n13315) );
  INV_X1 U16514 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13972) );
  INV_X1 U16515 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13310) );
  OAI22_X1 U16516 ( .A1(n13972), .A2(n19613), .B1(n19428), .B2(n13310), .ZN(
        n13314) );
  INV_X1 U16517 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13975) );
  INV_X1 U16518 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13312) );
  OAI22_X1 U16519 ( .A1(n13975), .A2(n19489), .B1(n13311), .B2(n13312), .ZN(
        n13313) );
  NOR3_X1 U16520 ( .A1(n13315), .A2(n13314), .A3(n13313), .ZN(n13316) );
  NAND4_X1 U16521 ( .A1(n13319), .A2(n13318), .A3(n13317), .A4(n13316), .ZN(
        n13322) );
  NAND2_X1 U16522 ( .A1(n13320), .A2(n10055), .ZN(n13321) );
  INV_X1 U16523 ( .A(n13352), .ZN(n13323) );
  NAND2_X1 U16524 ( .A1(n13535), .A2(n13543), .ZN(n13328) );
  INV_X1 U16525 ( .A(n13380), .ZN(n13327) );
  NAND2_X1 U16526 ( .A1(n13325), .A2(n13324), .ZN(n13326) );
  NAND2_X1 U16527 ( .A1(n13327), .A2(n13326), .ZN(n18908) );
  NAND2_X1 U16528 ( .A1(n13328), .A2(n18908), .ZN(n13349) );
  INV_X1 U16529 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15384) );
  XNOR2_X1 U16530 ( .A(n13349), .B(n15384), .ZN(n15376) );
  NAND2_X1 U16531 ( .A1(n15038), .A2(n13543), .ZN(n13331) );
  NAND2_X1 U16532 ( .A1(n13331), .A2(n13330), .ZN(n15031) );
  INV_X1 U16533 ( .A(n14693), .ZN(n13332) );
  NOR2_X1 U16534 ( .A1(n13333), .A2(n13332), .ZN(n13335) );
  NOR2_X1 U16535 ( .A1(n13335), .A2(n13334), .ZN(n13338) );
  XNOR2_X1 U16536 ( .A(n13338), .B(n13336), .ZN(n13650) );
  NAND2_X1 U16537 ( .A1(n13650), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13651) );
  INV_X1 U16538 ( .A(n13336), .ZN(n13337) );
  OR2_X1 U16539 ( .A1(n13338), .A2(n13337), .ZN(n13339) );
  INV_X1 U16540 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13631) );
  XNOR2_X1 U16541 ( .A(n13341), .B(n13340), .ZN(n19108) );
  INV_X1 U16542 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19123) );
  AND2_X1 U16543 ( .A1(n19108), .A2(n19123), .ZN(n13343) );
  AOI21_X1 U16544 ( .B1(n19107), .B2(n13631), .A(n13343), .ZN(n13342) );
  NAND2_X1 U16545 ( .A1(n15031), .A2(n13342), .ZN(n13348) );
  INV_X1 U16546 ( .A(n19107), .ZN(n13346) );
  INV_X1 U16547 ( .A(n13343), .ZN(n13344) );
  AND2_X1 U16548 ( .A1(n13344), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13345) );
  INV_X1 U16549 ( .A(n19108), .ZN(n18929) );
  AOI22_X1 U16550 ( .A1(n13346), .A2(n13345), .B1(n18929), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U16551 ( .A1(n13348), .A2(n13347), .ZN(n15375) );
  NAND2_X1 U16552 ( .A1(n15376), .A2(n15375), .ZN(n13351) );
  NAND2_X1 U16553 ( .A1(n13349), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13350) );
  NAND2_X1 U16554 ( .A1(n13351), .A2(n13350), .ZN(n15360) );
  INV_X1 U16555 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13993) );
  INV_X1 U16556 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13994) );
  OAI22_X1 U16557 ( .A1(n13993), .A2(n19358), .B1(n13305), .B2(n13994), .ZN(
        n13356) );
  INV_X1 U16558 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13997) );
  INV_X1 U16559 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13354) );
  OAI22_X1 U16560 ( .A1(n13997), .A2(n19246), .B1(n15435), .B2(n13354), .ZN(
        n13355) );
  NOR2_X1 U16561 ( .A1(n13356), .A2(n13355), .ZN(n13375) );
  INV_X1 U16562 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13358) );
  INV_X1 U16563 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13357) );
  OAI22_X1 U16564 ( .A1(n13358), .A2(n19578), .B1(n15454), .B2(n13357), .ZN(
        n13359) );
  INV_X1 U16565 ( .A(n13359), .ZN(n13374) );
  INV_X1 U16566 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13361) );
  INV_X1 U16567 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13360) );
  OAI22_X1 U16568 ( .A1(n13361), .A2(n19327), .B1(n19185), .B2(n13360), .ZN(
        n13365) );
  INV_X1 U16569 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13996) );
  INV_X1 U16570 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13362) );
  OAI22_X1 U16571 ( .A1(n13996), .A2(n19212), .B1(n13363), .B2(n13362), .ZN(
        n13364) );
  NOR2_X1 U16572 ( .A1(n13365), .A2(n13364), .ZN(n13373) );
  INV_X1 U16573 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14005) );
  INV_X1 U16574 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13366) );
  OAI22_X1 U16575 ( .A1(n14005), .A2(n19462), .B1(n19389), .B2(n13366), .ZN(
        n13371) );
  INV_X1 U16576 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14003) );
  INV_X1 U16577 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14007) );
  OAI22_X1 U16578 ( .A1(n14003), .A2(n19613), .B1(n19489), .B2(n14007), .ZN(
        n13370) );
  INV_X1 U16579 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13368) );
  INV_X1 U16580 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13367) );
  OAI22_X1 U16581 ( .A1(n13368), .A2(n19428), .B1(n13311), .B2(n13367), .ZN(
        n13369) );
  NOR3_X1 U16582 ( .A1(n13371), .A2(n13370), .A3(n13369), .ZN(n13372) );
  NAND4_X1 U16583 ( .A1(n13375), .A2(n13374), .A3(n13373), .A4(n13372), .ZN(
        n13378) );
  NAND2_X1 U16584 ( .A1(n13376), .A2(n10055), .ZN(n13377) );
  NOR2_X1 U16585 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  OR2_X1 U16586 ( .A1(n13386), .A2(n13381), .ZN(n18895) );
  INV_X1 U16587 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15366) );
  XNOR2_X1 U16588 ( .A(n13382), .B(n15366), .ZN(n15362) );
  NAND2_X1 U16589 ( .A1(n13382), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13383) );
  INV_X1 U16590 ( .A(n13384), .ZN(n13385) );
  XNOR2_X1 U16591 ( .A(n13386), .B(n13385), .ZN(n13393) );
  NOR2_X1 U16592 ( .A1(n13387), .A2(n13543), .ZN(n13391) );
  NAND2_X1 U16593 ( .A1(n13391), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15342) );
  AND2_X1 U16594 ( .A1(n13502), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13388) );
  MUX2_X1 U16595 ( .A(n11979), .B(n13388), .S(n13389), .Z(n13390) );
  NOR2_X1 U16596 ( .A1(n13390), .A2(n13396), .ZN(n18868) );
  NAND2_X1 U16597 ( .A1(n18868), .A2(n13510), .ZN(n13401) );
  INV_X1 U16598 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21038) );
  NAND2_X1 U16599 ( .A1(n13401), .A2(n21038), .ZN(n15329) );
  INV_X1 U16600 ( .A(n13391), .ZN(n13392) );
  INV_X1 U16601 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15354) );
  NAND2_X1 U16602 ( .A1(n13392), .A2(n15354), .ZN(n15341) );
  INV_X1 U16603 ( .A(n13393), .ZN(n18887) );
  INV_X1 U16604 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13394) );
  NAND2_X1 U16605 ( .A1(n18887), .A2(n13394), .ZN(n15021) );
  AND2_X1 U16606 ( .A1(n15341), .A2(n15021), .ZN(n15306) );
  NOR2_X1 U16607 ( .A1(n13396), .A2(n12743), .ZN(n13397) );
  NAND2_X1 U16608 ( .A1(n13502), .A2(n13397), .ZN(n13398) );
  AND2_X1 U16609 ( .A1(n13485), .A2(n13398), .ZN(n13399) );
  NAND2_X1 U16610 ( .A1(n13404), .A2(n13399), .ZN(n18862) );
  OR2_X1 U16611 ( .A1(n18862), .A2(n13543), .ZN(n13400) );
  INV_X1 U16612 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U16613 ( .A1(n13400), .A2(n15312), .ZN(n15305) );
  AND3_X1 U16614 ( .A1(n15329), .A2(n15306), .A3(n15305), .ZN(n13403) );
  OR2_X1 U16615 ( .A1(n13401), .A2(n21038), .ZN(n15330) );
  OR3_X1 U16616 ( .A1(n18862), .A2(n13543), .A3(n15312), .ZN(n15304) );
  NAND2_X1 U16617 ( .A1(n15330), .A2(n15304), .ZN(n13402) );
  AND3_X1 U16618 ( .A1(n13502), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n13404), .ZN(
        n13405) );
  OR2_X1 U16619 ( .A1(n13406), .A2(n13405), .ZN(n14685) );
  NOR2_X1 U16620 ( .A1(n14685), .A2(n13543), .ZN(n13435) );
  NAND2_X1 U16621 ( .A1(n13435), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15289) );
  NAND2_X1 U16622 ( .A1(n13502), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13407) );
  INV_X1 U16623 ( .A(n13407), .ZN(n13408) );
  NAND2_X1 U16624 ( .A1(n13408), .A2(n9842), .ZN(n13409) );
  NAND2_X1 U16625 ( .A1(n13424), .A2(n13409), .ZN(n18846) );
  XNOR2_X1 U16626 ( .A(n13439), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15269) );
  AND2_X1 U16627 ( .A1(n13502), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13423) );
  NAND2_X1 U16628 ( .A1(n18811), .A2(n18824), .ZN(n13411) );
  AND2_X1 U16629 ( .A1(n13502), .A2(n13411), .ZN(n13412) );
  NAND2_X1 U16630 ( .A1(n13502), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13416) );
  NAND2_X1 U16631 ( .A1(n13502), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13428) );
  NAND2_X1 U16632 ( .A1(n13502), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n13448) );
  AND2_X1 U16633 ( .A1(n13502), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13445) );
  NAND2_X1 U16634 ( .A1(n13502), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13413) );
  XNOR2_X1 U16635 ( .A(n13441), .B(n13413), .ZN(n18754) );
  NAND2_X1 U16636 ( .A1(n18754), .A2(n13510), .ZN(n13414) );
  INV_X1 U16637 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15172) );
  NAND2_X1 U16638 ( .A1(n13414), .A2(n15172), .ZN(n14948) );
  MUX2_X1 U16639 ( .A(n13416), .B(P2_EBX_REG_16__SCAN_IN), .S(n13415), .Z(
        n13417) );
  NAND2_X1 U16640 ( .A1(n13417), .A2(n13485), .ZN(n14674) );
  INV_X1 U16641 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15227) );
  OAI21_X1 U16642 ( .B1(n14674), .B2(n13543), .A(n15227), .ZN(n13420) );
  INV_X1 U16643 ( .A(n14674), .ZN(n13419) );
  AND2_X1 U16644 ( .A1(n13510), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13418) );
  NAND2_X1 U16645 ( .A1(n13419), .A2(n13418), .ZN(n14929) );
  NAND2_X1 U16646 ( .A1(n13502), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13421) );
  MUX2_X1 U16647 ( .A(n13502), .B(n13421), .S(n13426), .Z(n13422) );
  NAND2_X1 U16648 ( .A1(n13410), .A2(n18824), .ZN(n13432) );
  NAND2_X1 U16649 ( .A1(n13422), .A2(n13432), .ZN(n13457) );
  INV_X1 U16650 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15249) );
  OAI21_X1 U16651 ( .B1(n13457), .B2(n13543), .A(n15249), .ZN(n15244) );
  NAND2_X1 U16652 ( .A1(n13424), .A2(n13423), .ZN(n13425) );
  NAND2_X1 U16653 ( .A1(n13426), .A2(n13425), .ZN(n18837) );
  INV_X1 U16654 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13427) );
  OAI21_X1 U16655 ( .B1(n18837), .B2(n13543), .A(n13427), .ZN(n16131) );
  AND2_X1 U16656 ( .A1(n15244), .A2(n16131), .ZN(n14926) );
  NOR2_X1 U16657 ( .A1(n13429), .A2(n13428), .ZN(n13430) );
  NAND2_X1 U16658 ( .A1(n9843), .A2(n13510), .ZN(n13455) );
  INV_X1 U16659 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13431) );
  NAND2_X1 U16660 ( .A1(n13455), .A2(n13431), .ZN(n14987) );
  INV_X1 U16661 ( .A(n13415), .ZN(n13434) );
  NAND3_X1 U16662 ( .A1(n13432), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n13502), 
        .ZN(n13433) );
  NAND2_X1 U16663 ( .A1(n13434), .A2(n13433), .ZN(n18813) );
  INV_X1 U16664 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15209) );
  NAND2_X1 U16665 ( .A1(n13459), .A2(n15209), .ZN(n15008) );
  INV_X1 U16666 ( .A(n13435), .ZN(n13437) );
  INV_X1 U16667 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13436) );
  NAND2_X1 U16668 ( .A1(n13437), .A2(n13436), .ZN(n15288) );
  INV_X1 U16669 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13438) );
  NAND2_X1 U16670 ( .A1(n13439), .A2(n13438), .ZN(n14925) );
  AND4_X1 U16671 ( .A1(n14987), .A2(n15008), .A3(n15288), .A4(n14925), .ZN(
        n13440) );
  NAND4_X1 U16672 ( .A1(n14948), .A2(n14997), .A3(n14926), .A4(n13440), .ZN(
        n13452) );
  INV_X1 U16673 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14653) );
  NAND2_X1 U16674 ( .A1(n13443), .A2(n14653), .ZN(n13469) );
  NAND2_X1 U16675 ( .A1(n13469), .A2(n13485), .ZN(n13467) );
  NAND2_X1 U16676 ( .A1(n13502), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n13442) );
  NOR2_X1 U16677 ( .A1(n13443), .A2(n13442), .ZN(n13444) );
  INV_X1 U16678 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15111) );
  INV_X1 U16679 ( .A(n13445), .ZN(n13446) );
  XNOR2_X1 U16680 ( .A(n13447), .B(n13446), .ZN(n18772) );
  NAND2_X1 U16681 ( .A1(n18772), .A2(n13510), .ZN(n13463) );
  INV_X1 U16682 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15183) );
  NAND2_X1 U16683 ( .A1(n13463), .A2(n15183), .ZN(n14958) );
  XNOR2_X1 U16684 ( .A(n13449), .B(n10072), .ZN(n18785) );
  NAND2_X1 U16685 ( .A1(n18785), .A2(n13510), .ZN(n13450) );
  INV_X1 U16686 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14975) );
  NAND2_X1 U16687 ( .A1(n13450), .A2(n14975), .ZN(n14960) );
  AND2_X1 U16688 ( .A1(n14958), .A2(n14960), .ZN(n14946) );
  NAND2_X1 U16689 ( .A1(n14933), .A2(n14946), .ZN(n13451) );
  NOR2_X1 U16690 ( .A1(n13453), .A2(n15111), .ZN(n14935) );
  AND2_X1 U16691 ( .A1(n13510), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13454) );
  INV_X1 U16692 ( .A(n13455), .ZN(n13456) );
  NAND2_X1 U16693 ( .A1(n13456), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14930) );
  INV_X1 U16694 ( .A(n13457), .ZN(n18826) );
  AND2_X1 U16695 ( .A1(n13510), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13458) );
  NAND2_X1 U16696 ( .A1(n18826), .A2(n13458), .ZN(n15243) );
  INV_X1 U16697 ( .A(n13459), .ZN(n13460) );
  NAND2_X1 U16698 ( .A1(n13460), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14928) );
  INV_X1 U16699 ( .A(n18837), .ZN(n13462) );
  AND2_X1 U16700 ( .A1(n13510), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13461) );
  NAND2_X1 U16701 ( .A1(n13462), .A2(n13461), .ZN(n16130) );
  AND4_X1 U16702 ( .A1(n14930), .A2(n15243), .A3(n14928), .A4(n16130), .ZN(
        n13465) );
  AND2_X1 U16703 ( .A1(n13510), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13464) );
  NAND2_X1 U16704 ( .A1(n18785), .A2(n13464), .ZN(n14931) );
  NAND2_X1 U16705 ( .A1(n13502), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n13466) );
  INV_X1 U16706 ( .A(n13466), .ZN(n13470) );
  INV_X1 U16707 ( .A(n13472), .ZN(n13468) );
  AOI21_X1 U16708 ( .B1(n13470), .B2(n13469), .A(n13468), .ZN(n14639) );
  AOI21_X1 U16709 ( .B1(n14639), .B2(n13510), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14912) );
  NAND3_X1 U16710 ( .A1(n14639), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n13510), .ZN(n14913) );
  OAI21_X1 U16711 ( .B1(n14916), .B2(n14912), .A(n14913), .ZN(n14904) );
  AND2_X1 U16712 ( .A1(n13502), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U16713 ( .A1(n13472), .A2(n13471), .ZN(n13473) );
  NAND2_X1 U16714 ( .A1(n14594), .A2(n13473), .ZN(n14627) );
  OR2_X1 U16715 ( .A1(n14627), .A2(n13543), .ZN(n13474) );
  XNOR2_X1 U16716 ( .A(n13474), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14905) );
  INV_X1 U16717 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13573) );
  NOR3_X1 U16718 ( .A1(n14627), .A2(n13543), .A3(n13573), .ZN(n13475) );
  INV_X1 U16719 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15118) );
  NAND2_X1 U16720 ( .A1(n13485), .A2(n13510), .ZN(n14893) );
  INV_X1 U16721 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16085) );
  NOR2_X1 U16722 ( .A1(n13479), .A2(n16085), .ZN(n13476) );
  NAND2_X1 U16723 ( .A1(n13502), .A2(n13476), .ZN(n13477) );
  NAND2_X1 U16724 ( .A1(n13485), .A2(n13477), .ZN(n13478) );
  AOI21_X1 U16725 ( .B1(n13479), .B2(n16085), .A(n13478), .ZN(n16089) );
  AND2_X1 U16726 ( .A1(n16089), .A2(n13510), .ZN(n13496) );
  NOR2_X1 U16727 ( .A1(n13496), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14882) );
  NAND2_X1 U16728 ( .A1(n13479), .A2(n16085), .ZN(n13480) );
  AND2_X1 U16729 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n13480), .ZN(n13481) );
  AOI21_X1 U16730 ( .B1(n13502), .B2(n13481), .A(n13484), .ZN(n13482) );
  NAND2_X1 U16731 ( .A1(n13485), .A2(n13482), .ZN(n16074) );
  NOR2_X1 U16732 ( .A1(n16074), .A2(n13543), .ZN(n13483) );
  NAND2_X1 U16733 ( .A1(n13483), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13497) );
  OAI21_X1 U16734 ( .B1(n13483), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13497), .ZN(n14876) );
  INV_X1 U16735 ( .A(n13484), .ZN(n13487) );
  NAND2_X1 U16736 ( .A1(n13485), .A2(n13487), .ZN(n13506) );
  NAND2_X1 U16737 ( .A1(n13502), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n13486) );
  INV_X1 U16738 ( .A(n13486), .ZN(n13488) );
  NAND2_X1 U16739 ( .A1(n13488), .A2(n13487), .ZN(n13489) );
  NAND2_X1 U16740 ( .A1(n13490), .A2(n13489), .ZN(n14583) );
  NOR2_X1 U16741 ( .A1(n14583), .A2(n13543), .ZN(n14858) );
  AND2_X1 U16742 ( .A1(n13502), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13491) );
  AOI21_X1 U16743 ( .B1(n13491), .B2(n13490), .A(n13501), .ZN(n14576) );
  NAND2_X1 U16744 ( .A1(n14576), .A2(n13510), .ZN(n14859) );
  INV_X1 U16745 ( .A(n14859), .ZN(n13492) );
  OAI21_X1 U16746 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n13492), .ZN(n13493) );
  INV_X1 U16747 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15069) );
  NAND2_X1 U16748 ( .A1(n14859), .A2(n15069), .ZN(n13494) );
  NAND2_X1 U16749 ( .A1(n13495), .A2(n13494), .ZN(n13498) );
  NAND2_X1 U16750 ( .A1(n13496), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14883) );
  NAND2_X1 U16751 ( .A1(n14883), .A2(n13497), .ZN(n14855) );
  NAND2_X1 U16752 ( .A1(n13498), .A2(n10051), .ZN(n14847) );
  NAND2_X1 U16753 ( .A1(n13502), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13500) );
  INV_X1 U16754 ( .A(n13501), .ZN(n13499) );
  XOR2_X1 U16755 ( .A(n13500), .B(n13499), .Z(n13505) );
  INV_X1 U16756 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15060) );
  OAI21_X1 U16757 ( .B1(n13505), .B2(n13543), .A(n15060), .ZN(n14849) );
  NAND2_X1 U16758 ( .A1(n14847), .A2(n14849), .ZN(n14835) );
  NAND2_X1 U16759 ( .A1(n13501), .A2(n13500), .ZN(n13507) );
  NAND2_X1 U16760 ( .A1(n13502), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13503) );
  XNOR2_X1 U16761 ( .A(n13507), .B(n13503), .ZN(n13504) );
  AOI21_X1 U16762 ( .B1(n13504), .B2(n13510), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14838) );
  INV_X1 U16763 ( .A(n13504), .ZN(n16045) );
  INV_X1 U16764 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13643) );
  INV_X1 U16765 ( .A(n13505), .ZN(n16063) );
  NAND3_X1 U16766 ( .A1(n16063), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n13510), .ZN(n14848) );
  INV_X1 U16767 ( .A(n13506), .ZN(n13509) );
  NOR2_X1 U16768 ( .A1(n13507), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13508) );
  MUX2_X1 U16769 ( .A(n13509), .B(n13508), .S(n13502), .Z(n14564) );
  NAND2_X1 U16770 ( .A1(n14564), .A2(n13510), .ZN(n13511) );
  XNOR2_X1 U16771 ( .A(n13511), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13512) );
  XNOR2_X1 U16772 ( .A(n13513), .B(n13512), .ZN(n14834) );
  INV_X1 U16773 ( .A(n13514), .ZN(n13516) );
  NAND2_X1 U16774 ( .A1(n13516), .A2(n13515), .ZN(n13518) );
  NAND2_X1 U16775 ( .A1(n13518), .A2(n13517), .ZN(n13521) );
  XOR2_X1 U16776 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13521), .Z(
        n13660) );
  XOR2_X1 U16777 ( .A(n13520), .B(n13519), .Z(n13659) );
  NAND2_X1 U16778 ( .A1(n13660), .A2(n13659), .ZN(n13658) );
  NAND2_X1 U16779 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13521), .ZN(
        n13522) );
  NAND2_X1 U16780 ( .A1(n13658), .A2(n13522), .ZN(n13523) );
  XNOR2_X1 U16781 ( .A(n13523), .B(n13631), .ZN(n15037) );
  NAND2_X1 U16782 ( .A1(n13523), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13524) );
  NAND2_X1 U16783 ( .A1(n13525), .A2(n13524), .ZN(n13530) );
  NAND2_X1 U16784 ( .A1(n13527), .A2(n13526), .ZN(n13529) );
  XNOR2_X1 U16785 ( .A(n13529), .B(n13528), .ZN(n13531) );
  NAND2_X1 U16786 ( .A1(n13530), .A2(n13531), .ZN(n19111) );
  NAND2_X1 U16787 ( .A1(n19111), .A2(n19123), .ZN(n13534) );
  INV_X1 U16788 ( .A(n13530), .ZN(n13533) );
  INV_X1 U16789 ( .A(n13531), .ZN(n13532) );
  NAND2_X1 U16790 ( .A1(n13533), .A2(n13532), .ZN(n19112) );
  INV_X1 U16791 ( .A(n13535), .ZN(n13536) );
  NAND2_X1 U16792 ( .A1(n13536), .A2(n15384), .ZN(n15386) );
  NAND2_X1 U16793 ( .A1(n13535), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15387) );
  NAND2_X1 U16794 ( .A1(n9863), .A2(n15387), .ZN(n13537) );
  INV_X1 U16795 ( .A(n15387), .ZN(n15390) );
  NAND2_X1 U16796 ( .A1(n15390), .A2(n10037), .ZN(n13539) );
  NAND2_X1 U16797 ( .A1(n15371), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15370) );
  NAND2_X1 U16798 ( .A1(n15391), .A2(n15387), .ZN(n13540) );
  NAND2_X1 U16799 ( .A1(n13540), .A2(n9863), .ZN(n13541) );
  NAND2_X2 U16800 ( .A1(n15370), .A2(n13541), .ZN(n15020) );
  NAND2_X1 U16801 ( .A1(n13542), .A2(n13543), .ZN(n13544) );
  NAND2_X1 U16802 ( .A1(n13545), .A2(n13544), .ZN(n15018) );
  INV_X1 U16803 ( .A(n13545), .ZN(n13546) );
  NAND2_X1 U16804 ( .A1(n13546), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13547) );
  NAND2_X2 U16805 ( .A1(n15349), .A2(n13547), .ZN(n14992) );
  NAND2_X1 U16806 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15254) );
  NAND2_X1 U16807 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15293) );
  NOR2_X1 U16808 ( .A1(n15254), .A2(n15293), .ZN(n13548) );
  AND3_X1 U16809 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n13548), .ZN(n15203) );
  AND3_X1 U16810 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13549) );
  NAND2_X1 U16811 ( .A1(n15203), .A2(n13549), .ZN(n15195) );
  INV_X1 U16812 ( .A(n15195), .ZN(n13550) );
  AND2_X1 U16814 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15127) );
  NAND2_X1 U16815 ( .A1(n15127), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13628) );
  AND2_X1 U16816 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15090) );
  AOI22_X1 U16817 ( .A1(n13595), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n13553) );
  NAND2_X1 U16818 ( .A1(n9803), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13552) );
  OAI211_X1 U16819 ( .C1(n13574), .C2(n15227), .A(n13553), .B(n13552), .ZN(
        n14664) );
  INV_X1 U16820 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n18794) );
  NAND2_X1 U16821 ( .A1(n13595), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n13555) );
  NAND2_X1 U16822 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13554) );
  OAI211_X1 U16823 ( .C1(n13598), .C2(n18794), .A(n13555), .B(n13554), .ZN(
        n13556) );
  AOI21_X1 U16824 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n13556), .ZN(n14728) );
  OR2_X2 U16825 ( .A1(n14663), .A2(n14728), .ZN(n14977) );
  INV_X1 U16826 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18783) );
  INV_X1 U16827 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19717) );
  OR2_X1 U16828 ( .A1(n13585), .A2(n19717), .ZN(n13558) );
  NAND2_X1 U16829 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13557) );
  OAI211_X1 U16830 ( .C1(n13598), .C2(n18783), .A(n13558), .B(n13557), .ZN(
        n13559) );
  AOI21_X1 U16831 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n13559), .ZN(n14976) );
  AOI22_X1 U16832 ( .A1(n13595), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n13561) );
  NAND2_X1 U16833 ( .A1(n9803), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n13560) );
  OAI211_X1 U16834 ( .C1(n13574), .C2(n15183), .A(n13561), .B(n13560), .ZN(
        n13757) );
  AOI22_X1 U16835 ( .A1(n13595), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n13563) );
  NAND2_X1 U16836 ( .A1(n9803), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n13562) );
  OAI211_X1 U16837 ( .C1(n13574), .C2(n15172), .A(n13563), .B(n13562), .ZN(
        n14951) );
  INV_X1 U16838 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19723) );
  OR2_X1 U16839 ( .A1(n13585), .A2(n19723), .ZN(n13565) );
  NAND2_X1 U16840 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13564) );
  OAI211_X1 U16841 ( .C1(n13598), .C2(n14653), .A(n13565), .B(n13564), .ZN(
        n13566) );
  AOI21_X1 U16842 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n13566), .ZN(n14645) );
  INV_X1 U16843 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n13569) );
  INV_X1 U16844 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19725) );
  OR2_X1 U16845 ( .A1(n13585), .A2(n19725), .ZN(n13568) );
  NAND2_X1 U16846 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13567) );
  OAI211_X1 U16847 ( .C1(n13598), .C2(n13569), .A(n13568), .B(n13567), .ZN(
        n13570) );
  AOI21_X1 U16848 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n13570), .ZN(n14628) );
  AOI22_X1 U16849 ( .A1(n13595), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n13572) );
  NAND2_X1 U16850 ( .A1(n9803), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n13571) );
  OAI211_X1 U16851 ( .C1(n13574), .C2(n13573), .A(n13572), .B(n13571), .ZN(
        n14615) );
  AOI22_X1 U16853 ( .A1(n13595), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n13577) );
  NAND2_X1 U16854 ( .A1(n9803), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n13576) );
  OAI211_X1 U16855 ( .C1(n13574), .C2(n15118), .A(n13577), .B(n13576), .ZN(
        n13861) );
  NAND2_X1 U16856 ( .A1(n14617), .A2(n13861), .ZN(n13860) );
  INV_X1 U16857 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19731) );
  OR2_X1 U16858 ( .A1(n13585), .A2(n19731), .ZN(n13579) );
  NAND2_X1 U16859 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13578) );
  OAI211_X1 U16860 ( .C1(n13598), .C2(n16085), .A(n13579), .B(n13578), .ZN(
        n13580) );
  AOI21_X1 U16861 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n13580), .ZN(n13894) );
  OR2_X2 U16862 ( .A1(n13860), .A2(n13894), .ZN(n14713) );
  INV_X1 U16863 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n13583) );
  INV_X1 U16864 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19733) );
  OR2_X1 U16865 ( .A1(n13585), .A2(n19733), .ZN(n13582) );
  NAND2_X1 U16866 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13581) );
  OAI211_X1 U16867 ( .C1(n13598), .C2(n13583), .A(n13582), .B(n13581), .ZN(
        n13584) );
  AOI21_X1 U16868 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n13584), .ZN(n14714) );
  OR2_X2 U16869 ( .A1(n14713), .A2(n14714), .ZN(n14715) );
  INV_X1 U16870 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n14589) );
  INV_X1 U16871 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19736) );
  OR2_X1 U16872 ( .A1(n13585), .A2(n19736), .ZN(n13587) );
  NAND2_X1 U16873 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13586) );
  OAI211_X1 U16874 ( .C1(n13598), .C2(n14589), .A(n13587), .B(n13586), .ZN(
        n13588) );
  AOI21_X1 U16875 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n13588), .ZN(n13957) );
  NOR2_X2 U16876 ( .A1(n14715), .A2(n13957), .ZN(n13985) );
  AOI22_X1 U16877 ( .A1(n13595), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n13590) );
  NAND2_X1 U16878 ( .A1(n9803), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n13589) );
  OAI211_X1 U16879 ( .C1(n13574), .C2(n15069), .A(n13590), .B(n13589), .ZN(
        n13984) );
  AND2_X2 U16880 ( .A1(n13985), .A2(n13984), .ZN(n14705) );
  AOI22_X1 U16881 ( .A1(n13595), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n13592) );
  NAND2_X1 U16882 ( .A1(n9803), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13591) );
  OAI211_X1 U16883 ( .C1(n13574), .C2(n15060), .A(n13592), .B(n13591), .ZN(
        n14704) );
  AND2_X2 U16884 ( .A1(n14705), .A2(n14704), .ZN(n14707) );
  AOI22_X1 U16885 ( .A1(n13595), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n13594) );
  NAND2_X1 U16886 ( .A1(n9803), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13593) );
  OAI211_X1 U16887 ( .C1(n13574), .C2(n13643), .A(n13594), .B(n13593), .ZN(
        n14055) );
  NAND2_X1 U16888 ( .A1(n14707), .A2(n14055), .ZN(n13602) );
  NAND2_X1 U16889 ( .A1(n13595), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n13597) );
  NAND2_X1 U16890 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13596) );
  OAI211_X1 U16891 ( .C1(n13598), .C2(n16093), .A(n13597), .B(n13596), .ZN(
        n13599) );
  AOI21_X1 U16892 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13599), .ZN(n13601) );
  XNOR2_X2 U16893 ( .A(n13602), .B(n13601), .ZN(n16094) );
  INV_X1 U16894 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n15012) );
  NAND2_X1 U16895 ( .A1(n13604), .A2(n13603), .ZN(n13606) );
  AOI22_X1 U16896 ( .A1(n13625), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13605) );
  OAI211_X1 U16897 ( .C1(n12150), .C2(n15012), .A(n13606), .B(n13605), .ZN(
        n15230) );
  INV_X1 U16898 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19713) );
  AOI22_X1 U16899 ( .A1(n13625), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13607) );
  OAI21_X1 U16900 ( .B1(n12150), .B2(n19713), .A(n13607), .ZN(n14666) );
  INV_X1 U16901 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19715) );
  AOI22_X1 U16902 ( .A1(n13625), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13608) );
  OAI21_X1 U16903 ( .B1(n12150), .B2(n19715), .A(n13608), .ZN(n14818) );
  AOI22_X1 U16904 ( .A1(n13625), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13609) );
  OAI21_X1 U16905 ( .B1(n12150), .B2(n19717), .A(n13609), .ZN(n15189) );
  INV_X1 U16906 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19719) );
  AOI22_X1 U16907 ( .A1(n13625), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13610) );
  OAI21_X1 U16908 ( .B1(n12150), .B2(n19719), .A(n13610), .ZN(n14808) );
  INV_X1 U16909 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19721) );
  AOI22_X1 U16910 ( .A1(n13625), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13611) );
  OAI21_X1 U16911 ( .B1(n12150), .B2(n19721), .A(n13611), .ZN(n15163) );
  AOI22_X1 U16912 ( .A1(n13625), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13612) );
  OAI21_X1 U16913 ( .B1(n12150), .B2(n19723), .A(n13612), .ZN(n14650) );
  AOI22_X1 U16914 ( .A1(n13625), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13613) );
  OAI21_X1 U16915 ( .B1(n13621), .B2(n19725), .A(n13613), .ZN(n14631) );
  INV_X1 U16916 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19727) );
  AOI22_X1 U16917 ( .A1(n13625), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13614) );
  OAI21_X1 U16918 ( .B1(n12150), .B2(n19727), .A(n13614), .ZN(n14619) );
  INV_X1 U16919 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19729) );
  AOI22_X1 U16920 ( .A1(n13625), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13615) );
  OAI21_X1 U16921 ( .B1(n13621), .B2(n19729), .A(n13615), .ZN(n14602) );
  AOI22_X1 U16922 ( .A1(n13625), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13616) );
  OAI21_X1 U16923 ( .B1(n13621), .B2(n19731), .A(n13616), .ZN(n14768) );
  AOI22_X1 U16924 ( .A1(n13625), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13617) );
  OAI21_X1 U16925 ( .B1(n13621), .B2(n19733), .A(n13617), .ZN(n14757) );
  AOI22_X1 U16926 ( .A1(n13625), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13618) );
  OAI21_X1 U16927 ( .B1(n13621), .B2(n19736), .A(n13618), .ZN(n14584) );
  INV_X1 U16928 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19737) );
  AOI22_X1 U16929 ( .A1(n13625), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13619) );
  OAI21_X1 U16930 ( .B1(n13621), .B2(n19737), .A(n13619), .ZN(n14570) );
  INV_X1 U16931 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19739) );
  AOI22_X1 U16932 ( .A1(n13625), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13620) );
  OAI21_X1 U16933 ( .B1(n13621), .B2(n19739), .A(n13620), .ZN(n14735) );
  NAND2_X1 U16934 ( .A1(n14736), .A2(n14735), .ZN(n14734) );
  NAND2_X1 U16935 ( .A1(n13626), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13623) );
  AOI22_X1 U16936 ( .A1(n13625), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n13624), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13622) );
  AND2_X1 U16937 ( .A1(n13623), .A2(n13622), .ZN(n14047) );
  NOR2_X2 U16938 ( .A1(n14734), .A2(n14047), .ZN(n14046) );
  AOI222_X1 U16939 ( .A1(n13626), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n13625), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n13624), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13627) );
  NAND2_X1 U16940 ( .A1(n19132), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14826) );
  NOR2_X1 U16941 ( .A1(n15354), .A2(n13394), .ZN(n15353) );
  NOR2_X1 U16942 ( .A1(n15384), .A2(n19123), .ZN(n13634) );
  INV_X1 U16943 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13655) );
  NAND2_X1 U16944 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15401) );
  NOR2_X1 U16945 ( .A1(n13655), .A2(n15401), .ZN(n13664) );
  NAND2_X1 U16946 ( .A1(n13655), .A2(n15401), .ZN(n13632) );
  OAI211_X1 U16947 ( .C1(n13662), .C2(n13664), .A(n13632), .B(n15402), .ZN(
        n16218) );
  NOR2_X1 U16948 ( .A1(n13631), .A2(n16218), .ZN(n19124) );
  NAND2_X1 U16949 ( .A1(n13634), .A2(n19124), .ZN(n15369) );
  NOR2_X1 U16950 ( .A1(n15366), .A2(n15369), .ZN(n16201) );
  NAND2_X1 U16951 ( .A1(n15353), .A2(n16201), .ZN(n15250) );
  OR2_X1 U16952 ( .A1(n14975), .A2(n15195), .ZN(n13638) );
  NOR2_X1 U16953 ( .A1(n15250), .A2(n13638), .ZN(n15181) );
  NOR2_X1 U16954 ( .A1(n15172), .A2(n15183), .ZN(n13639) );
  NAND2_X1 U16955 ( .A1(n15181), .A2(n13639), .ZN(n15154) );
  INV_X1 U16956 ( .A(n13628), .ZN(n13629) );
  NAND2_X1 U16957 ( .A1(n13629), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13641) );
  NAND2_X1 U16958 ( .A1(n15090), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13630) );
  OR2_X1 U16959 ( .A1(n15103), .A2(n13630), .ZN(n15056) );
  NOR2_X1 U16960 ( .A1(n15056), .A2(n15069), .ZN(n15061) );
  NAND4_X1 U16961 ( .A1(n15061), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n13646), .ZN(n13647) );
  NAND3_X1 U16962 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13644) );
  INV_X1 U16963 ( .A(n15402), .ZN(n15252) );
  NAND2_X1 U16964 ( .A1(n15402), .A2(n13631), .ZN(n13633) );
  INV_X1 U16965 ( .A(n13632), .ZN(n13663) );
  NOR2_X1 U16966 ( .A1(n13654), .A2(n13664), .ZN(n13653) );
  AOI211_X1 U16967 ( .C1(n13662), .C2(n13663), .A(n13653), .B(n15399), .ZN(
        n16217) );
  NAND2_X1 U16968 ( .A1(n13633), .A2(n16217), .ZN(n19127) );
  INV_X1 U16969 ( .A(n13634), .ZN(n15378) );
  OR3_X1 U16970 ( .A1(n19127), .A2(n15378), .A3(n15366), .ZN(n13635) );
  NAND2_X1 U16971 ( .A1(n13645), .A2(n13635), .ZN(n16198) );
  INV_X1 U16972 ( .A(n15353), .ZN(n13636) );
  NAND2_X1 U16973 ( .A1(n15402), .A2(n13636), .ZN(n13637) );
  NAND2_X1 U16974 ( .A1(n16198), .A2(n13637), .ZN(n15334) );
  OAI21_X1 U16975 ( .B1(n15334), .B2(n13638), .A(n13645), .ZN(n15188) );
  INV_X1 U16976 ( .A(n13639), .ZN(n15169) );
  NAND2_X1 U16977 ( .A1(n13645), .A2(n15169), .ZN(n13640) );
  NAND2_X1 U16978 ( .A1(n15188), .A2(n13640), .ZN(n15157) );
  AND2_X1 U16979 ( .A1(n13645), .A2(n13641), .ZN(n13642) );
  NOR2_X1 U16980 ( .A1(n15157), .A2(n13642), .ZN(n15119) );
  OAI21_X1 U16981 ( .B1(n15090), .B2(n15252), .A(n15119), .ZN(n15082) );
  AOI211_X1 U16982 ( .C1(n15402), .C2(n13644), .A(n13643), .B(n15082), .ZN(
        n15043) );
  INV_X1 U16983 ( .A(n13645), .ZN(n15291) );
  OAI21_X1 U16984 ( .B1(n14834), .B2(n16192), .A(n13649), .ZN(P2_U3015) );
  NOR2_X1 U16985 ( .A1(n13650), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13679) );
  INV_X1 U16986 ( .A(n13651), .ZN(n13678) );
  NOR3_X1 U16987 ( .A1(n13679), .A2(n13678), .A3(n16192), .ZN(n13671) );
  INV_X1 U16988 ( .A(n15401), .ZN(n13652) );
  AND2_X1 U16989 ( .A1(n13653), .A2(n13652), .ZN(n13670) );
  INV_X1 U16990 ( .A(n13654), .ZN(n15208) );
  NAND2_X1 U16991 ( .A1(n15208), .A2(n15401), .ZN(n13656) );
  AOI21_X1 U16992 ( .B1(n13657), .B2(n13656), .A(n13655), .ZN(n13669) );
  OAI21_X1 U16993 ( .B1(n13660), .B2(n13659), .A(n13658), .ZN(n13661) );
  INV_X1 U16994 ( .A(n13661), .ZN(n13682) );
  NAND2_X1 U16995 ( .A1(n13682), .A2(n19129), .ZN(n13667) );
  NAND2_X1 U16996 ( .A1(n18885), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U16997 ( .A1(n19775), .A2(n19126), .ZN(n13666) );
  OAI21_X1 U16998 ( .B1(n13664), .B2(n13663), .A(n13662), .ZN(n13665) );
  NAND4_X1 U16999 ( .A1(n13667), .A2(n13675), .A3(n13666), .A4(n13665), .ZN(
        n13668) );
  NOR4_X1 U17000 ( .A1(n13671), .A2(n13670), .A3(n13669), .A4(n13668), .ZN(
        n13672) );
  OAI21_X1 U17001 ( .B1(n13691), .B2(n16191), .A(n13672), .ZN(P2_U3044) );
  INV_X1 U17002 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13677) );
  INV_X1 U17003 ( .A(n13673), .ZN(n13674) );
  NAND2_X1 U17004 ( .A1(n16178), .A2(n13674), .ZN(n13676) );
  OAI211_X1 U17005 ( .C1(n13677), .C2(n16186), .A(n13676), .B(n13675), .ZN(
        n13681) );
  NOR3_X1 U17006 ( .A1(n13679), .A2(n13678), .A3(n16179), .ZN(n13680) );
  AOI211_X1 U17007 ( .C1(n19115), .C2(n13682), .A(n13681), .B(n13680), .ZN(
        n13683) );
  OAI21_X1 U17008 ( .B1(n13691), .B2(n15430), .A(n13683), .ZN(P2_U3012) );
  INV_X2 U17009 ( .A(n19000), .ZN(n18996) );
  NOR2_X1 U17010 ( .A1(n18958), .A2(n18996), .ZN(n13684) );
  AOI21_X1 U17011 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n18996), .A(n13684), .ZN(
        n13685) );
  OAI21_X1 U17012 ( .B1(n19030), .B2(n18992), .A(n13685), .ZN(P2_U2887) );
  NAND2_X1 U17013 ( .A1(n13687), .A2(n13686), .ZN(n13688) );
  MUX2_X1 U17014 ( .A(n14697), .B(n14698), .S(n19000), .Z(n13690) );
  OAI21_X1 U17015 ( .B1(n19780), .B2(n18992), .A(n13690), .ZN(P2_U2886) );
  MUX2_X1 U17016 ( .A(n13691), .B(n12447), .S(n18996), .Z(n13692) );
  OAI21_X1 U17017 ( .B1(n19772), .B2(n18992), .A(n13692), .ZN(P2_U2885) );
  NOR2_X1 U17018 ( .A1(n13234), .A2(n18996), .ZN(n13693) );
  AOI21_X1 U17019 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n18996), .A(n13693), .ZN(
        n13694) );
  OAI21_X1 U17020 ( .B1(n19423), .B2(n18992), .A(n13694), .ZN(P2_U2884) );
  XOR2_X1 U17021 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n18934), .Z(n13700)
         );
  INV_X1 U17022 ( .A(n13695), .ZN(n13696) );
  AOI21_X1 U17023 ( .B1(n13697), .B2(n18938), .A(n13696), .ZN(n18915) );
  NOR2_X1 U17024 ( .A1(n19000), .A2(n12502), .ZN(n13698) );
  AOI21_X1 U17025 ( .B1(n18915), .B2(n19000), .A(n13698), .ZN(n13699) );
  OAI21_X1 U17026 ( .B1(n13700), .B2(n18992), .A(n13699), .ZN(P2_U2882) );
  XNOR2_X1 U17027 ( .A(n18991), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13705) );
  NOR2_X1 U17028 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  OR2_X1 U17029 ( .A1(n13027), .A2(n13703), .ZN(n18889) );
  MUX2_X1 U17030 ( .A(n18889), .B(n13047), .S(n18996), .Z(n13704) );
  OAI21_X1 U17031 ( .B1(n13705), .B2(n18992), .A(n13704), .ZN(P2_U2880) );
  CLKBUF_X1 U17032 ( .A(n13706), .Z(n18986) );
  XNOR2_X1 U17033 ( .A(n18986), .B(n18978), .ZN(n13711) );
  NAND2_X1 U17034 ( .A1(n13707), .A2(n15315), .ZN(n13709) );
  INV_X1 U17035 ( .A(n15275), .ZN(n13708) );
  AND2_X1 U17036 ( .A1(n13709), .A2(n13708), .ZN(n16150) );
  INV_X1 U17037 ( .A(n16150), .ZN(n15297) );
  MUX2_X1 U17038 ( .A(n12746), .B(n15297), .S(n19000), .Z(n13710) );
  OAI21_X1 U17039 ( .B1(n13711), .B2(n18992), .A(n13710), .ZN(P2_U2876) );
  AOI22_X1 U17040 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13836), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U17041 ( .A1(n12279), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U17042 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U17043 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13712) );
  NAND4_X1 U17044 ( .A1(n13715), .A2(n13714), .A3(n13713), .A4(n13712), .ZN(
        n13721) );
  AOI22_X1 U17045 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13719) );
  AOI22_X1 U17046 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13718) );
  AOI22_X1 U17047 ( .A1(n12205), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U17048 ( .A1(n12206), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13716) );
  NAND4_X1 U17049 ( .A1(n13719), .A2(n13718), .A3(n13717), .A4(n13716), .ZN(
        n13720) );
  NOR2_X1 U17050 ( .A1(n13721), .A2(n13720), .ZN(n18970) );
  AOI22_X1 U17051 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13836), .ZN(n13726) );
  AOI22_X1 U17052 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13725) );
  AOI22_X1 U17053 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13724) );
  AOI22_X1 U17054 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13723) );
  NAND4_X1 U17055 ( .A1(n13726), .A2(n13725), .A3(n13724), .A4(n13723), .ZN(
        n13732) );
  AOI22_X1 U17056 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13730) );
  AOI22_X1 U17057 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13729) );
  AOI22_X1 U17058 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11986), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13728) );
  AOI22_X1 U17059 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12654), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13727) );
  NAND4_X1 U17060 ( .A1(n13730), .A2(n13729), .A3(n13728), .A4(n13727), .ZN(
        n13731) );
  NOR2_X1 U17061 ( .A1(n13732), .A2(n13731), .ZN(n14731) );
  NOR2_X2 U17062 ( .A1(n14729), .A2(n14731), .ZN(n14730) );
  AOI22_X1 U17063 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n13836), .ZN(n13736) );
  AOI22_X1 U17064 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13735) );
  AOI22_X1 U17065 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13734) );
  AOI22_X1 U17066 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13733) );
  NAND4_X1 U17067 ( .A1(n13736), .A2(n13735), .A3(n13734), .A4(n13733), .ZN(
        n13742) );
  AOI22_X1 U17068 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13740) );
  AOI22_X1 U17069 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13739) );
  AOI22_X1 U17070 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11986), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13738) );
  AOI22_X1 U17071 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12654), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13737) );
  NAND4_X1 U17072 ( .A1(n13740), .A2(n13739), .A3(n13738), .A4(n13737), .ZN(
        n13741) );
  NOR2_X1 U17073 ( .A1(n13742), .A2(n13741), .ZN(n16106) );
  INV_X1 U17074 ( .A(n16106), .ZN(n13743) );
  AND2_X2 U17075 ( .A1(n14730), .A2(n13743), .ZN(n13754) );
  AOI22_X1 U17076 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n13836), .ZN(n13747) );
  AOI22_X1 U17077 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13746) );
  AOI22_X1 U17078 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13745) );
  AOI22_X1 U17079 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13744) );
  NAND4_X1 U17080 ( .A1(n13747), .A2(n13746), .A3(n13745), .A4(n13744), .ZN(
        n13753) );
  AOI22_X1 U17081 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13751) );
  AOI22_X1 U17082 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13750) );
  AOI22_X1 U17083 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11986), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13749) );
  AOI22_X1 U17084 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12654), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13748) );
  NAND4_X1 U17085 ( .A1(n13751), .A2(n13750), .A3(n13749), .A4(n13748), .ZN(
        n13752) );
  OR2_X1 U17086 ( .A1(n13753), .A2(n13752), .ZN(n13756) );
  INV_X1 U17087 ( .A(n9884), .ZN(n13755) );
  OAI21_X1 U17088 ( .B1(n13754), .B2(n13756), .A(n13755), .ZN(n14815) );
  NOR2_X1 U17089 ( .A1(n14978), .A2(n13757), .ZN(n13758) );
  OR2_X1 U17090 ( .A1(n14953), .A2(n13758), .ZN(n18773) );
  NOR2_X1 U17091 ( .A1(n18773), .A2(n18996), .ZN(n13759) );
  AOI21_X1 U17092 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n18996), .A(n13759), .ZN(
        n13760) );
  OAI21_X1 U17093 ( .B1(n14815), .B2(n18992), .A(n13760), .ZN(P2_U2868) );
  INV_X1 U17094 ( .A(n14035), .ZN(n13995) );
  INV_X1 U17095 ( .A(n14034), .ZN(n14004) );
  OAI22_X1 U17096 ( .A1(n13995), .A2(n13762), .B1(n14004), .B2(n13761), .ZN(
        n13766) );
  INV_X1 U17097 ( .A(n14036), .ZN(n14008) );
  INV_X1 U17098 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13764) );
  INV_X1 U17099 ( .A(n11946), .ZN(n14006) );
  OAI22_X1 U17100 ( .A1(n14008), .A2(n13764), .B1(n14006), .B2(n13763), .ZN(
        n13765) );
  NOR2_X1 U17101 ( .A1(n13766), .A2(n13765), .ZN(n13771) );
  AOI22_X1 U17102 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13770) );
  AOI22_X1 U17103 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13769) );
  XNOR2_X1 U17104 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14027) );
  NAND4_X1 U17105 ( .A1(n13771), .A2(n13770), .A3(n13769), .A4(n14027), .ZN(
        n13780) );
  OAI22_X1 U17106 ( .A1(n13995), .A2(n13772), .B1(n14004), .B2(n13272), .ZN(
        n13775) );
  OAI22_X1 U17107 ( .A1(n14008), .A2(n13773), .B1(n14006), .B2(n21044), .ZN(
        n13774) );
  NOR2_X1 U17108 ( .A1(n13775), .A2(n13774), .ZN(n13778) );
  INV_X1 U17109 ( .A(n14027), .ZN(n14032) );
  AOI22_X1 U17110 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13777) );
  AOI22_X1 U17111 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13776) );
  NAND4_X1 U17112 ( .A1(n13778), .A2(n14032), .A3(n13777), .A4(n13776), .ZN(
        n13779) );
  AND2_X1 U17113 ( .A1(n13780), .A2(n13779), .ZN(n13855) );
  NAND2_X1 U17114 ( .A1(n10055), .A2(n13855), .ZN(n13865) );
  AOI22_X1 U17115 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n13836), .ZN(n13784) );
  AOI22_X1 U17116 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13783) );
  AOI22_X1 U17117 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13782) );
  AOI22_X1 U17118 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13781) );
  NAND4_X1 U17119 ( .A1(n13784), .A2(n13783), .A3(n13782), .A4(n13781), .ZN(
        n13790) );
  AOI22_X1 U17120 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U17121 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U17122 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12205), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13786) );
  AOI22_X1 U17123 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12654), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13785) );
  NAND4_X1 U17124 ( .A1(n13788), .A2(n13787), .A3(n13786), .A4(n13785), .ZN(
        n13789) );
  OR2_X1 U17125 ( .A1(n13790), .A2(n13789), .ZN(n16103) );
  AOI22_X1 U17126 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13836), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13799) );
  AOI22_X1 U17127 ( .A1(n12279), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U17128 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13797) );
  INV_X1 U17129 ( .A(n13791), .ZN(n13793) );
  OAI22_X1 U17130 ( .A1(n13794), .A2(n13306), .B1(n13793), .B2(n13792), .ZN(
        n13795) );
  INV_X1 U17131 ( .A(n13795), .ZN(n13796) );
  NAND4_X1 U17132 ( .A1(n13799), .A2(n13798), .A3(n13797), .A4(n13796), .ZN(
        n13805) );
  AOI22_X1 U17133 ( .A1(n11984), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13803) );
  AOI22_X1 U17134 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13802) );
  AOI22_X1 U17135 ( .A1(n12205), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13801) );
  AOI22_X1 U17136 ( .A1(n12206), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12654), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13800) );
  NAND4_X1 U17137 ( .A1(n13803), .A2(n13802), .A3(n13801), .A4(n13800), .ZN(
        n13804) );
  NOR2_X1 U17138 ( .A1(n13805), .A2(n13804), .ZN(n14724) );
  AOI22_X1 U17139 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n13836), .ZN(n13809) );
  AOI22_X1 U17140 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U17141 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13807) );
  AOI22_X1 U17142 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13806) );
  NAND4_X1 U17143 ( .A1(n13809), .A2(n13808), .A3(n13807), .A4(n13806), .ZN(
        n13815) );
  AOI22_X1 U17144 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13813) );
  AOI22_X1 U17145 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13812) );
  AOI22_X1 U17146 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11986), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13811) );
  AOI22_X1 U17147 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12654), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13810) );
  NAND4_X1 U17148 ( .A1(n13813), .A2(n13812), .A3(n13811), .A4(n13810), .ZN(
        n13814) );
  OR2_X1 U17149 ( .A1(n13815), .A2(n13814), .ZN(n14792) );
  INV_X1 U17150 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13817) );
  INV_X1 U17151 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13816) );
  OAI22_X1 U17152 ( .A1(n13995), .A2(n13817), .B1(n14004), .B2(n13816), .ZN(
        n13821) );
  INV_X1 U17153 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13819) );
  INV_X1 U17154 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13818) );
  OAI22_X1 U17155 ( .A1(n14008), .A2(n13819), .B1(n14006), .B2(n13818), .ZN(
        n13820) );
  NOR2_X1 U17156 ( .A1(n13821), .A2(n13820), .ZN(n13824) );
  AOI22_X1 U17157 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11949), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13823) );
  AOI22_X1 U17158 ( .A1(n9786), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13822) );
  NAND4_X1 U17159 ( .A1(n13824), .A2(n13823), .A3(n13822), .A4(n14027), .ZN(
        n13835) );
  INV_X1 U17160 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13826) );
  INV_X1 U17161 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13825) );
  OAI22_X1 U17162 ( .A1(n11956), .A2(n13826), .B1(n14004), .B2(n13825), .ZN(
        n13830) );
  INV_X1 U17163 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13828) );
  INV_X1 U17164 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13827) );
  OAI22_X1 U17165 ( .A1(n14008), .A2(n13828), .B1(n14006), .B2(n13827), .ZN(
        n13829) );
  NOR2_X1 U17166 ( .A1(n13830), .A2(n13829), .ZN(n13833) );
  AOI22_X1 U17167 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U17168 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14035), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13831) );
  NAND4_X1 U17169 ( .A1(n13833), .A2(n14032), .A3(n13832), .A4(n13831), .ZN(
        n13834) );
  NAND2_X1 U17170 ( .A1(n13835), .A2(n13834), .ZN(n13866) );
  NOR2_X1 U17171 ( .A1(n10055), .A2(n13866), .ZN(n13849) );
  AOI22_X1 U17172 ( .A1(n12200), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13836), .ZN(n13842) );
  AOI22_X1 U17173 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12279), .B1(
        n13837), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13841) );
  AOI22_X1 U17174 ( .A1(n12151), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13838), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U17175 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13791), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13839) );
  NAND4_X1 U17176 ( .A1(n13842), .A2(n13841), .A3(n13840), .A4(n13839), .ZN(
        n13848) );
  AOI22_X1 U17177 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12152), .B1(
        n11984), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17178 ( .A1(n11985), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12170), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17179 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11986), .B1(
        n12205), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17180 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12654), .B1(
        n12206), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13843) );
  NAND4_X1 U17181 ( .A1(n13846), .A2(n13845), .A3(n13844), .A4(n13843), .ZN(
        n13847) );
  XNOR2_X1 U17182 ( .A(n13849), .B(n13854), .ZN(n13867) );
  INV_X1 U17183 ( .A(n13866), .ZN(n13853) );
  NAND2_X1 U17184 ( .A1(n10055), .A2(n13853), .ZN(n14785) );
  INV_X1 U17185 ( .A(n13867), .ZN(n13852) );
  AND2_X1 U17186 ( .A1(n13854), .A2(n13853), .ZN(n13856) );
  NAND2_X1 U17187 ( .A1(n13856), .A2(n13855), .ZN(n13868) );
  OAI211_X1 U17188 ( .C1(n13856), .C2(n13855), .A(n13948), .B(n13868), .ZN(
        n13857) );
  AOI21_X1 U17189 ( .B1(n13858), .B2(n13857), .A(n9849), .ZN(n13859) );
  XOR2_X1 U17190 ( .A(n13865), .B(n13859), .Z(n14783) );
  OR2_X1 U17191 ( .A1(n14617), .A2(n13861), .ZN(n13862) );
  NAND2_X1 U17192 ( .A1(n13860), .A2(n13862), .ZN(n14897) );
  NOR2_X1 U17193 ( .A1(n14897), .A2(n18996), .ZN(n13863) );
  AOI21_X1 U17194 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n18996), .A(n13863), .ZN(
        n13864) );
  OAI21_X1 U17195 ( .B1(n14783), .B2(n18992), .A(n13864), .ZN(P2_U2863) );
  INV_X1 U17196 ( .A(n13868), .ZN(n13889) );
  INV_X1 U17197 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13870) );
  INV_X1 U17198 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13869) );
  OAI22_X1 U17199 ( .A1(n13995), .A2(n13870), .B1(n14004), .B2(n13869), .ZN(
        n13874) );
  INV_X1 U17200 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13872) );
  INV_X1 U17201 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13871) );
  OAI22_X1 U17202 ( .A1(n14008), .A2(n13872), .B1(n14006), .B2(n13871), .ZN(
        n13873) );
  NOR2_X1 U17203 ( .A1(n13874), .A2(n13873), .ZN(n13877) );
  AOI22_X1 U17204 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U17205 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13875) );
  NAND4_X1 U17206 ( .A1(n13877), .A2(n13876), .A3(n13875), .A4(n14027), .ZN(
        n13888) );
  INV_X1 U17207 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13879) );
  INV_X1 U17208 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13878) );
  OAI22_X1 U17209 ( .A1(n13995), .A2(n13879), .B1(n14004), .B2(n13878), .ZN(
        n13883) );
  INV_X1 U17210 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13881) );
  INV_X1 U17211 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13880) );
  OAI22_X1 U17212 ( .A1(n14008), .A2(n13881), .B1(n14006), .B2(n13880), .ZN(
        n13882) );
  NOR2_X1 U17213 ( .A1(n13883), .A2(n13882), .ZN(n13886) );
  AOI22_X1 U17214 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U17215 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9786), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13884) );
  NAND4_X1 U17216 ( .A1(n13886), .A2(n14032), .A3(n13885), .A4(n13884), .ZN(
        n13887) );
  AND2_X1 U17217 ( .A1(n13888), .A2(n13887), .ZN(n13890) );
  NAND2_X1 U17218 ( .A1(n13889), .A2(n13890), .ZN(n13923) );
  OAI211_X1 U17219 ( .C1(n13889), .C2(n13890), .A(n13948), .B(n13923), .ZN(
        n13898) );
  INV_X1 U17220 ( .A(n13890), .ZN(n13891) );
  NOR2_X1 U17221 ( .A1(n14018), .A2(n13891), .ZN(n13892) );
  OAI21_X1 U17222 ( .B1(n13893), .B2(n13892), .A(n13901), .ZN(n14778) );
  NAND2_X1 U17223 ( .A1(n13860), .A2(n13894), .ZN(n13895) );
  NAND2_X1 U17224 ( .A1(n14713), .A2(n13895), .ZN(n15099) );
  MUX2_X1 U17225 ( .A(n16085), .B(n15099), .S(n19000), .Z(n13896) );
  OAI21_X1 U17226 ( .B1(n14778), .B2(n18992), .A(n13896), .ZN(P2_U2862) );
  OAI22_X1 U17227 ( .A1(n13995), .A2(n13903), .B1(n14004), .B2(n13902), .ZN(
        n13907) );
  OAI22_X1 U17228 ( .A1(n14008), .A2(n13905), .B1(n14006), .B2(n13904), .ZN(
        n13906) );
  NOR2_X1 U17229 ( .A1(n13907), .A2(n13906), .ZN(n13910) );
  AOI22_X1 U17230 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U17231 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13908) );
  NAND4_X1 U17232 ( .A1(n13910), .A2(n13909), .A3(n13908), .A4(n14027), .ZN(
        n13921) );
  OAI22_X1 U17233 ( .A1(n13995), .A2(n13912), .B1(n14004), .B2(n13911), .ZN(
        n13916) );
  OAI22_X1 U17234 ( .A1(n14008), .A2(n13914), .B1(n14006), .B2(n13913), .ZN(
        n13915) );
  NOR2_X1 U17235 ( .A1(n13916), .A2(n13915), .ZN(n13919) );
  AOI22_X1 U17236 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U17237 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9786), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13917) );
  NAND4_X1 U17238 ( .A1(n13919), .A2(n14032), .A3(n13918), .A4(n13917), .ZN(
        n13920) );
  NAND2_X1 U17239 ( .A1(n13921), .A2(n13920), .ZN(n13925) );
  AOI21_X1 U17240 ( .B1(n13923), .B2(n13925), .A(n13922), .ZN(n13924) );
  INV_X1 U17241 ( .A(n13925), .ZN(n13926) );
  NAND2_X1 U17242 ( .A1(n10055), .A2(n13926), .ZN(n14719) );
  NOR2_X2 U17243 ( .A1(n14720), .A2(n14719), .ZN(n14718) );
  INV_X1 U17244 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13929) );
  INV_X1 U17245 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13928) );
  OAI22_X1 U17246 ( .A1(n11956), .A2(n13929), .B1(n14004), .B2(n13928), .ZN(
        n13933) );
  INV_X1 U17247 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13931) );
  INV_X1 U17248 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13930) );
  OAI22_X1 U17249 ( .A1(n14008), .A2(n13931), .B1(n14006), .B2(n13930), .ZN(
        n13932) );
  NOR2_X1 U17250 ( .A1(n13933), .A2(n13932), .ZN(n13936) );
  AOI22_X1 U17251 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11949), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13935) );
  INV_X1 U17252 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n20945) );
  AOI22_X1 U17253 ( .A1(n14035), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13934) );
  NAND4_X1 U17254 ( .A1(n13936), .A2(n13935), .A3(n13934), .A4(n14027), .ZN(
        n13946) );
  INV_X1 U17255 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n19530) );
  INV_X1 U17256 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13937) );
  OAI22_X1 U17257 ( .A1(n13995), .A2(n19530), .B1(n14004), .B2(n13937), .ZN(
        n13941) );
  INV_X1 U17258 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13939) );
  INV_X1 U17259 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13938) );
  OAI22_X1 U17260 ( .A1(n14008), .A2(n13939), .B1(n14006), .B2(n13938), .ZN(
        n13940) );
  NOR2_X1 U17261 ( .A1(n13941), .A2(n13940), .ZN(n13944) );
  AOI22_X1 U17262 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13943) );
  INV_X1 U17263 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n20959) );
  AOI22_X1 U17264 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13942) );
  NAND4_X1 U17265 ( .A1(n13944), .A2(n14032), .A3(n13943), .A4(n13942), .ZN(
        n13945) );
  NAND2_X1 U17266 ( .A1(n13946), .A2(n13945), .ZN(n13954) );
  INV_X1 U17267 ( .A(n13954), .ZN(n13950) );
  INV_X1 U17268 ( .A(n13947), .ZN(n13949) );
  OR2_X1 U17269 ( .A1(n13947), .A2(n13954), .ZN(n13962) );
  OAI211_X1 U17270 ( .C1(n13950), .C2(n13949), .A(n13962), .B(n13948), .ZN(
        n13951) );
  NOR2_X1 U17271 ( .A1(n13952), .A2(n13951), .ZN(n13961) );
  NOR2_X1 U17272 ( .A1(n13271), .A2(n13954), .ZN(n13956) );
  NAND2_X1 U17273 ( .A1(n13955), .A2(n13956), .ZN(n13992) );
  OAI21_X1 U17274 ( .B1(n13955), .B2(n13956), .A(n13992), .ZN(n14755) );
  AND2_X1 U17275 ( .A1(n14715), .A2(n13957), .ZN(n13958) );
  OR2_X1 U17276 ( .A1(n13958), .A2(n13985), .ZN(n15078) );
  NOR2_X1 U17277 ( .A1(n15078), .A2(n18996), .ZN(n13959) );
  AOI21_X1 U17278 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n18996), .A(n13959), .ZN(
        n13960) );
  OAI21_X1 U17279 ( .B1(n14755), .B2(n18992), .A(n13960), .ZN(P2_U2860) );
  INV_X1 U17280 ( .A(n13962), .ZN(n14020) );
  NOR2_X1 U17281 ( .A1(n13961), .A2(n14020), .ZN(n13983) );
  OAI22_X1 U17282 ( .A1(n13995), .A2(n13964), .B1(n14004), .B2(n13963), .ZN(
        n13968) );
  OAI22_X1 U17283 ( .A1(n14008), .A2(n13966), .B1(n14006), .B2(n13965), .ZN(
        n13967) );
  NOR2_X1 U17284 ( .A1(n13968), .A2(n13967), .ZN(n13971) );
  AOI22_X1 U17285 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13970) );
  AOI22_X1 U17286 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13969) );
  NAND4_X1 U17287 ( .A1(n13971), .A2(n13970), .A3(n13969), .A4(n14027), .ZN(
        n13982) );
  OAI22_X1 U17288 ( .A1(n13995), .A2(n13973), .B1(n14004), .B2(n13972), .ZN(
        n13977) );
  OAI22_X1 U17289 ( .A1(n14008), .A2(n13975), .B1(n14006), .B2(n13974), .ZN(
        n13976) );
  NOR2_X1 U17290 ( .A1(n13977), .A2(n13976), .ZN(n13980) );
  AOI22_X1 U17291 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13979) );
  AOI22_X1 U17292 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9786), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13978) );
  NAND4_X1 U17293 ( .A1(n13980), .A2(n14032), .A3(n13979), .A4(n13978), .ZN(
        n13981) );
  NAND2_X1 U17294 ( .A1(n13982), .A2(n13981), .ZN(n14016) );
  XNOR2_X1 U17295 ( .A(n13983), .B(n14016), .ZN(n14749) );
  NOR2_X1 U17296 ( .A1(n15065), .A2(n18996), .ZN(n13986) );
  AOI21_X1 U17297 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n18996), .A(n13986), .ZN(
        n13987) );
  OAI21_X1 U17298 ( .B1(n14749), .B2(n18992), .A(n13987), .ZN(P2_U2859) );
  INV_X1 U17299 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16308) );
  NAND3_X1 U17300 ( .A1(n13988), .A2(n20091), .A3(n14271), .ZN(n13990) );
  AOI22_X1 U17301 ( .A1(n14265), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14235), .ZN(n13989) );
  OAI211_X1 U17302 ( .C1(n14239), .C2(n16308), .A(n13990), .B(n13989), .ZN(
        P1_U2873) );
  INV_X1 U17303 ( .A(n13961), .ZN(n13991) );
  AOI21_X2 U17304 ( .B1(n13992), .B2(n13991), .A(n14016), .ZN(n14709) );
  OAI22_X1 U17305 ( .A1(n13995), .A2(n13994), .B1(n14004), .B2(n13993), .ZN(
        n13999) );
  OAI22_X1 U17306 ( .A1(n14008), .A2(n13997), .B1(n14006), .B2(n13996), .ZN(
        n13998) );
  NOR2_X1 U17307 ( .A1(n13999), .A2(n13998), .ZN(n14002) );
  AOI22_X1 U17308 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U17309 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14000) );
  NAND4_X1 U17310 ( .A1(n14002), .A2(n14001), .A3(n14000), .A4(n14027), .ZN(
        n14015) );
  OAI22_X1 U17311 ( .A1(n11956), .A2(n13367), .B1(n14004), .B2(n14003), .ZN(
        n14010) );
  OAI22_X1 U17312 ( .A1(n14008), .A2(n14007), .B1(n14006), .B2(n14005), .ZN(
        n14009) );
  NOR2_X1 U17313 ( .A1(n14010), .A2(n14009), .ZN(n14013) );
  AOI22_X1 U17314 ( .A1(n11949), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14012) );
  AOI22_X1 U17315 ( .A1(n13768), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14035), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14011) );
  NAND4_X1 U17316 ( .A1(n14013), .A2(n14032), .A3(n14012), .A4(n14011), .ZN(
        n14014) );
  NAND2_X1 U17317 ( .A1(n14015), .A2(n14014), .ZN(n14022) );
  INV_X1 U17318 ( .A(n14016), .ZN(n14017) );
  AND2_X1 U17319 ( .A1(n14018), .A2(n14017), .ZN(n14019) );
  NAND2_X1 U17320 ( .A1(n14020), .A2(n14019), .ZN(n14021) );
  NOR2_X1 U17321 ( .A1(n14021), .A2(n14022), .ZN(n14023) );
  AOI21_X1 U17322 ( .B1(n14022), .B2(n14021), .A(n14023), .ZN(n14708) );
  NAND2_X1 U17323 ( .A1(n14709), .A2(n14708), .ZN(n14710) );
  INV_X1 U17324 ( .A(n14023), .ZN(n14024) );
  NAND2_X1 U17325 ( .A1(n14710), .A2(n14024), .ZN(n14045) );
  AOI22_X1 U17326 ( .A1(n14035), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14026) );
  AOI22_X1 U17327 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9784), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14025) );
  NAND2_X1 U17328 ( .A1(n14026), .A2(n14025), .ZN(n14042) );
  AOI22_X1 U17329 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9786), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14029) );
  AOI22_X1 U17330 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14028) );
  NAND3_X1 U17331 ( .A1(n14029), .A2(n14028), .A3(n14027), .ZN(n14041) );
  AOI22_X1 U17332 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11955), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U17333 ( .A1(n13767), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14030), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14031) );
  NAND3_X1 U17334 ( .A1(n14033), .A2(n14032), .A3(n14031), .ZN(n14040) );
  AOI22_X1 U17335 ( .A1(n14035), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14034), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14038) );
  AOI22_X1 U17336 ( .A1(n14036), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11946), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14037) );
  NAND2_X1 U17337 ( .A1(n14038), .A2(n14037), .ZN(n14039) );
  OAI22_X1 U17338 ( .A1(n14042), .A2(n14041), .B1(n14040), .B2(n14039), .ZN(
        n14043) );
  INV_X1 U17339 ( .A(n14043), .ZN(n14044) );
  XNOR2_X1 U17340 ( .A(n14045), .B(n14044), .ZN(n14058) );
  AOI21_X1 U17341 ( .B1(n14047), .B2(n14734), .A(n14046), .ZN(n16048) );
  NOR2_X2 U17342 ( .A1(n14049), .A2(n15431), .ZN(n19006) );
  INV_X1 U17343 ( .A(n19006), .ZN(n14765) );
  INV_X1 U17344 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U17345 ( .A1(n19005), .A2(n14048), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19056), .ZN(n14051) );
  NOR2_X2 U17346 ( .A1(n14049), .A2(n15429), .ZN(n19007) );
  NAND2_X1 U17347 ( .A1(n19007), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14050) );
  OAI211_X1 U17348 ( .C1(n14765), .C2(n14052), .A(n14051), .B(n14050), .ZN(
        n14053) );
  AOI21_X1 U17349 ( .B1(n16048), .B2(n19057), .A(n14053), .ZN(n14054) );
  OAI21_X1 U17350 ( .B1(n14058), .B2(n19061), .A(n14054), .ZN(P2_U2889) );
  XNOR2_X1 U17351 ( .A(n14707), .B(n14055), .ZN(n16046) );
  NOR2_X1 U17352 ( .A1(n16046), .A2(n18996), .ZN(n14056) );
  AOI21_X1 U17353 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n18996), .A(n14056), .ZN(
        n14057) );
  OAI21_X1 U17354 ( .B1(n14058), .B2(n18992), .A(n14057), .ZN(P2_U2857) );
  INV_X1 U17355 ( .A(n14060), .ZN(n14066) );
  INV_X1 U17356 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20690) );
  INV_X1 U17357 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14061) );
  OAI21_X1 U17358 ( .B1(n14075), .B2(n20690), .A(n14061), .ZN(n14063) );
  NAND2_X1 U17359 ( .A1(n14063), .A2(n14062), .ZN(n14065) );
  AOI22_X1 U17360 ( .A1(n19901), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19897), .ZN(n14064) );
  OAI211_X1 U17361 ( .C1(n14066), .C2(n19906), .A(n14065), .B(n14064), .ZN(
        n14067) );
  AOI21_X1 U17362 ( .B1(n11471), .B2(n19880), .A(n14067), .ZN(n14068) );
  OAI21_X1 U17363 ( .B1(n14069), .B2(n19847), .A(n14068), .ZN(P1_U2810) );
  AOI21_X1 U17364 ( .B1(n14072), .B2(n14071), .A(n14070), .ZN(n14279) );
  INV_X1 U17365 ( .A(n14279), .ZN(n14217) );
  AOI21_X1 U17366 ( .B1(n14074), .B2(n9839), .A(n14073), .ZN(n14404) );
  NOR2_X1 U17367 ( .A1(n14075), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U17368 ( .A1(n19901), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19897), .ZN(n14078) );
  NAND2_X1 U17369 ( .A1(n14076), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14077) );
  OAI211_X1 U17370 ( .C1(n19906), .C2(n14277), .A(n14078), .B(n14077), .ZN(
        n14079) );
  AOI211_X1 U17371 ( .C1(n14404), .C2(n19880), .A(n14080), .B(n14079), .ZN(
        n14081) );
  OAI21_X1 U17372 ( .B1(n14217), .B2(n19847), .A(n14081), .ZN(P1_U2811) );
  OR2_X1 U17373 ( .A1(n14097), .A2(n14082), .ZN(n14083) );
  NAND2_X1 U17374 ( .A1(n9853), .A2(n14083), .ZN(n14421) );
  AOI21_X1 U17375 ( .B1(n14086), .B2(n14084), .A(n14085), .ZN(n14300) );
  NAND2_X1 U17376 ( .A1(n14300), .A2(n19873), .ZN(n14094) );
  INV_X1 U17377 ( .A(n14298), .ZN(n14092) );
  INV_X1 U17378 ( .A(n14087), .ZN(n14088) );
  NAND2_X1 U17379 ( .A1(n19885), .A2(n14088), .ZN(n14101) );
  INV_X1 U17380 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20985) );
  AOI22_X1 U17381 ( .A1(n19901), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19897), .ZN(n14089) );
  OAI21_X1 U17382 ( .B1(n14101), .B2(n20985), .A(n14089), .ZN(n14091) );
  INV_X1 U17383 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20856) );
  NOR3_X1 U17384 ( .A1(n14102), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n20856), 
        .ZN(n14090) );
  AOI211_X1 U17385 ( .C1(n19838), .C2(n14092), .A(n14091), .B(n14090), .ZN(
        n14093) );
  OAI211_X1 U17386 ( .C1(n19892), .C2(n14421), .A(n14094), .B(n14093), .ZN(
        P1_U2813) );
  NOR2_X1 U17387 ( .A1(n14112), .A2(n14095), .ZN(n14096) );
  OR2_X1 U17388 ( .A1(n14097), .A2(n14096), .ZN(n14433) );
  INV_X1 U17389 ( .A(n14306), .ZN(n14100) );
  NAND2_X1 U17390 ( .A1(n14100), .A2(n19873), .ZN(n14106) );
  OAI22_X1 U17391 ( .A1(n19866), .A2(n14160), .B1(n14305), .B2(n15826), .ZN(
        n14104) );
  AOI21_X1 U17392 ( .B1(n14102), .B2(n20856), .A(n14101), .ZN(n14103) );
  AOI211_X1 U17393 ( .C1(n19838), .C2(n14309), .A(n14104), .B(n14103), .ZN(
        n14105) );
  OAI211_X1 U17394 ( .C1(n19892), .C2(n14433), .A(n14106), .B(n14105), .ZN(
        P1_U2814) );
  AOI21_X1 U17395 ( .B1(n14108), .B2(n14107), .A(n14098), .ZN(n14319) );
  INV_X1 U17396 ( .A(n14319), .ZN(n14228) );
  INV_X1 U17397 ( .A(n14124), .ZN(n14110) );
  OAI21_X1 U17398 ( .B1(n15751), .B2(n14110), .A(n14109), .ZN(n14111) );
  INV_X1 U17399 ( .A(n14111), .ZN(n14113) );
  OR2_X1 U17400 ( .A1(n14113), .A2(n14112), .ZN(n14441) );
  INV_X1 U17401 ( .A(n14441), .ZN(n14119) );
  INV_X1 U17402 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20683) );
  AOI21_X1 U17403 ( .B1(n19878), .B2(n14125), .A(n15758), .ZN(n15756) );
  OAI21_X1 U17404 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n19891), .A(n15756), 
        .ZN(n14115) );
  INV_X1 U17405 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14161) );
  OAI22_X1 U17406 ( .A1(n10976), .A2(n15826), .B1(n14161), .B2(n19866), .ZN(
        n14114) );
  AOI221_X1 U17407 ( .B1(n14116), .B2(n20683), .C1(n14115), .C2(
        P1_REIP_REG_25__SCAN_IN), .A(n14114), .ZN(n14117) );
  OAI21_X1 U17408 ( .B1(n14317), .B2(n19906), .A(n14117), .ZN(n14118) );
  AOI21_X1 U17409 ( .B1(n14119), .B2(n19880), .A(n14118), .ZN(n14120) );
  OAI21_X1 U17410 ( .B1(n14228), .B2(n19847), .A(n14120), .ZN(P1_U2815) );
  OAI21_X1 U17412 ( .B1(n14122), .B2(n14123), .A(n14107), .ZN(n14325) );
  XNOR2_X1 U17413 ( .A(n15751), .B(n14124), .ZN(n14461) );
  INV_X1 U17414 ( .A(n14328), .ZN(n14130) );
  NOR3_X1 U17415 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n19891), .A3(n14125), 
        .ZN(n14128) );
  OAI22_X1 U17416 ( .A1(n15756), .A2(n20681), .B1(n14126), .B2(n19866), .ZN(
        n14127) );
  AOI211_X1 U17417 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14128), .B(n14127), .ZN(n14129) );
  OAI21_X1 U17418 ( .B1(n14130), .B2(n19906), .A(n14129), .ZN(n14131) );
  AOI21_X1 U17419 ( .B1(n14461), .B2(n19880), .A(n14131), .ZN(n14132) );
  OAI21_X1 U17420 ( .B1(n14325), .B2(n19847), .A(n14132), .ZN(P1_U2816) );
  OAI21_X1 U17421 ( .B1(n14133), .B2(n14135), .A(n14191), .ZN(n15886) );
  INV_X1 U17422 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20669) );
  NAND2_X1 U17423 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15803) );
  NOR2_X1 U17424 ( .A1(n20669), .A2(n15803), .ZN(n14138) );
  OAI21_X1 U17425 ( .B1(n14136), .B2(n19832), .A(n19885), .ZN(n15822) );
  OAI21_X1 U17426 ( .B1(n14138), .B2(n14137), .A(n15822), .ZN(n15796) );
  NAND2_X1 U17427 ( .A1(n19878), .A2(n14139), .ZN(n15805) );
  OAI21_X1 U17428 ( .B1(n15803), .B2(n15805), .A(n20669), .ZN(n14141) );
  INV_X1 U17429 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14194) );
  OAI22_X1 U17430 ( .A1(n21018), .A2(n15826), .B1(n14194), .B2(n19866), .ZN(
        n14140) );
  AOI211_X1 U17431 ( .C1(n15796), .C2(n14141), .A(n19895), .B(n14140), .ZN(
        n14146) );
  NAND2_X1 U17432 ( .A1(n14201), .A2(n14142), .ZN(n14143) );
  AND2_X1 U17433 ( .A1(n14144), .A2(n14143), .ZN(n15944) );
  AOI22_X1 U17434 ( .A1(n19838), .A2(n15887), .B1(n19880), .B2(n15944), .ZN(
        n14145) );
  OAI211_X1 U17435 ( .C1(n15886), .C2(n19847), .A(n14146), .B(n14145), .ZN(
        P1_U2823) );
  INV_X1 U17436 ( .A(n14148), .ZN(n14149) );
  AOI21_X1 U17437 ( .B1(n14150), .B2(n14205), .A(n14149), .ZN(n15894) );
  INV_X1 U17438 ( .A(n15894), .ZN(n14270) );
  AND2_X1 U17439 ( .A1(n9878), .A2(n14151), .ZN(n14152) );
  OR2_X1 U17440 ( .A1(n14199), .A2(n14152), .ZN(n15958) );
  INV_X1 U17441 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14204) );
  OAI22_X1 U17442 ( .A1(n15958), .A2(n19892), .B1(n19866), .B2(n14204), .ZN(
        n14155) );
  INV_X1 U17443 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20665) );
  AOI21_X1 U17444 ( .B1(n19897), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n19895), .ZN(n14153) );
  OAI221_X1 U17445 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15805), .C1(n20665), 
        .C2(n15822), .A(n14153), .ZN(n14154) );
  AOI211_X1 U17446 ( .C1(n15893), .C2(n19838), .A(n14155), .B(n14154), .ZN(
        n14156) );
  OAI21_X1 U17447 ( .B1(n14270), .B2(n19847), .A(n14156), .ZN(P1_U2825) );
  OAI22_X1 U17448 ( .A1(n14393), .A2(n19912), .B1(n19919), .B2(n14157), .ZN(
        P1_U2841) );
  AOI22_X1 U17449 ( .A1(n14404), .A2(n19908), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14188), .ZN(n14158) );
  OAI21_X1 U17450 ( .B1(n14217), .B2(n9794), .A(n14158), .ZN(P1_U2843) );
  INV_X1 U17451 ( .A(n14300), .ZN(n14221) );
  INV_X1 U17452 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14159) );
  OAI222_X1 U17453 ( .A1(n9794), .A2(n14221), .B1(n14159), .B2(n19919), .C1(
        n14421), .C2(n19912), .ZN(P1_U2845) );
  OAI222_X1 U17454 ( .A1(n9794), .A2(n14228), .B1(n19919), .B2(n14161), .C1(
        n14441), .C2(n19912), .ZN(P1_U2847) );
  AOI22_X1 U17455 ( .A1(n14461), .A2(n19908), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n14188), .ZN(n14162) );
  OAI21_X1 U17456 ( .B1(n14325), .B2(n9794), .A(n14162), .ZN(P1_U2848) );
  INV_X1 U17457 ( .A(n14163), .ZN(n14164) );
  OAI21_X1 U17458 ( .B1(n14164), .B2(n9901), .A(n14233), .ZN(n15763) );
  OR2_X1 U17459 ( .A1(n9876), .A2(n14165), .ZN(n14166) );
  NAND2_X1 U17460 ( .A1(n15749), .A2(n14166), .ZN(n15762) );
  OAI22_X1 U17461 ( .A1(n15762), .A2(n19912), .B1(n15769), .B2(n19919), .ZN(
        n14167) );
  INV_X1 U17462 ( .A(n14167), .ZN(n14168) );
  OAI21_X1 U17463 ( .B1(n15763), .B2(n9794), .A(n14168), .ZN(P1_U2850) );
  OAI21_X1 U17464 ( .B1(n14175), .B2(n14169), .A(n14163), .ZN(n15774) );
  INV_X1 U17465 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14173) );
  INV_X1 U17466 ( .A(n14187), .ZN(n14171) );
  AOI21_X1 U17467 ( .B1(n14171), .B2(n14178), .A(n14170), .ZN(n14172) );
  OR2_X1 U17468 ( .A1(n14172), .A2(n9876), .ZN(n15706) );
  OAI222_X1 U17469 ( .A1(n9794), .A2(n15774), .B1(n14173), .B2(n19919), .C1(
        n15706), .C2(n19912), .ZN(P1_U2851) );
  INV_X1 U17470 ( .A(n14175), .ZN(n14176) );
  OAI21_X1 U17471 ( .B1(n14177), .B2(n14174), .A(n14176), .ZN(n15866) );
  INV_X1 U17472 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14179) );
  XNOR2_X1 U17473 ( .A(n14187), .B(n14178), .ZN(n15727) );
  INV_X1 U17474 ( .A(n15727), .ZN(n15778) );
  OAI222_X1 U17475 ( .A1(n9794), .A2(n15866), .B1(n19919), .B2(n14179), .C1(
        n19912), .C2(n15778), .ZN(P1_U2852) );
  INV_X1 U17476 ( .A(n14180), .ZN(n14182) );
  AND2_X1 U17477 ( .A1(n14182), .A2(n14181), .ZN(n14183) );
  OR2_X1 U17478 ( .A1(n14183), .A2(n14174), .ZN(n15787) );
  NAND2_X1 U17479 ( .A1(n14185), .A2(n14184), .ZN(n14186) );
  AND2_X1 U17480 ( .A1(n14187), .A2(n14186), .ZN(n15934) );
  AOI22_X1 U17481 ( .A1(n15934), .A2(n19908), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14188), .ZN(n14189) );
  OAI21_X1 U17482 ( .B1(n15787), .B2(n9794), .A(n14189), .ZN(P1_U2853) );
  XNOR2_X1 U17483 ( .A(n14191), .B(n14190), .ZN(n15797) );
  OAI22_X1 U17484 ( .A1(n15802), .A2(n19912), .B1(n15794), .B2(n19919), .ZN(
        n14192) );
  INV_X1 U17485 ( .A(n14192), .ZN(n14193) );
  OAI21_X1 U17486 ( .B1(n15797), .B2(n9794), .A(n14193), .ZN(P1_U2854) );
  INV_X1 U17487 ( .A(n15944), .ZN(n14195) );
  OAI222_X1 U17488 ( .A1(n14195), .A2(n19912), .B1(n19919), .B2(n14194), .C1(
        n15886), .C2(n9794), .ZN(P1_U2855) );
  AND2_X1 U17489 ( .A1(n14148), .A2(n14196), .ZN(n14197) );
  OR2_X1 U17490 ( .A1(n14197), .A2(n14133), .ZN(n15807) );
  OR2_X1 U17491 ( .A1(n14199), .A2(n14198), .ZN(n14200) );
  NAND2_X1 U17492 ( .A1(n14201), .A2(n14200), .ZN(n15952) );
  OAI22_X1 U17493 ( .A1(n15952), .A2(n19912), .B1(n15812), .B2(n19919), .ZN(
        n14202) );
  INV_X1 U17494 ( .A(n14202), .ZN(n14203) );
  OAI21_X1 U17495 ( .B1(n15807), .B2(n9794), .A(n14203), .ZN(P1_U2856) );
  OAI222_X1 U17496 ( .A1(n15958), .A2(n19912), .B1(n14204), .B2(n19919), .C1(
        n14270), .C2(n9794), .ZN(P1_U2857) );
  AOI21_X1 U17497 ( .B1(n14206), .B2(n13134), .A(n14147), .ZN(n15819) );
  OR2_X1 U17498 ( .A1(n14208), .A2(n14207), .ZN(n14209) );
  NAND2_X1 U17499 ( .A1(n9878), .A2(n14209), .ZN(n15814) );
  OAI22_X1 U17500 ( .A1(n15814), .A2(n19912), .B1(n15815), .B2(n19919), .ZN(
        n14210) );
  AOI21_X1 U17501 ( .B1(n15819), .B2(n19915), .A(n14210), .ZN(n14211) );
  INV_X1 U17502 ( .A(n14211), .ZN(P1_U2858) );
  OAI22_X1 U17503 ( .A1(n14262), .A2(n14213), .B1(n14271), .B2(n14212), .ZN(
        n14214) );
  AOI21_X1 U17504 ( .B1(n14264), .B2(BUF1_REG_29__SCAN_IN), .A(n14214), .ZN(
        n14216) );
  NAND2_X1 U17505 ( .A1(n14265), .A2(DATAI_29_), .ZN(n14215) );
  OAI211_X1 U17506 ( .C1(n14217), .C2(n14268), .A(n14216), .B(n14215), .ZN(
        P1_U2875) );
  INV_X1 U17507 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19156) );
  AOI22_X1 U17508 ( .A1(n14237), .A2(n19963), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n14235), .ZN(n14218) );
  OAI21_X1 U17509 ( .B1(n19156), .B2(n14239), .A(n14218), .ZN(n14219) );
  AOI21_X1 U17510 ( .B1(n14265), .B2(DATAI_27_), .A(n14219), .ZN(n14220) );
  OAI21_X1 U17511 ( .B1(n14221), .B2(n14268), .A(n14220), .ZN(P1_U2877) );
  OAI22_X1 U17512 ( .A1(n14262), .A2(n19960), .B1(n14271), .B2(n12144), .ZN(
        n14222) );
  AOI21_X1 U17513 ( .B1(n14264), .B2(BUF1_REG_26__SCAN_IN), .A(n14222), .ZN(
        n14224) );
  NAND2_X1 U17514 ( .A1(n14265), .A2(DATAI_26_), .ZN(n14223) );
  OAI211_X1 U17515 ( .C1(n14306), .C2(n14268), .A(n14224), .B(n14223), .ZN(
        P1_U2878) );
  INV_X1 U17516 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16317) );
  AOI22_X1 U17517 ( .A1(n14237), .A2(n19957), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n14235), .ZN(n14225) );
  OAI21_X1 U17518 ( .B1(n16317), .B2(n14239), .A(n14225), .ZN(n14226) );
  AOI21_X1 U17519 ( .B1(n14265), .B2(DATAI_25_), .A(n14226), .ZN(n14227) );
  OAI21_X1 U17520 ( .B1(n14228), .B2(n14268), .A(n14227), .ZN(P1_U2879) );
  OAI22_X1 U17521 ( .A1(n14262), .A2(n19954), .B1(n14271), .B2(n12129), .ZN(
        n14229) );
  AOI21_X1 U17522 ( .B1(n14264), .B2(BUF1_REG_24__SCAN_IN), .A(n14229), .ZN(
        n14231) );
  NAND2_X1 U17523 ( .A1(n14265), .A2(DATAI_24_), .ZN(n14230) );
  OAI211_X1 U17524 ( .C1(n14325), .C2(n14268), .A(n14231), .B(n14230), .ZN(
        P1_U2880) );
  AND2_X1 U17525 ( .A1(n14233), .A2(n14232), .ZN(n14234) );
  OR2_X1 U17526 ( .A1(n14234), .A2(n14122), .ZN(n15853) );
  INV_X1 U17527 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20970) );
  AOI22_X1 U17528 ( .A1(n14237), .A2(n14236), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n14235), .ZN(n14238) );
  OAI21_X1 U17529 ( .B1(n20970), .B2(n14239), .A(n14238), .ZN(n14240) );
  AOI21_X1 U17530 ( .B1(n14265), .B2(DATAI_23_), .A(n14240), .ZN(n14241) );
  OAI21_X1 U17531 ( .B1(n15853), .B2(n14268), .A(n14241), .ZN(P1_U2881) );
  OAI22_X1 U17532 ( .A1(n14262), .A2(n20087), .B1(n14271), .B2(n20884), .ZN(
        n14242) );
  AOI21_X1 U17533 ( .B1(n14264), .B2(BUF1_REG_22__SCAN_IN), .A(n14242), .ZN(
        n14244) );
  NAND2_X1 U17534 ( .A1(n14265), .A2(DATAI_22_), .ZN(n14243) );
  OAI211_X1 U17535 ( .C1(n15763), .C2(n14268), .A(n14244), .B(n14243), .ZN(
        P1_U2882) );
  OAI22_X1 U17536 ( .A1(n14262), .A2(n20084), .B1(n14271), .B2(n14245), .ZN(
        n14246) );
  AOI21_X1 U17537 ( .B1(n14264), .B2(BUF1_REG_21__SCAN_IN), .A(n14246), .ZN(
        n14248) );
  NAND2_X1 U17538 ( .A1(n14265), .A2(DATAI_21_), .ZN(n14247) );
  OAI211_X1 U17539 ( .C1(n15774), .C2(n14268), .A(n14248), .B(n14247), .ZN(
        P1_U2883) );
  OAI22_X1 U17540 ( .A1(n14262), .A2(n20080), .B1(n14271), .B2(n20828), .ZN(
        n14249) );
  AOI21_X1 U17541 ( .B1(n14264), .B2(BUF1_REG_20__SCAN_IN), .A(n14249), .ZN(
        n14251) );
  NAND2_X1 U17542 ( .A1(n14265), .A2(DATAI_20_), .ZN(n14250) );
  OAI211_X1 U17543 ( .C1(n15866), .C2(n14268), .A(n14251), .B(n14250), .ZN(
        P1_U2884) );
  OAI22_X1 U17544 ( .A1(n14262), .A2(n20076), .B1(n14271), .B2(n12136), .ZN(
        n14252) );
  AOI21_X1 U17545 ( .B1(n14264), .B2(BUF1_REG_19__SCAN_IN), .A(n14252), .ZN(
        n14254) );
  NAND2_X1 U17546 ( .A1(n14265), .A2(DATAI_19_), .ZN(n14253) );
  OAI211_X1 U17547 ( .C1(n15787), .C2(n14268), .A(n14254), .B(n14253), .ZN(
        P1_U2885) );
  OAI22_X1 U17548 ( .A1(n14262), .A2(n20071), .B1(n14271), .B2(n12146), .ZN(
        n14255) );
  AOI21_X1 U17549 ( .B1(n14264), .B2(BUF1_REG_18__SCAN_IN), .A(n14255), .ZN(
        n14257) );
  NAND2_X1 U17550 ( .A1(n14265), .A2(DATAI_18_), .ZN(n14256) );
  OAI211_X1 U17551 ( .C1(n15797), .C2(n14268), .A(n14257), .B(n14256), .ZN(
        P1_U2886) );
  OAI22_X1 U17552 ( .A1(n14262), .A2(n20067), .B1(n14271), .B2(n14258), .ZN(
        n14259) );
  AOI21_X1 U17553 ( .B1(n14264), .B2(BUF1_REG_17__SCAN_IN), .A(n14259), .ZN(
        n14261) );
  NAND2_X1 U17554 ( .A1(n14265), .A2(DATAI_17_), .ZN(n14260) );
  OAI211_X1 U17555 ( .C1(n15886), .C2(n14268), .A(n14261), .B(n14260), .ZN(
        P1_U2887) );
  OAI22_X1 U17556 ( .A1(n14262), .A2(n20058), .B1(n14271), .B2(n12138), .ZN(
        n14263) );
  AOI21_X1 U17557 ( .B1(n14264), .B2(BUF1_REG_16__SCAN_IN), .A(n14263), .ZN(
        n14267) );
  NAND2_X1 U17558 ( .A1(n14265), .A2(DATAI_16_), .ZN(n14266) );
  OAI211_X1 U17559 ( .C1(n15807), .C2(n14268), .A(n14267), .B(n14266), .ZN(
        P1_U2888) );
  OAI222_X1 U17560 ( .A1(n14268), .A2(n14270), .B1(n14273), .B2(n14269), .C1(
        n14271), .C2(n19926), .ZN(P1_U2889) );
  INV_X1 U17561 ( .A(n15819), .ZN(n14274) );
  INV_X1 U17562 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14272) );
  OAI222_X1 U17563 ( .A1(n14268), .A2(n14274), .B1(n19967), .B2(n14273), .C1(
        n14272), .C2(n14271), .ZN(P1_U2890) );
  XNOR2_X1 U17564 ( .A(n14275), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14409) );
  NOR2_X1 U17565 ( .A1(n20002), .A2(n20690), .ZN(n14403) );
  AOI21_X1 U17566 ( .B1(n19987), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14403), .ZN(n14276) );
  OAI21_X1 U17567 ( .B1(n14277), .B2(n19998), .A(n14276), .ZN(n14278) );
  AOI21_X1 U17568 ( .B1(n14279), .B2(n19993), .A(n14278), .ZN(n14280) );
  OAI21_X1 U17569 ( .B1(n19817), .B2(n14409), .A(n14280), .ZN(P1_U2970) );
  NAND2_X1 U17570 ( .A1(n11179), .A2(n14281), .ZN(n14302) );
  NAND2_X1 U17571 ( .A1(n15855), .A2(n14302), .ZN(n14285) );
  OAI21_X1 U17572 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14282), .A(
        n14285), .ZN(n14284) );
  INV_X1 U17573 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14426) );
  MUX2_X1 U17574 ( .A(n14426), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n11179), .Z(n14283) );
  OAI211_X1 U17575 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14285), .A(
        n14284), .B(n14283), .ZN(n14287) );
  XNOR2_X1 U17576 ( .A(n14287), .B(n14286), .ZN(n14419) );
  NAND2_X1 U17577 ( .A1(n20033), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14413) );
  OAI21_X1 U17578 ( .B1(n15871), .B2(n14288), .A(n14413), .ZN(n14291) );
  NOR2_X1 U17579 ( .A1(n14289), .A2(n20044), .ZN(n14290) );
  OAI21_X1 U17580 ( .B1(n19817), .B2(n14419), .A(n14293), .ZN(P1_U2971) );
  MUX2_X1 U17581 ( .A(n14295), .B(n14294), .S(n11189), .Z(n14296) );
  XNOR2_X1 U17582 ( .A(n14296), .B(n14426), .ZN(n14429) );
  NAND2_X1 U17583 ( .A1(n20033), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14420) );
  NAND2_X1 U17584 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14297) );
  OAI211_X1 U17585 ( .C1(n14298), .C2(n19998), .A(n14420), .B(n14297), .ZN(
        n14299) );
  AOI21_X1 U17586 ( .B1(n14300), .B2(n19993), .A(n14299), .ZN(n14301) );
  OAI21_X1 U17587 ( .B1(n19817), .B2(n14429), .A(n14301), .ZN(P1_U2972) );
  OAI211_X1 U17588 ( .C1(n11189), .C2(n15855), .A(n14303), .B(n14302), .ZN(
        n14304) );
  XNOR2_X1 U17589 ( .A(n14304), .B(n14430), .ZN(n14438) );
  NAND2_X1 U17590 ( .A1(n20033), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14432) );
  OAI21_X1 U17591 ( .B1(n15871), .B2(n14305), .A(n14432), .ZN(n14308) );
  NOR2_X1 U17592 ( .A1(n14306), .A2(n20044), .ZN(n14307) );
  OAI21_X1 U17593 ( .B1(n19817), .B2(n14438), .A(n14310), .ZN(P1_U2973) );
  INV_X1 U17594 ( .A(n15855), .ZN(n14311) );
  NAND3_X1 U17595 ( .A1(n14311), .A2(n21047), .A3(n14457), .ZN(n14314) );
  NAND2_X1 U17596 ( .A1(n14321), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14313) );
  MUX2_X1 U17597 ( .A(n14314), .B(n14313), .S(n11179), .Z(n14315) );
  XNOR2_X1 U17598 ( .A(n14315), .B(n20954), .ZN(n14446) );
  NAND2_X1 U17599 ( .A1(n20033), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14440) );
  NAND2_X1 U17600 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14316) );
  OAI211_X1 U17601 ( .C1(n14317), .C2(n19998), .A(n14440), .B(n14316), .ZN(
        n14318) );
  AOI21_X1 U17602 ( .B1(n14319), .B2(n19993), .A(n14318), .ZN(n14320) );
  OAI21_X1 U17603 ( .B1(n19817), .B2(n14446), .A(n14320), .ZN(P1_U2974) );
  NOR2_X1 U17604 ( .A1(n14321), .A2(n15855), .ZN(n14322) );
  MUX2_X1 U17605 ( .A(n14322), .B(n14321), .S(n11179), .Z(n14323) );
  XNOR2_X1 U17606 ( .A(n14323), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14463) );
  NAND2_X1 U17607 ( .A1(n20033), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14449) );
  OAI21_X1 U17608 ( .B1(n15871), .B2(n14324), .A(n14449), .ZN(n14327) );
  NOR2_X1 U17609 ( .A1(n14325), .A2(n20044), .ZN(n14326) );
  AOI211_X1 U17610 ( .C1(n15899), .C2(n14328), .A(n14327), .B(n14326), .ZN(
        n14329) );
  OAI21_X1 U17611 ( .B1(n19817), .B2(n14463), .A(n14329), .ZN(P1_U2975) );
  NAND2_X1 U17612 ( .A1(n14331), .A2(n14330), .ZN(n14332) );
  XNOR2_X1 U17613 ( .A(n14332), .B(n14447), .ZN(n14476) );
  NAND2_X1 U17614 ( .A1(n20033), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14471) );
  OAI21_X1 U17615 ( .B1(n15871), .B2(n10926), .A(n14471), .ZN(n14334) );
  NOR2_X1 U17616 ( .A1(n15763), .A2(n20044), .ZN(n14333) );
  AOI211_X1 U17617 ( .C1(n15899), .C2(n15766), .A(n14334), .B(n14333), .ZN(
        n14335) );
  OAI21_X1 U17618 ( .B1(n19817), .B2(n14476), .A(n14335), .ZN(P1_U2977) );
  OAI22_X1 U17619 ( .A1(n15871), .A2(n14336), .B1(n20002), .B2(n20671), .ZN(
        n14338) );
  NOR2_X1 U17620 ( .A1(n15797), .A2(n20044), .ZN(n14337) );
  AOI211_X1 U17621 ( .C1(n15899), .C2(n15798), .A(n14338), .B(n14337), .ZN(
        n14339) );
  OAI21_X1 U17622 ( .B1(n19817), .B2(n14340), .A(n14339), .ZN(P1_U2981) );
  NAND2_X1 U17623 ( .A1(n14341), .A2(n14342), .ZN(n14363) );
  INV_X1 U17624 ( .A(n14343), .ZN(n14344) );
  NAND2_X1 U17625 ( .A1(n14363), .A2(n14344), .ZN(n14347) );
  INV_X1 U17626 ( .A(n14345), .ZN(n14346) );
  NAND2_X1 U17627 ( .A1(n14347), .A2(n14346), .ZN(n15892) );
  NOR2_X1 U17628 ( .A1(n11179), .A2(n15961), .ZN(n14348) );
  NAND2_X1 U17629 ( .A1(n15880), .A2(n14349), .ZN(n14350) );
  NAND2_X1 U17630 ( .A1(n14350), .A2(n14352), .ZN(n14354) );
  AND2_X1 U17631 ( .A1(n11179), .A2(n15961), .ZN(n14351) );
  NOR2_X1 U17632 ( .A1(n14352), .A2(n14351), .ZN(n14353) );
  NAND2_X1 U17633 ( .A1(n15880), .A2(n14353), .ZN(n15881) );
  NAND2_X1 U17634 ( .A1(n15954), .A2(n19994), .ZN(n14359) );
  INV_X1 U17635 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14355) );
  OAI22_X1 U17636 ( .A1(n15871), .A2(n14356), .B1(n20002), .B2(n14355), .ZN(
        n14357) );
  AOI21_X1 U17637 ( .B1(n15809), .B2(n15899), .A(n14357), .ZN(n14358) );
  OAI211_X1 U17638 ( .C1(n20044), .C2(n15807), .A(n14359), .B(n14358), .ZN(
        P1_U2983) );
  INV_X1 U17639 ( .A(n14360), .ZN(n14361) );
  AOI21_X1 U17640 ( .B1(n14363), .B2(n14362), .A(n14361), .ZN(n14365) );
  XNOR2_X1 U17641 ( .A(n11179), .B(n20982), .ZN(n14364) );
  XNOR2_X1 U17642 ( .A(n14365), .B(n14364), .ZN(n14486) );
  INV_X1 U17643 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14366) );
  NOR2_X1 U17644 ( .A1(n20002), .A2(n14366), .ZN(n14483) );
  AOI21_X1 U17645 ( .B1(n19987), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n14483), .ZN(n14367) );
  OAI21_X1 U17646 ( .B1(n19998), .B2(n15817), .A(n14367), .ZN(n14368) );
  AOI21_X1 U17647 ( .B1(n15819), .B2(n19993), .A(n14368), .ZN(n14369) );
  OAI21_X1 U17648 ( .B1(n14486), .B2(n19817), .A(n14369), .ZN(P1_U2985) );
  INV_X1 U17649 ( .A(n14341), .ZN(n15903) );
  INV_X1 U17650 ( .A(n14370), .ZN(n14371) );
  AOI22_X1 U17651 ( .A1(n15903), .A2(n14372), .B1(n11189), .B2(n14371), .ZN(
        n14496) );
  INV_X1 U17652 ( .A(n14374), .ZN(n14373) );
  AOI21_X1 U17653 ( .B1(n11189), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14373), .ZN(n14495) );
  NAND2_X1 U17654 ( .A1(n14496), .A2(n14495), .ZN(n14494) );
  NAND2_X1 U17655 ( .A1(n14494), .A2(n14374), .ZN(n14376) );
  XNOR2_X1 U17656 ( .A(n14376), .B(n14375), .ZN(n15975) );
  AOI22_X1 U17657 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20033), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14377) );
  OAI21_X1 U17658 ( .B1(n19998), .B2(n14378), .A(n14377), .ZN(n14379) );
  AOI21_X1 U17659 ( .B1(n14380), .B2(n19993), .A(n14379), .ZN(n14381) );
  OAI21_X1 U17660 ( .B1(n15975), .B2(n19817), .A(n14381), .ZN(P1_U2986) );
  NAND2_X1 U17661 ( .A1(n14382), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14384) );
  XNOR2_X1 U17662 ( .A(n14341), .B(n14385), .ZN(n14383) );
  MUX2_X1 U17663 ( .A(n14384), .B(n14383), .S(n11179), .Z(n14387) );
  INV_X1 U17664 ( .A(n14382), .ZN(n14386) );
  NAND3_X1 U17665 ( .A1(n14386), .A2(n11189), .A3(n14385), .ZN(n15904) );
  NAND2_X1 U17666 ( .A1(n14387), .A2(n15904), .ZN(n15997) );
  NAND2_X1 U17667 ( .A1(n15997), .A2(n19994), .ZN(n14392) );
  INV_X1 U17668 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14388) );
  OAI22_X1 U17669 ( .A1(n15871), .A2(n14389), .B1(n20002), .B2(n14388), .ZN(
        n14390) );
  AOI21_X1 U17670 ( .B1(n15847), .B2(n15899), .A(n14390), .ZN(n14391) );
  OAI211_X1 U17671 ( .C1(n20044), .C2(n15845), .A(n14392), .B(n14391), .ZN(
        P1_U2989) );
  AND3_X1 U17672 ( .A1(n14394), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16012), .ZN(n14399) );
  NOR3_X1 U17673 ( .A1(n14396), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14395), .ZN(n14397) );
  NOR3_X1 U17674 ( .A1(n14410), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14401), .ZN(n14402) );
  AOI211_X1 U17675 ( .C1(n14404), .C2(n20027), .A(n14403), .B(n14402), .ZN(
        n14408) );
  INV_X1 U17676 ( .A(n14405), .ZN(n14406) );
  NAND2_X1 U17677 ( .A1(n14406), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14407) );
  OAI211_X1 U17678 ( .C1(n14409), .C2(n15966), .A(n14408), .B(n14407), .ZN(
        P1_U3002) );
  INV_X1 U17679 ( .A(n14410), .ZN(n14427) );
  NOR2_X1 U17680 ( .A1(n14412), .A2(n14411), .ZN(n14417) );
  AND3_X1 U17681 ( .A1(n14436), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16012), .ZN(n14416) );
  OAI21_X1 U17682 ( .B1(n14414), .B2(n20003), .A(n14413), .ZN(n14415) );
  AOI211_X1 U17683 ( .C1(n14427), .C2(n14417), .A(n14416), .B(n14415), .ZN(
        n14418) );
  OAI21_X1 U17684 ( .B1(n14419), .B2(n15966), .A(n14418), .ZN(P1_U3003) );
  OAI21_X1 U17685 ( .B1(n14421), .B2(n20003), .A(n14420), .ZN(n14425) );
  INV_X1 U17686 ( .A(n14436), .ZN(n14423) );
  NOR3_X1 U17687 ( .A1(n14423), .A2(n14422), .A3(n14426), .ZN(n14424) );
  AOI211_X1 U17688 ( .C1(n14427), .C2(n14426), .A(n14425), .B(n14424), .ZN(
        n14428) );
  OAI21_X1 U17689 ( .B1(n14429), .B2(n15966), .A(n14428), .ZN(P1_U3004) );
  INV_X1 U17690 ( .A(n14444), .ZN(n14431) );
  OAI21_X1 U17691 ( .B1(n14431), .B2(n20954), .A(n14430), .ZN(n14435) );
  OAI21_X1 U17692 ( .B1(n14433), .B2(n20003), .A(n14432), .ZN(n14434) );
  AOI21_X1 U17693 ( .B1(n14436), .B2(n14435), .A(n14434), .ZN(n14437) );
  OAI21_X1 U17694 ( .B1(n14438), .B2(n15966), .A(n14437), .ZN(P1_U3005) );
  NOR2_X1 U17695 ( .A1(n14439), .A2(n20954), .ZN(n14443) );
  OAI21_X1 U17696 ( .B1(n14441), .B2(n20003), .A(n14440), .ZN(n14442) );
  AOI211_X1 U17697 ( .C1(n14444), .C2(n20954), .A(n14443), .B(n14442), .ZN(
        n14445) );
  OAI21_X1 U17698 ( .B1(n14446), .B2(n15966), .A(n14445), .ZN(P1_U3006) );
  NOR4_X1 U17699 ( .A1(n14451), .A2(n21047), .A3(n14447), .A4(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14448) );
  NAND2_X1 U17700 ( .A1(n14453), .A2(n14448), .ZN(n14450) );
  OAI21_X1 U17701 ( .B1(n15942), .B2(n14450), .A(n14449), .ZN(n14460) );
  INV_X1 U17702 ( .A(n14451), .ZN(n14452) );
  NAND4_X1 U17703 ( .A1(n14453), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14452), .A4(n21047), .ZN(n14454) );
  NOR2_X1 U17704 ( .A1(n14455), .A2(n14454), .ZN(n15926) );
  AOI21_X1 U17705 ( .B1(n14487), .B2(n15926), .A(n14456), .ZN(n14458) );
  NOR2_X1 U17706 ( .A1(n14458), .A2(n14457), .ZN(n14459) );
  AOI211_X1 U17707 ( .C1(n20027), .C2(n14461), .A(n14460), .B(n14459), .ZN(
        n14462) );
  OAI21_X1 U17708 ( .B1(n14463), .B2(n15966), .A(n14462), .ZN(P1_U3007) );
  NAND2_X1 U17709 ( .A1(n15990), .A2(n14477), .ZN(n15968) );
  NOR3_X1 U17710 ( .A1(n20023), .A2(n14464), .A3(n15968), .ZN(n14465) );
  AOI21_X1 U17711 ( .B1(n14466), .B2(n14491), .A(n14465), .ZN(n14480) );
  NOR2_X1 U17712 ( .A1(n14480), .A2(n14467), .ZN(n15937) );
  INV_X1 U17713 ( .A(n15937), .ZN(n15728) );
  OAI21_X1 U17714 ( .B1(n15969), .B2(n14468), .A(n15728), .ZN(n15731) );
  NAND2_X1 U17715 ( .A1(n14469), .A2(n15731), .ZN(n15709) );
  AOI21_X1 U17716 ( .B1(n11186), .B2(n14447), .A(n15709), .ZN(n14473) );
  NAND2_X1 U17717 ( .A1(n15703), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14470) );
  OAI211_X1 U17718 ( .C1(n15762), .C2(n20003), .A(n14471), .B(n14470), .ZN(
        n14472) );
  AOI21_X1 U17719 ( .B1(n14474), .B2(n14473), .A(n14472), .ZN(n14475) );
  OAI21_X1 U17720 ( .B1(n14476), .B2(n15966), .A(n14475), .ZN(P1_U3009) );
  INV_X1 U17721 ( .A(n15814), .ZN(n14484) );
  OAI22_X1 U17722 ( .A1(n14477), .A2(n20024), .B1(n15970), .B2(n15969), .ZN(
        n14478) );
  AOI211_X1 U17723 ( .C1(n14479), .C2(n15968), .A(n15992), .B(n14478), .ZN(
        n15981) );
  NOR2_X1 U17724 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14480), .ZN(
        n15971) );
  NOR2_X1 U17725 ( .A1(n20982), .A2(n15971), .ZN(n14481) );
  AOI22_X1 U17726 ( .A1(n15942), .A2(n20982), .B1(n15981), .B2(n14481), .ZN(
        n14482) );
  AOI211_X1 U17727 ( .C1(n20027), .C2(n14484), .A(n14483), .B(n14482), .ZN(
        n14485) );
  OAI21_X1 U17728 ( .B1(n14486), .B2(n15966), .A(n14485), .ZN(P1_U3017) );
  INV_X1 U17729 ( .A(n14487), .ZN(n14492) );
  NAND2_X1 U17730 ( .A1(n15988), .A2(n14488), .ZN(n15983) );
  AOI21_X1 U17731 ( .B1(n15990), .B2(n14488), .A(n20001), .ZN(n14489) );
  AOI211_X1 U17732 ( .C1(n14491), .C2(n14490), .A(n14489), .B(n15992), .ZN(
        n15989) );
  OAI21_X1 U17733 ( .B1(n14492), .B2(n15983), .A(n15989), .ZN(n14500) );
  NAND2_X1 U17734 ( .A1(n14493), .A2(n16014), .ZN(n14498) );
  OAI21_X1 U17735 ( .B1(n14496), .B2(n14495), .A(n14494), .ZN(n14497) );
  INV_X1 U17736 ( .A(n14497), .ZN(n15902) );
  OAI22_X1 U17737 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14498), .B1(
        n15902), .B2(n15966), .ZN(n14499) );
  AOI21_X1 U17738 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14500), .A(
        n14499), .ZN(n14502) );
  NAND2_X1 U17739 ( .A1(n19986), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14501) );
  OAI211_X1 U17740 ( .C1(n20003), .C2(n15825), .A(n14502), .B(n14501), .ZN(
        P1_U3019) );
  NAND3_X1 U17741 ( .A1(n14503), .A2(n12276), .A3(n20031), .ZN(n14514) );
  INV_X1 U17742 ( .A(n14504), .ZN(n14510) );
  INV_X1 U17743 ( .A(n14505), .ZN(n14509) );
  AOI21_X1 U17744 ( .B1(n14507), .B2(n14506), .A(n20022), .ZN(n14508) );
  AOI211_X1 U17745 ( .C1(n20027), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        n14513) );
  NAND3_X1 U17746 ( .A1(n14511), .A2(n20022), .A3(n20034), .ZN(n14512) );
  NAND3_X1 U17747 ( .A1(n14514), .A2(n14513), .A3(n14512), .ZN(P1_U3030) );
  INV_X1 U17748 ( .A(n14515), .ZN(n14518) );
  INV_X1 U17749 ( .A(n14516), .ZN(n14517) );
  NAND2_X1 U17750 ( .A1(n14518), .A2(n14517), .ZN(n14524) );
  INV_X1 U17751 ( .A(n12799), .ZN(n20517) );
  INV_X1 U17752 ( .A(n15669), .ZN(n14519) );
  OAI22_X1 U17753 ( .A1(n14519), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n14524), .B2(n15667), .ZN(n14520) );
  AOI21_X1 U17754 ( .B1(n20517), .B2(n14521), .A(n14520), .ZN(n15671) );
  INV_X1 U17755 ( .A(n20708), .ZN(n14522) );
  OAI222_X1 U17756 ( .A1(n14524), .A2(n20706), .B1(n20714), .B2(n15671), .C1(
        n14523), .C2(n14522), .ZN(n14525) );
  MUX2_X1 U17757 ( .A(n14525), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n20711), .Z(P1_U3473) );
  AOI22_X1 U17758 ( .A1(n11907), .A2(n19574), .B1(n19681), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14528) );
  INV_X1 U17759 ( .A(n14526), .ZN(n16221) );
  OAI21_X1 U17760 ( .B1(n19680), .B2(n19390), .A(n16221), .ZN(n14527) );
  OAI21_X1 U17761 ( .B1(n14528), .B2(n11897), .A(n14527), .ZN(n14532) );
  AOI22_X1 U17762 ( .A1(n19097), .A2(n15735), .B1(n19616), .B2(n14529), .ZN(
        n14530) );
  NAND2_X1 U17763 ( .A1(n14530), .A2(n18730), .ZN(n14531) );
  MUX2_X1 U17764 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n14532), .S(n14531), 
        .Z(P2_U3610) );
  NAND2_X1 U17765 ( .A1(n18916), .A2(n18912), .ZN(n18800) );
  INV_X1 U17766 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16060) );
  INV_X1 U17767 ( .A(n14534), .ZN(n14533) );
  AOI21_X1 U17768 ( .B1(n16060), .B2(n14533), .A(n14561), .ZN(n16059) );
  INV_X1 U17769 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14536) );
  INV_X1 U17770 ( .A(n14538), .ZN(n14535) );
  AOI21_X1 U17771 ( .B1(n14536), .B2(n14535), .A(n14534), .ZN(n14862) );
  AND2_X1 U17772 ( .A1(n14541), .A2(n14868), .ZN(n14537) );
  NOR2_X1 U17773 ( .A1(n14538), .A2(n14537), .ZN(n14871) );
  INV_X1 U17774 ( .A(n14871), .ZN(n14580) );
  NAND2_X1 U17775 ( .A1(n14542), .A2(n14539), .ZN(n14540) );
  NAND2_X1 U17776 ( .A1(n14541), .A2(n14540), .ZN(n16073) );
  INV_X1 U17777 ( .A(n14542), .ZN(n14543) );
  AOI21_X1 U17778 ( .B1(n14887), .B2(n14560), .A(n14543), .ZN(n16084) );
  AOI21_X1 U17779 ( .B1(n14906), .B2(n14557), .A(n9897), .ZN(n14908) );
  INV_X1 U17780 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14940) );
  AOI21_X1 U17781 ( .B1(n14556), .B2(n14940), .A(n14558), .ZN(n14942) );
  AOI21_X1 U17782 ( .B1(n14965), .B2(n14554), .A(n9896), .ZN(n18768) );
  INV_X1 U17783 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18793) );
  AOI21_X1 U17784 ( .B1(n14552), .B2(n18793), .A(n14555), .ZN(n18803) );
  AOI21_X1 U17785 ( .B1(n18812), .B2(n14550), .A(n14551), .ZN(n18810) );
  AOI21_X1 U17786 ( .B1(n16138), .B2(n14548), .A(n9871), .ZN(n18841) );
  AOI21_X1 U17787 ( .B1(n16153), .B2(n14546), .A(n14549), .ZN(n16146) );
  AOI21_X1 U17788 ( .B1(n18869), .B2(n14544), .A(n14547), .ZN(n18875) );
  NAND2_X1 U17789 ( .A1(n14545), .A2(n16170), .ZN(n18873) );
  NOR2_X1 U17790 ( .A1(n18875), .A2(n18873), .ZN(n18857) );
  OAI21_X1 U17791 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n14547), .A(
        n14546), .ZN(n18859) );
  NAND2_X1 U17792 ( .A1(n18857), .A2(n18859), .ZN(n14676) );
  NOR2_X1 U17793 ( .A1(n16146), .A2(n14676), .ZN(n14675) );
  OAI21_X1 U17794 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n14549), .A(
        n14548), .ZN(n18852) );
  NAND2_X1 U17795 ( .A1(n14675), .A2(n18852), .ZN(n18833) );
  NOR2_X1 U17796 ( .A1(n18841), .A2(n18833), .ZN(n18821) );
  OAI21_X1 U17797 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9871), .A(
        n14550), .ZN(n18822) );
  NAND2_X1 U17798 ( .A1(n18821), .A2(n18822), .ZN(n18808) );
  NOR2_X1 U17799 ( .A1(n18810), .A2(n18808), .ZN(n14660) );
  OR2_X1 U17800 ( .A1(n14551), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14553) );
  NAND2_X1 U17801 ( .A1(n14553), .A2(n14552), .ZN(n15000) );
  NAND2_X1 U17802 ( .A1(n14660), .A2(n15000), .ZN(n18802) );
  NOR2_X1 U17803 ( .A1(n18803), .A2(n18802), .ZN(n18801) );
  OAI21_X1 U17804 ( .B1(n14555), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14554), .ZN(n18779) );
  NAND2_X1 U17805 ( .A1(n18801), .A2(n18779), .ZN(n18766) );
  NOR2_X1 U17806 ( .A1(n18768), .A2(n18766), .ZN(n18758) );
  OAI21_X1 U17807 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9896), .A(
        n14556), .ZN(n18757) );
  NAND2_X1 U17808 ( .A1(n18758), .A2(n18757), .ZN(n14641) );
  NOR2_X1 U17809 ( .A1(n14942), .A2(n14641), .ZN(n14633) );
  OAI21_X1 U17810 ( .B1(n14558), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14557), .ZN(n14920) );
  NAND2_X1 U17811 ( .A1(n14633), .A2(n14920), .ZN(n14611) );
  NOR2_X1 U17812 ( .A1(n14908), .A2(n14611), .ZN(n14595) );
  OR2_X1 U17813 ( .A1(n9897), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14559) );
  AND2_X1 U17814 ( .A1(n14560), .A2(n14559), .ZN(n14598) );
  INV_X1 U17815 ( .A(n14598), .ZN(n14899) );
  AOI21_X1 U17816 ( .B1(n14595), .B2(n14899), .A(n18941), .ZN(n16083) );
  NOR2_X1 U17817 ( .A1(n16084), .A2(n16083), .ZN(n16082) );
  OR2_X1 U17818 ( .A1(n18941), .A2(n16082), .ZN(n16072) );
  NAND2_X1 U17819 ( .A1(n16073), .A2(n16072), .ZN(n16071) );
  NAND2_X1 U17820 ( .A1(n18912), .A2(n16071), .ZN(n14579) );
  OAI21_X1 U17821 ( .B1(n18941), .B2(n14580), .A(n14579), .ZN(n14568) );
  NOR2_X1 U17822 ( .A1(n14862), .A2(n14568), .ZN(n14567) );
  NOR2_X1 U17823 ( .A1(n18941), .A2(n14567), .ZN(n16058) );
  AOI21_X1 U17824 ( .B1(n16059), .B2(n18912), .A(n16058), .ZN(n16051) );
  XNOR2_X1 U17825 ( .A(n14561), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16050) );
  NAND2_X1 U17826 ( .A1(n16051), .A2(n16050), .ZN(n16049) );
  AOI22_X1 U17827 ( .A1(n18950), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n18949), .ZN(n14562) );
  OAI21_X1 U17828 ( .B1(n18800), .B2(n16049), .A(n14562), .ZN(n14563) );
  AOI21_X1 U17829 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18928), .A(
        n14563), .ZN(n14566) );
  AOI22_X1 U17830 ( .A1(n19001), .A2(n18952), .B1(n14564), .B2(n18954), .ZN(
        n14565) );
  OAI211_X1 U17831 ( .C1(n16094), .C2(n18957), .A(n14566), .B(n14565), .ZN(
        P2_U2824) );
  AOI211_X1 U17832 ( .C1(n14568), .C2(n14862), .A(n18967), .B(n14567), .ZN(
        n14569) );
  INV_X1 U17833 ( .A(n14569), .ZN(n14578) );
  INV_X1 U17834 ( .A(n18949), .ZN(n18926) );
  OAI22_X1 U17835 ( .A1(n14536), .A2(n18961), .B1(n19737), .B2(n18926), .ZN(
        n14575) );
  NOR2_X1 U17836 ( .A1(n14586), .A2(n14570), .ZN(n14571) );
  NOR2_X1 U17837 ( .A1(n14736), .A2(n14571), .ZN(n15067) );
  INV_X1 U17838 ( .A(n15067), .ZN(n14573) );
  INV_X1 U17839 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n14572) );
  OAI22_X1 U17840 ( .A1(n14573), .A2(n18920), .B1(n14572), .B2(n18925), .ZN(
        n14574) );
  AOI211_X1 U17841 ( .C1(n18954), .C2(n14576), .A(n14575), .B(n14574), .ZN(
        n14577) );
  OAI211_X1 U17842 ( .C1(n18957), .C2(n15065), .A(n14578), .B(n14577), .ZN(
        P2_U2827) );
  INV_X1 U17843 ( .A(n14579), .ZN(n14581) );
  AOI221_X1 U17844 ( .B1(n14871), .B2(n14581), .C1(n14580), .C2(n14579), .A(
        n18967), .ZN(n14582) );
  INV_X1 U17845 ( .A(n14582), .ZN(n14593) );
  INV_X1 U17846 ( .A(n14583), .ZN(n14591) );
  NOR2_X1 U17847 ( .A1(n14759), .A2(n14584), .ZN(n14585) );
  NOR2_X1 U17848 ( .A1(n14586), .A2(n14585), .ZN(n15075) );
  NAND2_X1 U17849 ( .A1(n15075), .A2(n18952), .ZN(n14588) );
  AOI22_X1 U17850 ( .A1(n18949), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18928), .ZN(n14587) );
  OAI211_X1 U17851 ( .C1(n14589), .C2(n18925), .A(n14588), .B(n14587), .ZN(
        n14590) );
  AOI21_X1 U17852 ( .B1(n14591), .B2(n18954), .A(n14590), .ZN(n14592) );
  OAI211_X1 U17853 ( .C1(n18957), .C2(n15078), .A(n14593), .B(n14592), .ZN(
        P2_U2828) );
  XNOR2_X1 U17854 ( .A(n14594), .B(P2_EBX_REG_24__SCAN_IN), .ZN(n14610) );
  NOR2_X1 U17855 ( .A1(n18941), .A2(n14595), .ZN(n14597) );
  OAI21_X1 U17856 ( .B1(n14598), .B2(n14597), .A(n18916), .ZN(n14596) );
  AOI21_X1 U17857 ( .B1(n14598), .B2(n14597), .A(n14596), .ZN(n14599) );
  INV_X1 U17858 ( .A(n14599), .ZN(n14609) );
  INV_X1 U17859 ( .A(n14897), .ZN(n15116) );
  INV_X1 U17860 ( .A(n14600), .ZN(n14770) );
  INV_X1 U17861 ( .A(n14601), .ZN(n14622) );
  INV_X1 U17862 ( .A(n14602), .ZN(n14603) );
  NAND2_X1 U17863 ( .A1(n14622), .A2(n14603), .ZN(n14604) );
  NAND2_X1 U17864 ( .A1(n14770), .A2(n14604), .ZN(n15114) );
  AOI22_X1 U17865 ( .A1(n18949), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18928), .ZN(n14606) );
  NAND2_X1 U17866 ( .A1(n18950), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n14605) );
  OAI211_X1 U17867 ( .C1(n15114), .C2(n18920), .A(n14606), .B(n14605), .ZN(
        n14607) );
  AOI21_X1 U17868 ( .B1(n15116), .B2(n18939), .A(n14607), .ZN(n14608) );
  OAI211_X1 U17869 ( .C1(n14610), .C2(n18907), .A(n14609), .B(n14608), .ZN(
        P2_U2831) );
  NAND2_X1 U17870 ( .A1(n18912), .A2(n14611), .ZN(n14612) );
  XNOR2_X1 U17871 ( .A(n14908), .B(n14612), .ZN(n14613) );
  AOI22_X1 U17872 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18928), .B1(
        n18916), .B2(n14613), .ZN(n14626) );
  NOR2_X1 U17873 ( .A1(n14614), .A2(n14615), .ZN(n14616) );
  OR2_X1 U17874 ( .A1(n14617), .A2(n14616), .ZN(n15126) );
  INV_X1 U17875 ( .A(n15126), .ZN(n16095) );
  INV_X1 U17876 ( .A(n14618), .ZN(n14630) );
  INV_X1 U17877 ( .A(n14619), .ZN(n14620) );
  NAND2_X1 U17878 ( .A1(n14630), .A2(n14620), .ZN(n14621) );
  NAND2_X1 U17879 ( .A1(n14622), .A2(n14621), .ZN(n15131) );
  AOI22_X1 U17880 ( .A1(n18950), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18949), .ZN(n14623) );
  OAI21_X1 U17881 ( .B1(n15131), .B2(n18920), .A(n14623), .ZN(n14624) );
  AOI21_X1 U17882 ( .B1(n16095), .B2(n18939), .A(n14624), .ZN(n14625) );
  OAI211_X1 U17883 ( .C1(n14627), .C2(n18907), .A(n14626), .B(n14625), .ZN(
        P2_U2832) );
  AND2_X1 U17884 ( .A1(n14648), .A2(n14628), .ZN(n14629) );
  OR2_X1 U17885 ( .A1(n14629), .A2(n14614), .ZN(n16101) );
  OAI21_X1 U17886 ( .B1(n14652), .B2(n14631), .A(n14630), .ZN(n15139) );
  INV_X1 U17887 ( .A(n15139), .ZN(n14797) );
  AOI22_X1 U17888 ( .A1(n14797), .A2(n18952), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18928), .ZN(n14632) );
  OAI21_X1 U17889 ( .B1(n16101), .B2(n18957), .A(n14632), .ZN(n14638) );
  NOR2_X1 U17890 ( .A1(n18941), .A2(n14633), .ZN(n14634) );
  XOR2_X1 U17891 ( .A(n14920), .B(n14634), .Z(n14636) );
  AOI22_X1 U17892 ( .A1(n18950), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18949), .ZN(n14635) );
  OAI21_X1 U17893 ( .B1(n18967), .B2(n14636), .A(n14635), .ZN(n14637) );
  AOI211_X1 U17894 ( .C1(n18954), .C2(n14639), .A(n14638), .B(n14637), .ZN(
        n14640) );
  INV_X1 U17895 ( .A(n14640), .ZN(P2_U2833) );
  AND2_X1 U17896 ( .A1(n18912), .A2(n14641), .ZN(n14643) );
  OAI21_X1 U17897 ( .B1(n14942), .B2(n14643), .A(n18916), .ZN(n14642) );
  AOI21_X1 U17898 ( .B1(n14643), .B2(n14942), .A(n14642), .ZN(n14659) );
  NOR2_X1 U17899 ( .A1(n14644), .A2(n18907), .ZN(n14658) );
  NAND2_X1 U17900 ( .A1(n14646), .A2(n14645), .ZN(n14647) );
  NAND2_X1 U17901 ( .A1(n14648), .A2(n14647), .ZN(n15153) );
  NOR2_X1 U17902 ( .A1(n14649), .A2(n14650), .ZN(n14651) );
  NOR2_X1 U17903 ( .A1(n14652), .A2(n14651), .ZN(n15150) );
  OAI22_X1 U17904 ( .A1(n14940), .A2(n18961), .B1(n19723), .B2(n18926), .ZN(
        n14655) );
  NOR2_X1 U17905 ( .A1(n18925), .A2(n14653), .ZN(n14654) );
  AOI211_X1 U17906 ( .C1(n15150), .C2(n18952), .A(n14655), .B(n14654), .ZN(
        n14656) );
  OAI21_X1 U17907 ( .B1(n15153), .B2(n18957), .A(n14656), .ZN(n14657) );
  OR3_X1 U17908 ( .A1(n14659), .A2(n14658), .A3(n14657), .ZN(P2_U2834) );
  NOR2_X1 U17909 ( .A1(n18941), .A2(n14660), .ZN(n14661) );
  XNOR2_X1 U17910 ( .A(n14661), .B(n15000), .ZN(n14662) );
  NAND2_X1 U17911 ( .A1(n14662), .A2(n18916), .ZN(n14673) );
  OAI21_X1 U17912 ( .B1(n14665), .B2(n14664), .A(n14663), .ZN(n18972) );
  INV_X1 U17913 ( .A(n18972), .ZN(n15002) );
  NOR2_X1 U17914 ( .A1(n14667), .A2(n14666), .ZN(n14668) );
  NOR2_X1 U17915 ( .A1(n14820), .A2(n14668), .ZN(n19008) );
  AOI22_X1 U17916 ( .A1(n19008), .A2(n18952), .B1(n18950), .B2(
        P2_EBX_REG_16__SCAN_IN), .ZN(n14670) );
  AOI21_X1 U17917 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18928), .A(
        n18885), .ZN(n14669) );
  OAI211_X1 U17918 ( .C1(n19713), .C2(n18926), .A(n14670), .B(n14669), .ZN(
        n14671) );
  AOI21_X1 U17919 ( .B1(n15002), .B2(n18939), .A(n14671), .ZN(n14672) );
  OAI211_X1 U17920 ( .C1(n18907), .C2(n14674), .A(n14673), .B(n14672), .ZN(
        P2_U2839) );
  OR2_X1 U17921 ( .A1(n18941), .A2(n14675), .ZN(n18851) );
  AOI211_X1 U17922 ( .C1(n14676), .C2(n16146), .A(n18967), .B(n18851), .ZN(
        n14677) );
  INV_X1 U17923 ( .A(n14677), .ZN(n14684) );
  INV_X1 U17924 ( .A(n16146), .ZN(n14681) );
  NAND2_X1 U17925 ( .A1(n18941), .A2(n18916), .ZN(n18960) );
  AOI22_X1 U17926 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n18950), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n18949), .ZN(n14678) );
  OAI211_X1 U17927 ( .C1(n15298), .C2(n18920), .A(n14678), .B(n18905), .ZN(
        n14679) );
  AOI21_X1 U17928 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18928), .A(
        n14679), .ZN(n14680) );
  OAI21_X1 U17929 ( .B1(n14681), .B2(n18960), .A(n14680), .ZN(n14682) );
  AOI21_X1 U17930 ( .B1(n16150), .B2(n18939), .A(n14682), .ZN(n14683) );
  OAI211_X1 U17931 ( .C1(n14685), .C2(n18907), .A(n14684), .B(n14683), .ZN(
        P2_U2844) );
  AOI211_X1 U17932 ( .C1(n15407), .C2(n14687), .A(n18941), .B(n14686), .ZN(
        n15415) );
  NAND2_X1 U17933 ( .A1(n15415), .A2(n18916), .ZN(n14702) );
  INV_X1 U17934 ( .A(n14688), .ZN(n14690) );
  NAND2_X1 U17935 ( .A1(n14690), .A2(n14689), .ZN(n14691) );
  NAND2_X1 U17936 ( .A1(n14692), .A2(n14691), .ZN(n19785) );
  NAND2_X1 U17937 ( .A1(n18954), .A2(n14693), .ZN(n14696) );
  INV_X1 U17938 ( .A(n18960), .ZN(n18840) );
  MUX2_X1 U17939 ( .A(n18840), .B(n18928), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14694) );
  AOI21_X1 U17940 ( .B1(n18949), .B2(P2_REIP_REG_1__SCAN_IN), .A(n14694), .ZN(
        n14695) );
  OAI211_X1 U17941 ( .C1(n18925), .C2(n14697), .A(n14696), .B(n14695), .ZN(
        n14700) );
  NOR2_X1 U17942 ( .A1(n14698), .A2(n18957), .ZN(n14699) );
  AOI211_X1 U17943 ( .C1(n18952), .C2(n19785), .A(n14700), .B(n14699), .ZN(
        n14701) );
  OAI211_X1 U17944 ( .C1(n19780), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        P2_U2854) );
  OR2_X2 U17945 ( .A1(n14707), .A2(n14706), .ZN(n15052) );
  OR2_X1 U17946 ( .A1(n14709), .A2(n14708), .ZN(n14737) );
  NAND3_X1 U17947 ( .A1(n14737), .A2(n14710), .A3(n18998), .ZN(n14712) );
  NAND2_X1 U17948 ( .A1(n18996), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14711) );
  OAI211_X1 U17949 ( .C1(n18996), .C2(n15052), .A(n14712), .B(n14711), .ZN(
        P2_U2858) );
  INV_X1 U17950 ( .A(n14713), .ZN(n14717) );
  INV_X1 U17951 ( .A(n14714), .ZN(n14716) );
  OAI21_X1 U17952 ( .B1(n14717), .B2(n14716), .A(n14715), .ZN(n16068) );
  AOI21_X1 U17953 ( .B1(n14720), .B2(n14719), .A(n14718), .ZN(n14756) );
  NAND2_X1 U17954 ( .A1(n14756), .A2(n18998), .ZN(n14722) );
  NAND2_X1 U17955 ( .A1(n18996), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14721) );
  OAI211_X1 U17956 ( .C1(n16068), .C2(n18996), .A(n14722), .B(n14721), .ZN(
        P2_U2861) );
  AOI21_X1 U17957 ( .B1(n14724), .B2(n16102), .A(n14723), .ZN(n14801) );
  NAND2_X1 U17958 ( .A1(n14801), .A2(n18998), .ZN(n14726) );
  NAND2_X1 U17959 ( .A1(n18996), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n14725) );
  OAI211_X1 U17960 ( .C1(n15153), .C2(n18996), .A(n14726), .B(n14725), .ZN(
        P2_U2866) );
  INV_X1 U17961 ( .A(n14977), .ZN(n14727) );
  AOI21_X1 U17962 ( .B1(n14728), .B2(n14663), .A(n14727), .ZN(n14991) );
  INV_X1 U17963 ( .A(n14991), .ZN(n18798) );
  AOI21_X1 U17964 ( .B1(n14731), .B2(n18968), .A(n14730), .ZN(n14816) );
  NAND2_X1 U17965 ( .A1(n14816), .A2(n18998), .ZN(n14733) );
  NAND2_X1 U17966 ( .A1(n18996), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14732) );
  OAI211_X1 U17967 ( .C1(n18798), .C2(n18996), .A(n14733), .B(n14732), .ZN(
        P2_U2870) );
  INV_X1 U17968 ( .A(n19057), .ZN(n16117) );
  OAI21_X1 U17969 ( .B1(n14736), .B2(n14735), .A(n14734), .ZN(n16067) );
  NAND3_X1 U17970 ( .A1(n14737), .A2(n14710), .A3(n19038), .ZN(n14743) );
  INV_X1 U17971 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n14740) );
  AOI22_X1 U17972 ( .A1(n19005), .A2(n14738), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19056), .ZN(n14739) );
  OAI21_X1 U17973 ( .B1(n14765), .B2(n14740), .A(n14739), .ZN(n14741) );
  AOI21_X1 U17974 ( .B1(n19007), .B2(BUF1_REG_29__SCAN_IN), .A(n14741), .ZN(
        n14742) );
  OAI211_X1 U17975 ( .C1(n16117), .C2(n16067), .A(n14743), .B(n14742), .ZN(
        P2_U2890) );
  INV_X1 U17976 ( .A(n19007), .ZN(n14766) );
  AOI22_X1 U17977 ( .A1(n19005), .A2(n19016), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19056), .ZN(n14745) );
  NAND2_X1 U17978 ( .A1(n19006), .A2(BUF2_REG_28__SCAN_IN), .ZN(n14744) );
  OAI211_X1 U17979 ( .C1(n14766), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14747) );
  AOI21_X1 U17980 ( .B1(n15067), .B2(n19057), .A(n14747), .ZN(n14748) );
  OAI21_X1 U17981 ( .B1(n14749), .B2(n19061), .A(n14748), .ZN(P2_U2891) );
  AOI22_X1 U17982 ( .A1(n19005), .A2(n14750), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n19056), .ZN(n14752) );
  NAND2_X1 U17983 ( .A1(n19006), .A2(BUF2_REG_27__SCAN_IN), .ZN(n14751) );
  OAI211_X1 U17984 ( .C1(n14766), .C2(n19156), .A(n14752), .B(n14751), .ZN(
        n14753) );
  AOI21_X1 U17985 ( .B1(n15075), .B2(n19057), .A(n14753), .ZN(n14754) );
  OAI21_X1 U17986 ( .B1(n14755), .B2(n19061), .A(n14754), .ZN(P2_U2892) );
  NAND2_X1 U17987 ( .A1(n14756), .A2(n19038), .ZN(n14763) );
  AOI22_X1 U17988 ( .A1(n19005), .A2(n19019), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19056), .ZN(n14762) );
  AOI22_X1 U17989 ( .A1(n19007), .A2(BUF1_REG_26__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14761) );
  NOR2_X1 U17990 ( .A1(n14767), .A2(n14757), .ZN(n14758) );
  NOR2_X1 U17991 ( .A1(n14759), .A2(n14758), .ZN(n16069) );
  NAND2_X1 U17992 ( .A1(n16069), .A2(n19057), .ZN(n14760) );
  NAND4_X1 U17993 ( .A1(n14763), .A2(n14762), .A3(n14761), .A4(n14760), .ZN(
        P2_U2893) );
  INV_X1 U17994 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n14764) );
  OAI22_X1 U17995 ( .A1(n14766), .A2(n16317), .B1(n14765), .B2(n14764), .ZN(
        n14775) );
  INV_X1 U17996 ( .A(n14767), .ZN(n14772) );
  INV_X1 U17997 ( .A(n14768), .ZN(n14769) );
  NAND2_X1 U17998 ( .A1(n14770), .A2(n14769), .ZN(n14771) );
  NAND2_X1 U17999 ( .A1(n14772), .A2(n14771), .ZN(n16092) );
  OAI22_X1 U18000 ( .A1(n16092), .A2(n16117), .B1(n14810), .B2(n14773), .ZN(
        n14774) );
  AOI211_X1 U18001 ( .C1(n19005), .C2(n14776), .A(n14775), .B(n14774), .ZN(
        n14777) );
  OAI21_X1 U18002 ( .B1(n14778), .B2(n19061), .A(n14777), .ZN(P2_U2894) );
  OAI22_X1 U18003 ( .A1(n15114), .A2(n16117), .B1(n14810), .B2(n11871), .ZN(
        n14779) );
  AOI21_X1 U18004 ( .B1(n19005), .B2(n14780), .A(n14779), .ZN(n14782) );
  AOI22_X1 U18005 ( .A1(n19007), .A2(BUF1_REG_24__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n14781) );
  OAI211_X1 U18006 ( .C1(n14783), .C2(n19061), .A(n14782), .B(n14781), .ZN(
        P2_U2895) );
  AOI21_X1 U18007 ( .B1(n14786), .B2(n14785), .A(n14784), .ZN(n16096) );
  AOI22_X1 U18008 ( .A1(n19005), .A2(n14787), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n19056), .ZN(n14789) );
  AOI22_X1 U18009 ( .A1(n19007), .A2(BUF1_REG_23__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n14788) );
  OAI211_X1 U18010 ( .C1(n15131), .C2(n16117), .A(n14789), .B(n14788), .ZN(
        n14790) );
  AOI21_X1 U18011 ( .B1(n16096), .B2(n19038), .A(n14790), .ZN(n14791) );
  INV_X1 U18012 ( .A(n14791), .ZN(P2_U2896) );
  INV_X1 U18013 ( .A(n14792), .ZN(n14794) );
  AOI21_X1 U18014 ( .B1(n14794), .B2(n10303), .A(n14793), .ZN(n16099) );
  INV_X1 U18015 ( .A(n16099), .ZN(n14800) );
  OAI22_X1 U18016 ( .A1(n19176), .A2(n14811), .B1(n14810), .B2(n14795), .ZN(
        n14796) );
  AOI21_X1 U18017 ( .B1(n14797), .B2(n19057), .A(n14796), .ZN(n14799) );
  AOI22_X1 U18018 ( .A1(n19007), .A2(BUF1_REG_22__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n14798) );
  OAI211_X1 U18019 ( .C1(n14800), .C2(n19061), .A(n14799), .B(n14798), .ZN(
        P2_U2897) );
  NAND2_X1 U18020 ( .A1(n14801), .A2(n19038), .ZN(n14806) );
  AOI22_X1 U18021 ( .A1(n19005), .A2(n14802), .B1(n19056), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U18022 ( .A1(n19007), .A2(BUF1_REG_21__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n14804) );
  NAND2_X1 U18023 ( .A1(n15150), .A2(n19057), .ZN(n14803) );
  NAND4_X1 U18024 ( .A1(n14806), .A2(n14805), .A3(n14804), .A4(n14803), .ZN(
        P2_U2898) );
  INV_X1 U18025 ( .A(n15164), .ZN(n14807) );
  OAI21_X1 U18026 ( .B1(n15192), .B2(n14808), .A(n14807), .ZN(n15178) );
  INV_X1 U18027 ( .A(n15178), .ZN(n18774) );
  OAI22_X1 U18028 ( .A1(n19158), .A2(n14811), .B1(n14810), .B2(n14809), .ZN(
        n14812) );
  AOI21_X1 U18029 ( .B1(n18774), .B2(n19057), .A(n14812), .ZN(n14814) );
  AOI22_X1 U18030 ( .A1(n19007), .A2(BUF1_REG_19__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n14813) );
  OAI211_X1 U18031 ( .C1(n14815), .C2(n19061), .A(n14814), .B(n14813), .ZN(
        P2_U2900) );
  NAND2_X1 U18032 ( .A1(n14816), .A2(n19038), .ZN(n14824) );
  AOI22_X1 U18033 ( .A1(n19005), .A2(n14817), .B1(n19056), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n14823) );
  AOI22_X1 U18034 ( .A1(n19007), .A2(BUF1_REG_17__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n14822) );
  INV_X1 U18035 ( .A(n14818), .ZN(n14819) );
  XNOR2_X1 U18036 ( .A(n14820), .B(n14819), .ZN(n18805) );
  NAND2_X1 U18037 ( .A1(n19057), .A2(n18805), .ZN(n14821) );
  NAND4_X1 U18038 ( .A1(n14824), .A2(n14823), .A3(n14822), .A4(n14821), .ZN(
        P2_U2902) );
  INV_X1 U18039 ( .A(n14825), .ZN(n14829) );
  OAI21_X1 U18040 ( .B1(n16186), .B2(n14827), .A(n14826), .ZN(n14828) );
  AOI21_X1 U18041 ( .B1(n16178), .B2(n14829), .A(n14828), .ZN(n14830) );
  OAI21_X1 U18042 ( .B1(n16094), .B2(n15430), .A(n14830), .ZN(n14831) );
  AOI21_X1 U18043 ( .B1(n14832), .B2(n19115), .A(n14831), .ZN(n14833) );
  OAI21_X1 U18044 ( .B1(n14834), .B2(n16179), .A(n14833), .ZN(P2_U2983) );
  NAND2_X1 U18045 ( .A1(n14835), .A2(n14848), .ZN(n14840) );
  INV_X1 U18046 ( .A(n14836), .ZN(n14837) );
  NOR2_X1 U18047 ( .A1(n14838), .A2(n14837), .ZN(n14839) );
  XNOR2_X1 U18048 ( .A(n14840), .B(n14839), .ZN(n15050) );
  NOR2_X1 U18049 ( .A1(n16046), .A2(n15430), .ZN(n14843) );
  NAND2_X1 U18050 ( .A1(n18885), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15044) );
  NAND2_X1 U18051 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14841) );
  OAI211_X1 U18052 ( .C1(n19120), .C2(n16050), .A(n15044), .B(n14841), .ZN(
        n14842) );
  OAI21_X1 U18053 ( .B1(n15050), .B2(n16179), .A(n14844), .ZN(P2_U2984) );
  OAI21_X1 U18054 ( .B1(n14845), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14846), .ZN(n15064) );
  NAND2_X1 U18055 ( .A1(n14849), .A2(n14848), .ZN(n14850) );
  NAND2_X1 U18056 ( .A1(n15051), .A2(n19116), .ZN(n14854) );
  NAND2_X1 U18057 ( .A1(n18885), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15053) );
  OAI21_X1 U18058 ( .B1(n16186), .B2(n16060), .A(n15053), .ZN(n14852) );
  NOR2_X1 U18059 ( .A1(n15052), .A2(n15430), .ZN(n14851) );
  AOI211_X1 U18060 ( .C1(n16178), .C2(n16059), .A(n14852), .B(n14851), .ZN(
        n14853) );
  OAI211_X1 U18061 ( .C1(n16181), .C2(n15064), .A(n14854), .B(n14853), .ZN(
        P2_U2985) );
  XNOR2_X1 U18062 ( .A(n14856), .B(n14858), .ZN(n14867) );
  INV_X1 U18063 ( .A(n14856), .ZN(n14857) );
  AOI22_X1 U18064 ( .A1(n14867), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14858), .B2(n14857), .ZN(n14861) );
  XNOR2_X1 U18065 ( .A(n14859), .B(n15069), .ZN(n14860) );
  XNOR2_X1 U18066 ( .A(n14861), .B(n14860), .ZN(n15074) );
  AOI21_X1 U18067 ( .B1(n15069), .B2(n15083), .A(n14845), .ZN(n15072) );
  NOR2_X1 U18068 ( .A1(n18905), .A2(n19737), .ZN(n15066) );
  AOI21_X1 U18069 ( .B1(n19104), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15066), .ZN(n14864) );
  NAND2_X1 U18070 ( .A1(n16178), .A2(n14862), .ZN(n14863) );
  OAI211_X1 U18071 ( .C1(n15065), .C2(n15430), .A(n14864), .B(n14863), .ZN(
        n14865) );
  AOI21_X1 U18072 ( .B1(n15072), .B2(n19115), .A(n14865), .ZN(n14866) );
  OAI21_X1 U18073 ( .B1(n15074), .B2(n16179), .A(n14866), .ZN(P2_U2986) );
  XNOR2_X1 U18074 ( .A(n14867), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15087) );
  NAND2_X1 U18075 ( .A1(n18885), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15077) );
  OAI21_X1 U18076 ( .B1(n16186), .B2(n14868), .A(n15077), .ZN(n14870) );
  NOR2_X1 U18077 ( .A1(n15078), .A2(n15430), .ZN(n14869) );
  AOI211_X1 U18078 ( .C1(n16178), .C2(n14871), .A(n14870), .B(n14869), .ZN(
        n14874) );
  INV_X1 U18079 ( .A(n14877), .ZN(n14872) );
  INV_X1 U18080 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15055) );
  NAND2_X1 U18081 ( .A1(n14872), .A2(n15055), .ZN(n15084) );
  NAND3_X1 U18082 ( .A1(n15084), .A2(n19115), .A3(n15083), .ZN(n14873) );
  OAI211_X1 U18083 ( .C1(n15087), .C2(n16179), .A(n14874), .B(n14873), .ZN(
        P2_U2987) );
  AOI21_X1 U18084 ( .B1(n14886), .B2(n14883), .A(n14882), .ZN(n14875) );
  XOR2_X1 U18085 ( .A(n14876), .B(n14875), .Z(n15098) );
  INV_X1 U18086 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15092) );
  NAND2_X1 U18087 ( .A1(n14896), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15106) );
  AOI21_X1 U18088 ( .B1(n15092), .B2(n15106), .A(n14877), .ZN(n15095) );
  NOR2_X1 U18089 ( .A1(n18905), .A2(n19733), .ZN(n15088) );
  NOR2_X1 U18090 ( .A1(n19120), .A2(n16073), .ZN(n14878) );
  AOI211_X1 U18091 ( .C1(n19104), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15088), .B(n14878), .ZN(n14879) );
  OAI21_X1 U18092 ( .B1(n16068), .B2(n15430), .A(n14879), .ZN(n14880) );
  AOI21_X1 U18093 ( .B1(n15095), .B2(n19115), .A(n14880), .ZN(n14881) );
  OAI21_X1 U18094 ( .B1(n15098), .B2(n16179), .A(n14881), .ZN(P2_U2988) );
  INV_X1 U18095 ( .A(n14882), .ZN(n14884) );
  NAND2_X1 U18096 ( .A1(n14884), .A2(n14883), .ZN(n14885) );
  XNOR2_X1 U18097 ( .A(n14886), .B(n14885), .ZN(n15110) );
  NAND2_X1 U18098 ( .A1(n18885), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15100) );
  OAI21_X1 U18099 ( .B1(n16186), .B2(n14887), .A(n15100), .ZN(n14889) );
  NOR2_X1 U18100 ( .A1(n15099), .A2(n15430), .ZN(n14888) );
  AOI211_X1 U18101 ( .C1(n16178), .C2(n16084), .A(n14889), .B(n14888), .ZN(
        n14892) );
  INV_X1 U18102 ( .A(n14896), .ZN(n14890) );
  INV_X1 U18103 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15091) );
  NAND2_X1 U18104 ( .A1(n14890), .A2(n15091), .ZN(n15107) );
  NAND3_X1 U18105 ( .A1(n15107), .A2(n19115), .A3(n15106), .ZN(n14891) );
  OAI211_X1 U18106 ( .C1(n15110), .C2(n16179), .A(n14892), .B(n14891), .ZN(
        P2_U2989) );
  XOR2_X1 U18107 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14893), .Z(
        n14894) );
  XNOR2_X1 U18108 ( .A(n14895), .B(n14894), .ZN(n15123) );
  INV_X1 U18109 ( .A(n14918), .ZN(n14939) );
  NAND2_X1 U18110 ( .A1(n14939), .A2(n15127), .ZN(n14903) );
  AOI21_X1 U18111 ( .B1(n15118), .B2(n14903), .A(n14896), .ZN(n15121) );
  NOR2_X1 U18112 ( .A1(n14897), .A2(n15430), .ZN(n14901) );
  NAND2_X1 U18113 ( .A1(n18885), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15113) );
  NAND2_X1 U18114 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14898) );
  OAI211_X1 U18115 ( .C1(n19120), .C2(n14899), .A(n15113), .B(n14898), .ZN(
        n14900) );
  AOI211_X1 U18116 ( .C1(n15121), .C2(n19115), .A(n14901), .B(n14900), .ZN(
        n14902) );
  OAI21_X1 U18117 ( .B1(n15123), .B2(n16179), .A(n14902), .ZN(P2_U2990) );
  INV_X1 U18118 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15143) );
  NOR2_X1 U18119 ( .A1(n14918), .A2(n15143), .ZN(n14917) );
  OAI21_X1 U18120 ( .B1(n14917), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14903), .ZN(n15136) );
  XOR2_X1 U18121 ( .A(n14905), .B(n14904), .Z(n15124) );
  NAND2_X1 U18122 ( .A1(n18885), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15130) );
  OAI21_X1 U18123 ( .B1(n16186), .B2(n14906), .A(n15130), .ZN(n14907) );
  AOI21_X1 U18124 ( .B1(n16178), .B2(n14908), .A(n14907), .ZN(n14909) );
  OAI21_X1 U18125 ( .B1(n15126), .B2(n15430), .A(n14909), .ZN(n14910) );
  AOI21_X1 U18126 ( .B1(n15124), .B2(n19116), .A(n14910), .ZN(n14911) );
  OAI21_X1 U18127 ( .B1(n16181), .B2(n15136), .A(n14911), .ZN(P2_U2991) );
  INV_X1 U18128 ( .A(n14912), .ZN(n14914) );
  NAND2_X1 U18129 ( .A1(n14914), .A2(n14913), .ZN(n14915) );
  XNOR2_X1 U18130 ( .A(n14916), .B(n14915), .ZN(n15149) );
  INV_X1 U18131 ( .A(n14917), .ZN(n15138) );
  NAND2_X1 U18132 ( .A1(n14918), .A2(n15143), .ZN(n15137) );
  NAND3_X1 U18133 ( .A1(n15138), .A2(n19115), .A3(n15137), .ZN(n14924) );
  INV_X1 U18134 ( .A(n16101), .ZN(n14922) );
  NOR2_X1 U18135 ( .A1(n18905), .A2(n19725), .ZN(n15141) );
  AOI21_X1 U18136 ( .B1(n19104), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15141), .ZN(n14919) );
  OAI21_X1 U18137 ( .B1(n19120), .B2(n14920), .A(n14919), .ZN(n14921) );
  AOI21_X1 U18138 ( .B1(n14922), .B2(n19114), .A(n14921), .ZN(n14923) );
  OAI211_X1 U18139 ( .C1(n15149), .C2(n16179), .A(n14924), .B(n14923), .ZN(
        P2_U2992) );
  NAND2_X1 U18140 ( .A1(n15270), .A2(n15269), .ZN(n15268) );
  INV_X1 U18141 ( .A(n14926), .ZN(n14927) );
  NAND2_X1 U18142 ( .A1(n15006), .A2(n14928), .ZN(n14996) );
  NAND2_X1 U18143 ( .A1(n14996), .A2(n14997), .ZN(n15223) );
  NAND2_X1 U18144 ( .A1(n15223), .A2(n14929), .ZN(n14986) );
  INV_X1 U18145 ( .A(n14931), .ZN(n14970) );
  NAND3_X1 U18146 ( .A1(n14947), .A2(n14946), .A3(n14948), .ZN(n14932) );
  NAND2_X1 U18147 ( .A1(n14932), .A2(n9895), .ZN(n14937) );
  INV_X1 U18148 ( .A(n14933), .ZN(n14934) );
  NOR2_X1 U18149 ( .A1(n14935), .A2(n14934), .ZN(n14936) );
  XNOR2_X1 U18150 ( .A(n14937), .B(n14936), .ZN(n15161) );
  AOI21_X1 U18151 ( .B1(n15111), .B2(n14938), .A(n14939), .ZN(n15158) );
  NAND2_X1 U18152 ( .A1(n18885), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15152) );
  OAI21_X1 U18153 ( .B1(n16186), .B2(n14940), .A(n15152), .ZN(n14941) );
  AOI21_X1 U18154 ( .B1(n16178), .B2(n14942), .A(n14941), .ZN(n14943) );
  OAI21_X1 U18155 ( .B1(n15153), .B2(n15430), .A(n14943), .ZN(n14944) );
  AOI21_X1 U18156 ( .B1(n15158), .B2(n19115), .A(n14944), .ZN(n14945) );
  OAI21_X1 U18157 ( .B1(n15161), .B2(n16179), .A(n14945), .ZN(P2_U2993) );
  NAND2_X1 U18158 ( .A1(n14947), .A2(n14946), .ZN(n14950) );
  NAND2_X1 U18159 ( .A1(n9895), .A2(n14948), .ZN(n14949) );
  XNOR2_X1 U18160 ( .A(n14950), .B(n14949), .ZN(n15176) );
  INV_X1 U18161 ( .A(n14951), .ZN(n14952) );
  XNOR2_X1 U18162 ( .A(n14953), .B(n14952), .ZN(n18756) );
  NOR2_X1 U18163 ( .A1(n18905), .A2(n19721), .ZN(n15168) );
  AOI21_X1 U18164 ( .B1(n19104), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15168), .ZN(n14954) );
  OAI21_X1 U18165 ( .B1(n19120), .B2(n18757), .A(n14954), .ZN(n14956) );
  OAI21_X1 U18166 ( .B1(n14964), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14938), .ZN(n15162) );
  NOR2_X1 U18167 ( .A1(n15162), .A2(n16181), .ZN(n14955) );
  AOI211_X1 U18168 ( .C1(n19114), .C2(n18756), .A(n14956), .B(n14955), .ZN(
        n14957) );
  OAI21_X1 U18169 ( .B1(n15176), .B2(n16179), .A(n14957), .ZN(P2_U2994) );
  NAND2_X1 U18170 ( .A1(n14959), .A2(n14958), .ZN(n14963) );
  INV_X1 U18171 ( .A(n14960), .ZN(n14971) );
  NOR2_X1 U18172 ( .A1(n14961), .A2(n14971), .ZN(n14962) );
  XOR2_X1 U18173 ( .A(n14963), .B(n14962), .Z(n15187) );
  AOI21_X1 U18174 ( .B1(n15183), .B2(n14973), .A(n14964), .ZN(n15185) );
  NAND2_X1 U18175 ( .A1(n18885), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15177) );
  OAI21_X1 U18176 ( .B1(n16186), .B2(n14965), .A(n15177), .ZN(n14966) );
  AOI21_X1 U18177 ( .B1(n16178), .B2(n18768), .A(n14966), .ZN(n14967) );
  OAI21_X1 U18178 ( .B1(n18773), .B2(n15430), .A(n14967), .ZN(n14968) );
  AOI21_X1 U18179 ( .B1(n15185), .B2(n19115), .A(n14968), .ZN(n14969) );
  OAI21_X1 U18180 ( .B1(n15187), .B2(n16179), .A(n14969), .ZN(P2_U2995) );
  NOR2_X1 U18181 ( .A1(n14971), .A2(n14970), .ZN(n14972) );
  XNOR2_X1 U18182 ( .A(n14984), .B(n14972), .ZN(n15202) );
  INV_X1 U18183 ( .A(n14973), .ZN(n14974) );
  AOI21_X1 U18184 ( .B1(n14975), .B2(n14993), .A(n14974), .ZN(n15199) );
  AND2_X1 U18185 ( .A1(n14977), .A2(n14976), .ZN(n14979) );
  OR2_X1 U18186 ( .A1(n14979), .A2(n14978), .ZN(n18787) );
  NOR2_X1 U18187 ( .A1(n18787), .A2(n15430), .ZN(n14982) );
  NAND2_X1 U18188 ( .A1(n18885), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U18189 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14980) );
  OAI211_X1 U18190 ( .C1(n19120), .C2(n18779), .A(n15194), .B(n14980), .ZN(
        n14981) );
  AOI211_X1 U18191 ( .C1(n15199), .C2(n19115), .A(n14982), .B(n14981), .ZN(
        n14983) );
  OAI21_X1 U18192 ( .B1(n15202), .B2(n16179), .A(n14983), .ZN(P2_U2996) );
  INV_X1 U18193 ( .A(n14984), .ZN(n14988) );
  AOI22_X1 U18194 ( .A1(n14988), .A2(n14987), .B1(n14986), .B2(n14985), .ZN(
        n15218) );
  NAND2_X1 U18195 ( .A1(n16178), .A2(n18803), .ZN(n14989) );
  NAND2_X1 U18196 ( .A1(n18885), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15213) );
  OAI211_X1 U18197 ( .C1(n16186), .C2(n18793), .A(n14989), .B(n15213), .ZN(
        n14990) );
  AOI21_X1 U18198 ( .B1(n14991), .B2(n19114), .A(n14990), .ZN(n14995) );
  NAND2_X1 U18199 ( .A1(n15248), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15010) );
  NOR2_X1 U18200 ( .A1(n15010), .A2(n15227), .ZN(n15205) );
  OAI211_X1 U18201 ( .C1(n15205), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19115), .B(n14993), .ZN(n14994) );
  OAI211_X1 U18202 ( .C1(n15218), .C2(n16179), .A(n14995), .B(n14994), .ZN(
        P2_U2997) );
  XNOR2_X1 U18203 ( .A(n15010), .B(n15227), .ZN(n15005) );
  INV_X1 U18204 ( .A(n14996), .ZN(n15009) );
  INV_X1 U18205 ( .A(n14997), .ZN(n14998) );
  NAND2_X1 U18206 ( .A1(n15009), .A2(n14998), .ZN(n15224) );
  NAND3_X1 U18207 ( .A1(n15224), .A2(n19116), .A3(n15223), .ZN(n15004) );
  NAND2_X1 U18208 ( .A1(n18885), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15219) );
  NAND2_X1 U18209 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14999) );
  OAI211_X1 U18210 ( .C1(n15000), .C2(n19120), .A(n15219), .B(n14999), .ZN(
        n15001) );
  AOI21_X1 U18211 ( .B1(n15002), .B2(n19114), .A(n15001), .ZN(n15003) );
  OAI211_X1 U18212 ( .C1(n16181), .C2(n15005), .A(n15004), .B(n15003), .ZN(
        P2_U2998) );
  AOI22_X1 U18213 ( .A1(n15009), .A2(n15008), .B1(n15007), .B2(n15006), .ZN(
        n15240) );
  INV_X1 U18214 ( .A(n15248), .ZN(n15011) );
  INV_X1 U18215 ( .A(n15010), .ZN(n15211) );
  AOI21_X1 U18216 ( .B1(n15209), .B2(n15011), .A(n15211), .ZN(n15238) );
  INV_X1 U18217 ( .A(n18817), .ZN(n15015) );
  NOR2_X1 U18218 ( .A1(n18905), .A2(n15012), .ZN(n15233) );
  AOI21_X1 U18219 ( .B1(n19104), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15233), .ZN(n15014) );
  NAND2_X1 U18220 ( .A1(n18810), .A2(n16178), .ZN(n15013) );
  OAI211_X1 U18221 ( .C1(n15015), .C2(n15430), .A(n15014), .B(n15013), .ZN(
        n15016) );
  AOI21_X1 U18222 ( .B1(n15238), .B2(n19115), .A(n15016), .ZN(n15017) );
  OAI21_X1 U18223 ( .B1(n15240), .B2(n16179), .A(n15017), .ZN(P2_U2999) );
  XNOR2_X1 U18224 ( .A(n15018), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15019) );
  XNOR2_X1 U18225 ( .A(n15020), .B(n15019), .ZN(n16206) );
  INV_X1 U18226 ( .A(n15344), .ZN(n15025) );
  INV_X1 U18227 ( .A(n15021), .ZN(n15343) );
  OAI21_X1 U18228 ( .B1(n15023), .B2(n15343), .A(n15022), .ZN(n15024) );
  OAI21_X1 U18229 ( .B1(n15025), .B2(n15343), .A(n15024), .ZN(n16203) );
  OAI22_X1 U18230 ( .A1(n16186), .A2(n15026), .B1(n19703), .B2(n18905), .ZN(
        n15027) );
  AOI21_X1 U18231 ( .B1(n16178), .B2(n18882), .A(n15027), .ZN(n15028) );
  OAI21_X1 U18232 ( .B1(n18889), .B2(n15430), .A(n15028), .ZN(n15029) );
  AOI21_X1 U18233 ( .B1(n16203), .B2(n19116), .A(n15029), .ZN(n15030) );
  OAI21_X1 U18234 ( .B1(n16181), .B2(n16206), .A(n15030), .ZN(P2_U3007) );
  NOR2_X1 U18235 ( .A1(n15031), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19105) );
  INV_X1 U18236 ( .A(n19105), .ZN(n15032) );
  NAND2_X1 U18237 ( .A1(n15031), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19106) );
  NAND2_X1 U18238 ( .A1(n15032), .A2(n19106), .ZN(n15033) );
  XNOR2_X1 U18239 ( .A(n15033), .B(n19107), .ZN(n16207) );
  NAND2_X1 U18240 ( .A1(n16178), .A2(n15034), .ZN(n15035) );
  NAND2_X1 U18241 ( .A1(n19132), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16208) );
  OAI211_X1 U18242 ( .C1(n15036), .C2(n16186), .A(n15035), .B(n16208), .ZN(
        n15040) );
  XNOR2_X1 U18243 ( .A(n15038), .B(n15037), .ZN(n16213) );
  NOR2_X1 U18244 ( .A1(n16213), .A2(n16181), .ZN(n15039) );
  AOI211_X1 U18245 ( .C1(n19114), .C2(n13263), .A(n15040), .B(n15039), .ZN(
        n15041) );
  OAI21_X1 U18246 ( .B1(n16207), .B2(n16179), .A(n15041), .ZN(P2_U3011) );
  AOI21_X1 U18247 ( .B1(n15061), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15042) );
  NOR2_X1 U18248 ( .A1(n15043), .A2(n15042), .ZN(n15047) );
  NAND2_X1 U18249 ( .A1(n16048), .A2(n19126), .ZN(n15045) );
  OAI211_X1 U18250 ( .C1(n16046), .C2(n16191), .A(n15045), .B(n15044), .ZN(
        n15046) );
  OAI21_X1 U18251 ( .B1(n15050), .B2(n16192), .A(n15049), .ZN(P2_U3016) );
  NAND2_X1 U18252 ( .A1(n15051), .A2(n19130), .ZN(n15063) );
  INV_X1 U18253 ( .A(n15052), .ZN(n16064) );
  NAND2_X1 U18254 ( .A1(n16064), .A2(n19121), .ZN(n15054) );
  OAI211_X1 U18255 ( .C1(n16067), .C2(n16209), .A(n15054), .B(n15053), .ZN(
        n15059) );
  AOI21_X1 U18256 ( .B1(n15055), .B2(n15402), .A(n15082), .ZN(n15070) );
  INV_X1 U18257 ( .A(n15056), .ZN(n15057) );
  NAND2_X1 U18258 ( .A1(n15057), .A2(n15069), .ZN(n15068) );
  AOI21_X1 U18259 ( .B1(n15070), .B2(n15068), .A(n15060), .ZN(n15058) );
  OAI211_X1 U18260 ( .C1(n15064), .C2(n16212), .A(n15063), .B(n15062), .ZN(
        P2_U3017) );
  AOI21_X1 U18261 ( .B1(n15072), .B2(n19129), .A(n15071), .ZN(n15073) );
  OAI21_X1 U18262 ( .B1(n15074), .B2(n16192), .A(n15073), .ZN(P2_U3018) );
  NAND2_X1 U18263 ( .A1(n15075), .A2(n19126), .ZN(n15076) );
  OAI211_X1 U18264 ( .C1(n15078), .C2(n16191), .A(n15077), .B(n15076), .ZN(
        n15081) );
  INV_X1 U18265 ( .A(n15090), .ZN(n15079) );
  NOR3_X1 U18266 ( .A1(n15103), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15079), .ZN(n15080) );
  AOI211_X1 U18267 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15082), .A(
        n15081), .B(n15080), .ZN(n15086) );
  NAND3_X1 U18268 ( .A1(n15084), .A2(n19129), .A3(n15083), .ZN(n15085) );
  OAI211_X1 U18269 ( .C1(n15087), .C2(n16192), .A(n15086), .B(n15085), .ZN(
        P2_U3019) );
  INV_X1 U18270 ( .A(n15119), .ZN(n15105) );
  AOI21_X1 U18271 ( .B1(n16069), .B2(n19126), .A(n15088), .ZN(n15089) );
  OAI21_X1 U18272 ( .B1(n16068), .B2(n16191), .A(n15089), .ZN(n15094) );
  AOI211_X1 U18273 ( .C1(n15092), .C2(n15091), .A(n15090), .B(n15103), .ZN(
        n15093) );
  AOI211_X1 U18274 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n15105), .A(
        n15094), .B(n15093), .ZN(n15097) );
  NAND2_X1 U18275 ( .A1(n15095), .A2(n19129), .ZN(n15096) );
  OAI211_X1 U18276 ( .C1(n15098), .C2(n16192), .A(n15097), .B(n15096), .ZN(
        P2_U3020) );
  INV_X1 U18277 ( .A(n15099), .ZN(n16088) );
  OAI21_X1 U18278 ( .B1(n16092), .B2(n16209), .A(n15100), .ZN(n15101) );
  AOI21_X1 U18279 ( .B1(n16088), .B2(n19121), .A(n15101), .ZN(n15102) );
  OAI21_X1 U18280 ( .B1(n15103), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15102), .ZN(n15104) );
  AOI21_X1 U18281 ( .B1(n15105), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15104), .ZN(n15109) );
  NAND3_X1 U18282 ( .A1(n15107), .A2(n19129), .A3(n15106), .ZN(n15108) );
  OAI211_X1 U18283 ( .C1(n15110), .C2(n16192), .A(n15109), .B(n15108), .ZN(
        P2_U3021) );
  NOR2_X1 U18284 ( .A1(n15111), .A2(n15154), .ZN(n15142) );
  NAND3_X1 U18285 ( .A1(n15127), .A2(n15118), .A3(n15142), .ZN(n15112) );
  OAI211_X1 U18286 ( .C1(n15114), .C2(n16209), .A(n15113), .B(n15112), .ZN(
        n15115) );
  AOI21_X1 U18287 ( .B1(n15116), .B2(n19121), .A(n15115), .ZN(n15117) );
  OAI21_X1 U18288 ( .B1(n15119), .B2(n15118), .A(n15117), .ZN(n15120) );
  AOI21_X1 U18289 ( .B1(n15121), .B2(n19129), .A(n15120), .ZN(n15122) );
  OAI21_X1 U18290 ( .B1(n15123), .B2(n16192), .A(n15122), .ZN(P2_U3022) );
  NAND2_X1 U18291 ( .A1(n15124), .A2(n19130), .ZN(n15135) );
  INV_X1 U18292 ( .A(n15157), .ZN(n15125) );
  OAI21_X1 U18293 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15250), .A(
        n15125), .ZN(n15146) );
  NOR2_X1 U18294 ( .A1(n15126), .A2(n16191), .ZN(n15133) );
  INV_X1 U18295 ( .A(n15127), .ZN(n15128) );
  OAI211_X1 U18296 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15128), .B(n15142), .ZN(
        n15129) );
  OAI211_X1 U18297 ( .C1(n15131), .C2(n16209), .A(n15130), .B(n15129), .ZN(
        n15132) );
  AOI211_X1 U18298 ( .C1(n15146), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15133), .B(n15132), .ZN(n15134) );
  OAI211_X1 U18299 ( .C1(n15136), .C2(n16212), .A(n15135), .B(n15134), .ZN(
        P2_U3023) );
  NAND3_X1 U18300 ( .A1(n15138), .A2(n19129), .A3(n15137), .ZN(n15148) );
  NOR2_X1 U18301 ( .A1(n15139), .A2(n16209), .ZN(n15140) );
  AOI211_X1 U18302 ( .C1(n15143), .C2(n15142), .A(n15141), .B(n15140), .ZN(
        n15144) );
  OAI21_X1 U18303 ( .B1(n16101), .B2(n16191), .A(n15144), .ZN(n15145) );
  AOI21_X1 U18304 ( .B1(n15146), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15145), .ZN(n15147) );
  OAI211_X1 U18305 ( .C1(n15149), .C2(n16192), .A(n15148), .B(n15147), .ZN(
        P2_U3024) );
  NAND2_X1 U18306 ( .A1(n15150), .A2(n19126), .ZN(n15151) );
  OAI211_X1 U18307 ( .C1(n15153), .C2(n16191), .A(n15152), .B(n15151), .ZN(
        n15156) );
  NOR2_X1 U18308 ( .A1(n15154), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15155) );
  AOI211_X1 U18309 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15157), .A(
        n15156), .B(n15155), .ZN(n15160) );
  NAND2_X1 U18310 ( .A1(n15158), .A2(n19129), .ZN(n15159) );
  OAI211_X1 U18311 ( .C1(n15161), .C2(n16192), .A(n15160), .B(n15159), .ZN(
        P2_U3025) );
  INV_X1 U18312 ( .A(n15162), .ZN(n15174) );
  NOR2_X1 U18313 ( .A1(n15164), .A2(n15163), .ZN(n15165) );
  NOR2_X1 U18314 ( .A1(n14649), .A2(n15165), .ZN(n18755) );
  INV_X1 U18315 ( .A(n18756), .ZN(n15166) );
  NOR2_X1 U18316 ( .A1(n15166), .A2(n16191), .ZN(n15167) );
  AOI211_X1 U18317 ( .C1(n19126), .C2(n18755), .A(n15168), .B(n15167), .ZN(
        n15171) );
  OAI211_X1 U18318 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15181), .B(n15169), .ZN(
        n15170) );
  OAI211_X1 U18319 ( .C1(n15188), .C2(n15172), .A(n15171), .B(n15170), .ZN(
        n15173) );
  AOI21_X1 U18320 ( .B1(n15174), .B2(n19129), .A(n15173), .ZN(n15175) );
  OAI21_X1 U18321 ( .B1(n15176), .B2(n16192), .A(n15175), .ZN(P2_U3026) );
  NOR2_X1 U18322 ( .A1(n18773), .A2(n16191), .ZN(n15180) );
  OAI21_X1 U18323 ( .B1(n16209), .B2(n15178), .A(n15177), .ZN(n15179) );
  AOI211_X1 U18324 ( .C1(n15181), .C2(n15183), .A(n15180), .B(n15179), .ZN(
        n15182) );
  OAI21_X1 U18325 ( .B1(n15188), .B2(n15183), .A(n15182), .ZN(n15184) );
  AOI21_X1 U18326 ( .B1(n15185), .B2(n19129), .A(n15184), .ZN(n15186) );
  OAI21_X1 U18327 ( .B1(n15187), .B2(n16192), .A(n15186), .ZN(P2_U3027) );
  INV_X1 U18328 ( .A(n15188), .ZN(n15198) );
  NOR2_X1 U18329 ( .A1(n15190), .A2(n15189), .ZN(n15191) );
  NOR2_X1 U18330 ( .A1(n15192), .A2(n15191), .ZN(n16116) );
  NAND2_X1 U18331 ( .A1(n19126), .A2(n16116), .ZN(n15193) );
  OAI211_X1 U18332 ( .C1(n18787), .C2(n16191), .A(n15194), .B(n15193), .ZN(
        n15197) );
  NOR3_X1 U18333 ( .A1(n15250), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15195), .ZN(n15196) );
  AOI211_X1 U18334 ( .C1(n15198), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15197), .B(n15196), .ZN(n15201) );
  NAND2_X1 U18335 ( .A1(n15199), .A2(n19129), .ZN(n15200) );
  OAI211_X1 U18336 ( .C1(n15202), .C2(n16192), .A(n15201), .B(n15200), .ZN(
        P2_U3028) );
  INV_X1 U18337 ( .A(n15203), .ZN(n15229) );
  AND2_X1 U18338 ( .A1(n15402), .A2(n15229), .ZN(n15204) );
  OR2_X1 U18339 ( .A1(n15334), .A2(n15204), .ZN(n15232) );
  AOI21_X1 U18340 ( .B1(n16212), .B2(n15206), .A(n15205), .ZN(n15207) );
  AOI211_X1 U18341 ( .C1(n15208), .C2(n15209), .A(n15232), .B(n15207), .ZN(
        n15228) );
  OAI21_X1 U18342 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15252), .A(
        n15228), .ZN(n15216) );
  NOR3_X1 U18343 ( .A1(n15250), .A2(n15229), .A3(n15209), .ZN(n15210) );
  AOI21_X1 U18344 ( .B1(n15211), .B2(n19129), .A(n15210), .ZN(n15220) );
  NOR3_X1 U18345 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15227), .ZN(n15215) );
  NAND2_X1 U18346 ( .A1(n19126), .A2(n18805), .ZN(n15212) );
  OAI211_X1 U18347 ( .C1(n18798), .C2(n16191), .A(n15213), .B(n15212), .ZN(
        n15214) );
  AOI211_X1 U18348 ( .C1(n15216), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15215), .B(n15214), .ZN(n15217) );
  OAI21_X1 U18349 ( .B1(n15218), .B2(n16192), .A(n15217), .ZN(P2_U3029) );
  OAI21_X1 U18350 ( .B1(n18972), .B2(n16191), .A(n15219), .ZN(n15222) );
  NOR2_X1 U18351 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15221) );
  AOI211_X1 U18352 ( .C1(n19126), .C2(n19008), .A(n15222), .B(n15221), .ZN(
        n15226) );
  NAND3_X1 U18353 ( .A1(n15224), .A2(n19130), .A3(n15223), .ZN(n15225) );
  OAI211_X1 U18354 ( .C1(n15228), .C2(n15227), .A(n15226), .B(n15225), .ZN(
        P2_U3030) );
  NOR3_X1 U18355 ( .A1(n15250), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n15229), .ZN(n15237) );
  XNOR2_X1 U18356 ( .A(n15231), .B(n15230), .ZN(n18816) );
  NAND2_X1 U18357 ( .A1(n15232), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15235) );
  AOI21_X1 U18358 ( .B1(n18817), .B2(n19121), .A(n15233), .ZN(n15234) );
  OAI211_X1 U18359 ( .C1(n18816), .C2(n16209), .A(n15235), .B(n15234), .ZN(
        n15236) );
  AOI211_X1 U18360 ( .C1(n15238), .C2(n19129), .A(n15237), .B(n15236), .ZN(
        n15239) );
  OAI21_X1 U18361 ( .B1(n15240), .B2(n16192), .A(n15239), .ZN(P2_U3031) );
  INV_X1 U18362 ( .A(n16131), .ZN(n15241) );
  AND2_X1 U18363 ( .A1(n15244), .A2(n15243), .ZN(n15245) );
  XNOR2_X1 U18364 ( .A(n15246), .B(n15245), .ZN(n16123) );
  INV_X1 U18365 ( .A(n16123), .ZN(n15267) );
  NAND2_X1 U18366 ( .A1(n14992), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15328) );
  INV_X1 U18367 ( .A(n15286), .ZN(n15282) );
  INV_X1 U18368 ( .A(n15254), .ZN(n15247) );
  NAND2_X1 U18369 ( .A1(n15282), .A2(n15247), .ZN(n16134) );
  AOI21_X1 U18370 ( .B1(n16134), .B2(n15249), .A(n15248), .ZN(n16124) );
  INV_X1 U18371 ( .A(n15250), .ZN(n15335) );
  NAND2_X1 U18372 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15335), .ZN(
        n15319) );
  NOR2_X1 U18373 ( .A1(n15293), .A2(n15319), .ZN(n16187) );
  INV_X1 U18374 ( .A(n16187), .ZN(n15251) );
  NOR2_X1 U18375 ( .A1(n15254), .A2(n15251), .ZN(n15256) );
  NOR2_X1 U18376 ( .A1(n21038), .A2(n15293), .ZN(n15253) );
  INV_X1 U18377 ( .A(n15334), .ZN(n15292) );
  OAI21_X1 U18378 ( .B1(n15253), .B2(n15252), .A(n15292), .ZN(n15274) );
  AOI21_X1 U18379 ( .B1(n16187), .B2(n15254), .A(n15274), .ZN(n16189) );
  INV_X1 U18380 ( .A(n16189), .ZN(n15255) );
  MUX2_X1 U18381 ( .A(n15256), .B(n15255), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n15265) );
  NAND2_X1 U18382 ( .A1(n15258), .A2(n15257), .ZN(n15259) );
  NAND2_X1 U18383 ( .A1(n15260), .A2(n15259), .ZN(n18976) );
  NAND2_X1 U18384 ( .A1(n19126), .A2(n15261), .ZN(n15263) );
  NAND2_X1 U18385 ( .A1(n18885), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n15262) );
  OAI211_X1 U18386 ( .C1(n18976), .C2(n16191), .A(n15263), .B(n15262), .ZN(
        n15264) );
  AOI211_X1 U18387 ( .C1(n16124), .C2(n19129), .A(n15265), .B(n15264), .ZN(
        n15266) );
  OAI21_X1 U18388 ( .B1(n16192), .B2(n15267), .A(n15266), .ZN(P2_U3032) );
  OAI21_X1 U18389 ( .B1(n15270), .B2(n15269), .A(n15268), .ZN(n16143) );
  XNOR2_X1 U18390 ( .A(n15272), .B(n15271), .ZN(n19018) );
  NOR2_X1 U18391 ( .A1(n12628), .A2(n18905), .ZN(n15273) );
  AOI221_X1 U18392 ( .B1(n16187), .B2(n13438), .C1(n15274), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15273), .ZN(n15281) );
  OR2_X1 U18393 ( .A1(n15276), .A2(n15275), .ZN(n15277) );
  NAND2_X1 U18394 ( .A1(n15278), .A2(n15277), .ZN(n18983) );
  INV_X1 U18395 ( .A(n18983), .ZN(n15279) );
  NAND2_X1 U18396 ( .A1(n19121), .A2(n15279), .ZN(n15280) );
  OAI211_X1 U18397 ( .C1(n16209), .C2(n19018), .A(n15281), .B(n15280), .ZN(
        n15284) );
  NOR2_X1 U18398 ( .A1(n15282), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16140) );
  NOR2_X1 U18399 ( .A1(n13438), .A2(n15286), .ZN(n16139) );
  NOR3_X1 U18400 ( .A1(n16140), .A2(n16139), .A3(n16212), .ZN(n15283) );
  AOI211_X1 U18401 ( .C1(n19130), .C2(n16143), .A(n15284), .B(n15283), .ZN(
        n15285) );
  INV_X1 U18402 ( .A(n15285), .ZN(P2_U3034) );
  NOR2_X1 U18403 ( .A1(n15328), .A2(n15312), .ZN(n15311) );
  OAI21_X1 U18404 ( .B1(n15311), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15286), .ZN(n16148) );
  NAND2_X1 U18405 ( .A1(n15289), .A2(n15288), .ZN(n15290) );
  XNOR2_X1 U18406 ( .A(n15287), .B(n15290), .ZN(n16147) );
  AOI21_X1 U18407 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15292), .A(
        n15291), .ZN(n15325) );
  INV_X1 U18408 ( .A(n15293), .ZN(n15294) );
  AOI211_X1 U18409 ( .C1(n15312), .C2(n13436), .A(n15294), .B(n15319), .ZN(
        n15296) );
  INV_X1 U18410 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20894) );
  NOR2_X1 U18411 ( .A1(n20894), .A2(n18905), .ZN(n15295) );
  AOI211_X1 U18412 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15325), .A(
        n15296), .B(n15295), .ZN(n15301) );
  OAI22_X1 U18413 ( .A1(n15298), .A2(n16209), .B1(n16191), .B2(n15297), .ZN(
        n15299) );
  INV_X1 U18414 ( .A(n15299), .ZN(n15300) );
  OAI211_X1 U18415 ( .C1(n16147), .C2(n16192), .A(n15301), .B(n15300), .ZN(
        n15302) );
  INV_X1 U18416 ( .A(n15302), .ZN(n15303) );
  OAI21_X1 U18417 ( .B1(n16148), .B2(n16212), .A(n15303), .ZN(P2_U3035) );
  NAND2_X1 U18418 ( .A1(n15305), .A2(n15304), .ZN(n15310) );
  NAND2_X1 U18419 ( .A1(n15307), .A2(n15306), .ZN(n15332) );
  INV_X1 U18420 ( .A(n15329), .ZN(n15308) );
  OAI21_X1 U18421 ( .B1(n15332), .B2(n15308), .A(n15330), .ZN(n15309) );
  XOR2_X1 U18422 ( .A(n15310), .B(n15309), .Z(n16154) );
  AOI21_X1 U18423 ( .B1(n15312), .B2(n15328), .A(n15311), .ZN(n16156) );
  NAND2_X1 U18424 ( .A1(n16156), .A2(n19129), .ZN(n15327) );
  OR2_X1 U18425 ( .A1(n15314), .A2(n15313), .ZN(n15316) );
  NAND2_X1 U18426 ( .A1(n15316), .A2(n15315), .ZN(n18985) );
  XNOR2_X1 U18427 ( .A(n15318), .B(n15317), .ZN(n19022) );
  INV_X1 U18428 ( .A(n19022), .ZN(n15322) );
  NOR2_X1 U18429 ( .A1(n12540), .A2(n18905), .ZN(n15321) );
  NOR2_X1 U18430 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15319), .ZN(
        n15320) );
  AOI211_X1 U18431 ( .C1(n19126), .C2(n15322), .A(n15321), .B(n15320), .ZN(
        n15323) );
  OAI21_X1 U18432 ( .B1(n16191), .B2(n18985), .A(n15323), .ZN(n15324) );
  AOI21_X1 U18433 ( .B1(n15325), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15324), .ZN(n15326) );
  OAI211_X1 U18434 ( .C1(n16154), .C2(n16192), .A(n15327), .B(n15326), .ZN(
        P2_U3036) );
  OAI21_X1 U18435 ( .B1(n14992), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15328), .ZN(n16160) );
  NAND2_X1 U18436 ( .A1(n15330), .A2(n15329), .ZN(n15331) );
  XNOR2_X1 U18437 ( .A(n15332), .B(n15331), .ZN(n16159) );
  NOR2_X1 U18438 ( .A1(n12364), .A2(n18905), .ZN(n15333) );
  AOI221_X1 U18439 ( .B1(n15335), .B2(n21038), .C1(n15334), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15333), .ZN(n15338) );
  INV_X1 U18440 ( .A(n18880), .ZN(n15336) );
  AOI22_X1 U18441 ( .A1(n19121), .A2(n18876), .B1(n19126), .B2(n15336), .ZN(
        n15337) );
  OAI211_X1 U18442 ( .C1(n16159), .C2(n16192), .A(n15338), .B(n15337), .ZN(
        n15339) );
  INV_X1 U18443 ( .A(n15339), .ZN(n15340) );
  OAI21_X1 U18444 ( .B1(n16160), .B2(n16212), .A(n15340), .ZN(P2_U3037) );
  NAND2_X1 U18445 ( .A1(n15342), .A2(n15341), .ZN(n15346) );
  NOR2_X1 U18446 ( .A1(n15344), .A2(n15343), .ZN(n15345) );
  XOR2_X1 U18447 ( .A(n15346), .B(n15345), .Z(n16165) );
  NOR2_X1 U18448 ( .A1(n15348), .A2(n15347), .ZN(n16164) );
  INV_X1 U18449 ( .A(n16164), .ZN(n15350) );
  NAND3_X1 U18450 ( .A1(n15350), .A2(n19129), .A3(n15349), .ZN(n15359) );
  INV_X1 U18451 ( .A(n18997), .ZN(n15357) );
  OAI22_X1 U18452 ( .A1(n16209), .A2(n15351), .B1(n12293), .B2(n18905), .ZN(
        n15356) );
  OAI21_X1 U18453 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16201), .ZN(n15352) );
  OAI22_X1 U18454 ( .A1(n16198), .A2(n15354), .B1(n15353), .B2(n15352), .ZN(
        n15355) );
  AOI211_X1 U18455 ( .C1(n15357), .C2(n19121), .A(n15356), .B(n15355), .ZN(
        n15358) );
  OAI211_X1 U18456 ( .C1(n16165), .C2(n16192), .A(n15359), .B(n15358), .ZN(
        P2_U3038) );
  INV_X1 U18457 ( .A(n15360), .ZN(n15361) );
  XNOR2_X1 U18458 ( .A(n15362), .B(n15361), .ZN(n16171) );
  INV_X1 U18459 ( .A(n18904), .ZN(n15364) );
  NOR2_X1 U18460 ( .A1(n19702), .A2(n18905), .ZN(n15363) );
  AOI21_X1 U18461 ( .B1(n19126), .B2(n15364), .A(n15363), .ZN(n15365) );
  OAI21_X1 U18462 ( .B1(n16198), .B2(n15366), .A(n15365), .ZN(n15367) );
  AOI21_X1 U18463 ( .B1(n9894), .B2(n19121), .A(n15367), .ZN(n15368) );
  OAI21_X1 U18464 ( .B1(n15369), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15368), .ZN(n15373) );
  OAI21_X1 U18465 ( .B1(n15371), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15370), .ZN(n16174) );
  NOR2_X1 U18466 ( .A1(n16174), .A2(n16212), .ZN(n15372) );
  AOI211_X1 U18467 ( .C1(n16171), .C2(n19130), .A(n15373), .B(n15372), .ZN(
        n15374) );
  INV_X1 U18468 ( .A(n15374), .ZN(P2_U3040) );
  XNOR2_X1 U18469 ( .A(n15376), .B(n15375), .ZN(n16180) );
  INV_X1 U18470 ( .A(n19127), .ZN(n15385) );
  XNOR2_X1 U18471 ( .A(n15377), .B(n18922), .ZN(n19024) );
  INV_X1 U18472 ( .A(n19024), .ZN(n15382) );
  OAI211_X1 U18473 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n19124), .B(n15378), .ZN(n15379) );
  OAI21_X1 U18474 ( .B1(n18905), .B2(n15380), .A(n15379), .ZN(n15381) );
  AOI21_X1 U18475 ( .B1(n19126), .B2(n15382), .A(n15381), .ZN(n15383) );
  OAI21_X1 U18476 ( .B1(n15385), .B2(n15384), .A(n15383), .ZN(n15393) );
  AND2_X1 U18477 ( .A1(n15387), .A2(n15386), .ZN(n15388) );
  OAI22_X1 U18478 ( .A1(n15391), .A2(n15390), .B1(n15389), .B2(n15388), .ZN(
        n16182) );
  NOR2_X1 U18479 ( .A1(n16182), .A2(n16212), .ZN(n15392) );
  AOI211_X1 U18480 ( .C1(n19121), .C2(n18915), .A(n15393), .B(n15392), .ZN(
        n15394) );
  OAI21_X1 U18481 ( .B1(n16192), .B2(n16180), .A(n15394), .ZN(P2_U3041) );
  NOR2_X1 U18482 ( .A1(n16212), .A2(n15395), .ZN(n15396) );
  AOI211_X1 U18483 ( .C1(n15398), .C2(n19130), .A(n15397), .B(n15396), .ZN(
        n15406) );
  AOI22_X1 U18484 ( .A1(n15399), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19126), .B2(n19785), .ZN(n15405) );
  NAND2_X1 U18485 ( .A1(n15400), .A2(n19121), .ZN(n15404) );
  OAI211_X1 U18486 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15402), .B(n15401), .ZN(n15403) );
  NAND4_X1 U18487 ( .A1(n15406), .A2(n15405), .A3(n15404), .A4(n15403), .ZN(
        P2_U3045) );
  INV_X1 U18488 ( .A(n15416), .ZN(n19759) );
  NAND2_X1 U18489 ( .A1(n18912), .A2(n15407), .ZN(n18966) );
  OAI21_X1 U18490 ( .B1(n18912), .B2(n15408), .A(n18966), .ZN(n15414) );
  OAI22_X1 U18491 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19616), .B1(n15411), 
        .B2(n18734), .ZN(n15412) );
  AOI21_X1 U18492 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15739), .A(n15412), .ZN(
        n19760) );
  INV_X1 U18493 ( .A(n19760), .ZN(n15483) );
  MUX2_X1 U18494 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15413), .S(
        n15483), .Z(P2_U3601) );
  NAND2_X1 U18495 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15414), .ZN(n19757) );
  INV_X1 U18496 ( .A(n19757), .ZN(n15417) );
  AOI21_X1 U18497 ( .B1(n18941), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15415), .ZN(n19758) );
  AOI222_X1 U18498 ( .A1(n15418), .A2(n19764), .B1(n15417), .B2(n19758), .C1(
        n19783), .C2(n15416), .ZN(n15420) );
  NAND2_X1 U18499 ( .A1(n19760), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15419) );
  OAI21_X1 U18500 ( .B1(n15420), .B2(n19760), .A(n15419), .ZN(P2_U3600) );
  OAI22_X1 U18501 ( .A1(n15421), .A2(n19756), .B1(n19423), .B2(n19759), .ZN(
        n15422) );
  MUX2_X1 U18502 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15422), .S(
        n15483), .Z(P2_U3596) );
  NAND2_X1 U18503 ( .A1(n19423), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19362) );
  OR2_X1 U18504 ( .A1(n19362), .A2(n15428), .ZN(n15423) );
  NAND2_X1 U18505 ( .A1(n15423), .A2(n19771), .ZN(n15438) );
  INV_X1 U18506 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19770) );
  NAND3_X1 U18507 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19770), .A3(
        n19787), .ZN(n19275) );
  INV_X1 U18508 ( .A(n19275), .ZN(n15424) );
  OR2_X1 U18509 ( .A1(n15438), .A2(n15424), .ZN(n15427) );
  NOR2_X1 U18510 ( .A1(n19794), .A2(n19275), .ZN(n19330) );
  INV_X1 U18511 ( .A(n19330), .ZN(n15445) );
  OAI211_X1 U18512 ( .C1(n15435), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n15445), 
        .B(n19762), .ZN(n15425) );
  AND2_X1 U18513 ( .A1(n15425), .A2(n19624), .ZN(n15426) );
  NAND2_X1 U18514 ( .A1(n15427), .A2(n15426), .ZN(n19319) );
  INV_X1 U18515 ( .A(n19319), .ZN(n19309) );
  INV_X1 U18516 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15442) );
  AOI22_X1 U18517 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19173), .ZN(n19629) );
  INV_X1 U18518 ( .A(n19629), .ZN(n19573) );
  INV_X1 U18519 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18058) );
  INV_X1 U18520 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16319) );
  OAI22_X2 U18521 ( .A1(n18058), .A2(n19169), .B1(n16319), .B2(n19171), .ZN(
        n19626) );
  INV_X1 U18522 ( .A(n19175), .ZN(n15432) );
  NAND2_X1 U18523 ( .A1(n15433), .A2(n15432), .ZN(n19137) );
  OAI22_X1 U18524 ( .A1(n19587), .A2(n19322), .B1(n15445), .B2(n19137), .ZN(
        n15434) );
  AOI21_X1 U18525 ( .B1(n19353), .B2(n19573), .A(n15434), .ZN(n15441) );
  INV_X1 U18526 ( .A(n15435), .ZN(n15436) );
  OAI21_X1 U18527 ( .B1(n15436), .B2(n19330), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15437) );
  NOR2_X2 U18528 ( .A1(n15439), .A2(n19281), .ZN(n19619) );
  NAND2_X1 U18529 ( .A1(n19318), .A2(n19619), .ZN(n15440) );
  OAI211_X1 U18530 ( .C1(n19309), .C2(n15442), .A(n15441), .B(n15440), .ZN(
        P2_U3088) );
  INV_X1 U18531 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15449) );
  INV_X1 U18532 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16326) );
  INV_X1 U18533 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18067) );
  OAI22_X1 U18534 ( .A1(n16326), .A2(n19171), .B1(n18067), .B2(n19169), .ZN(
        n19523) );
  AOI22_X1 U18535 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19173), .ZN(n19500) );
  NOR2_X2 U18536 ( .A1(n15443), .A2(n19175), .ZN(n19636) );
  INV_X1 U18537 ( .A(n19636), .ZN(n15444) );
  OAI22_X1 U18538 ( .A1(n19500), .A2(n19322), .B1(n15445), .B2(n15444), .ZN(
        n15446) );
  AOI21_X1 U18539 ( .B1(n19353), .B2(n19523), .A(n15446), .ZN(n15448) );
  INV_X1 U18540 ( .A(n16115), .ZN(n19055) );
  NOR2_X2 U18541 ( .A1(n19055), .A2(n19281), .ZN(n19637) );
  NAND2_X1 U18542 ( .A1(n19318), .A2(n19637), .ZN(n15447) );
  OAI211_X1 U18543 ( .C1(n19309), .C2(n15449), .A(n15448), .B(n15447), .ZN(
        P2_U3090) );
  NOR2_X2 U18544 ( .A1(n19421), .A2(n19491), .ZN(n19536) );
  OAI21_X1 U18545 ( .B1(n19567), .B2(n19536), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15456) );
  NOR2_X1 U18546 ( .A1(n15451), .A2(n15450), .ZN(n19274) );
  NAND2_X1 U18547 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19274), .ZN(
        n15457) );
  NAND3_X1 U18548 ( .A1(n19787), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19547) );
  NOR2_X1 U18549 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19547), .ZN(
        n19534) );
  INV_X1 U18550 ( .A(n19534), .ZN(n15452) );
  AND2_X1 U18551 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15452), .ZN(n15453) );
  NAND2_X1 U18552 ( .A1(n15454), .A2(n15453), .ZN(n15459) );
  OAI211_X1 U18553 ( .C1(n19534), .C2(n19616), .A(n15459), .B(n19624), .ZN(
        n15455) );
  INV_X1 U18554 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15463) );
  INV_X1 U18555 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18098) );
  OAI22_X2 U18556 ( .A1(n16308), .A2(n19171), .B1(n18098), .B2(n19169), .ZN(
        n19672) );
  INV_X1 U18557 ( .A(n19678), .ZN(n19512) );
  AOI22_X1 U18558 ( .A1(n19536), .A2(n19672), .B1(n19567), .B2(n19512), .ZN(
        n15462) );
  OAI21_X1 U18559 ( .B1(n15457), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19390), 
        .ZN(n15458) );
  AND2_X1 U18560 ( .A1(n15459), .A2(n15458), .ZN(n19535) );
  NOR2_X2 U18561 ( .A1(n15460), .A2(n19281), .ZN(n19670) );
  AOI22_X1 U18562 ( .A1(n19535), .A2(n19670), .B1(n19668), .B2(n19534), .ZN(
        n15461) );
  OAI211_X1 U18563 ( .C1(n19539), .C2(n15463), .A(n15462), .B(n15461), .ZN(
        P2_U3151) );
  AOI22_X1 U18564 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15467) );
  AOI22_X1 U18565 ( .A1(n9790), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15466) );
  AOI22_X1 U18566 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15465) );
  AOI22_X1 U18567 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15464) );
  NAND4_X1 U18568 ( .A1(n15467), .A2(n15466), .A3(n15465), .A4(n15464), .ZN(
        n15473) );
  AOI22_X1 U18569 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15471) );
  AOI22_X1 U18570 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U18571 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15469) );
  AOI22_X1 U18572 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15468) );
  NAND4_X1 U18573 ( .A1(n15471), .A2(n15470), .A3(n15469), .A4(n15468), .ZN(
        n15472) );
  NOR2_X1 U18574 ( .A1(n15473), .A2(n15472), .ZN(n17176) );
  INV_X1 U18575 ( .A(n17076), .ZN(n17079) );
  NOR2_X1 U18576 ( .A1(n17079), .A2(n17057), .ZN(n17061) );
  INV_X1 U18577 ( .A(n17061), .ZN(n17062) );
  NOR2_X1 U18578 ( .A1(n15474), .A2(n17062), .ZN(n15475) );
  NAND2_X1 U18579 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n15475), .ZN(n16964) );
  OAI21_X1 U18580 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n15475), .A(n16964), .ZN(
        n15476) );
  AOI22_X1 U18581 ( .A1(n17080), .A2(n17176), .B1(n15476), .B2(n17075), .ZN(
        P3_U2690) );
  NOR4_X1 U18582 ( .A1(n15479), .A2(n15478), .A3(n15477), .A4(n19756), .ZN(
        n15480) );
  NAND2_X1 U18583 ( .A1(n15483), .A2(n15480), .ZN(n15481) );
  OAI21_X1 U18584 ( .B1(n15483), .B2(n15482), .A(n15481), .ZN(P2_U3595) );
  INV_X1 U18585 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16298) );
  AOI22_X1 U18586 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15484) );
  OAI21_X1 U18587 ( .B1(n15485), .B2(n21015), .A(n15484), .ZN(n15491) );
  AOI22_X1 U18588 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11493), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U18589 ( .A1(n9791), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15489) );
  AOI22_X1 U18590 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9793), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15488) );
  AOI22_X1 U18591 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11510), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15487) );
  AOI22_X1 U18592 ( .A1(n11525), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15493) );
  INV_X1 U18593 ( .A(n15493), .ZN(n15496) );
  AOI22_X1 U18594 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15494) );
  INV_X1 U18595 ( .A(n15494), .ZN(n15495) );
  INV_X1 U18596 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18668) );
  NOR2_X1 U18597 ( .A1(n17232), .A2(n18668), .ZN(n15508) );
  AOI22_X1 U18598 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15507) );
  AOI22_X1 U18599 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U18600 ( .A1(n15486), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15498) );
  OAI21_X1 U18601 ( .B1(n11567), .B2(n18061), .A(n15498), .ZN(n15504) );
  AOI22_X1 U18602 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9791), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15502) );
  AOI22_X1 U18603 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15501) );
  AOI22_X1 U18604 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11493), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18605 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11510), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15499) );
  NAND4_X1 U18606 ( .A1(n15502), .A2(n15501), .A3(n15500), .A4(n15499), .ZN(
        n15503) );
  AOI211_X1 U18607 ( .C1(n17016), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n15504), .B(n15503), .ZN(n15505) );
  NAND3_X1 U18608 ( .A1(n15507), .A2(n15506), .A3(n15505), .ZN(n17706) );
  NAND2_X1 U18609 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17706), .ZN(
        n17705) );
  XNOR2_X1 U18610 ( .A(n15620), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17700) );
  NOR2_X1 U18611 ( .A1(n17705), .A2(n17700), .ZN(n17699) );
  NOR2_X1 U18612 ( .A1(n15508), .A2(n17699), .ZN(n17691) );
  INV_X1 U18613 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U18614 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n16971), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15516) );
  AOI22_X1 U18615 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12889), .B1(
        P3_INSTQUEUE_REG_8__2__SCAN_IN), .B2(n11493), .ZN(n15515) );
  AOI22_X1 U18616 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9789), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15509) );
  OAI21_X1 U18617 ( .B1(n11567), .B2(n18072), .A(n15509), .ZN(n15514) );
  AOI22_X1 U18618 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n17036), .B1(
        P3_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n15546), .ZN(n15513) );
  AOI22_X1 U18619 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n17020), .B1(
        P3_INSTQUEUE_REG_10__2__SCAN_IN), .B2(n17004), .ZN(n15512) );
  AOI22_X1 U18620 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n9793), .B1(n9798), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U18621 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n9787), .B1(
        P3_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n11496), .ZN(n15510) );
  XNOR2_X1 U18622 ( .A(n18005), .B(n15517), .ZN(n17690) );
  NOR2_X1 U18623 ( .A1(n17691), .A2(n17690), .ZN(n15519) );
  NOR2_X1 U18624 ( .A1(n18005), .A2(n15517), .ZN(n15518) );
  INV_X1 U18625 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17983) );
  AOI22_X1 U18626 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15523) );
  AOI22_X1 U18627 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U18628 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15521) );
  AOI22_X1 U18629 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15520) );
  NAND4_X1 U18630 ( .A1(n15523), .A2(n15522), .A3(n15521), .A4(n15520), .ZN(
        n15529) );
  AOI22_X1 U18631 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U18632 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15526) );
  AOI22_X1 U18633 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15525) );
  AOI22_X1 U18634 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15524) );
  NAND4_X1 U18635 ( .A1(n15527), .A2(n15526), .A3(n15525), .A4(n15524), .ZN(
        n15528) );
  INV_X1 U18636 ( .A(n17219), .ZN(n15612) );
  XOR2_X1 U18637 ( .A(n15532), .B(n15612), .Z(n17674) );
  NOR2_X1 U18638 ( .A1(n15530), .A2(n17983), .ZN(n15531) );
  AOI22_X1 U18639 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U18640 ( .A1(n9790), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15541) );
  AOI22_X1 U18641 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15533) );
  OAI21_X1 U18642 ( .B1(n11567), .B2(n18083), .A(n15533), .ZN(n15539) );
  AOI22_X1 U18643 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15537) );
  AOI22_X1 U18644 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15536) );
  AOI22_X1 U18645 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15535) );
  AOI22_X1 U18646 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15534) );
  NAND4_X1 U18647 ( .A1(n15537), .A2(n15536), .A3(n15535), .A4(n15534), .ZN(
        n15538) );
  AOI211_X1 U18648 ( .C1(n16924), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n15539), .B(n15538), .ZN(n15540) );
  NAND3_X1 U18649 ( .A1(n15542), .A2(n15541), .A3(n15540), .ZN(n15613) );
  INV_X1 U18650 ( .A(n15613), .ZN(n17216) );
  XNOR2_X1 U18651 ( .A(n15545), .B(n17216), .ZN(n15543) );
  XNOR2_X1 U18652 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n15543), .ZN(
        n17665) );
  AND2_X1 U18653 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15543), .ZN(
        n15544) );
  AOI22_X1 U18654 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17003), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15550) );
  AOI22_X1 U18655 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15549) );
  AOI22_X1 U18656 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9787), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15548) );
  AOI22_X1 U18657 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15547) );
  NAND4_X1 U18658 ( .A1(n15550), .A2(n15549), .A3(n15548), .A4(n15547), .ZN(
        n15557) );
  AOI22_X1 U18659 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15555) );
  AOI22_X1 U18660 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15554) );
  AOI22_X1 U18661 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15553) );
  AOI22_X1 U18662 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15552) );
  NAND4_X1 U18663 ( .A1(n15555), .A2(n15554), .A3(n15553), .A4(n15552), .ZN(
        n15556) );
  INV_X1 U18664 ( .A(n17211), .ZN(n15614) );
  XOR2_X1 U18665 ( .A(n15558), .B(n15614), .Z(n17649) );
  AOI22_X1 U18666 ( .A1(n9790), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U18667 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15567) );
  AOI22_X1 U18668 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15559) );
  OAI21_X1 U18669 ( .B1(n15575), .B2(n20973), .A(n15559), .ZN(n15565) );
  AOI22_X1 U18670 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U18671 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U18672 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15561) );
  AOI22_X1 U18673 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15560) );
  NAND4_X1 U18674 ( .A1(n15563), .A2(n15562), .A3(n15561), .A4(n15560), .ZN(
        n15564) );
  AOI211_X1 U18675 ( .C1(n17003), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n15565), .B(n15564), .ZN(n15566) );
  NAND3_X1 U18676 ( .A1(n15568), .A2(n15567), .A3(n15566), .ZN(n15631) );
  INV_X1 U18677 ( .A(n15631), .ZN(n17208) );
  XNOR2_X1 U18678 ( .A(n15570), .B(n17208), .ZN(n15569) );
  XNOR2_X1 U18679 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15569), .ZN(
        n17635) );
  NAND2_X1 U18680 ( .A1(n15570), .A2(n15631), .ZN(n16290) );
  AOI22_X1 U18681 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U18682 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U18683 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U18684 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9788), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15571) );
  NAND4_X1 U18685 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15581) );
  AOI22_X1 U18686 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15579) );
  AOI22_X1 U18687 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15578) );
  AOI22_X1 U18688 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15577) );
  AOI22_X1 U18689 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15576) );
  NAND4_X1 U18690 ( .A1(n15579), .A2(n15578), .A3(n15577), .A4(n15576), .ZN(
        n15580) );
  INV_X1 U18691 ( .A(n15582), .ZN(n15647) );
  AOI21_X1 U18692 ( .B1(n16290), .B2(n17204), .A(n15582), .ZN(n15583) );
  INV_X1 U18693 ( .A(n15583), .ZN(n15584) );
  INV_X1 U18694 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17962) );
  NOR2_X1 U18695 ( .A1(n15585), .A2(n15584), .ZN(n15586) );
  NOR2_X2 U18696 ( .A1(n17624), .A2(n15586), .ZN(n15646) );
  INV_X1 U18697 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17948) );
  NOR2_X2 U18698 ( .A1(n15646), .A2(n17948), .ZN(n17916) );
  INV_X1 U18699 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17903) );
  NAND2_X1 U18700 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17922) );
  INV_X1 U18701 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17574) );
  NOR2_X1 U18702 ( .A1(n17922), .A2(n17574), .ZN(n17906) );
  NAND3_X1 U18703 ( .A1(n17906), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17521) );
  NOR2_X1 U18704 ( .A1(n17903), .A2(n17521), .ZN(n17524) );
  NAND2_X1 U18705 ( .A1(n17524), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15648) );
  INV_X1 U18706 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17848) );
  INV_X1 U18707 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17837) );
  NOR2_X1 U18708 ( .A1(n17848), .A2(n17837), .ZN(n17827) );
  INV_X1 U18709 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17830) );
  INV_X1 U18710 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17783) );
  NAND2_X1 U18711 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17452) );
  NOR3_X1 U18712 ( .A1(n17830), .A2(n17783), .A3(n17452), .ZN(n17785) );
  NAND2_X1 U18713 ( .A1(n17827), .A2(n17785), .ZN(n17779) );
  NAND2_X1 U18714 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17732) );
  NOR2_X1 U18715 ( .A1(n17779), .A2(n17732), .ZN(n15650) );
  NAND2_X1 U18716 ( .A1(n17856), .A2(n15650), .ZN(n17762) );
  INV_X1 U18717 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17765) );
  NOR2_X1 U18718 ( .A1(n17762), .A2(n17765), .ZN(n17388) );
  NAND2_X1 U18719 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17388), .ZN(
        n17387) );
  INV_X1 U18720 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17735) );
  INV_X1 U18721 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17730) );
  NOR3_X1 U18722 ( .A1(n16298), .A2(n17723), .A3(n17730), .ZN(n16264) );
  INV_X1 U18723 ( .A(n15591), .ZN(n15592) );
  NAND3_X1 U18724 ( .A1(n15592), .A2(n18708), .A3(n18514), .ZN(n15593) );
  NAND2_X1 U18725 ( .A1(n15594), .A2(n15593), .ZN(n18507) );
  XOR2_X1 U18726 ( .A(n18069), .B(n18062), .Z(n15596) );
  INV_X1 U18727 ( .A(n17204), .ZN(n16288) );
  NAND2_X1 U18728 ( .A1(n15595), .A2(n18496), .ZN(n15608) );
  OAI21_X1 U18729 ( .B1(n18707), .B2(n15596), .A(n18702), .ZN(n16398) );
  INV_X1 U18730 ( .A(n18080), .ZN(n15597) );
  OAI21_X1 U18731 ( .B1(n15598), .B2(n15597), .A(n18498), .ZN(n15607) );
  NOR2_X1 U18732 ( .A1(n18062), .A2(n15599), .ZN(n15605) );
  INV_X1 U18733 ( .A(n15600), .ZN(n15603) );
  OAI21_X1 U18734 ( .B1(n15603), .B2(n15602), .A(n15601), .ZN(n18500) );
  NAND3_X1 U18735 ( .A1(n15605), .A2(n15604), .A3(n18500), .ZN(n15606) );
  OAI211_X1 U18736 ( .C1(n15608), .C2(n16398), .A(n15607), .B(n15606), .ZN(
        n15609) );
  OAI21_X2 U18737 ( .B1(n15610), .B2(n15609), .A(n18706), .ZN(n18022) );
  NOR2_X1 U18738 ( .A1(n17915), .A2(n18022), .ZN(n17888) );
  NAND2_X1 U18739 ( .A1(n17232), .A2(n17706), .ZN(n15618) );
  NAND2_X1 U18740 ( .A1(n10128), .A2(n15618), .ZN(n15617) );
  AND2_X1 U18741 ( .A1(n15613), .A2(n15627), .ZN(n15615) );
  NAND2_X1 U18742 ( .A1(n15615), .A2(n15614), .ZN(n15630) );
  NOR2_X1 U18743 ( .A1(n17208), .A2(n15630), .ZN(n15635) );
  NAND2_X1 U18744 ( .A1(n15635), .A2(n16288), .ZN(n15636) );
  XNOR2_X1 U18745 ( .A(n17211), .B(n15615), .ZN(n15616) );
  AND2_X1 U18746 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15616), .ZN(
        n15629) );
  XNOR2_X1 U18747 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n15616), .ZN(
        n17653) );
  XOR2_X1 U18748 ( .A(n17219), .B(n15617), .Z(n15625) );
  NOR2_X1 U18749 ( .A1(n17983), .A2(n15625), .ZN(n15626) );
  XOR2_X1 U18750 ( .A(n10128), .B(n15618), .Z(n15619) );
  NOR2_X1 U18751 ( .A1(n15619), .A2(n18005), .ZN(n15624) );
  XNOR2_X1 U18752 ( .A(n18005), .B(n15619), .ZN(n17689) );
  INV_X1 U18753 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18031) );
  NOR2_X1 U18754 ( .A1(n15620), .A2(n18031), .ZN(n15623) );
  INV_X1 U18755 ( .A(n17706), .ZN(n15622) );
  NAND3_X1 U18756 ( .A1(n15622), .A2(n15620), .A3(n18031), .ZN(n15621) );
  OAI221_X1 U18757 ( .B1(n15623), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n15622), .C2(n15620), .A(n15621), .ZN(n17688) );
  NOR2_X1 U18758 ( .A1(n17689), .A2(n17688), .ZN(n17687) );
  NOR2_X1 U18759 ( .A1(n15624), .A2(n17687), .ZN(n17680) );
  XNOR2_X1 U18760 ( .A(n17983), .B(n15625), .ZN(n17679) );
  NOR2_X1 U18761 ( .A1(n17680), .A2(n17679), .ZN(n17678) );
  NOR2_X1 U18762 ( .A1(n15626), .A2(n17678), .ZN(n17660) );
  XOR2_X1 U18763 ( .A(n17216), .B(n15627), .Z(n17661) );
  NOR2_X1 U18764 ( .A1(n17660), .A2(n17661), .ZN(n15628) );
  NAND2_X1 U18765 ( .A1(n17660), .A2(n17661), .ZN(n17659) );
  OAI21_X1 U18766 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15628), .A(
        n17659), .ZN(n17652) );
  NOR2_X1 U18767 ( .A1(n17653), .A2(n17652), .ZN(n17651) );
  NOR2_X1 U18768 ( .A1(n15629), .A2(n17651), .ZN(n15632) );
  XOR2_X1 U18769 ( .A(n15631), .B(n15630), .Z(n15633) );
  NOR2_X1 U18770 ( .A1(n15632), .A2(n15633), .ZN(n15634) );
  INV_X1 U18771 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17641) );
  XNOR2_X1 U18772 ( .A(n15633), .B(n15632), .ZN(n17640) );
  NOR2_X1 U18773 ( .A1(n17641), .A2(n17640), .ZN(n17639) );
  NOR2_X1 U18774 ( .A1(n15634), .A2(n17639), .ZN(n15637) );
  XNOR2_X1 U18775 ( .A(n16288), .B(n15635), .ZN(n15638) );
  NAND2_X1 U18776 ( .A1(n15637), .A2(n15638), .ZN(n17626) );
  NAND2_X1 U18777 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17626), .ZN(
        n15640) );
  NOR2_X1 U18778 ( .A1(n15636), .A2(n15640), .ZN(n15642) );
  INV_X1 U18779 ( .A(n15636), .ZN(n15641) );
  OR2_X1 U18780 ( .A1(n15638), .A2(n15637), .ZN(n17627) );
  OAI21_X1 U18781 ( .B1(n15641), .B2(n15640), .A(n17627), .ZN(n15639) );
  AOI21_X1 U18782 ( .B1(n15641), .B2(n15640), .A(n15639), .ZN(n17614) );
  NOR2_X2 U18783 ( .A1(n17529), .A2(n15648), .ZN(n17867) );
  NAND2_X1 U18784 ( .A1(n15650), .A2(n17867), .ZN(n17758) );
  NOR2_X1 U18785 ( .A1(n17765), .A2(n17758), .ZN(n17397) );
  NAND2_X1 U18786 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17397), .ZN(
        n17396) );
  NOR2_X1 U18787 ( .A1(n17735), .A2(n17396), .ZN(n17721) );
  NAND3_X1 U18788 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n17721), .ZN(n16291) );
  NAND2_X1 U18789 ( .A1(n17785), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16297) );
  INV_X1 U18790 ( .A(n16297), .ZN(n17744) );
  NAND2_X1 U18791 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17746) );
  NAND2_X1 U18792 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17719) );
  NOR2_X1 U18793 ( .A1(n17746), .A2(n17719), .ZN(n15658) );
  INV_X1 U18794 ( .A(n15658), .ZN(n17715) );
  NOR2_X1 U18795 ( .A1(n17730), .A2(n17715), .ZN(n15660) );
  INV_X1 U18796 ( .A(n15660), .ZN(n17351) );
  NOR2_X1 U18797 ( .A1(n18022), .A2(n17351), .ZN(n16299) );
  INV_X1 U18798 ( .A(n18506), .ZN(n18524) );
  AOI21_X1 U18799 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17945) );
  NAND4_X1 U18800 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17961) );
  NOR2_X1 U18801 ( .A1(n17962), .A2(n17961), .ZN(n17952) );
  NAND2_X1 U18802 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17952), .ZN(
        n17821) );
  NOR2_X1 U18803 ( .A1(n17945), .A2(n17821), .ZN(n17874) );
  INV_X1 U18804 ( .A(n15648), .ZN(n17823) );
  AND2_X1 U18805 ( .A1(n17823), .A2(n17827), .ZN(n16296) );
  NAND2_X1 U18806 ( .A1(n17874), .A2(n16296), .ZN(n17829) );
  INV_X1 U18807 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17862) );
  NAND2_X1 U18808 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17944) );
  NOR2_X1 U18809 ( .A1(n17821), .A2(n17944), .ZN(n17912) );
  NAND2_X1 U18810 ( .A1(n17524), .A2(n17912), .ZN(n17875) );
  NOR2_X1 U18811 ( .A1(n17862), .A2(n17875), .ZN(n17844) );
  NAND2_X1 U18812 ( .A1(n17827), .A2(n17844), .ZN(n15657) );
  NAND2_X1 U18813 ( .A1(n18531), .A2(n18031), .ZN(n18025) );
  NAND2_X1 U18814 ( .A1(n18531), .A2(n18516), .ZN(n18003) );
  NAND2_X1 U18815 ( .A1(n18025), .A2(n18003), .ZN(n18008) );
  OAI22_X1 U18816 ( .A1(n18524), .A2(n17829), .B1(n15657), .B2(n18008), .ZN(
        n17743) );
  NAND4_X1 U18817 ( .A1(n17744), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n16299), .A4(n17743), .ZN(n16277) );
  OAI21_X1 U18818 ( .B1(n18039), .B2(n16291), .A(n16277), .ZN(n15643) );
  AOI21_X1 U18819 ( .B1(n16264), .B2(n17888), .A(n15643), .ZN(n15716) );
  INV_X1 U18820 ( .A(n18499), .ZN(n15644) );
  INV_X1 U18821 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17814) );
  NAND2_X1 U18822 ( .A1(n17486), .A2(n17814), .ZN(n15645) );
  NOR2_X1 U18823 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15645), .ZN(
        n17450) );
  NAND2_X1 U18824 ( .A1(n17450), .A2(n17783), .ZN(n17432) );
  NOR2_X2 U18825 ( .A1(n15648), .A2(n17519), .ZN(n15651) );
  NOR2_X2 U18826 ( .A1(n15649), .A2(n17617), .ZN(n17595) );
  NOR2_X1 U18827 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17581) );
  NAND2_X1 U18828 ( .A1(n17595), .A2(n17581), .ZN(n17573) );
  NOR2_X2 U18829 ( .A1(n17573), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17559) );
  INV_X1 U18830 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17558) );
  NAND2_X1 U18831 ( .A1(n17559), .A2(n17558), .ZN(n17520) );
  NOR2_X1 U18832 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17860) );
  NAND2_X1 U18833 ( .A1(n17827), .A2(n15651), .ZN(n17449) );
  NAND2_X1 U18834 ( .A1(n17415), .A2(n17449), .ZN(n17487) );
  INV_X1 U18835 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17429) );
  NOR3_X2 U18836 ( .A1(n17408), .A2(n17416), .A3(n17429), .ZN(n17399) );
  INV_X1 U18837 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17753) );
  NAND2_X1 U18838 ( .A1(n17617), .A2(n17753), .ZN(n15652) );
  OAI211_X2 U18839 ( .C1(n17399), .C2(n17753), .A(n17398), .B(n15652), .ZN(
        n17380) );
  NOR2_X2 U18840 ( .A1(n17380), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17379) );
  NOR2_X1 U18841 ( .A1(n17379), .A2(n15654), .ZN(n15655) );
  OR2_X2 U18842 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15655), .ZN(
        n16301) );
  NAND2_X1 U18843 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15655), .ZN(
        n16289) );
  NOR2_X1 U18844 ( .A1(n15715), .A2(n15714), .ZN(n15656) );
  XNOR2_X1 U18845 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n15656), .ZN(
        n16268) );
  NOR2_X1 U18846 ( .A1(n16297), .A2(n15657), .ZN(n15659) );
  AOI21_X1 U18847 ( .B1(n15658), .B2(n15659), .A(n18531), .ZN(n15662) );
  NOR2_X1 U18848 ( .A1(n17829), .A2(n16297), .ZN(n17763) );
  AOI21_X1 U18849 ( .B1(n17763), .B2(n15658), .A(n18524), .ZN(n17718) );
  AND2_X1 U18850 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15659), .ZN(
        n17716) );
  AOI21_X1 U18851 ( .B1(n17716), .B2(n15660), .A(n18516), .ZN(n15661) );
  NOR4_X1 U18852 ( .A1(n15662), .A2(n17718), .A3(n15661), .A4(n18022), .ZN(
        n15712) );
  OAI21_X1 U18853 ( .B1(n17930), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15712), .ZN(n16295) );
  AOI21_X1 U18854 ( .B1(n16298), .B2(n15710), .A(n16295), .ZN(n15663) );
  NAND3_X1 U18855 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16254) );
  NOR2_X1 U18856 ( .A1(n17723), .A2(n16254), .ZN(n16248) );
  INV_X1 U18857 ( .A(n16248), .ZN(n16253) );
  INV_X1 U18858 ( .A(n17721), .ZN(n17359) );
  NOR2_X1 U18859 ( .A1(n17359), .A2(n16254), .ZN(n16246) );
  INV_X1 U18860 ( .A(n16246), .ZN(n16252) );
  AOI22_X1 U18861 ( .A1(n17888), .A2(n16253), .B1(n18019), .B2(n16252), .ZN(
        n15719) );
  OAI21_X1 U18862 ( .B1(n18035), .B2(n15663), .A(n15719), .ZN(n15664) );
  AOI22_X1 U18863 ( .A1(n17955), .A2(n16268), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15664), .ZN(n15665) );
  NAND2_X1 U18864 ( .A1(n18035), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16274) );
  OAI211_X1 U18865 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15716), .A(
        n15665), .B(n16274), .ZN(P3_U2833) );
  INV_X1 U18866 ( .A(n15666), .ZN(n15679) );
  OAI22_X1 U18867 ( .A1(n20166), .A2(n15668), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15667), .ZN(n20705) );
  NAND2_X1 U18868 ( .A1(n15669), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n20713) );
  INV_X1 U18869 ( .A(n20713), .ZN(n15670) );
  NOR3_X1 U18870 ( .A1(n20705), .A2(n15670), .A3(n20489), .ZN(n15675) );
  AOI211_X1 U18871 ( .C1(n15675), .C2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15672), .B(n15671), .ZN(n15673) );
  INV_X1 U18872 ( .A(n15673), .ZN(n15674) );
  OAI21_X1 U18873 ( .B1(n15675), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15674), .ZN(n15676) );
  AOI222_X1 U18874 ( .A1(n15677), .A2(n20375), .B1(n15677), .B2(n15676), .C1(
        n20375), .C2(n15676), .ZN(n15678) );
  AOI222_X1 U18875 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15679), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15678), .C1(n15679), 
        .C2(n15678), .ZN(n15688) );
  NAND2_X1 U18876 ( .A1(n15680), .A2(n9932), .ZN(n15684) );
  OAI21_X1 U18877 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15681), .ZN(n15682) );
  NAND4_X1 U18878 ( .A1(n15685), .A2(n15684), .A3(n15683), .A4(n15682), .ZN(
        n15686) );
  AOI211_X1 U18879 ( .C1(n15688), .C2(n20042), .A(n15687), .B(n15686), .ZN(
        n15702) );
  INV_X1 U18880 ( .A(n15689), .ZN(n15692) );
  NAND3_X1 U18881 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20635), .A3(n10081), 
        .ZN(n15690) );
  AOI22_X1 U18882 ( .A1(n15693), .A2(n15692), .B1(n15691), .B2(n15690), .ZN(
        n16038) );
  OAI221_X1 U18883 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15702), 
        .A(n16038), .ZN(n16044) );
  AND2_X1 U18884 ( .A1(n15694), .A2(n15696), .ZN(n15695) );
  NOR2_X1 U18885 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15695), .ZN(n15700) );
  AOI211_X1 U18886 ( .C1(n20635), .C2(n10613), .A(n15697), .B(n15696), .ZN(
        n15698) );
  NAND2_X1 U18887 ( .A1(n16044), .A2(n15698), .ZN(n15699) );
  AOI22_X1 U18888 ( .A1(n16044), .A2(n15700), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15699), .ZN(n15701) );
  OAI21_X1 U18889 ( .B1(n15702), .B2(n19811), .A(n15701), .ZN(P1_U3161) );
  AOI22_X1 U18890 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15703), .B1(
        n19986), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15708) );
  NOR2_X1 U18891 ( .A1(n15704), .A2(n11179), .ZN(n15724) );
  NOR3_X1 U18892 ( .A1(n13163), .A2(n11189), .A3(n15874), .ZN(n15725) );
  MUX2_X1 U18893 ( .A(n15724), .B(n15725), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n15705) );
  XNOR2_X1 U18894 ( .A(n15705), .B(n11186), .ZN(n15861) );
  INV_X1 U18895 ( .A(n15706), .ZN(n15775) );
  AOI22_X1 U18896 ( .A1(n15861), .A2(n20031), .B1(n20027), .B2(n15775), .ZN(
        n15707) );
  OAI211_X1 U18897 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15709), .A(
        n15708), .B(n15707), .ZN(P1_U3010) );
  INV_X1 U18898 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16278) );
  NAND2_X1 U18899 ( .A1(n18032), .A2(n15710), .ZN(n17974) );
  INV_X1 U18900 ( .A(n17974), .ZN(n18026) );
  INV_X1 U18901 ( .A(n15712), .ZN(n15713) );
  AOI22_X1 U18902 ( .A1(n18026), .A2(n16254), .B1(n9800), .B2(n15713), .ZN(
        n16276) );
  INV_X1 U18903 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16279) );
  INV_X1 U18904 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18643) );
  NOR2_X1 U18905 ( .A1(n9800), .A2(n18643), .ZN(n16255) );
  NOR3_X1 U18906 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15716), .A3(
        n16279), .ZN(n15717) );
  AOI211_X1 U18907 ( .C1(n17955), .C2(n16261), .A(n16255), .B(n15717), .ZN(
        n15718) );
  INV_X1 U18908 ( .A(HOLD), .ZN(n20742) );
  INV_X1 U18909 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n15721) );
  NAND2_X1 U18910 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15721), .ZN(n20634) );
  INV_X1 U18911 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20630) );
  INV_X1 U18912 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20636) );
  NOR2_X1 U18913 ( .A1(n20630), .A2(n20636), .ZN(n20639) );
  AOI221_X1 U18914 ( .B1(n15721), .B2(n20639), .C1(n20742), .C2(n20639), .A(
        n15720), .ZN(n15723) );
  NAND2_X1 U18915 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20635), .ZN(n15722) );
  OAI211_X1 U18916 ( .C1(n20742), .C2(n20634), .A(n15723), .B(n15722), .ZN(
        P1_U3195) );
  INV_X1 U18917 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16386) );
  NOR2_X1 U18918 ( .A1(n19925), .A2(n16386), .ZN(P1_U2905) );
  NOR2_X1 U18919 ( .A1(n15725), .A2(n15724), .ZN(n15726) );
  XNOR2_X1 U18920 ( .A(n15726), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15868) );
  AOI22_X1 U18921 ( .A1(n15868), .A2(n20031), .B1(n20027), .B2(n15727), .ZN(
        n15734) );
  AOI21_X1 U18922 ( .B1(n15969), .B2(n15728), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15936) );
  INV_X1 U18923 ( .A(n15729), .ZN(n15933) );
  OAI21_X1 U18924 ( .B1(n15936), .B2(n15933), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15733) );
  NAND2_X1 U18925 ( .A1(n19986), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15869) );
  NAND3_X1 U18926 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15731), .A3(
        n15730), .ZN(n15732) );
  NAND4_X1 U18927 ( .A1(n15734), .A2(n15733), .A3(n15869), .A4(n15732), .ZN(
        P1_U3011) );
  NOR3_X1 U18928 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15737) );
  NOR2_X1 U18929 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15736) );
  NOR3_X1 U18930 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12943), .A3(n15735), 
        .ZN(n16222) );
  NOR4_X1 U18931 ( .A1(n15737), .A2(n15736), .A3(n16222), .A4(n15739), .ZN(
        P2_U3178) );
  AOI221_X1 U18932 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15739), .C1(n15738), .C2(
        n15739), .A(n19624), .ZN(n19795) );
  INV_X1 U18933 ( .A(n19795), .ZN(n19792) );
  NOR2_X1 U18934 ( .A1(n15740), .A2(n19792), .ZN(P2_U3047) );
  NAND3_X1 U18935 ( .A1(n18706), .A2(n18496), .A3(n18702), .ZN(n17278) );
  NAND2_X1 U18936 ( .A1(n18097), .A2(n17230), .ZN(n17222) );
  INV_X1 U18937 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17313) );
  NOR2_X1 U18938 ( .A1(n17215), .A2(n18530), .ZN(n17234) );
  NAND2_X1 U18939 ( .A1(n18530), .A2(n17230), .ZN(n17226) );
  AOI22_X1 U18940 ( .A1(n17234), .A2(BUF2_REG_0__SCAN_IN), .B1(n17233), .B2(
        n17706), .ZN(n15744) );
  OAI221_X1 U18941 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17222), .C1(n17313), 
        .C2(n17230), .A(n15744), .ZN(P3_U2735) );
  NOR4_X1 U18942 ( .A1(n19891), .A2(n20672), .A3(n20671), .A4(n15788), .ZN(
        n15760) );
  AOI21_X1 U18943 ( .B1(n15745), .B2(n15760), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15755) );
  OAI22_X1 U18944 ( .A1(n15746), .A2(n15826), .B1(n15859), .B2(n19906), .ZN(
        n15747) );
  AOI21_X1 U18945 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(n19901), .A(n15747), .ZN(
        n15754) );
  NAND2_X1 U18946 ( .A1(n15749), .A2(n15748), .ZN(n15750) );
  NAND2_X1 U18947 ( .A1(n15751), .A2(n15750), .ZN(n15927) );
  OAI22_X1 U18948 ( .A1(n15853), .A2(n19847), .B1(n15927), .B2(n19892), .ZN(
        n15752) );
  INV_X1 U18949 ( .A(n15752), .ZN(n15753) );
  OAI211_X1 U18950 ( .C1(n15756), .C2(n15755), .A(n15754), .B(n15753), .ZN(
        P1_U2817) );
  NAND2_X1 U18951 ( .A1(n15757), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15770) );
  AOI21_X1 U18952 ( .B1(n19878), .B2(n15770), .A(n15758), .ZN(n15783) );
  OAI21_X1 U18953 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n19891), .A(n15783), 
        .ZN(n15759) );
  AOI22_X1 U18954 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19897), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n15759), .ZN(n15768) );
  INV_X1 U18955 ( .A(n15760), .ZN(n15782) );
  NOR3_X1 U18956 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15761), .A3(n15782), 
        .ZN(n15765) );
  OAI22_X1 U18957 ( .A1(n15763), .A2(n19847), .B1(n15762), .B2(n19892), .ZN(
        n15764) );
  AOI211_X1 U18958 ( .C1(n19838), .C2(n15766), .A(n15765), .B(n15764), .ZN(
        n15767) );
  OAI211_X1 U18959 ( .C1(n15769), .C2(n19866), .A(n15768), .B(n15767), .ZN(
        P1_U2818) );
  NOR3_X1 U18960 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19891), .A3(n15770), 
        .ZN(n15773) );
  INV_X1 U18961 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20676) );
  INV_X1 U18962 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15771) );
  OAI22_X1 U18963 ( .A1(n15783), .A2(n20676), .B1(n15771), .B2(n15826), .ZN(
        n15772) );
  AOI211_X1 U18964 ( .C1(n19901), .C2(P1_EBX_REG_21__SCAN_IN), .A(n15773), .B(
        n15772), .ZN(n15777) );
  INV_X1 U18965 ( .A(n15774), .ZN(n15860) );
  AOI22_X1 U18966 ( .A1(n15860), .A2(n19873), .B1(n15775), .B2(n19880), .ZN(
        n15776) );
  OAI211_X1 U18967 ( .C1(n15864), .C2(n19906), .A(n15777), .B(n15776), .ZN(
        P1_U2819) );
  INV_X1 U18968 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20674) );
  OAI22_X1 U18969 ( .A1(n15872), .A2(n15826), .B1(n15865), .B2(n19906), .ZN(
        n15780) );
  OAI22_X1 U18970 ( .A1(n15866), .A2(n19847), .B1(n15778), .B2(n19892), .ZN(
        n15779) );
  AOI211_X1 U18971 ( .C1(P1_EBX_REG_20__SCAN_IN), .C2(n19901), .A(n15780), .B(
        n15779), .ZN(n15781) );
  OAI221_X1 U18972 ( .B1(n15783), .B2(n20674), .C1(n15783), .C2(n15782), .A(
        n15781), .ZN(P1_U2820) );
  NOR3_X1 U18973 ( .A1(n19891), .A2(n20671), .A3(n15788), .ZN(n15784) );
  AOI22_X1 U18974 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n19901), .B1(n15784), 
        .B2(n20672), .ZN(n15785) );
  OAI21_X1 U18975 ( .B1(n15879), .B2(n19906), .A(n15785), .ZN(n15786) );
  AOI211_X1 U18976 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19895), .B(n15786), .ZN(n15791) );
  INV_X1 U18977 ( .A(n15787), .ZN(n15876) );
  AOI22_X1 U18978 ( .A1(n15876), .A2(n19873), .B1(n15934), .B2(n19880), .ZN(
        n15790) );
  NOR3_X1 U18979 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n19891), .A3(n15788), 
        .ZN(n15792) );
  OAI21_X1 U18980 ( .B1(n15792), .B2(n15796), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15789) );
  NAND3_X1 U18981 ( .A1(n15791), .A2(n15790), .A3(n15789), .ZN(P1_U2821) );
  AOI211_X1 U18982 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15792), .B(n19895), .ZN(n15793) );
  OAI21_X1 U18983 ( .B1(n15794), .B2(n19866), .A(n15793), .ZN(n15795) );
  AOI21_X1 U18984 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15796), .A(n15795), 
        .ZN(n15801) );
  INV_X1 U18985 ( .A(n15797), .ZN(n15799) );
  AOI22_X1 U18986 ( .A1(n15799), .A2(n19873), .B1(n15798), .B2(n19838), .ZN(
        n15800) );
  OAI211_X1 U18987 ( .C1(n19892), .C2(n15802), .A(n15801), .B(n15800), .ZN(
        P1_U2822) );
  OAI21_X1 U18988 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15803), .ZN(n15804) );
  OAI22_X1 U18989 ( .A1(n14355), .A2(n15822), .B1(n15805), .B2(n15804), .ZN(
        n15806) );
  AOI211_X1 U18990 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19895), .B(n15806), .ZN(n15811) );
  OAI22_X1 U18991 ( .A1(n15807), .A2(n19847), .B1(n19892), .B2(n15952), .ZN(
        n15808) );
  AOI21_X1 U18992 ( .B1(n15809), .B2(n19838), .A(n15808), .ZN(n15810) );
  OAI211_X1 U18993 ( .C1(n15812), .C2(n19866), .A(n15811), .B(n15810), .ZN(
        P1_U2824) );
  AOI21_X1 U18994 ( .B1(n15813), .B2(n15840), .A(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n15823) );
  OAI22_X1 U18995 ( .A1(n15815), .A2(n19866), .B1(n19892), .B2(n15814), .ZN(
        n15816) );
  AOI211_X1 U18996 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n19895), .B(n15816), .ZN(n15821) );
  INV_X1 U18997 ( .A(n15817), .ZN(n15818) );
  AOI22_X1 U18998 ( .A1(n15819), .A2(n19873), .B1(n15818), .B2(n19838), .ZN(
        n15820) );
  OAI211_X1 U18999 ( .C1(n15823), .C2(n15822), .A(n15821), .B(n15820), .ZN(
        P1_U2826) );
  INV_X1 U19000 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20659) );
  NAND2_X1 U19001 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15834) );
  NOR2_X1 U19002 ( .A1(n20659), .A2(n15834), .ZN(n15824) );
  AOI21_X1 U19003 ( .B1(n15824), .B2(n15840), .A(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n15833) );
  OAI22_X1 U19004 ( .A1(n15827), .A2(n15826), .B1(n19892), .B2(n15825), .ZN(
        n15828) );
  AOI211_X1 U19005 ( .C1(n19901), .C2(P1_EBX_REG_12__SCAN_IN), .A(n19895), .B(
        n15828), .ZN(n15831) );
  INV_X1 U19006 ( .A(n15829), .ZN(n15897) );
  AOI22_X1 U19007 ( .A1(n15898), .A2(n19838), .B1(n19873), .B2(n15897), .ZN(
        n15830) );
  OAI211_X1 U19008 ( .C1(n15833), .C2(n15832), .A(n15831), .B(n15830), .ZN(
        P1_U2828) );
  OAI21_X1 U19009 ( .B1(n15834), .B2(n19832), .A(n19885), .ZN(n15849) );
  AOI22_X1 U19010 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n19901), .B1(n19880), 
        .B2(n15982), .ZN(n15837) );
  NOR3_X1 U19011 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15834), .A3(n19834), 
        .ZN(n15835) );
  AOI211_X1 U19012 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19895), .B(n15835), .ZN(n15836) );
  OAI211_X1 U19013 ( .C1(n15910), .C2(n19906), .A(n15837), .B(n15836), .ZN(
        n15838) );
  AOI21_X1 U19014 ( .B1(n19873), .B2(n15907), .A(n15838), .ZN(n15839) );
  OAI21_X1 U19015 ( .B1(n20659), .B2(n15849), .A(n15839), .ZN(P1_U2829) );
  NAND3_X1 U19016 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15840), .A3(n14388), 
        .ZN(n15844) );
  OAI22_X1 U19017 ( .A1(n15841), .A2(n19866), .B1(n19892), .B2(n15994), .ZN(
        n15842) );
  AOI211_X1 U19018 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19895), .B(n15842), .ZN(n15843) );
  OAI211_X1 U19019 ( .C1(n15845), .C2(n19847), .A(n15844), .B(n15843), .ZN(
        n15846) );
  AOI21_X1 U19020 ( .B1(n15847), .B2(n19838), .A(n15846), .ZN(n15848) );
  OAI21_X1 U19021 ( .B1(n14388), .B2(n15849), .A(n15848), .ZN(P1_U2830) );
  OAI22_X1 U19022 ( .A1(n15853), .A2(n9794), .B1(n15927), .B2(n19912), .ZN(
        n15850) );
  INV_X1 U19023 ( .A(n15850), .ZN(n15851) );
  OAI21_X1 U19024 ( .B1(n19919), .B2(n15852), .A(n15851), .ZN(P1_U2849) );
  AOI22_X1 U19025 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20033), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15858) );
  INV_X1 U19026 ( .A(n15853), .ZN(n15856) );
  XNOR2_X1 U19027 ( .A(n11179), .B(n21047), .ZN(n15854) );
  XNOR2_X1 U19028 ( .A(n15855), .B(n15854), .ZN(n15929) );
  AOI22_X1 U19029 ( .A1(n15856), .A2(n19993), .B1(n19994), .B2(n15929), .ZN(
        n15857) );
  OAI211_X1 U19030 ( .C1(n19998), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        P1_U2976) );
  AOI22_X1 U19031 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20033), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15863) );
  AOI22_X1 U19032 ( .A1(n15861), .A2(n19994), .B1(n19993), .B2(n15860), .ZN(
        n15862) );
  OAI211_X1 U19033 ( .C1(n19998), .C2(n15864), .A(n15863), .B(n15862), .ZN(
        P1_U2978) );
  OAI22_X1 U19034 ( .A1(n15866), .A2(n20044), .B1(n15865), .B2(n19998), .ZN(
        n15867) );
  AOI21_X1 U19035 ( .B1(n19994), .B2(n15868), .A(n15867), .ZN(n15870) );
  OAI211_X1 U19036 ( .C1(n15872), .C2(n15871), .A(n15870), .B(n15869), .ZN(
        P1_U2979) );
  AOI22_X1 U19037 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20033), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15878) );
  NOR2_X1 U19038 ( .A1(n11179), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15873) );
  MUX2_X1 U19039 ( .A(n11179), .B(n15873), .S(n13163), .Z(n15875) );
  XNOR2_X1 U19040 ( .A(n15875), .B(n15874), .ZN(n15935) );
  AOI22_X1 U19041 ( .A1(n15935), .A2(n19994), .B1(n19993), .B2(n15876), .ZN(
        n15877) );
  OAI211_X1 U19042 ( .C1(n19998), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        P1_U2980) );
  INV_X1 U19043 ( .A(n15880), .ZN(n15884) );
  INV_X1 U19044 ( .A(n15881), .ZN(n15883) );
  MUX2_X1 U19045 ( .A(n15884), .B(n15883), .S(n15882), .Z(n15885) );
  XNOR2_X1 U19046 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n15885), .ZN(
        n15949) );
  AOI22_X1 U19047 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20033), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15890) );
  INV_X1 U19048 ( .A(n15886), .ZN(n15888) );
  AOI22_X1 U19049 ( .A1(n15888), .A2(n19993), .B1(n15899), .B2(n15887), .ZN(
        n15889) );
  OAI211_X1 U19050 ( .C1(n19817), .C2(n15949), .A(n15890), .B(n15889), .ZN(
        P1_U2982) );
  XNOR2_X1 U19051 ( .A(n11179), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15891) );
  XNOR2_X1 U19052 ( .A(n15892), .B(n15891), .ZN(n15967) );
  AOI22_X1 U19053 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20033), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15896) );
  AOI22_X1 U19054 ( .A1(n15894), .A2(n19993), .B1(n15899), .B2(n15893), .ZN(
        n15895) );
  OAI211_X1 U19055 ( .C1(n15967), .C2(n19817), .A(n15896), .B(n15895), .ZN(
        P1_U2984) );
  AOI22_X1 U19056 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19986), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15901) );
  AOI22_X1 U19057 ( .A1(n15899), .A2(n15898), .B1(n19993), .B2(n15897), .ZN(
        n15900) );
  OAI211_X1 U19058 ( .C1(n15902), .C2(n19817), .A(n15901), .B(n15900), .ZN(
        P1_U2987) );
  AOI22_X1 U19059 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19986), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15909) );
  NAND3_X1 U19060 ( .A1(n15903), .A2(n11179), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15905) );
  NAND2_X1 U19061 ( .A1(n15905), .A2(n15904), .ZN(n15906) );
  XNOR2_X1 U19062 ( .A(n15906), .B(n15988), .ZN(n15985) );
  AOI22_X1 U19063 ( .A1(n19994), .A2(n15985), .B1(n19993), .B2(n15907), .ZN(
        n15908) );
  OAI211_X1 U19064 ( .C1(n19998), .C2(n15910), .A(n15909), .B(n15908), .ZN(
        P1_U2988) );
  AOI22_X1 U19065 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19986), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15916) );
  NAND2_X1 U19066 ( .A1(n15912), .A2(n15911), .ZN(n15913) );
  XNOR2_X1 U19067 ( .A(n15914), .B(n15913), .ZN(n16021) );
  AOI22_X1 U19068 ( .A1(n16021), .A2(n19994), .B1(n19993), .B2(n19861), .ZN(
        n15915) );
  OAI211_X1 U19069 ( .C1(n19998), .C2(n19859), .A(n15916), .B(n15915), .ZN(
        P1_U2992) );
  AOI22_X1 U19070 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19986), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15919) );
  AOI22_X1 U19071 ( .A1(n15917), .A2(n19994), .B1(n19993), .B2(n19874), .ZN(
        n15918) );
  OAI211_X1 U19072 ( .C1(n19998), .C2(n19876), .A(n15919), .B(n15918), .ZN(
        P1_U2993) );
  AOI22_X1 U19073 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19986), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15925) );
  OAI21_X1 U19074 ( .B1(n15922), .B2(n15921), .A(n15920), .ZN(n15923) );
  INV_X1 U19075 ( .A(n15923), .ZN(n16032) );
  AOI22_X1 U19076 ( .A1(n16032), .A2(n19994), .B1(n19993), .B2(n19916), .ZN(
        n15924) );
  OAI211_X1 U19077 ( .C1(n19998), .C2(n19889), .A(n15925), .B(n15924), .ZN(
        P1_U2994) );
  AOI22_X1 U19078 ( .A1(n20033), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n16014), 
        .B2(n15926), .ZN(n15931) );
  INV_X1 U19079 ( .A(n15927), .ZN(n15928) );
  AOI22_X1 U19080 ( .A1(n15929), .A2(n20031), .B1(n20027), .B2(n15928), .ZN(
        n15930) );
  OAI211_X1 U19081 ( .C1(n15932), .C2(n21047), .A(n15931), .B(n15930), .ZN(
        P1_U3008) );
  AOI22_X1 U19082 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15933), .B1(
        n20033), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15941) );
  AOI22_X1 U19083 ( .A1(n15935), .A2(n20031), .B1(n20027), .B2(n15934), .ZN(
        n15940) );
  OAI21_X1 U19084 ( .B1(n15938), .B2(n15937), .A(n15936), .ZN(n15939) );
  NAND3_X1 U19085 ( .A1(n15941), .A2(n15940), .A3(n15939), .ZN(P1_U3012) );
  OR2_X1 U19086 ( .A1(n20982), .A2(n15942), .ZN(n15962) );
  OAI21_X1 U19087 ( .B1(n15950), .B2(n15962), .A(n15943), .ZN(n15946) );
  AOI22_X1 U19088 ( .A1(n15946), .A2(n15945), .B1(n20027), .B2(n15944), .ZN(
        n15948) );
  NAND2_X1 U19089 ( .A1(n20033), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15947) );
  OAI211_X1 U19090 ( .C1(n15949), .C2(n15966), .A(n15948), .B(n15947), .ZN(
        P1_U3014) );
  INV_X1 U19091 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15957) );
  OAI21_X1 U19092 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15950), .ZN(n15951) );
  OAI22_X1 U19093 ( .A1(n15952), .A2(n20003), .B1(n15951), .B2(n15962), .ZN(
        n15953) );
  AOI21_X1 U19094 ( .B1(n20031), .B2(n15954), .A(n15953), .ZN(n15956) );
  NAND2_X1 U19095 ( .A1(n19986), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15955) );
  OAI211_X1 U19096 ( .C1(n15960), .C2(n15957), .A(n15956), .B(n15955), .ZN(
        P1_U3015) );
  INV_X1 U19097 ( .A(n15958), .ZN(n15964) );
  NAND2_X1 U19098 ( .A1(n19986), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15959) );
  OAI221_X1 U19099 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15962), 
        .C1(n15961), .C2(n15960), .A(n15959), .ZN(n15963) );
  AOI21_X1 U19100 ( .B1(n15964), .B2(n20027), .A(n15963), .ZN(n15965) );
  OAI21_X1 U19101 ( .B1(n15967), .B2(n15966), .A(n15965), .ZN(P1_U3016) );
  INV_X1 U19102 ( .A(n15968), .ZN(n15974) );
  NOR2_X1 U19103 ( .A1(n15970), .A2(n15969), .ZN(n15973) );
  NOR2_X1 U19104 ( .A1(n20002), .A2(n20662), .ZN(n15972) );
  AOI211_X1 U19105 ( .C1(n15974), .C2(n15973), .A(n15972), .B(n15971), .ZN(
        n15979) );
  INV_X1 U19106 ( .A(n15975), .ZN(n15977) );
  AOI22_X1 U19107 ( .A1(n15977), .A2(n20031), .B1(n20027), .B2(n15976), .ZN(
        n15978) );
  OAI211_X1 U19108 ( .C1(n15981), .C2(n15980), .A(n15979), .B(n15978), .ZN(
        P1_U3018) );
  AOI22_X1 U19109 ( .A1(n15982), .A2(n20027), .B1(n20033), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15987) );
  INV_X1 U19110 ( .A(n15983), .ZN(n15984) );
  AOI22_X1 U19111 ( .A1(n20031), .A2(n15985), .B1(n16014), .B2(n15984), .ZN(
        n15986) );
  OAI211_X1 U19112 ( .C1(n15989), .C2(n15988), .A(n15987), .B(n15986), .ZN(
        P1_U3020) );
  OAI21_X1 U19113 ( .B1(n20001), .B2(n15990), .A(n15993), .ZN(n15991) );
  OAI21_X1 U19114 ( .B1(n15992), .B2(n15991), .A(n16012), .ZN(n16009) );
  NAND2_X1 U19115 ( .A1(n15993), .A2(n16014), .ZN(n16005) );
  AOI221_X1 U19116 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14385), .C2(n16010), .A(
        n16005), .ZN(n15996) );
  OAI22_X1 U19117 ( .A1(n15994), .A2(n20003), .B1(n14388), .B2(n20002), .ZN(
        n15995) );
  AOI211_X1 U19118 ( .C1(n15997), .C2(n20031), .A(n15996), .B(n15995), .ZN(
        n15998) );
  OAI21_X1 U19119 ( .B1(n14385), .B2(n16009), .A(n15998), .ZN(P1_U3021) );
  INV_X1 U19120 ( .A(n15999), .ZN(n16007) );
  AND2_X1 U19121 ( .A1(n16001), .A2(n16000), .ZN(n16002) );
  NOR2_X1 U19122 ( .A1(n16003), .A2(n16002), .ZN(n19907) );
  AOI22_X1 U19123 ( .A1(n19907), .A2(n20027), .B1(n20033), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n16004) );
  OAI21_X1 U19124 ( .B1(n16005), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16004), .ZN(n16006) );
  AOI21_X1 U19125 ( .B1(n16007), .B2(n20031), .A(n16006), .ZN(n16008) );
  OAI21_X1 U19126 ( .B1(n16010), .B2(n16009), .A(n16008), .ZN(P1_U3022) );
  INV_X1 U19127 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16019) );
  NAND2_X1 U19128 ( .A1(n16012), .A2(n16011), .ZN(n16023) );
  INV_X1 U19129 ( .A(n16013), .ZN(n16017) );
  INV_X1 U19130 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16024) );
  NAND2_X1 U19131 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16014), .ZN(
        n16025) );
  AOI221_X1 U19132 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16019), .C2(n16024), .A(
        n16025), .ZN(n16016) );
  INV_X1 U19133 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21024) );
  OAI22_X1 U19134 ( .A1(n19844), .A2(n20003), .B1(n21024), .B2(n20002), .ZN(
        n16015) );
  AOI211_X1 U19135 ( .C1(n16017), .C2(n20031), .A(n16016), .B(n16015), .ZN(
        n16018) );
  OAI21_X1 U19136 ( .B1(n16019), .B2(n16023), .A(n16018), .ZN(P1_U3023) );
  INV_X1 U19137 ( .A(n19855), .ZN(n16020) );
  AOI222_X1 U19138 ( .A1(n16021), .A2(n20031), .B1(n20027), .B2(n16020), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(n19986), .ZN(n16022) );
  OAI221_X1 U19139 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16025), .C1(
        n16024), .C2(n16023), .A(n16022), .ZN(P1_U3024) );
  NOR2_X1 U19140 ( .A1(n16027), .A2(n16026), .ZN(n16028) );
  OR2_X1 U19141 ( .A1(n16029), .A2(n16028), .ZN(n19913) );
  INV_X1 U19142 ( .A(n19913), .ZN(n19879) );
  AOI22_X1 U19143 ( .A1(n19879), .A2(n20027), .B1(n20033), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16034) );
  INV_X1 U19144 ( .A(n16030), .ZN(n16031) );
  AOI22_X1 U19145 ( .A1(n16032), .A2(n20031), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16031), .ZN(n16033) );
  OAI211_X1 U19146 ( .C1(n20014), .C2(n16035), .A(n16034), .B(n16033), .ZN(
        P1_U3026) );
  AOI21_X1 U19147 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16044), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16042) );
  NAND4_X1 U19148 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n10613), .A4(n20726), .ZN(n16036) );
  AND2_X1 U19149 ( .A1(n16037), .A2(n16036), .ZN(n20628) );
  AOI21_X1 U19150 ( .B1(n20628), .B2(n16039), .A(n16038), .ZN(n16041) );
  AOI21_X1 U19151 ( .B1(n20704), .B2(n20726), .A(n20730), .ZN(n16040) );
  NOR3_X1 U19152 ( .A1(n16042), .A2(n16041), .A3(n16040), .ZN(P1_U3162) );
  OAI221_X1 U19153 ( .B1(n20704), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20704), 
        .C2(n16044), .A(n16043), .ZN(P1_U3466) );
  AOI22_X1 U19154 ( .A1(n18950), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18949), .ZN(n16055) );
  OAI22_X1 U19155 ( .A1(n16046), .A2(n18957), .B1(n16045), .B2(n18907), .ZN(
        n16047) );
  AOI21_X1 U19156 ( .B1(n16048), .B2(n18952), .A(n16047), .ZN(n16054) );
  OAI211_X1 U19157 ( .C1(n16051), .C2(n16050), .A(n18916), .B(n16049), .ZN(
        n16053) );
  NAND2_X1 U19158 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18928), .ZN(
        n16052) );
  NAND4_X1 U19159 ( .A1(n16055), .A2(n16054), .A3(n16053), .A4(n16052), .ZN(
        P2_U2825) );
  INV_X1 U19160 ( .A(n16059), .ZN(n16057) );
  INV_X1 U19161 ( .A(n16058), .ZN(n16056) );
  AOI221_X1 U19162 ( .B1(n16059), .B2(n16058), .C1(n16057), .C2(n16056), .A(
        n18967), .ZN(n16062) );
  INV_X1 U19163 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n20938) );
  OAI22_X1 U19164 ( .A1(n18925), .A2(n20938), .B1(n16060), .B2(n18961), .ZN(
        n16061) );
  AOI211_X1 U19165 ( .C1(n18949), .C2(P2_REIP_REG_29__SCAN_IN), .A(n16062), 
        .B(n16061), .ZN(n16066) );
  AOI22_X1 U19166 ( .A1(n16064), .A2(n18939), .B1(n18954), .B2(n16063), .ZN(
        n16065) );
  INV_X1 U19167 ( .A(n16068), .ZN(n16070) );
  AOI22_X1 U19168 ( .A1(n16070), .A2(n18939), .B1(n16069), .B2(n18952), .ZN(
        n16081) );
  OAI211_X1 U19169 ( .C1(n16073), .C2(n16072), .A(n18916), .B(n16071), .ZN(
        n16079) );
  AOI22_X1 U19170 ( .A1(n18949), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18928), .ZN(n16078) );
  NAND2_X1 U19171 ( .A1(n18950), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16077) );
  INV_X1 U19172 ( .A(n16074), .ZN(n16075) );
  NAND2_X1 U19173 ( .A1(n16075), .A2(n18954), .ZN(n16076) );
  AND4_X1 U19174 ( .A1(n16079), .A2(n16078), .A3(n16077), .A4(n16076), .ZN(
        n16080) );
  NAND2_X1 U19175 ( .A1(n16081), .A2(n16080), .ZN(P2_U2829) );
  AOI211_X1 U19176 ( .C1(n16084), .C2(n16083), .A(n16082), .B(n18967), .ZN(
        n16087) );
  OAI22_X1 U19177 ( .A1(n18926), .A2(n19731), .B1(n16085), .B2(n18925), .ZN(
        n16086) );
  AOI211_X1 U19178 ( .C1(n18928), .C2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16087), .B(n16086), .ZN(n16091) );
  AOI22_X1 U19179 ( .A1(n16089), .A2(n18954), .B1(n16088), .B2(n18939), .ZN(
        n16090) );
  OAI211_X1 U19180 ( .C1(n16092), .C2(n18920), .A(n16091), .B(n16090), .ZN(
        P2_U2830) );
  AOI22_X1 U19181 ( .A1(n19000), .A2(n16094), .B1(n16093), .B2(n18996), .ZN(
        P2_U2856) );
  INV_X1 U19182 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16098) );
  AOI22_X1 U19183 ( .A1(n16096), .A2(n18998), .B1(n19000), .B2(n16095), .ZN(
        n16097) );
  OAI21_X1 U19184 ( .B1(n19000), .B2(n16098), .A(n16097), .ZN(P2_U2864) );
  AOI22_X1 U19185 ( .A1(n16099), .A2(n18998), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n18996), .ZN(n16100) );
  OAI21_X1 U19186 ( .B1(n18996), .B2(n16101), .A(n16100), .ZN(P2_U2865) );
  OAI21_X1 U19187 ( .B1(n9884), .B2(n16103), .A(n16102), .ZN(n16104) );
  INV_X1 U19188 ( .A(n16104), .ZN(n16111) );
  AOI22_X1 U19189 ( .A1(n16111), .A2(n18998), .B1(n19000), .B2(n18756), .ZN(
        n16105) );
  OAI21_X1 U19190 ( .B1(n19000), .B2(n10070), .A(n16105), .ZN(P2_U2867) );
  AND2_X1 U19191 ( .A1(n16107), .A2(n16106), .ZN(n16108) );
  OR2_X1 U19192 ( .A1(n16108), .A2(n13754), .ZN(n16118) );
  OAI22_X1 U19193 ( .A1(n16118), .A2(n18992), .B1(n19000), .B2(n18783), .ZN(
        n16109) );
  INV_X1 U19194 ( .A(n16109), .ZN(n16110) );
  OAI21_X1 U19195 ( .B1(n18996), .B2(n18787), .A(n16110), .ZN(P2_U2869) );
  AOI22_X1 U19196 ( .A1(n19005), .A2(n19028), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19056), .ZN(n16114) );
  AOI22_X1 U19197 ( .A1(n19007), .A2(BUF1_REG_20__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16113) );
  AOI22_X1 U19198 ( .A1(n16111), .A2(n19038), .B1(n19057), .B2(n18755), .ZN(
        n16112) );
  NAND3_X1 U19199 ( .A1(n16114), .A2(n16113), .A3(n16112), .ZN(P2_U2899) );
  AOI22_X1 U19200 ( .A1(n19005), .A2(n16115), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19056), .ZN(n16122) );
  AOI22_X1 U19201 ( .A1(n19007), .A2(BUF1_REG_18__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16121) );
  INV_X1 U19202 ( .A(n16116), .ZN(n18786) );
  OAI22_X1 U19203 ( .A1(n16118), .A2(n19061), .B1(n16117), .B2(n18786), .ZN(
        n16119) );
  INV_X1 U19204 ( .A(n16119), .ZN(n16120) );
  NAND3_X1 U19205 ( .A1(n16122), .A2(n16121), .A3(n16120), .ZN(P2_U2901) );
  AOI22_X1 U19206 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19132), .ZN(n16129) );
  NAND2_X1 U19207 ( .A1(n16123), .A2(n19116), .ZN(n16126) );
  NAND2_X1 U19208 ( .A1(n16124), .A2(n19115), .ZN(n16125) );
  OAI211_X1 U19209 ( .C1(n15430), .C2(n18976), .A(n16126), .B(n16125), .ZN(
        n16127) );
  INV_X1 U19210 ( .A(n16127), .ZN(n16128) );
  OAI211_X1 U19211 ( .C1(n19120), .C2(n18822), .A(n16129), .B(n16128), .ZN(
        P2_U3000) );
  AOI22_X1 U19212 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19132), .B1(n16178), 
        .B2(n18841), .ZN(n16137) );
  NAND2_X1 U19213 ( .A1(n16131), .A2(n16130), .ZN(n16132) );
  XNOR2_X1 U19214 ( .A(n16133), .B(n16132), .ZN(n16193) );
  OAI21_X1 U19215 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16139), .A(
        n16134), .ZN(n16197) );
  OAI22_X1 U19216 ( .A1(n16193), .A2(n16179), .B1(n16197), .B2(n16181), .ZN(
        n16135) );
  AOI21_X1 U19217 ( .B1(n19114), .B2(n18842), .A(n16135), .ZN(n16136) );
  OAI211_X1 U19218 ( .C1(n16186), .C2(n16138), .A(n16137), .B(n16136), .ZN(
        P2_U3001) );
  AOI22_X1 U19219 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19132), .ZN(n16145) );
  NOR2_X1 U19220 ( .A1(n18983), .A2(n15430), .ZN(n16142) );
  NOR3_X1 U19221 ( .A1(n16140), .A2(n16139), .A3(n16181), .ZN(n16141) );
  AOI211_X1 U19222 ( .C1(n19116), .C2(n16143), .A(n16142), .B(n16141), .ZN(
        n16144) );
  OAI211_X1 U19223 ( .C1(n19120), .C2(n18852), .A(n16145), .B(n16144), .ZN(
        P2_U3002) );
  AOI22_X1 U19224 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19132), .B1(n16178), 
        .B2(n16146), .ZN(n16152) );
  OAI22_X1 U19225 ( .A1(n16148), .A2(n16181), .B1(n16147), .B2(n16179), .ZN(
        n16149) );
  AOI21_X1 U19226 ( .B1(n19114), .B2(n16150), .A(n16149), .ZN(n16151) );
  OAI211_X1 U19227 ( .C1(n16186), .C2(n16153), .A(n16152), .B(n16151), .ZN(
        P2_U3003) );
  AOI22_X1 U19228 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18885), .ZN(n16158) );
  OAI22_X1 U19229 ( .A1(n16154), .A2(n16179), .B1(n15430), .B2(n18985), .ZN(
        n16155) );
  AOI21_X1 U19230 ( .B1(n16156), .B2(n19115), .A(n16155), .ZN(n16157) );
  OAI211_X1 U19231 ( .C1(n19120), .C2(n18859), .A(n16158), .B(n16157), .ZN(
        P2_U3004) );
  AOI22_X1 U19232 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19132), .B1(n16178), 
        .B2(n18875), .ZN(n16163) );
  OAI22_X1 U19233 ( .A1(n16160), .A2(n16181), .B1(n16179), .B2(n16159), .ZN(
        n16161) );
  AOI21_X1 U19234 ( .B1(n19114), .B2(n18876), .A(n16161), .ZN(n16162) );
  OAI211_X1 U19235 ( .C1(n16186), .C2(n18869), .A(n16163), .B(n16162), .ZN(
        P2_U3005) );
  AOI22_X1 U19236 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19132), .ZN(n16169) );
  NOR2_X1 U19237 ( .A1(n16164), .A2(n16181), .ZN(n16167) );
  OAI22_X1 U19238 ( .A1(n16165), .A2(n16179), .B1(n15430), .B2(n18997), .ZN(
        n16166) );
  AOI21_X1 U19239 ( .B1(n16167), .B2(n15349), .A(n16166), .ZN(n16168) );
  OAI211_X1 U19240 ( .C1(n19120), .C2(n16170), .A(n16169), .B(n16168), .ZN(
        P2_U3006) );
  AOI22_X1 U19241 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19132), .ZN(n16177) );
  NAND2_X1 U19242 ( .A1(n16171), .A2(n19116), .ZN(n16173) );
  NAND2_X1 U19243 ( .A1(n9894), .A2(n19114), .ZN(n16172) );
  OAI211_X1 U19244 ( .C1(n16174), .C2(n16181), .A(n16173), .B(n16172), .ZN(
        n16175) );
  INV_X1 U19245 ( .A(n16175), .ZN(n16176) );
  OAI211_X1 U19246 ( .C1(n19120), .C2(n18899), .A(n16177), .B(n16176), .ZN(
        P2_U3008) );
  AOI22_X1 U19247 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19132), .B1(n16178), 
        .B2(n18914), .ZN(n16185) );
  OAI22_X1 U19248 ( .A1(n16182), .A2(n16181), .B1(n16180), .B2(n16179), .ZN(
        n16183) );
  AOI21_X1 U19249 ( .B1(n19114), .B2(n18915), .A(n16183), .ZN(n16184) );
  OAI211_X1 U19250 ( .C1(n16186), .C2(n18906), .A(n16185), .B(n16184), .ZN(
        P2_U3009) );
  AOI21_X1 U19251 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16187), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16188) );
  OAI22_X1 U19252 ( .A1(n16189), .A2(n16188), .B1(n16209), .B2(n18845), .ZN(
        n16195) );
  INV_X1 U19253 ( .A(n18842), .ZN(n16190) );
  OAI22_X1 U19254 ( .A1(n16193), .A2(n16192), .B1(n16191), .B2(n16190), .ZN(
        n16194) );
  AOI211_X1 U19255 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18885), .A(n16195), 
        .B(n16194), .ZN(n16196) );
  OAI21_X1 U19256 ( .B1(n16212), .B2(n16197), .A(n16196), .ZN(P2_U3033) );
  NOR2_X1 U19257 ( .A1(n19703), .A2(n18905), .ZN(n16200) );
  OAI22_X1 U19258 ( .A1(n16198), .A2(n13394), .B1(n16209), .B2(n18888), .ZN(
        n16199) );
  AOI211_X1 U19259 ( .C1(n16201), .C2(n13394), .A(n16200), .B(n16199), .ZN(
        n16205) );
  INV_X1 U19260 ( .A(n18889), .ZN(n16202) );
  AOI22_X1 U19261 ( .A1(n16203), .A2(n19130), .B1(n19121), .B2(n16202), .ZN(
        n16204) );
  OAI211_X1 U19262 ( .C1(n16212), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        P2_U3039) );
  INV_X1 U19263 ( .A(n16207), .ZN(n16215) );
  OAI21_X1 U19264 ( .B1(n16209), .B2(n19033), .A(n16208), .ZN(n16210) );
  AOI21_X1 U19265 ( .B1(n13263), .B2(n19121), .A(n16210), .ZN(n16211) );
  OAI21_X1 U19266 ( .B1(n16213), .B2(n16212), .A(n16211), .ZN(n16214) );
  AOI21_X1 U19267 ( .B1(n16215), .B2(n19130), .A(n16214), .ZN(n16216) );
  OAI221_X1 U19268 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16218), .C1(
        n13631), .C2(n16217), .A(n16216), .ZN(P2_U3043) );
  NAND2_X1 U19269 ( .A1(n19759), .A2(n12943), .ZN(n16220) );
  AOI21_X1 U19270 ( .B1(n16221), .B2(n16220), .A(n16219), .ZN(n16223) );
  NOR3_X1 U19271 ( .A1(n16224), .A2(n16223), .A3(n16222), .ZN(n16229) );
  NOR2_X1 U19272 ( .A1(n16226), .A2(n16225), .ZN(n19788) );
  OAI21_X1 U19273 ( .B1(n16227), .B2(n19788), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16228) );
  OAI211_X1 U19274 ( .C1(n16230), .C2(n18734), .A(n16229), .B(n16228), .ZN(
        P2_U3176) );
  INV_X1 U19275 ( .A(n18500), .ZN(n16232) );
  NOR2_X1 U19276 ( .A1(n15582), .A2(n16233), .ZN(n16241) );
  OAI21_X1 U19277 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17617), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16234) );
  OAI221_X1 U19278 ( .B1(n16278), .B2(n16235), .C1(n17617), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16234), .ZN(n16240) );
  OAI21_X1 U19279 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16278), .A(
        n16235), .ZN(n16238) );
  NAND2_X1 U19280 ( .A1(n17617), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16236) );
  OAI22_X1 U19281 ( .A1(n15582), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n16236), .B2(n16278), .ZN(n16237) );
  OAI21_X1 U19282 ( .B1(n16241), .B2(n16238), .A(n16237), .ZN(n16239) );
  OAI21_X1 U19283 ( .B1(n16241), .B2(n16240), .A(n16239), .ZN(n16287) );
  INV_X1 U19284 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18645) );
  NOR2_X1 U19285 ( .A1(n9800), .A2(n18645), .ZN(n16280) );
  NOR2_X1 U19286 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18720), .ZN(n17546) );
  NAND2_X2 U19287 ( .A1(n18315), .A2(n18364), .ZN(n18132) );
  OAI21_X1 U19288 ( .B1(n17457), .B2(n21011), .A(n18132), .ZN(n17561) );
  INV_X1 U19289 ( .A(n17561), .ZN(n17472) );
  OR2_X1 U19290 ( .A1(n16242), .A2(n17472), .ZN(n16258) );
  XOR2_X1 U19291 ( .A(n10110), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16244) );
  NOR2_X1 U19292 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17457), .ZN(
        n16269) );
  NOR2_X1 U19293 ( .A1(n21011), .A2(n17352), .ZN(n16421) );
  NAND3_X1 U19294 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(n16421), .ZN(n16418) );
  AOI22_X1 U19295 ( .A1(n17546), .A2(n16418), .B1(n18442), .B2(n16242), .ZN(
        n16243) );
  NAND2_X1 U19296 ( .A1(n16243), .A2(n17708), .ZN(n16270) );
  NOR2_X1 U19297 ( .A1(n16269), .A2(n16270), .ZN(n16257) );
  OAI22_X1 U19298 ( .A1(n16258), .A2(n16244), .B1(n16257), .B2(n10110), .ZN(
        n16245) );
  AOI211_X1 U19299 ( .C1(n17565), .C2(n16733), .A(n16280), .B(n16245), .ZN(
        n16251) );
  NOR2_X2 U19300 ( .A1(n18708), .A2(n16402), .ZN(n17698) );
  NAND2_X1 U19301 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16246), .ZN(
        n16247) );
  XNOR2_X1 U19302 ( .A(n16247), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16284) );
  NAND2_X1 U19303 ( .A1(n16248), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16249) );
  XNOR2_X1 U19304 ( .A(n16249), .B(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16283) );
  AOI22_X1 U19305 ( .A1(n17698), .A2(n16284), .B1(n17543), .B2(n16283), .ZN(
        n16250) );
  OAI211_X1 U19306 ( .C1(n17606), .C2(n16287), .A(n16251), .B(n16250), .ZN(
        P3_U2799) );
  NAND2_X1 U19307 ( .A1(n9792), .A2(n16252), .ZN(n16263) );
  NAND2_X1 U19308 ( .A1(n17543), .A2(n16253), .ZN(n16265) );
  NAND2_X1 U19309 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17378), .ZN(
        n17430) );
  NOR4_X1 U19310 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16254), .A3(
        n17715), .A4(n17430), .ZN(n16260) );
  XOR2_X1 U19311 ( .A(n9909), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(n16438) );
  AOI21_X1 U19312 ( .B1(n17565), .B2(n16438), .A(n16255), .ZN(n16256) );
  OAI221_X1 U19313 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16258), .C1(
        n10111), .C2(n16257), .A(n16256), .ZN(n16259) );
  AOI211_X1 U19314 ( .C1(n17618), .C2(n16261), .A(n16260), .B(n16259), .ZN(
        n16262) );
  AOI21_X1 U19315 ( .B1(n16291), .B2(n16279), .A(n16263), .ZN(n16267) );
  INV_X1 U19316 ( .A(n16264), .ZN(n16292) );
  AOI21_X1 U19317 ( .B1(n16292), .B2(n16279), .A(n16265), .ZN(n16266) );
  AOI211_X1 U19318 ( .C1(n17618), .C2(n16268), .A(n16267), .B(n16266), .ZN(
        n16275) );
  AOI21_X1 U19319 ( .B1(n10109), .B2(n16418), .A(n9909), .ZN(n16449) );
  OAI21_X1 U19320 ( .B1(n17565), .B2(n16269), .A(n16449), .ZN(n16273) );
  OAI221_X1 U19321 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16271), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18442), .A(n16270), .ZN(
        n16272) );
  NAND4_X1 U19322 ( .A1(n16275), .A2(n16274), .A3(n16273), .A4(n16272), .ZN(
        P3_U2801) );
  OAI21_X1 U19323 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17974), .A(
        n16276), .ZN(n16282) );
  NOR4_X1 U19324 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16279), .A3(
        n16278), .A4(n16277), .ZN(n16281) );
  AOI211_X1 U19325 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16282), .A(
        n16281), .B(n16280), .ZN(n16286) );
  AOI22_X1 U19326 ( .A1(n16284), .A2(n18019), .B1(n16283), .B2(n17888), .ZN(
        n16285) );
  OAI211_X1 U19327 ( .C1(n17942), .C2(n16287), .A(n16286), .B(n16285), .ZN(
        P3_U2831) );
  NAND2_X1 U19328 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18035), .ZN(n17355) );
  NAND2_X1 U19329 ( .A1(n17617), .A2(n17366), .ZN(n17365) );
  AOI22_X1 U19330 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17617), .B1(
        n15647), .B2(n16298), .ZN(n17348) );
  AOI22_X1 U19331 ( .A1(n17894), .A2(n16292), .B1(n18494), .B2(n16291), .ZN(
        n16293) );
  OAI211_X1 U19332 ( .C1(n16295), .C2(n16294), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n9800), .ZN(n16304) );
  AND2_X1 U19333 ( .A1(n17617), .A2(n17346), .ZN(n16300) );
  OAI22_X1 U19334 ( .A1(n17529), .A2(n17914), .B1(n17915), .B2(n9952), .ZN(
        n17820) );
  AOI21_X1 U19335 ( .B1(n16296), .B2(n17820), .A(n17743), .ZN(n17801) );
  NOR2_X1 U19336 ( .A1(n17801), .A2(n16297), .ZN(n17773) );
  OAI211_X1 U19337 ( .C1(n16300), .C2(n17773), .A(n16299), .B(n16298), .ZN(
        n16303) );
  OR3_X1 U19338 ( .A1(n16301), .A2(n17942), .A3(n17348), .ZN(n16302) );
  NAND4_X1 U19339 ( .A1(n17355), .A2(n16304), .A3(n16303), .A4(n16302), .ZN(
        P3_U2834) );
  NOR3_X1 U19340 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16306) );
  NOR4_X1 U19341 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16305) );
  NAND4_X1 U19342 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16306), .A3(n16305), .A4(
        U215), .ZN(U213) );
  INV_X1 U19343 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19066) );
  INV_X2 U19344 ( .A(U214), .ZN(n16349) );
  NOR2_X2 U19345 ( .A1(n16349), .A2(n16307), .ZN(n16341) );
  OAI222_X1 U19346 ( .A1(U212), .A2(n19066), .B1(n16352), .B2(n16308), .C1(
        U214), .C2(n16386), .ZN(U216) );
  INV_X1 U19347 ( .A(U212), .ZN(n16350) );
  AOI222_X1 U19348 ( .A1(n16349), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16341), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16350), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n16309) );
  INV_X1 U19349 ( .A(n16309), .ZN(U217) );
  INV_X1 U19350 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16311) );
  AOI22_X1 U19351 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16349), .ZN(n16310) );
  OAI21_X1 U19352 ( .B1(n16311), .B2(n16352), .A(n16310), .ZN(U218) );
  AOI22_X1 U19353 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16349), .ZN(n16312) );
  OAI21_X1 U19354 ( .B1(n14746), .B2(n16352), .A(n16312), .ZN(U219) );
  AOI22_X1 U19355 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16349), .ZN(n16313) );
  OAI21_X1 U19356 ( .B1(n19156), .B2(n16352), .A(n16313), .ZN(U220) );
  INV_X1 U19357 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16315) );
  AOI22_X1 U19358 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16349), .ZN(n16314) );
  OAI21_X1 U19359 ( .B1(n16315), .B2(n16352), .A(n16314), .ZN(U221) );
  AOI22_X1 U19360 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16349), .ZN(n16316) );
  OAI21_X1 U19361 ( .B1(n16317), .B2(n16352), .A(n16316), .ZN(U222) );
  AOI22_X1 U19362 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16349), .ZN(n16318) );
  OAI21_X1 U19363 ( .B1(n16319), .B2(n16352), .A(n16318), .ZN(U223) );
  AOI22_X1 U19364 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16349), .ZN(n16320) );
  OAI21_X1 U19365 ( .B1(n20970), .B2(n16352), .A(n16320), .ZN(U224) );
  INV_X1 U19366 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19172) );
  AOI22_X1 U19367 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16349), .ZN(n16321) );
  OAI21_X1 U19368 ( .B1(n19172), .B2(n16352), .A(n16321), .ZN(U225) );
  AOI222_X1 U19369 ( .A1(n16349), .A2(P1_DATAO_REG_21__SCAN_IN), .B1(n16341), 
        .B2(BUF1_REG_21__SCAN_IN), .C1(n16350), .C2(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n16322) );
  INV_X1 U19370 ( .A(n16322), .ZN(U226) );
  AOI222_X1 U19371 ( .A1(n16349), .A2(P1_DATAO_REG_20__SCAN_IN), .B1(n16341), 
        .B2(BUF1_REG_20__SCAN_IN), .C1(n16350), .C2(P2_DATAO_REG_20__SCAN_IN), 
        .ZN(n16323) );
  INV_X1 U19372 ( .A(n16323), .ZN(U227) );
  INV_X1 U19373 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n20853) );
  AOI22_X1 U19374 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n16341), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16349), .ZN(n16324) );
  OAI21_X1 U19375 ( .B1(n20853), .B2(U212), .A(n16324), .ZN(U228) );
  AOI22_X1 U19376 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16349), .ZN(n16325) );
  OAI21_X1 U19377 ( .B1(n16326), .B2(n16352), .A(n16325), .ZN(U229) );
  AOI222_X1 U19378 ( .A1(n16349), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n16341), 
        .B2(BUF1_REG_17__SCAN_IN), .C1(n16350), .C2(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n16327) );
  INV_X1 U19379 ( .A(n16327), .ZN(U230) );
  INV_X1 U19380 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16329) );
  AOI22_X1 U19381 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16349), .ZN(n16328) );
  OAI21_X1 U19382 ( .B1(n16329), .B2(n16352), .A(n16328), .ZN(U231) );
  INV_X1 U19383 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n19924) );
  AOI22_X1 U19384 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16341), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16350), .ZN(n16330) );
  OAI21_X1 U19385 ( .B1(n19924), .B2(U214), .A(n16330), .ZN(U232) );
  INV_X1 U19386 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16368) );
  AOI22_X1 U19387 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16341), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16349), .ZN(n16331) );
  OAI21_X1 U19388 ( .B1(n16368), .B2(U212), .A(n16331), .ZN(U233) );
  INV_X1 U19389 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16366) );
  AOI22_X1 U19390 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16341), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16349), .ZN(n16332) );
  OAI21_X1 U19391 ( .B1(n16366), .B2(U212), .A(n16332), .ZN(U234) );
  INV_X1 U19392 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n16333) );
  INV_X1 U19393 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20968) );
  INV_X1 U19394 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n20869) );
  OAI222_X1 U19395 ( .A1(U214), .A2(n16333), .B1(n16352), .B2(n20968), .C1(
        U212), .C2(n20869), .ZN(U235) );
  INV_X1 U19396 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16365) );
  AOI22_X1 U19397 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16341), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16349), .ZN(n16334) );
  OAI21_X1 U19398 ( .B1(n16365), .B2(U212), .A(n16334), .ZN(U236) );
  AOI22_X1 U19399 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16349), .ZN(n16335) );
  OAI21_X1 U19400 ( .B1(n21043), .B2(n16352), .A(n16335), .ZN(U237) );
  INV_X1 U19401 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16362) );
  AOI22_X1 U19402 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16341), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16349), .ZN(n16336) );
  OAI21_X1 U19403 ( .B1(n16362), .B2(U212), .A(n16336), .ZN(U238) );
  AOI22_X1 U19404 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16349), .ZN(n16337) );
  OAI21_X1 U19405 ( .B1(n16338), .B2(n16352), .A(n16337), .ZN(U239) );
  INV_X1 U19406 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n21027) );
  AOI22_X1 U19407 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16341), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16349), .ZN(n16339) );
  OAI21_X1 U19408 ( .B1(n21027), .B2(U212), .A(n16339), .ZN(U240) );
  INV_X1 U19409 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16359) );
  AOI22_X1 U19410 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16341), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16349), .ZN(n16340) );
  OAI21_X1 U19411 ( .B1(n16359), .B2(U212), .A(n16340), .ZN(U241) );
  INV_X1 U19412 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16358) );
  AOI22_X1 U19413 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16341), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16349), .ZN(n16342) );
  OAI21_X1 U19414 ( .B1(n16358), .B2(U212), .A(n16342), .ZN(U242) );
  AOI22_X1 U19415 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16349), .ZN(n16343) );
  OAI21_X1 U19416 ( .B1(n16344), .B2(n16352), .A(n16343), .ZN(U243) );
  INV_X1 U19417 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n20811) );
  INV_X1 U19418 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16345) );
  INV_X1 U19419 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n20956) );
  OAI222_X1 U19420 ( .A1(U214), .A2(n20811), .B1(n16352), .B2(n16345), .C1(
        U212), .C2(n20956), .ZN(U244) );
  AOI22_X1 U19421 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16349), .ZN(n16346) );
  OAI21_X1 U19422 ( .B1(n16347), .B2(n16352), .A(n16346), .ZN(U245) );
  INV_X1 U19423 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20881) );
  AOI22_X1 U19424 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16349), .ZN(n16348) );
  OAI21_X1 U19425 ( .B1(n20881), .B2(n16352), .A(n16348), .ZN(U246) );
  AOI22_X1 U19426 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16350), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16349), .ZN(n16351) );
  OAI21_X1 U19427 ( .B1(n16353), .B2(n16352), .A(n16351), .ZN(U247) );
  INV_X1 U19428 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16354) );
  AOI22_X1 U19429 ( .A1(n16384), .A2(n16354), .B1(n18054), .B2(U215), .ZN(U251) );
  OAI22_X1 U19430 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16384), .ZN(n16355) );
  INV_X1 U19431 ( .A(n16355), .ZN(U252) );
  INV_X1 U19432 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16356) );
  AOI22_X1 U19433 ( .A1(n16384), .A2(n16356), .B1(n18068), .B2(U215), .ZN(U253) );
  INV_X1 U19434 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U19435 ( .A1(n16384), .A2(n20956), .B1(n18074), .B2(U215), .ZN(U254) );
  INV_X1 U19436 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16357) );
  AOI22_X1 U19437 ( .A1(n16384), .A2(n16357), .B1(n18079), .B2(U215), .ZN(U255) );
  INV_X1 U19438 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18084) );
  AOI22_X1 U19439 ( .A1(n16384), .A2(n16358), .B1(n18084), .B2(U215), .ZN(U256) );
  INV_X1 U19440 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18090) );
  AOI22_X1 U19441 ( .A1(n16384), .A2(n16359), .B1(n18090), .B2(U215), .ZN(U257) );
  INV_X1 U19442 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20841) );
  AOI22_X1 U19443 ( .A1(n16384), .A2(n21027), .B1(n20841), .B2(U215), .ZN(U258) );
  INV_X1 U19444 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16360) );
  INV_X1 U19445 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U19446 ( .A1(n16384), .A2(n16360), .B1(n17203), .B2(U215), .ZN(U259) );
  INV_X1 U19447 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n16361) );
  AOI22_X1 U19448 ( .A1(n16378), .A2(n16362), .B1(n16361), .B2(U215), .ZN(U260) );
  INV_X1 U19449 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16363) );
  INV_X1 U19450 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U19451 ( .A1(n16378), .A2(n16363), .B1(n17193), .B2(U215), .ZN(U261) );
  INV_X1 U19452 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n16364) );
  AOI22_X1 U19453 ( .A1(n16384), .A2(n16365), .B1(n16364), .B2(U215), .ZN(U262) );
  INV_X1 U19454 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U19455 ( .A1(n16384), .A2(n20869), .B1(n17184), .B2(U215), .ZN(U263) );
  INV_X1 U19456 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U19457 ( .A1(n16384), .A2(n16366), .B1(n17179), .B2(U215), .ZN(U264) );
  INV_X1 U19458 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19459 ( .A1(n16378), .A2(n16368), .B1(n16367), .B2(U215), .ZN(U265) );
  OAI22_X1 U19460 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16384), .ZN(n16369) );
  INV_X1 U19461 ( .A(n16369), .ZN(U266) );
  OAI22_X1 U19462 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16378), .ZN(n16370) );
  INV_X1 U19463 ( .A(n16370), .ZN(U267) );
  INV_X1 U19464 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n20906) );
  INV_X1 U19465 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18063) );
  AOI22_X1 U19466 ( .A1(n16384), .A2(n20906), .B1(n18063), .B2(U215), .ZN(U268) );
  INV_X1 U19467 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n16371) );
  AOI22_X1 U19468 ( .A1(n16378), .A2(n16371), .B1(n18067), .B2(U215), .ZN(U269) );
  INV_X1 U19469 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18073) );
  AOI22_X1 U19470 ( .A1(n16384), .A2(n20853), .B1(n18073), .B2(U215), .ZN(U270) );
  OAI22_X1 U19471 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16384), .ZN(n16372) );
  INV_X1 U19472 ( .A(n16372), .ZN(U271) );
  OAI22_X1 U19473 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16378), .ZN(n16373) );
  INV_X1 U19474 ( .A(n16373), .ZN(U272) );
  INV_X1 U19475 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16374) );
  INV_X1 U19476 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19170) );
  AOI22_X1 U19477 ( .A1(n16378), .A2(n16374), .B1(n19170), .B2(U215), .ZN(U273) );
  OAI22_X1 U19478 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16378), .ZN(n16375) );
  INV_X1 U19479 ( .A(n16375), .ZN(U274) );
  INV_X1 U19480 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n16376) );
  AOI22_X1 U19481 ( .A1(n16378), .A2(n16376), .B1(n18058), .B2(U215), .ZN(U275) );
  INV_X1 U19482 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16377) );
  AOI22_X1 U19483 ( .A1(n16384), .A2(n16377), .B1(n14764), .B2(U215), .ZN(U276) );
  OAI22_X1 U19484 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16378), .ZN(n16379) );
  INV_X1 U19485 ( .A(n16379), .ZN(U277) );
  INV_X1 U19486 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16380) );
  INV_X1 U19487 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19155) );
  AOI22_X1 U19488 ( .A1(n16384), .A2(n16380), .B1(n19155), .B2(U215), .ZN(U278) );
  INV_X1 U19489 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16381) );
  INV_X1 U19490 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19161) );
  AOI22_X1 U19491 ( .A1(n16384), .A2(n16381), .B1(n19161), .B2(U215), .ZN(U279) );
  OAI22_X1 U19492 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16384), .ZN(n16382) );
  INV_X1 U19493 ( .A(n16382), .ZN(U280) );
  OAI22_X1 U19494 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16384), .ZN(n16383) );
  INV_X1 U19495 ( .A(n16383), .ZN(U281) );
  AOI22_X1 U19496 ( .A1(n16384), .A2(n19066), .B1(n18098), .B2(U215), .ZN(U282) );
  INV_X1 U19497 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16385) );
  AOI222_X1 U19498 ( .A1(n19066), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16386), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16385), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16387) );
  INV_X2 U19499 ( .A(n16389), .ZN(n16388) );
  INV_X1 U19500 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18605) );
  INV_X1 U19501 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19707) );
  AOI22_X1 U19502 ( .A1(n16388), .A2(n18605), .B1(n19707), .B2(n16389), .ZN(
        U347) );
  INV_X1 U19503 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18603) );
  INV_X1 U19504 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19706) );
  AOI22_X1 U19505 ( .A1(n16388), .A2(n18603), .B1(n19706), .B2(n16389), .ZN(
        U348) );
  INV_X1 U19506 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18600) );
  INV_X1 U19507 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19705) );
  AOI22_X1 U19508 ( .A1(n16388), .A2(n18600), .B1(n19705), .B2(n16389), .ZN(
        U349) );
  INV_X1 U19509 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18599) );
  INV_X1 U19510 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19704) );
  AOI22_X1 U19511 ( .A1(n16388), .A2(n18599), .B1(n19704), .B2(n16389), .ZN(
        U350) );
  INV_X1 U19512 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18597) );
  INV_X1 U19513 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20918) );
  AOI22_X1 U19514 ( .A1(n16388), .A2(n18597), .B1(n20918), .B2(n16389), .ZN(
        U351) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18594) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19701) );
  AOI22_X1 U19517 ( .A1(n16388), .A2(n18594), .B1(n19701), .B2(n16389), .ZN(
        U352) );
  INV_X1 U19518 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18593) );
  INV_X1 U19519 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19700) );
  AOI22_X1 U19520 ( .A1(n16388), .A2(n18593), .B1(n19700), .B2(n16389), .ZN(
        U353) );
  INV_X1 U19521 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18590) );
  AOI22_X1 U19522 ( .A1(n16388), .A2(n18590), .B1(n19699), .B2(n16389), .ZN(
        U354) );
  INV_X1 U19523 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18644) );
  INV_X1 U19524 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19742) );
  AOI22_X1 U19525 ( .A1(n16388), .A2(n18644), .B1(n19742), .B2(n16389), .ZN(
        U355) );
  INV_X1 U19526 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18641) );
  INV_X1 U19527 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19740) );
  AOI22_X1 U19528 ( .A1(n16388), .A2(n18641), .B1(n19740), .B2(n16389), .ZN(
        U356) );
  INV_X1 U19529 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18638) );
  INV_X1 U19530 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19738) );
  AOI22_X1 U19531 ( .A1(n16388), .A2(n18638), .B1(n19738), .B2(n16389), .ZN(
        U357) );
  INV_X1 U19532 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20983) );
  INV_X1 U19533 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19735) );
  AOI22_X1 U19534 ( .A1(n16388), .A2(n20983), .B1(n19735), .B2(n16389), .ZN(
        U358) );
  INV_X1 U19535 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18634) );
  INV_X1 U19536 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19734) );
  AOI22_X1 U19537 ( .A1(n16388), .A2(n18634), .B1(n19734), .B2(n16389), .ZN(
        U359) );
  INV_X1 U19538 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18632) );
  INV_X1 U19539 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19732) );
  AOI22_X1 U19540 ( .A1(n16388), .A2(n18632), .B1(n19732), .B2(n16389), .ZN(
        U360) );
  INV_X1 U19541 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18631) );
  INV_X1 U19542 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19730) );
  AOI22_X1 U19543 ( .A1(n16388), .A2(n18631), .B1(n19730), .B2(n16389), .ZN(
        U361) );
  INV_X1 U19544 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18628) );
  INV_X1 U19545 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19728) );
  AOI22_X1 U19546 ( .A1(n16388), .A2(n18628), .B1(n19728), .B2(n16389), .ZN(
        U362) );
  INV_X1 U19547 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18627) );
  INV_X1 U19548 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19726) );
  AOI22_X1 U19549 ( .A1(n16388), .A2(n18627), .B1(n19726), .B2(n16389), .ZN(
        U363) );
  INV_X1 U19550 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18625) );
  INV_X1 U19551 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19724) );
  AOI22_X1 U19552 ( .A1(n16388), .A2(n18625), .B1(n19724), .B2(n16389), .ZN(
        U364) );
  INV_X1 U19553 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18589) );
  INV_X1 U19554 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19698) );
  AOI22_X1 U19555 ( .A1(n16388), .A2(n18589), .B1(n19698), .B2(n16389), .ZN(
        U365) );
  INV_X1 U19556 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18624) );
  INV_X1 U19557 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19722) );
  AOI22_X1 U19558 ( .A1(n16388), .A2(n18624), .B1(n19722), .B2(n16389), .ZN(
        U366) );
  INV_X1 U19559 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18621) );
  INV_X1 U19560 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19720) );
  AOI22_X1 U19561 ( .A1(n16388), .A2(n18621), .B1(n19720), .B2(n16389), .ZN(
        U367) );
  INV_X1 U19562 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18620) );
  INV_X1 U19563 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19718) );
  AOI22_X1 U19564 ( .A1(n16388), .A2(n18620), .B1(n19718), .B2(n16389), .ZN(
        U368) );
  INV_X1 U19565 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18617) );
  INV_X1 U19566 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19716) );
  AOI22_X1 U19567 ( .A1(n16388), .A2(n18617), .B1(n19716), .B2(n16389), .ZN(
        U369) );
  INV_X1 U19568 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18616) );
  INV_X1 U19569 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19714) );
  AOI22_X1 U19570 ( .A1(n16388), .A2(n18616), .B1(n19714), .B2(n16389), .ZN(
        U370) );
  INV_X1 U19571 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18614) );
  INV_X1 U19572 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19712) );
  AOI22_X1 U19573 ( .A1(n16388), .A2(n18614), .B1(n19712), .B2(n16389), .ZN(
        U371) );
  INV_X1 U19574 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18611) );
  INV_X1 U19575 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19711) );
  AOI22_X1 U19576 ( .A1(n16388), .A2(n18611), .B1(n19711), .B2(n16389), .ZN(
        U372) );
  INV_X1 U19577 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18610) );
  INV_X1 U19578 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19710) );
  AOI22_X1 U19579 ( .A1(n16388), .A2(n18610), .B1(n19710), .B2(n16389), .ZN(
        U373) );
  INV_X1 U19580 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18608) );
  INV_X1 U19581 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19709) );
  AOI22_X1 U19582 ( .A1(n16388), .A2(n18608), .B1(n19709), .B2(n16389), .ZN(
        U374) );
  INV_X1 U19583 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18607) );
  INV_X1 U19584 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19708) );
  AOI22_X1 U19585 ( .A1(n16388), .A2(n18607), .B1(n19708), .B2(n16389), .ZN(
        U375) );
  INV_X1 U19586 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18588) );
  INV_X1 U19587 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19695) );
  AOI22_X1 U19588 ( .A1(n16388), .A2(n18588), .B1(n19695), .B2(n16389), .ZN(
        U376) );
  INV_X1 U19589 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16391) );
  INV_X1 U19590 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18586) );
  NAND2_X1 U19591 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18586), .ZN(n16390) );
  AOI22_X1 U19592 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n16390), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18584), .ZN(n18656) );
  OAI21_X1 U19593 ( .B1(n18584), .B2(n16391), .A(n18570), .ZN(P3_U2633) );
  NOR2_X1 U19594 ( .A1(n17281), .A2(n16392), .ZN(n16399) );
  OAI21_X1 U19595 ( .B1(n16399), .B2(n17277), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16393) );
  OAI21_X1 U19596 ( .B1(n16394), .B2(n18559), .A(n16393), .ZN(P3_U2634) );
  AOI21_X1 U19597 ( .B1(n18584), .B2(n18586), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16395) );
  AOI22_X1 U19598 ( .A1(n18652), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16395), 
        .B2(n18718), .ZN(P3_U2635) );
  OAI21_X1 U19599 ( .B1(n16396), .B2(BS16), .A(n18656), .ZN(n18654) );
  OAI21_X1 U19600 ( .B1(n18656), .B2(n16397), .A(n18654), .ZN(P3_U2636) );
  INV_X1 U19601 ( .A(n16398), .ZN(n16400) );
  NOR3_X1 U19602 ( .A1(n16401), .A2(n16400), .A3(n16399), .ZN(n18501) );
  INV_X1 U19603 ( .A(n18706), .ZN(n18550) );
  NOR2_X1 U19604 ( .A1(n18501), .A2(n18550), .ZN(n18700) );
  OAI21_X1 U19605 ( .B1(n18700), .B2(n16403), .A(n16402), .ZN(P3_U2637) );
  NOR4_X1 U19606 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16407) );
  NOR4_X1 U19607 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_14__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16406) );
  NOR4_X1 U19608 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16405) );
  NOR4_X1 U19609 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16404) );
  NAND4_X1 U19610 ( .A1(n16407), .A2(n16406), .A3(n16405), .A4(n16404), .ZN(
        n16413) );
  NOR4_X1 U19611 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16411) );
  AOI211_X1 U19612 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_27__SCAN_IN), .B(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16410) );
  NOR4_X1 U19613 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n16409) );
  NOR4_X1 U19614 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n16408) );
  NAND4_X1 U19615 ( .A1(n16411), .A2(n16410), .A3(n16409), .A4(n16408), .ZN(
        n16412) );
  NOR2_X1 U19616 ( .A1(n16413), .A2(n16412), .ZN(n18699) );
  INV_X1 U19617 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18650) );
  NOR3_X1 U19618 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16415) );
  OAI21_X1 U19619 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16415), .A(n18699), .ZN(
        n16414) );
  OAI21_X1 U19620 ( .B1(n18699), .B2(n18650), .A(n16414), .ZN(P3_U2638) );
  INV_X1 U19621 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18647) );
  NOR2_X1 U19622 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18693) );
  OAI21_X1 U19623 ( .B1(n16415), .B2(n18693), .A(n18699), .ZN(n16416) );
  OAI21_X1 U19624 ( .B1(n18699), .B2(n18647), .A(n16416), .ZN(P3_U2639) );
  INV_X1 U19625 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20842) );
  NAND3_X1 U19626 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(P3_REIP_REG_22__SCAN_IN), .ZN(n16431) );
  NAND2_X1 U19627 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16507), .ZN(n16499) );
  NOR2_X1 U19628 ( .A1(n20842), .A2(n16499), .ZN(n16476) );
  NAND2_X1 U19629 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16476), .ZN(n16475) );
  INV_X1 U19630 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18637) );
  INV_X1 U19631 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18635) );
  NOR2_X1 U19632 ( .A1(n18637), .A2(n18635), .ZN(n16457) );
  INV_X1 U19633 ( .A(n16457), .ZN(n16417) );
  NOR2_X1 U19634 ( .A1(n16475), .A2(n16417), .ZN(n16454) );
  NAND2_X1 U19635 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16454), .ZN(n16436) );
  NAND2_X1 U19636 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18645), .ZN(n16435) );
  NAND2_X1 U19637 ( .A1(n16518), .A2(n16517), .ZN(n16516) );
  NOR2_X1 U19638 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16516), .ZN(n16489) );
  NAND2_X1 U19639 ( .A1(n16489), .A2(n16496), .ZN(n16478) );
  NOR2_X1 U19640 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16478), .ZN(n16477) );
  INV_X1 U19641 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16472) );
  NAND2_X1 U19642 ( .A1(n16477), .A2(n16472), .ZN(n16471) );
  NOR2_X1 U19643 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16471), .ZN(n16458) );
  INV_X1 U19644 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16811) );
  NAND2_X1 U19645 ( .A1(n16458), .A2(n16811), .ZN(n16439) );
  NOR2_X1 U19646 ( .A1(n16770), .A2(n16439), .ZN(n16442) );
  INV_X1 U19647 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16430) );
  INV_X1 U19648 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17367) );
  INV_X1 U19649 ( .A(n16421), .ZN(n16420) );
  NOR2_X1 U19650 ( .A1(n17367), .A2(n16420), .ZN(n16419) );
  OAI21_X1 U19651 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16419), .A(
        n16418), .ZN(n17356) );
  INV_X1 U19652 ( .A(n17356), .ZN(n16461) );
  AOI21_X1 U19653 ( .B1(n17367), .B2(n16420), .A(n16419), .ZN(n17364) );
  INV_X1 U19654 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16422) );
  INV_X1 U19655 ( .A(n17392), .ZN(n17390) );
  NAND2_X1 U19656 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17390), .ZN(
        n16425) );
  NOR2_X1 U19657 ( .A1(n17393), .A2(n16425), .ZN(n17349) );
  INV_X1 U19658 ( .A(n17349), .ZN(n16423) );
  AOI21_X1 U19659 ( .B1(n16422), .B2(n16423), .A(n16421), .ZN(n17377) );
  INV_X1 U19660 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17406) );
  NOR2_X1 U19661 ( .A1(n17406), .A2(n16425), .ZN(n16424) );
  OAI21_X1 U19662 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16424), .A(
        n16423), .ZN(n17395) );
  INV_X1 U19663 ( .A(n17395), .ZN(n16493) );
  AOI21_X1 U19664 ( .B1(n17406), .B2(n16425), .A(n16424), .ZN(n17404) );
  OAI21_X1 U19665 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17389), .A(
        n16425), .ZN(n17420) );
  INV_X1 U19666 ( .A(n17420), .ZN(n16512) );
  NOR2_X1 U19667 ( .A1(n16426), .A2(n16764), .ZN(n16511) );
  NOR2_X1 U19668 ( .A1(n16512), .A2(n16511), .ZN(n16510) );
  NOR2_X1 U19669 ( .A1(n16510), .A2(n16764), .ZN(n16502) );
  NOR2_X1 U19670 ( .A1(n17404), .A2(n16502), .ZN(n16501) );
  NOR2_X1 U19671 ( .A1(n16501), .A2(n16764), .ZN(n16492) );
  NOR2_X1 U19672 ( .A1(n16493), .A2(n16492), .ZN(n16491) );
  NOR2_X1 U19673 ( .A1(n16491), .A2(n16764), .ZN(n16480) );
  NOR2_X1 U19674 ( .A1(n17377), .A2(n16480), .ZN(n16479) );
  NOR2_X1 U19675 ( .A1(n16479), .A2(n16764), .ZN(n16468) );
  NOR2_X1 U19676 ( .A1(n17364), .A2(n16468), .ZN(n16467) );
  NOR2_X1 U19677 ( .A1(n16467), .A2(n16764), .ZN(n16460) );
  NOR2_X1 U19678 ( .A1(n16461), .A2(n16460), .ZN(n16459) );
  NOR2_X1 U19679 ( .A1(n16459), .A2(n16764), .ZN(n16448) );
  NOR2_X1 U19680 ( .A1(n16449), .A2(n16448), .ZN(n16447) );
  NOR2_X1 U19681 ( .A1(n16447), .A2(n16764), .ZN(n16437) );
  NOR4_X1 U19682 ( .A1(n16438), .A2(n16437), .A3(n16764), .A4(n18565), .ZN(
        n16429) );
  INV_X1 U19683 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16427) );
  OAI22_X1 U19684 ( .A1(n10110), .A2(n16745), .B1(n16427), .B2(n16767), .ZN(
        n16428) );
  AOI211_X1 U19685 ( .C1(n16442), .C2(n16430), .A(n16429), .B(n16428), .ZN(
        n16434) );
  NOR2_X1 U19686 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16436), .ZN(n16441) );
  NOR2_X1 U19687 ( .A1(n16431), .A2(n16536), .ZN(n16500) );
  NAND2_X1 U19688 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16500), .ZN(n16490) );
  NAND2_X1 U19689 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16432) );
  OAI21_X1 U19690 ( .B1(n16490), .B2(n16432), .A(n16777), .ZN(n16485) );
  OAI221_X1 U19691 ( .B1(n16581), .B2(n16457), .C1(n16581), .C2(
        P3_REIP_REG_29__SCAN_IN), .A(n16485), .ZN(n16446) );
  OAI21_X1 U19692 ( .B1(n16441), .B2(n16446), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16433) );
  OAI211_X1 U19693 ( .C1(n16436), .C2(n16435), .A(n16434), .B(n16433), .ZN(
        P3_U2640) );
  XNOR2_X1 U19694 ( .A(n16438), .B(n16437), .ZN(n16445) );
  NAND2_X1 U19695 ( .A1(n16749), .A2(n16439), .ZN(n16450) );
  OAI22_X1 U19696 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16450), .B1(n10111), 
        .B2(n16745), .ZN(n16440) );
  AOI211_X1 U19697 ( .C1(P3_REIP_REG_30__SCAN_IN), .C2(n16446), .A(n16441), 
        .B(n16440), .ZN(n16444) );
  OAI21_X1 U19698 ( .B1(n16722), .B2(n16442), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16443) );
  OAI211_X1 U19699 ( .C1(n18565), .C2(n16445), .A(n16444), .B(n16443), .ZN(
        P3_U2641) );
  AOI22_X1 U19700 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16446), .B1(n16722), 
        .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16456) );
  INV_X1 U19701 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18640) );
  AOI211_X1 U19702 ( .C1(n16449), .C2(n16448), .A(n16447), .B(n18565), .ZN(
        n16453) );
  INV_X1 U19703 ( .A(n16458), .ZN(n16451) );
  AOI21_X1 U19704 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16451), .A(n16450), .ZN(
        n16452) );
  AOI211_X1 U19705 ( .C1(n16454), .C2(n18640), .A(n16453), .B(n16452), .ZN(
        n16455) );
  OAI211_X1 U19706 ( .C1(n10109), .C2(n16745), .A(n16456), .B(n16455), .ZN(
        P3_U2642) );
  AOI22_X1 U19707 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16765), .B1(
        n16722), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16466) );
  AOI211_X1 U19708 ( .C1(n18637), .C2(n18635), .A(n16457), .B(n16475), .ZN(
        n16464) );
  AOI211_X1 U19709 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16471), .A(n16458), .B(
        n16770), .ZN(n16463) );
  AOI211_X1 U19710 ( .C1(n16461), .C2(n16460), .A(n16459), .B(n18565), .ZN(
        n16462) );
  NOR3_X1 U19711 ( .A1(n16464), .A2(n16463), .A3(n16462), .ZN(n16465) );
  OAI211_X1 U19712 ( .C1(n18637), .C2(n16485), .A(n16466), .B(n16465), .ZN(
        P3_U2643) );
  AOI211_X1 U19713 ( .C1(n17364), .C2(n16468), .A(n16467), .B(n18565), .ZN(
        n16470) );
  OAI22_X1 U19714 ( .A1(n18635), .A2(n16485), .B1(n16767), .B2(n16472), .ZN(
        n16469) );
  AOI211_X1 U19715 ( .C1(n16765), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16470), .B(n16469), .ZN(n16474) );
  OAI211_X1 U19716 ( .C1(n16477), .C2(n16472), .A(n16749), .B(n16471), .ZN(
        n16473) );
  OAI211_X1 U19717 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16475), .A(n16474), 
        .B(n16473), .ZN(P3_U2644) );
  NOR2_X1 U19718 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16476), .ZN(n16486) );
  AOI22_X1 U19719 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16765), .B1(
        n16722), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16484) );
  AOI211_X1 U19720 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16478), .A(n16477), .B(
        n16770), .ZN(n16482) );
  AOI211_X1 U19721 ( .C1(n17377), .C2(n16480), .A(n16479), .B(n18565), .ZN(
        n16481) );
  NOR2_X1 U19722 ( .A1(n16482), .A2(n16481), .ZN(n16483) );
  OAI211_X1 U19723 ( .C1(n16486), .C2(n16485), .A(n16484), .B(n16483), .ZN(
        P3_U2645) );
  INV_X1 U19724 ( .A(n16489), .ZN(n16487) );
  OAI21_X1 U19725 ( .B1(n16770), .B2(n16487), .A(n16767), .ZN(n16488) );
  AOI22_X1 U19726 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16765), .B1(
        P3_EBX_REG_25__SCAN_IN), .B2(n16488), .ZN(n16498) );
  NOR2_X1 U19727 ( .A1(n16489), .A2(n16770), .ZN(n16503) );
  AND3_X1 U19728 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16777), .A3(n16490), 
        .ZN(n16495) );
  AOI211_X1 U19729 ( .C1(n16493), .C2(n16492), .A(n16491), .B(n18565), .ZN(
        n16494) );
  AOI211_X1 U19730 ( .C1(n16503), .C2(n16496), .A(n16495), .B(n16494), .ZN(
        n16497) );
  OAI211_X1 U19731 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16499), .A(n16498), 
        .B(n16497), .ZN(P3_U2646) );
  NOR2_X1 U19732 ( .A1(n16581), .A2(n16500), .ZN(n16515) );
  AOI22_X1 U19733 ( .A1(n16722), .A2(P3_EBX_REG_24__SCAN_IN), .B1(
        P3_REIP_REG_24__SCAN_IN), .B2(n16515), .ZN(n16509) );
  INV_X1 U19734 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18630) );
  AOI211_X1 U19735 ( .C1(n17404), .C2(n16502), .A(n16501), .B(n18565), .ZN(
        n16506) );
  INV_X1 U19736 ( .A(n16503), .ZN(n16504) );
  AOI21_X1 U19737 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16516), .A(n16504), .ZN(
        n16505) );
  AOI211_X1 U19738 ( .C1(n16507), .C2(n18630), .A(n16506), .B(n16505), .ZN(
        n16508) );
  OAI211_X1 U19739 ( .C1(n17406), .C2(n16745), .A(n16509), .B(n16508), .ZN(
        P3_U2647) );
  AOI22_X1 U19740 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16765), .B1(
        n16722), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16521) );
  INV_X1 U19741 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20836) );
  NOR3_X1 U19742 ( .A1(n18626), .A2(n16532), .A3(n20836), .ZN(n16514) );
  INV_X1 U19743 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18629) );
  AOI211_X1 U19744 ( .C1(n16512), .C2(n16511), .A(n16510), .B(n18565), .ZN(
        n16513) );
  AOI221_X1 U19745 ( .B1(n16515), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n16514), 
        .C2(n18629), .A(n16513), .ZN(n16520) );
  OAI211_X1 U19746 ( .C1(n16518), .C2(n16517), .A(n16749), .B(n16516), .ZN(
        n16519) );
  NAND3_X1 U19747 ( .A1(n16521), .A2(n16520), .A3(n16519), .ZN(P3_U2648) );
  INV_X1 U19748 ( .A(n16534), .ZN(n16522) );
  AOI21_X1 U19749 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16522), .A(n16770), .ZN(
        n16530) );
  AOI211_X1 U19750 ( .C1(n16525), .C2(n16524), .A(n16523), .B(n18565), .ZN(
        n16528) );
  INV_X1 U19751 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17447) );
  OAI22_X1 U19752 ( .A1(n17447), .A2(n16745), .B1(n16767), .B2(n16526), .ZN(
        n16527) );
  AOI211_X1 U19753 ( .C1(n16530), .C2(n16529), .A(n16528), .B(n16527), .ZN(
        n16531) );
  OAI221_X1 U19754 ( .B1(n16533), .B2(n18626), .C1(n16533), .C2(n16532), .A(
        n16531), .ZN(P3_U2650) );
  AOI211_X1 U19755 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16553), .A(n16534), .B(
        n16770), .ZN(n16535) );
  AOI21_X1 U19756 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16722), .A(n16535), .ZN(
        n16543) );
  AND2_X1 U19757 ( .A1(n16777), .A2(n16536), .ZN(n16541) );
  INV_X1 U19758 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18623) );
  AOI211_X1 U19759 ( .C1(n17461), .C2(n16538), .A(n16537), .B(n18565), .ZN(
        n16539) );
  AOI221_X1 U19760 ( .B1(n16541), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n16540), 
        .C2(n18623), .A(n16539), .ZN(n16542) );
  OAI211_X1 U19761 ( .C1(n10097), .C2(n16745), .A(n16543), .B(n16542), .ZN(
        P3_U2651) );
  NAND2_X1 U19762 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17470), .ZN(
        n16557) );
  INV_X1 U19763 ( .A(n16557), .ZN(n16545) );
  OAI21_X1 U19764 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16545), .A(
        n16544), .ZN(n17476) );
  NAND2_X1 U19765 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17562), .ZN(
        n17545) );
  INV_X1 U19766 ( .A(n17545), .ZN(n16639) );
  AND2_X1 U19767 ( .A1(n17504), .A2(n16639), .ZN(n17507) );
  NAND2_X1 U19768 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17507), .ZN(
        n16589) );
  OAI21_X1 U19769 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16589), .A(
        n16733), .ZN(n16591) );
  OAI21_X1 U19770 ( .B1(n16545), .B2(n16764), .A(n16591), .ZN(n16546) );
  XNOR2_X1 U19771 ( .A(n17476), .B(n16546), .ZN(n16552) );
  OAI21_X1 U19772 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), 
        .A(n16547), .ZN(n16550) );
  NOR2_X1 U19773 ( .A1(n16581), .A2(n16548), .ZN(n16567) );
  AOI22_X1 U19774 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16765), .B1(
        P3_REIP_REG_19__SCAN_IN), .B2(n16567), .ZN(n16549) );
  OAI211_X1 U19775 ( .C1(n16561), .C2(n16550), .A(n16549), .B(n9800), .ZN(
        n16551) );
  AOI21_X1 U19776 ( .B1(n16552), .B2(n16753), .A(n16551), .ZN(n16555) );
  OAI211_X1 U19777 ( .C1(n16559), .C2(n16556), .A(n16749), .B(n16553), .ZN(
        n16554) );
  OAI211_X1 U19778 ( .C1(n16556), .C2(n16767), .A(n16555), .B(n16554), .ZN(
        P3_U2652) );
  OAI21_X1 U19779 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17470), .A(
        n16557), .ZN(n17481) );
  OAI21_X1 U19780 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16568), .A(
        n16733), .ZN(n16558) );
  XNOR2_X1 U19781 ( .A(n17481), .B(n16558), .ZN(n16565) );
  AOI211_X1 U19782 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16574), .A(n16559), .B(
        n16770), .ZN(n16563) );
  AOI22_X1 U19783 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16765), .B1(
        P3_REIP_REG_18__SCAN_IN), .B2(n16567), .ZN(n16560) );
  OAI211_X1 U19784 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(n16561), .A(n16560), 
        .B(n9800), .ZN(n16562) );
  AOI211_X1 U19785 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16722), .A(n16563), .B(
        n16562), .ZN(n16564) );
  OAI21_X1 U19786 ( .B1(n18565), .B2(n16565), .A(n16564), .ZN(P3_U2653) );
  INV_X1 U19787 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18613) );
  NOR2_X1 U19788 ( .A1(n16566), .A2(n18613), .ZN(n16584) );
  AOI21_X1 U19789 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16584), .A(
        P3_REIP_REG_17__SCAN_IN), .ZN(n16572) );
  INV_X1 U19790 ( .A(n16567), .ZN(n16571) );
  AOI21_X1 U19791 ( .B1(n17491), .B2(n16754), .A(n16764), .ZN(n16569) );
  AND2_X1 U19792 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17491), .ZN(
        n16582) );
  OAI21_X1 U19793 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16582), .A(
        n16568), .ZN(n17492) );
  XOR2_X1 U19794 ( .A(n16569), .B(n17492), .Z(n16570) );
  OAI22_X1 U19795 ( .A1(n16572), .A2(n16571), .B1(n18565), .B2(n16570), .ZN(
        n16573) );
  AOI211_X1 U19796 ( .C1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n16765), .A(
        n18035), .B(n16573), .ZN(n16576) );
  OAI211_X1 U19797 ( .C1(n16578), .C2(n16577), .A(n16749), .B(n16574), .ZN(
        n16575) );
  OAI211_X1 U19798 ( .C1(n16577), .C2(n16767), .A(n16576), .B(n16575), .ZN(
        P3_U2654) );
  AOI211_X1 U19799 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16597), .A(n16578), .B(
        n16770), .ZN(n16579) );
  AOI21_X1 U19800 ( .B1(n16765), .B2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16579), .ZN(n16588) );
  INV_X1 U19801 ( .A(n16580), .ZN(n16607) );
  AOI21_X1 U19802 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16607), .A(n16581), 
        .ZN(n16595) );
  AOI22_X1 U19803 ( .A1(n16722), .A2(P3_EBX_REG_16__SCAN_IN), .B1(
        P3_REIP_REG_16__SCAN_IN), .B2(n16595), .ZN(n16587) );
  INV_X1 U19804 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16583) );
  AOI21_X1 U19805 ( .B1(n16583), .B2(n16589), .A(n16582), .ZN(n17508) );
  XNOR2_X1 U19806 ( .A(n17508), .B(n16591), .ZN(n16585) );
  INV_X1 U19807 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18615) );
  AOI22_X1 U19808 ( .A1(n16585), .A2(n16753), .B1(n16584), .B2(n18615), .ZN(
        n16586) );
  NAND4_X1 U19809 ( .A1(n16588), .A2(n16587), .A3(n16586), .A4(n9800), .ZN(
        P3_U2655) );
  AOI21_X1 U19810 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n16765), .A(
        n18035), .ZN(n16602) );
  NAND2_X1 U19811 ( .A1(n16753), .A2(n16764), .ZN(n16757) );
  OAI21_X1 U19812 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17507), .A(
        n16589), .ZN(n17515) );
  NAND2_X1 U19813 ( .A1(n16733), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16590) );
  NAND2_X1 U19814 ( .A1(n16753), .A2(n16590), .ZN(n16776) );
  AOI211_X1 U19815 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16757), .A(
        n17515), .B(n16776), .ZN(n16594) );
  INV_X1 U19816 ( .A(n17515), .ZN(n16592) );
  NOR3_X1 U19817 ( .A1(n16592), .A2(n18565), .A3(n16591), .ZN(n16593) );
  AOI211_X1 U19818 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16722), .A(n16594), .B(
        n16593), .ZN(n16601) );
  OAI21_X1 U19819 ( .B1(n16596), .B2(P3_REIP_REG_15__SCAN_IN), .A(n16595), 
        .ZN(n16600) );
  OAI211_X1 U19820 ( .C1(n16603), .C2(n16598), .A(n16749), .B(n16597), .ZN(
        n16599) );
  NAND4_X1 U19821 ( .A1(n16602), .A2(n16601), .A3(n16600), .A4(n16599), .ZN(
        P3_U2656) );
  INV_X1 U19822 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16923) );
  AOI211_X1 U19823 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16619), .A(n16603), .B(
        n16770), .ZN(n16609) );
  NOR2_X1 U19824 ( .A1(n16768), .A2(n16604), .ZN(n16613) );
  AOI22_X1 U19825 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16777), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(n16613), .ZN(n16606) );
  INV_X1 U19826 ( .A(n17534), .ZN(n17551) );
  NAND2_X1 U19827 ( .A1(n17551), .A2(n16639), .ZN(n16612) );
  AOI21_X1 U19828 ( .B1(n17533), .B2(n16612), .A(n17507), .ZN(n17536) );
  OAI21_X1 U19829 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16612), .A(
        n16733), .ZN(n16611) );
  XOR2_X1 U19830 ( .A(n17536), .B(n16611), .Z(n16605) );
  OAI22_X1 U19831 ( .A1(n16607), .A2(n16606), .B1(n18565), .B2(n16605), .ZN(
        n16608) );
  AOI211_X1 U19832 ( .C1(n16765), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16609), .B(n16608), .ZN(n16610) );
  OAI211_X1 U19833 ( .C1(n16767), .C2(n16923), .A(n16610), .B(n9800), .ZN(
        P3_U2657) );
  INV_X1 U19834 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16623) );
  NOR2_X1 U19835 ( .A1(n16611), .A2(n18565), .ZN(n16618) );
  INV_X1 U19836 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16629) );
  NOR2_X1 U19837 ( .A1(n16629), .A2(n17545), .ZN(n16628) );
  OAI21_X1 U19838 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16628), .A(
        n16612), .ZN(n17548) );
  AOI211_X1 U19839 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16733), .A(
        n17548), .B(n16776), .ZN(n16617) );
  INV_X1 U19840 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20904) );
  OAI21_X1 U19841 ( .B1(n16768), .B2(n16625), .A(n16779), .ZN(n16637) );
  AOI21_X1 U19842 ( .B1(n16761), .B2(n20904), .A(n16637), .ZN(n16615) );
  AOI22_X1 U19843 ( .A1(n16722), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n16613), 
        .B2(n18609), .ZN(n16614) );
  OAI211_X1 U19844 ( .C1(n16615), .C2(n18609), .A(n16614), .B(n9800), .ZN(
        n16616) );
  AOI211_X1 U19845 ( .C1(n16618), .C2(n17548), .A(n16617), .B(n16616), .ZN(
        n16622) );
  OAI211_X1 U19846 ( .C1(n16626), .C2(n16620), .A(n16749), .B(n16619), .ZN(
        n16621) );
  OAI211_X1 U19847 ( .C1(n16745), .C2(n16623), .A(n16622), .B(n16621), .ZN(
        P3_U2658) );
  NOR2_X1 U19848 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16768), .ZN(n16624) );
  AOI22_X1 U19849 ( .A1(n16722), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16625), 
        .B2(n16624), .ZN(n16634) );
  AOI211_X1 U19850 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16646), .A(n16626), .B(
        n16770), .ZN(n16627) );
  AOI211_X1 U19851 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n16765), .A(
        n18035), .B(n16627), .ZN(n16633) );
  AOI21_X1 U19852 ( .B1(n16629), .B2(n17545), .A(n16628), .ZN(n17564) );
  NAND3_X1 U19853 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17623), .A3(
        n16754), .ZN(n16655) );
  NAND2_X1 U19854 ( .A1(n16733), .A2(n16655), .ZN(n16679) );
  OAI21_X1 U19855 ( .B1(n9912), .B2(n16764), .A(n16679), .ZN(n16630) );
  XOR2_X1 U19856 ( .A(n17564), .B(n16630), .Z(n16631) );
  AOI22_X1 U19857 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16637), .B1(n16753), 
        .B2(n16631), .ZN(n16632) );
  NAND3_X1 U19858 ( .A1(n16634), .A2(n16633), .A3(n16632), .ZN(P3_U2659) );
  INV_X1 U19859 ( .A(n16635), .ZN(n16636) );
  NOR3_X1 U19860 ( .A1(n16768), .A2(n16707), .A3(n16652), .ZN(n16704) );
  AOI21_X1 U19861 ( .B1(n16636), .B2(n16704), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16644) );
  INV_X1 U19862 ( .A(n16637), .ZN(n16643) );
  INV_X1 U19863 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20917) );
  INV_X1 U19864 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17587) );
  NAND2_X1 U19865 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16638) );
  NOR2_X1 U19866 ( .A1(n21011), .A2(n17637), .ZN(n16708) );
  INV_X1 U19867 ( .A(n16708), .ZN(n16699) );
  NOR2_X1 U19868 ( .A1(n17645), .A2(n16699), .ZN(n16698) );
  NAND2_X1 U19869 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16698), .ZN(
        n16685) );
  OR2_X1 U19870 ( .A1(n16638), .A2(n16685), .ZN(n16663) );
  NOR2_X1 U19871 ( .A1(n17587), .A2(n16663), .ZN(n16654) );
  INV_X1 U19872 ( .A(n16654), .ZN(n16640) );
  AOI21_X1 U19873 ( .B1(n20917), .B2(n16640), .A(n16639), .ZN(n17572) );
  OAI21_X1 U19874 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16640), .A(
        n16733), .ZN(n16641) );
  XOR2_X1 U19875 ( .A(n17572), .B(n16641), .Z(n16642) );
  OAI22_X1 U19876 ( .A1(n16644), .A2(n16643), .B1(n18565), .B2(n16642), .ZN(
        n16645) );
  AOI211_X1 U19877 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n16765), .A(
        n18035), .B(n16645), .ZN(n16648) );
  OAI211_X1 U19878 ( .C1(n16649), .C2(n16997), .A(n16749), .B(n16646), .ZN(
        n16647) );
  OAI211_X1 U19879 ( .C1(n16997), .C2(n16767), .A(n16648), .B(n16647), .ZN(
        P3_U2660) );
  AOI211_X1 U19880 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16650), .A(n16649), .B(
        n16770), .ZN(n16651) );
  AOI211_X1 U19881 ( .C1(n16722), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18035), .B(
        n16651), .ZN(n16660) );
  OR2_X1 U19882 ( .A1(n16707), .A2(n16773), .ZN(n16723) );
  OAI21_X1 U19883 ( .B1(n16652), .B2(n16723), .A(n16777), .ZN(n16711) );
  OAI21_X1 U19884 ( .B1(n16653), .B2(n16768), .A(n16711), .ZN(n16681) );
  INV_X1 U19885 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18604) );
  INV_X1 U19886 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18602) );
  NAND2_X1 U19887 ( .A1(n16653), .A2(n16704), .ZN(n16662) );
  AOI221_X1 U19888 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n18604), .C2(n18602), .A(n16662), .ZN(n16658) );
  AOI21_X1 U19889 ( .B1(n17587), .B2(n16663), .A(n16654), .ZN(n17590) );
  INV_X1 U19890 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17611) );
  NOR2_X1 U19891 ( .A1(n17611), .A2(n16655), .ZN(n16666) );
  AOI21_X1 U19892 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16666), .A(
        n16764), .ZN(n16665) );
  OAI21_X1 U19893 ( .B1(n17590), .B2(n16665), .A(n16753), .ZN(n16656) );
  AOI21_X1 U19894 ( .B1(n17590), .B2(n16665), .A(n16656), .ZN(n16657) );
  AOI211_X1 U19895 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16681), .A(n16658), 
        .B(n16657), .ZN(n16659) );
  OAI211_X1 U19896 ( .C1(n17587), .C2(n16745), .A(n16660), .B(n16659), .ZN(
        P3_U2661) );
  NOR3_X1 U19897 ( .A1(n16668), .A2(n16661), .A3(n16667), .ZN(n16676) );
  AOI22_X1 U19898 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16765), .B1(
        n16676), .B2(n16995), .ZN(n16674) );
  INV_X1 U19899 ( .A(n16662), .ZN(n16672) );
  NOR2_X1 U19900 ( .A1(n17611), .A2(n16685), .ZN(n16664) );
  OAI21_X1 U19901 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16664), .A(
        n16663), .ZN(n17601) );
  OAI211_X1 U19902 ( .C1(n16666), .C2(n17601), .A(n16753), .B(n16665), .ZN(
        n16670) );
  NAND2_X1 U19903 ( .A1(n16767), .A2(n16770), .ZN(n16778) );
  OAI211_X1 U19904 ( .C1(n16668), .C2(n16667), .A(P3_EBX_REG_9__SCAN_IN), .B(
        n16778), .ZN(n16669) );
  OAI211_X1 U19905 ( .C1(n16757), .C2(n17601), .A(n16670), .B(n16669), .ZN(
        n16671) );
  AOI221_X1 U19906 ( .B1(n16672), .B2(n18602), .C1(n16681), .C2(
        P3_REIP_REG_9__SCAN_IN), .A(n16671), .ZN(n16673) );
  NAND3_X1 U19907 ( .A1(n16674), .A2(n16673), .A3(n9800), .ZN(P3_U2662) );
  NAND2_X1 U19908 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16693), .ZN(n16675) );
  AOI22_X1 U19909 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16765), .B1(
        n16676), .B2(n16675), .ZN(n16684) );
  NOR2_X1 U19910 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16688), .ZN(n16677) );
  AOI22_X1 U19911 ( .A1(n16722), .A2(P3_EBX_REG_8__SCAN_IN), .B1(n16704), .B2(
        n16677), .ZN(n16683) );
  INV_X1 U19912 ( .A(n16685), .ZN(n16678) );
  AOI22_X1 U19913 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16685), .B1(
        n16678), .B2(n17611), .ZN(n17608) );
  XOR2_X1 U19914 ( .A(n17608), .B(n16679), .Z(n16680) );
  AOI22_X1 U19915 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16681), .B1(n16753), 
        .B2(n16680), .ZN(n16682) );
  NAND4_X1 U19916 ( .A1(n16684), .A2(n16683), .A3(n16682), .A4(n9800), .ZN(
        P3_U2663) );
  INV_X1 U19917 ( .A(n16711), .ZN(n16692) );
  OAI21_X1 U19918 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16698), .A(
        n16685), .ZN(n17629) );
  INV_X1 U19919 ( .A(n17623), .ZN(n17607) );
  INV_X1 U19920 ( .A(n16754), .ZN(n16686) );
  OAI21_X1 U19921 ( .B1(n17607), .B2(n16686), .A(n16733), .ZN(n16700) );
  OAI21_X1 U19922 ( .B1(n17629), .B2(n16700), .A(n16753), .ZN(n16687) );
  AOI21_X1 U19923 ( .B1(n17629), .B2(n16700), .A(n16687), .ZN(n16691) );
  OAI211_X1 U19924 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16704), .B(n16688), .ZN(n16689) );
  OAI211_X1 U19925 ( .C1(n10100), .C2(n16745), .A(n9800), .B(n16689), .ZN(
        n16690) );
  AOI211_X1 U19926 ( .C1(n16692), .C2(P3_REIP_REG_7__SCAN_IN), .A(n16691), .B(
        n16690), .ZN(n16695) );
  OAI211_X1 U19927 ( .C1(n16696), .C2(n16969), .A(n16749), .B(n16693), .ZN(
        n16694) );
  OAI211_X1 U19928 ( .C1(n16969), .C2(n16767), .A(n16695), .B(n16694), .ZN(
        P3_U2664) );
  INV_X1 U19929 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18596) );
  AOI211_X1 U19930 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16714), .A(n16696), .B(
        n16770), .ZN(n16697) );
  AOI211_X1 U19931 ( .C1(n16722), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18035), .B(
        n16697), .ZN(n16706) );
  AOI21_X1 U19932 ( .B1(n17645), .B2(n16699), .A(n16698), .ZN(n17642) );
  NOR3_X1 U19933 ( .A1(n17642), .A2(n18565), .A3(n16700), .ZN(n16703) );
  OAI21_X1 U19934 ( .B1(n16708), .B2(n16764), .A(n17642), .ZN(n16701) );
  OAI22_X1 U19935 ( .A1(n17645), .A2(n16745), .B1(n16776), .B2(n16701), .ZN(
        n16702) );
  AOI211_X1 U19936 ( .C1(n16704), .C2(n18596), .A(n16703), .B(n16702), .ZN(
        n16705) );
  OAI211_X1 U19937 ( .C1(n18596), .C2(n16711), .A(n16706), .B(n16705), .ZN(
        P3_U2665) );
  NOR2_X1 U19938 ( .A1(n16768), .A2(n16707), .ZN(n16726) );
  AOI21_X1 U19939 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16726), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16712) );
  INV_X1 U19940 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16709) );
  NAND2_X1 U19941 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17646), .ZN(
        n16718) );
  AOI21_X1 U19942 ( .B1(n16709), .B2(n16718), .A(n16708), .ZN(n17654) );
  OAI21_X1 U19943 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16718), .A(
        n16733), .ZN(n16717) );
  XOR2_X1 U19944 ( .A(n17654), .B(n16717), .Z(n16710) );
  OAI22_X1 U19945 ( .A1(n16712), .A2(n16711), .B1(n18565), .B2(n16710), .ZN(
        n16713) );
  AOI211_X1 U19946 ( .C1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n16765), .A(
        n18035), .B(n16713), .ZN(n16716) );
  OAI211_X1 U19947 ( .C1(n16724), .C2(n17060), .A(n16749), .B(n16714), .ZN(
        n16715) );
  OAI211_X1 U19948 ( .C1(n17060), .C2(n16767), .A(n16716), .B(n16715), .ZN(
        P3_U2666) );
  NOR2_X1 U19949 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17666), .ZN(
        n17663) );
  INV_X1 U19950 ( .A(n16717), .ZN(n16719) );
  NOR2_X1 U19951 ( .A1(n21011), .A2(n17666), .ZN(n16730) );
  OAI21_X1 U19952 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16730), .A(
        n16718), .ZN(n17669) );
  AOI22_X1 U19953 ( .A1(n16754), .A2(n17663), .B1(n16719), .B2(n17669), .ZN(
        n16729) );
  NAND2_X1 U19954 ( .A1(n18057), .A2(n18723), .ZN(n16782) );
  OAI221_X1 U19955 ( .B1(n16782), .B2(n11567), .C1(n16782), .C2(n18504), .A(
        n9800), .ZN(n16721) );
  OAI22_X1 U19956 ( .A1(n17668), .A2(n16745), .B1(n17669), .B2(n16757), .ZN(
        n16720) );
  AOI211_X1 U19957 ( .C1(n16722), .C2(P3_EBX_REG_4__SCAN_IN), .A(n16721), .B(
        n16720), .ZN(n16728) );
  AND2_X1 U19958 ( .A1(n16777), .A2(n16723), .ZN(n16739) );
  INV_X1 U19959 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18592) );
  AOI211_X1 U19960 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16740), .A(n16724), .B(
        n16770), .ZN(n16725) );
  AOI221_X1 U19961 ( .B1(n16739), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n16726), 
        .C2(n18592), .A(n16725), .ZN(n16727) );
  OAI211_X1 U19962 ( .C1(n16729), .C2(n18565), .A(n16728), .B(n16727), .ZN(
        P3_U2667) );
  NAND2_X1 U19963 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n16760) );
  INV_X1 U19964 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18591) );
  OAI21_X1 U19965 ( .B1(n16768), .B2(n16760), .A(n18591), .ZN(n16738) );
  INV_X1 U19966 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16731) );
  NAND2_X1 U19967 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16746) );
  AOI21_X1 U19968 ( .B1(n16731), .B2(n16746), .A(n16730), .ZN(n16732) );
  INV_X1 U19969 ( .A(n16732), .ZN(n17686) );
  OAI21_X1 U19970 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16746), .A(
        n16733), .ZN(n16751) );
  OAI21_X1 U19971 ( .B1(n17686), .B2(n16751), .A(n16753), .ZN(n16734) );
  AOI21_X1 U19972 ( .B1(n17686), .B2(n16751), .A(n16734), .ZN(n16737) );
  INV_X1 U19973 ( .A(n16782), .ZN(n18725) );
  NOR2_X1 U19974 ( .A1(n18675), .A2(n11599), .ZN(n18519) );
  NAND2_X1 U19975 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18519), .ZN(
        n18511) );
  AOI21_X1 U19976 ( .B1(n18665), .B2(n18511), .A(n17046), .ZN(n18662) );
  AOI22_X1 U19977 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16765), .B1(
        n18725), .B2(n18662), .ZN(n16735) );
  INV_X1 U19978 ( .A(n16735), .ZN(n16736) );
  AOI211_X1 U19979 ( .C1(n16739), .C2(n16738), .A(n16737), .B(n16736), .ZN(
        n16742) );
  OAI211_X1 U19980 ( .C1(n16747), .C2(n16743), .A(n16749), .B(n16740), .ZN(
        n16741) );
  OAI211_X1 U19981 ( .C1(n16743), .C2(n16767), .A(n16742), .B(n16741), .ZN(
        P3_U2668) );
  INV_X1 U19982 ( .A(n18511), .ZN(n16744) );
  AOI21_X1 U19983 ( .B1(n18675), .B2(n18526), .A(n16744), .ZN(n18673) );
  INV_X1 U19984 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17696) );
  INV_X1 U19985 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20808) );
  OAI22_X1 U19986 ( .A1(n17696), .A2(n16745), .B1(n20808), .B2(n16779), .ZN(
        n16759) );
  OAI21_X1 U19987 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16746), .ZN(n17692) );
  NOR2_X1 U19988 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16750) );
  INV_X1 U19989 ( .A(n16747), .ZN(n16748) );
  OAI211_X1 U19990 ( .C1(n16750), .C2(n17068), .A(n16749), .B(n16748), .ZN(
        n16756) );
  INV_X1 U19991 ( .A(n16751), .ZN(n16752) );
  OAI211_X1 U19992 ( .C1(n16754), .C2(n17692), .A(n16753), .B(n16752), .ZN(
        n16755) );
  OAI211_X1 U19993 ( .C1(n16757), .C2(n17692), .A(n16756), .B(n16755), .ZN(
        n16758) );
  AOI211_X1 U19994 ( .C1(n18673), .C2(n18725), .A(n16759), .B(n16758), .ZN(
        n16763) );
  OAI211_X1 U19995 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n16761), .B(n16760), .ZN(n16762) );
  OAI211_X1 U19996 ( .C1(n17068), .C2(n16767), .A(n16763), .B(n16762), .ZN(
        P3_U2669) );
  NOR2_X1 U19997 ( .A1(n16764), .A2(n18565), .ZN(n16766) );
  AOI21_X1 U19998 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16766), .A(
        n16765), .ZN(n16775) );
  INV_X1 U19999 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17077) );
  OAI22_X1 U20000 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16768), .B1(n16767), 
        .B2(n17077), .ZN(n16772) );
  OAI21_X1 U20001 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17071), .ZN(n17078) );
  NAND2_X1 U20002 ( .A1(n16769), .A2(n18526), .ZN(n18676) );
  OAI22_X1 U20003 ( .A1(n16770), .A2(n17078), .B1(n18676), .B2(n16782), .ZN(
        n16771) );
  AOI211_X1 U20004 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n16773), .A(n16772), .B(
        n16771), .ZN(n16774) );
  OAI221_X1 U20005 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16776), .C1(
        n21011), .C2(n16775), .A(n16774), .ZN(P3_U2670) );
  AOI22_X1 U20006 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16778), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16777), .ZN(n16781) );
  NAND3_X1 U20007 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18670), .A3(
        n16779), .ZN(n16780) );
  OAI211_X1 U20008 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16782), .A(
        n16781), .B(n16780), .ZN(P3_U2671) );
  AOI22_X1 U20009 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16786) );
  AOI22_X1 U20010 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16785) );
  AOI22_X1 U20011 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16784) );
  AOI22_X1 U20012 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16783) );
  NAND4_X1 U20013 ( .A1(n16786), .A2(n16785), .A3(n16784), .A4(n16783), .ZN(
        n16792) );
  AOI22_X1 U20014 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16790) );
  AOI22_X1 U20015 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16789) );
  AOI22_X1 U20016 ( .A1(n9787), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16788) );
  AOI22_X1 U20017 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16787) );
  NAND4_X1 U20018 ( .A1(n16790), .A2(n16789), .A3(n16788), .A4(n16787), .ZN(
        n16791) );
  NOR2_X1 U20019 ( .A1(n16792), .A2(n16791), .ZN(n16803) );
  AOI22_X1 U20020 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16802) );
  AOI22_X1 U20021 ( .A1(n17004), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U20022 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16793) );
  OAI21_X1 U20023 ( .B1(n9841), .B2(n20973), .A(n16793), .ZN(n16799) );
  AOI22_X1 U20024 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16797) );
  AOI22_X1 U20025 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16796) );
  AOI22_X1 U20026 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16795) );
  AOI22_X1 U20027 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9788), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16794) );
  NAND4_X1 U20028 ( .A1(n16797), .A2(n16796), .A3(n16795), .A4(n16794), .ZN(
        n16798) );
  AOI211_X1 U20029 ( .C1(n16924), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n16799), .B(n16798), .ZN(n16800) );
  NAND3_X1 U20030 ( .A1(n16802), .A2(n16801), .A3(n16800), .ZN(n16808) );
  NAND2_X1 U20031 ( .A1(n16809), .A2(n16808), .ZN(n16807) );
  XNOR2_X1 U20032 ( .A(n16803), .B(n16807), .ZN(n17092) );
  NOR2_X1 U20033 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16804), .ZN(n16806) );
  OAI22_X1 U20034 ( .A1(n17092), .A2(n17075), .B1(n16806), .B2(n16805), .ZN(
        P3_U2673) );
  OAI21_X1 U20035 ( .B1(n16809), .B2(n16808), .A(n16807), .ZN(n17096) );
  NOR2_X1 U20036 ( .A1(n16824), .A2(n16810), .ZN(n16812) );
  AOI22_X1 U20037 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16813), .B1(n16812), 
        .B2(n16811), .ZN(n16814) );
  OAI21_X1 U20038 ( .B1(n17096), .B2(n17075), .A(n16814), .ZN(P3_U2674) );
  OAI21_X1 U20039 ( .B1(n16819), .B2(n16816), .A(n16815), .ZN(n17105) );
  NAND3_X1 U20040 ( .A1(n16818), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17075), 
        .ZN(n16817) );
  OAI221_X1 U20041 ( .B1(n16818), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17075), 
        .C2(n17105), .A(n16817), .ZN(P3_U2676) );
  AOI21_X1 U20042 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17075), .A(n16828), .ZN(
        n16822) );
  AOI21_X1 U20043 ( .B1(n16820), .B2(n16825), .A(n16819), .ZN(n17106) );
  INV_X1 U20044 ( .A(n17106), .ZN(n16821) );
  OAI22_X1 U20045 ( .A1(n16823), .A2(n16822), .B1(n17075), .B2(n16821), .ZN(
        P3_U2677) );
  INV_X1 U20046 ( .A(n16824), .ZN(n16833) );
  AOI21_X1 U20047 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17075), .A(n16833), .ZN(
        n16827) );
  OAI21_X1 U20048 ( .B1(n16829), .B2(n16826), .A(n16825), .ZN(n17115) );
  OAI22_X1 U20049 ( .A1(n16828), .A2(n16827), .B1(n17075), .B2(n17115), .ZN(
        P3_U2678) );
  AOI21_X1 U20050 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17075), .A(n16839), .ZN(
        n16832) );
  AOI21_X1 U20051 ( .B1(n16830), .B2(n16835), .A(n16829), .ZN(n17116) );
  INV_X1 U20052 ( .A(n17116), .ZN(n16831) );
  OAI22_X1 U20053 ( .A1(n16833), .A2(n16832), .B1(n17075), .B2(n16831), .ZN(
        P3_U2679) );
  INV_X1 U20054 ( .A(n16834), .ZN(n16854) );
  AOI21_X1 U20055 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17075), .A(n16854), .ZN(
        n16838) );
  OAI21_X1 U20056 ( .B1(n16837), .B2(n16836), .A(n16835), .ZN(n17125) );
  OAI22_X1 U20057 ( .A1(n16839), .A2(n16838), .B1(n17075), .B2(n17125), .ZN(
        P3_U2680) );
  AOI21_X1 U20058 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17075), .A(n16840), .ZN(
        n16853) );
  AOI22_X1 U20059 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16851) );
  AOI22_X1 U20060 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16850) );
  AOI22_X1 U20061 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16841) );
  OAI21_X1 U20062 ( .B1(n16842), .B2(n20973), .A(n16841), .ZN(n16848) );
  AOI22_X1 U20063 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16846) );
  AOI22_X1 U20064 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16845) );
  AOI22_X1 U20065 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16844) );
  AOI22_X1 U20066 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16843) );
  NAND4_X1 U20067 ( .A1(n16846), .A2(n16845), .A3(n16844), .A4(n16843), .ZN(
        n16847) );
  AOI211_X1 U20068 ( .C1(n17035), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n16848), .B(n16847), .ZN(n16849) );
  NAND3_X1 U20069 ( .A1(n16851), .A2(n16850), .A3(n16849), .ZN(n17126) );
  INV_X1 U20070 ( .A(n17126), .ZN(n16852) );
  OAI22_X1 U20071 ( .A1(n16854), .A2(n16853), .B1(n16852), .B2(n17075), .ZN(
        P3_U2681) );
  NOR2_X1 U20072 ( .A1(n17080), .A2(n16855), .ZN(n16879) );
  AOI22_X1 U20073 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20074 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16858) );
  AOI22_X1 U20075 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16857) );
  AOI22_X1 U20076 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16856) );
  NAND4_X1 U20077 ( .A1(n16859), .A2(n16858), .A3(n16857), .A4(n16856), .ZN(
        n16865) );
  AOI22_X1 U20078 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16863) );
  AOI22_X1 U20079 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16862) );
  AOI22_X1 U20080 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20081 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16860) );
  NAND4_X1 U20082 ( .A1(n16863), .A2(n16862), .A3(n16861), .A4(n16860), .ZN(
        n16864) );
  NOR2_X1 U20083 ( .A1(n16865), .A2(n16864), .ZN(n17132) );
  INV_X1 U20084 ( .A(n17132), .ZN(n16866) );
  AOI22_X1 U20085 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16879), .B1(n17080), 
        .B2(n16866), .ZN(n16867) );
  OAI21_X1 U20086 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16868), .A(n16867), .ZN(
        P3_U2682) );
  AOI22_X1 U20087 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16878) );
  AOI22_X1 U20088 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16877) );
  AOI22_X1 U20089 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16869) );
  OAI21_X1 U20090 ( .B1(n16899), .B2(n18083), .A(n16869), .ZN(n16875) );
  AOI22_X1 U20091 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16873) );
  AOI22_X1 U20092 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16872) );
  AOI22_X1 U20093 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16871) );
  AOI22_X1 U20094 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16870) );
  NAND4_X1 U20095 ( .A1(n16873), .A2(n16872), .A3(n16871), .A4(n16870), .ZN(
        n16874) );
  AOI211_X1 U20096 ( .C1(n17016), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n16875), .B(n16874), .ZN(n16876) );
  NAND3_X1 U20097 ( .A1(n16878), .A2(n16877), .A3(n16876), .ZN(n17136) );
  INV_X1 U20098 ( .A(n17136), .ZN(n16882) );
  OAI21_X1 U20099 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16880), .A(n16879), .ZN(
        n16881) );
  OAI21_X1 U20100 ( .B1(n16882), .B2(n17075), .A(n16881), .ZN(P3_U2683) );
  AOI22_X1 U20101 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16886) );
  AOI22_X1 U20102 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16885) );
  AOI22_X1 U20103 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16884) );
  AOI22_X1 U20104 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16883) );
  NAND4_X1 U20105 ( .A1(n16886), .A2(n16885), .A3(n16884), .A4(n16883), .ZN(
        n16892) );
  AOI22_X1 U20106 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16890) );
  AOI22_X1 U20107 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20108 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U20109 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16887) );
  NAND4_X1 U20110 ( .A1(n16890), .A2(n16889), .A3(n16888), .A4(n16887), .ZN(
        n16891) );
  NOR2_X1 U20111 ( .A1(n16892), .A2(n16891), .ZN(n17144) );
  OAI21_X1 U20112 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16895), .A(n16893), .ZN(
        n16894) );
  AOI22_X1 U20113 ( .A1(n17080), .A2(n17144), .B1(n16894), .B2(n17075), .ZN(
        P3_U2684) );
  AOI21_X1 U20114 ( .B1(n16897), .B2(n16896), .A(n16895), .ZN(n16909) );
  AOI22_X1 U20115 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n15486), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16908) );
  AOI22_X1 U20116 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n9790), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16907) );
  AOI22_X1 U20117 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16898) );
  OAI21_X1 U20118 ( .B1(n16899), .B2(n18072), .A(n16898), .ZN(n16905) );
  AOI22_X1 U20119 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n17004), .ZN(n16903) );
  AOI22_X1 U20120 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__2__SCAN_IN), .B2(n17021), .ZN(n16902) );
  AOI22_X1 U20121 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n15546), .B1(
        P3_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n16971), .ZN(n16901) );
  AOI22_X1 U20122 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n9788), .ZN(n16900) );
  NAND4_X1 U20123 ( .A1(n16903), .A2(n16902), .A3(n16901), .A4(n16900), .ZN(
        n16904) );
  AOI211_X1 U20124 ( .C1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .C2(n17039), .A(
        n16905), .B(n16904), .ZN(n16906) );
  NAND3_X1 U20125 ( .A1(n16908), .A2(n16907), .A3(n16906), .ZN(n17145) );
  MUX2_X1 U20126 ( .A(n16909), .B(n17145), .S(n17080), .Z(P3_U2685) );
  AOI22_X1 U20127 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20128 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20129 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16911) );
  AOI22_X1 U20130 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9787), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16910) );
  NAND4_X1 U20131 ( .A1(n16913), .A2(n16912), .A3(n16911), .A4(n16910), .ZN(
        n16919) );
  AOI22_X1 U20132 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20133 ( .A1(n15486), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16916) );
  AOI22_X1 U20134 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16915) );
  AOI22_X1 U20135 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16914) );
  NAND4_X1 U20136 ( .A1(n16917), .A2(n16916), .A3(n16915), .A4(n16914), .ZN(
        n16918) );
  NOR2_X1 U20137 ( .A1(n16919), .A2(n16918), .ZN(n17155) );
  INV_X1 U20138 ( .A(n17082), .ZN(n17064) );
  OR2_X1 U20139 ( .A1(n17163), .A2(n16921), .ZN(n16938) );
  NAND3_X1 U20140 ( .A1(n17076), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n16938), 
        .ZN(n16920) );
  OAI221_X1 U20141 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16921), .C1(
        P3_EBX_REG_17__SCAN_IN), .C2(n17064), .A(n16920), .ZN(n16922) );
  OAI21_X1 U20142 ( .B1(n17155), .B2(n17075), .A(n16922), .ZN(P3_U2686) );
  NOR2_X1 U20143 ( .A1(n16923), .A2(n16964), .ZN(n16967) );
  NAND2_X1 U20144 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16967), .ZN(n16937) );
  AOI22_X1 U20145 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16928) );
  AOI22_X1 U20146 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U20147 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16926) );
  AOI22_X1 U20148 ( .A1(n9788), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16925) );
  NAND4_X1 U20149 ( .A1(n16928), .A2(n16927), .A3(n16926), .A4(n16925), .ZN(
        n16935) );
  AOI22_X1 U20150 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20151 ( .A1(n15486), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20152 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U20153 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16930) );
  NAND4_X1 U20154 ( .A1(n16933), .A2(n16932), .A3(n16931), .A4(n16930), .ZN(
        n16934) );
  NOR2_X1 U20155 ( .A1(n16935), .A2(n16934), .ZN(n17162) );
  INV_X1 U20156 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16936) );
  NAND2_X1 U20157 ( .A1(n17075), .A2(n16937), .ZN(n16949) );
  OAI222_X1 U20158 ( .A1(n16938), .A2(n16937), .B1(n17075), .B2(n17162), .C1(
        n16936), .C2(n16949), .ZN(P3_U2687) );
  AOI22_X1 U20159 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20160 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20161 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16939) );
  OAI21_X1 U20162 ( .B1(n9801), .B2(n21017), .A(n16939), .ZN(n16945) );
  AOI22_X1 U20163 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20164 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17039), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20165 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20166 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16940) );
  NAND4_X1 U20167 ( .A1(n16943), .A2(n16942), .A3(n16941), .A4(n16940), .ZN(
        n16944) );
  AOI211_X1 U20168 ( .C1(n17046), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n16945), .B(n16944), .ZN(n16946) );
  NAND3_X1 U20169 ( .A1(n16948), .A2(n16947), .A3(n16946), .ZN(n17165) );
  INV_X1 U20170 ( .A(n17165), .ZN(n16951) );
  NOR2_X1 U20171 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16967), .ZN(n16950) );
  OAI22_X1 U20172 ( .A1(n16951), .A2(n17075), .B1(n16950), .B2(n16949), .ZN(
        P3_U2688) );
  AOI22_X1 U20173 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20174 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20175 ( .A1(n9790), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16952) );
  OAI21_X1 U20176 ( .B1(n16953), .B2(n20973), .A(n16952), .ZN(n16960) );
  AOI22_X1 U20177 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n16954), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U20178 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20179 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16956) );
  AOI22_X1 U20180 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9788), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16955) );
  NAND4_X1 U20181 ( .A1(n16958), .A2(n16957), .A3(n16956), .A4(n16955), .ZN(
        n16959) );
  NAND3_X1 U20182 ( .A1(n16963), .A2(n16962), .A3(n16961), .ZN(n17171) );
  INV_X1 U20183 ( .A(n17171), .ZN(n16968) );
  INV_X1 U20184 ( .A(n16964), .ZN(n16965) );
  OAI21_X1 U20185 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16965), .A(n17075), .ZN(
        n16966) );
  OAI22_X1 U20186 ( .A1(n16968), .A2(n17075), .B1(n16967), .B2(n16966), .ZN(
        P3_U2689) );
  NOR3_X1 U20187 ( .A1(n16969), .A2(n17054), .A3(n17062), .ZN(n16994) );
  NAND2_X1 U20188 ( .A1(n18097), .A2(n16994), .ZN(n17050) );
  NOR2_X1 U20189 ( .A1(n16970), .A2(n17050), .ZN(n17013) );
  NAND3_X1 U20190 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n17013), .ZN(n16983) );
  AOI22_X1 U20191 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20192 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20193 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9798), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20194 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16972) );
  NAND4_X1 U20195 ( .A1(n16975), .A2(n16974), .A3(n16973), .A4(n16972), .ZN(
        n16981) );
  AOI22_X1 U20196 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20197 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16978) );
  AOI22_X1 U20198 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20199 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16976) );
  NAND4_X1 U20200 ( .A1(n16979), .A2(n16978), .A3(n16977), .A4(n16976), .ZN(
        n16980) );
  NOR2_X1 U20201 ( .A1(n16981), .A2(n16980), .ZN(n17181) );
  NAND3_X1 U20202 ( .A1(n16983), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17075), 
        .ZN(n16982) );
  OAI221_X1 U20203 ( .B1(n16983), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17075), 
        .C2(n17181), .A(n16982), .ZN(P3_U2691) );
  AOI22_X1 U20204 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17004), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20205 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20206 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17003), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20207 ( .A1(n17046), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16984) );
  NAND4_X1 U20208 ( .A1(n16987), .A2(n16986), .A3(n16985), .A4(n16984), .ZN(
        n16993) );
  AOI22_X1 U20209 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16991) );
  AOI22_X1 U20210 ( .A1(n9793), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20211 ( .A1(n12889), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20212 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16988) );
  NAND4_X1 U20213 ( .A1(n16991), .A2(n16990), .A3(n16989), .A4(n16988), .ZN(
        n16992) );
  NOR2_X1 U20214 ( .A1(n16993), .A2(n16992), .ZN(n17185) );
  NAND2_X1 U20215 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16994), .ZN(n17051) );
  NOR2_X1 U20216 ( .A1(n16995), .A2(n17051), .ZN(n17011) );
  NAND2_X1 U20217 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17011), .ZN(n16996) );
  XNOR2_X1 U20218 ( .A(n16997), .B(n16996), .ZN(n16998) );
  AOI22_X1 U20219 ( .A1(n17080), .A2(n17185), .B1(n16998), .B2(n17075), .ZN(
        P3_U2692) );
  AOI22_X1 U20220 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n9798), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20221 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n17036), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20222 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20223 ( .A1(n9789), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9788), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16999) );
  NAND4_X1 U20224 ( .A1(n17002), .A2(n17001), .A3(n17000), .A4(n16999), .ZN(
        n17010) );
  AOI22_X1 U20225 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n9793), .B1(
        P3_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n17003), .ZN(n17008) );
  AOI22_X1 U20226 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n17039), .B1(
        P3_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n15486), .ZN(n17007) );
  AOI22_X1 U20227 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n17004), .ZN(n17006) );
  AOI22_X1 U20228 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__2__SCAN_IN), .B2(n15546), .ZN(n17005) );
  NAND4_X1 U20229 ( .A1(n17008), .A2(n17007), .A3(n17006), .A4(n17005), .ZN(
        n17009) );
  NOR2_X1 U20230 ( .A1(n17010), .A2(n17009), .ZN(n17190) );
  NOR2_X1 U20231 ( .A1(n17080), .A2(n17011), .ZN(n17031) );
  AOI22_X1 U20232 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17031), .B1(n17013), 
        .B2(n17012), .ZN(n17014) );
  OAI21_X1 U20233 ( .B1(n17190), .B2(n17075), .A(n17014), .ZN(P3_U2693) );
  AOI22_X1 U20234 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17015), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20235 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15546), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20236 ( .A1(n17036), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17017) );
  OAI21_X1 U20237 ( .B1(n17018), .B2(n21015), .A(n17017), .ZN(n17027) );
  AOI22_X1 U20238 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16971), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20239 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15486), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20240 ( .A1(n17021), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9793), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20241 ( .A1(n16924), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9787), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17022) );
  NAND4_X1 U20242 ( .A1(n17025), .A2(n17024), .A3(n17023), .A4(n17022), .ZN(
        n17026) );
  AOI211_X1 U20243 ( .C1(n17035), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n17027), .B(n17026), .ZN(n17028) );
  NAND3_X1 U20244 ( .A1(n17030), .A2(n17029), .A3(n17028), .ZN(n17194) );
  INV_X1 U20245 ( .A(n17194), .ZN(n17034) );
  INV_X1 U20246 ( .A(n17051), .ZN(n17032) );
  OAI21_X1 U20247 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17032), .A(n17031), .ZN(
        n17033) );
  OAI21_X1 U20248 ( .B1(n17034), .B2(n17075), .A(n17033), .ZN(P3_U2694) );
  AOI22_X1 U20249 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17020), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20250 ( .A1(n12878), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17036), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20251 ( .A1(n17003), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15551), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17037) );
  OAI21_X1 U20252 ( .B1(n9801), .B2(n18061), .A(n17037), .ZN(n17045) );
  AOI22_X1 U20253 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17019), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20254 ( .A1(n17039), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17021), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20255 ( .A1(n16971), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15492), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20256 ( .A1(n9798), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9793), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17040) );
  NAND4_X1 U20257 ( .A1(n17043), .A2(n17042), .A3(n17041), .A4(n17040), .ZN(
        n17044) );
  AOI211_X1 U20258 ( .C1(n17046), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17045), .B(n17044), .ZN(n17047) );
  NAND3_X1 U20259 ( .A1(n17049), .A2(n17048), .A3(n17047), .ZN(n17201) );
  INV_X1 U20260 ( .A(n17201), .ZN(n17053) );
  INV_X1 U20261 ( .A(n17050), .ZN(n17056) );
  OAI21_X1 U20262 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17056), .A(n17051), .ZN(
        n17052) );
  AOI22_X1 U20263 ( .A1(n17080), .A2(n17053), .B1(n17052), .B2(n17075), .ZN(
        P3_U2695) );
  OAI21_X1 U20264 ( .B1(n17054), .B2(n17062), .A(n17075), .ZN(n17058) );
  OAI22_X1 U20265 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17058), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17075), .ZN(n17055) );
  NOR2_X1 U20266 ( .A1(n17056), .A2(n17055), .ZN(P3_U2696) );
  NOR2_X1 U20267 ( .A1(n17057), .A2(n17082), .ZN(n17067) );
  AOI21_X1 U20268 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17067), .A(
        P3_EBX_REG_6__SCAN_IN), .ZN(n17059) );
  INV_X1 U20269 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18094) );
  OAI22_X1 U20270 ( .A1(n17059), .A2(n17058), .B1(n18094), .B2(n17075), .ZN(
        P3_U2697) );
  INV_X1 U20271 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18089) );
  AOI22_X1 U20272 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17062), .B1(n17061), .B2(
        n17060), .ZN(n17063) );
  AOI22_X1 U20273 ( .A1(n17080), .A2(n18089), .B1(n17063), .B2(n17075), .ZN(
        P3_U2698) );
  AND2_X1 U20274 ( .A1(n17065), .A2(n17064), .ZN(n17070) );
  AOI21_X1 U20275 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17075), .A(n17070), .ZN(
        n17066) );
  OAI22_X1 U20276 ( .A1(n17067), .A2(n17066), .B1(n18083), .B2(n17075), .ZN(
        P3_U2699) );
  NOR3_X1 U20277 ( .A1(n17068), .A2(n17071), .A3(n17082), .ZN(n17074) );
  AOI21_X1 U20278 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17075), .A(n17074), .ZN(
        n17069) );
  INV_X1 U20279 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18078) );
  OAI22_X1 U20280 ( .A1(n17070), .A2(n17069), .B1(n18078), .B2(n17075), .ZN(
        P3_U2700) );
  NOR2_X1 U20281 ( .A1(n17071), .A2(n17082), .ZN(n17072) );
  AOI21_X1 U20282 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17075), .A(n17072), .ZN(
        n17073) );
  OAI22_X1 U20283 ( .A1(n17074), .A2(n17073), .B1(n18072), .B2(n17075), .ZN(
        P3_U2701) );
  INV_X1 U20284 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18066) );
  OAI222_X1 U20285 ( .A1(n17078), .A2(n17082), .B1(n17077), .B2(n17076), .C1(
        n18066), .C2(n17075), .ZN(P3_U2702) );
  AOI22_X1 U20286 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17080), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17079), .ZN(n17081) );
  OAI21_X1 U20287 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17082), .A(n17081), .ZN(
        P3_U2703) );
  INV_X1 U20288 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17307) );
  INV_X1 U20289 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17302) );
  INV_X1 U20290 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20940) );
  INV_X1 U20291 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17329) );
  NAND2_X1 U20292 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17223) );
  INV_X1 U20293 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17319) );
  INV_X1 U20294 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17327) );
  NAND4_X1 U20295 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17083) );
  NOR4_X1 U20296 ( .A1(n17223), .A2(n17319), .A3(n17327), .A4(n17083), .ZN(
        n17168) );
  INV_X1 U20297 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17340) );
  INV_X1 U20298 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17333) );
  INV_X1 U20299 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17338) );
  INV_X1 U20300 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17336) );
  NOR4_X1 U20301 ( .A1(n17340), .A2(n17333), .A3(n17338), .A4(n17336), .ZN(
        n17170) );
  INV_X1 U20302 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20845) );
  INV_X1 U20303 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17294) );
  NAND4_X1 U20304 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17084)
         );
  NOR4_X2 U20305 ( .A1(n17158), .A2(n20845), .A3(n17294), .A4(n17084), .ZN(
        n17122) );
  NAND2_X1 U20306 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17122), .ZN(n17121) );
  NAND2_X1 U20307 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17118), .ZN(n17117) );
  NAND2_X1 U20308 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17098), .ZN(n17093) );
  NAND2_X1 U20309 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17089), .ZN(n17088) );
  NAND3_X1 U20310 ( .A1(n17225), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17088), 
        .ZN(n17086) );
  NOR2_X2 U20311 ( .A1(n18091), .A2(n17215), .ZN(n17156) );
  NAND2_X1 U20312 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17156), .ZN(n17085) );
  OAI211_X1 U20313 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17088), .A(n17086), .B(
        n17085), .ZN(P3_U2704) );
  NOR2_X1 U20314 ( .A1(n17087), .A2(n17215), .ZN(n17157) );
  AOI22_X1 U20315 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17157), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17156), .ZN(n17091) );
  OAI211_X1 U20316 ( .C1(n17089), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17215), .B(
        n17088), .ZN(n17090) );
  OAI211_X1 U20317 ( .C1(n17092), .C2(n17226), .A(n17091), .B(n17090), .ZN(
        P3_U2705) );
  AOI22_X1 U20318 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17157), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17156), .ZN(n17095) );
  OAI211_X1 U20319 ( .C1(n17098), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17215), .B(
        n17093), .ZN(n17094) );
  OAI211_X1 U20320 ( .C1(n17096), .C2(n17226), .A(n17095), .B(n17094), .ZN(
        P3_U2706) );
  INV_X1 U20321 ( .A(n17156), .ZN(n17131) );
  AOI22_X1 U20322 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17157), .B1(n17233), .B2(
        n17097), .ZN(n17101) );
  AOI211_X1 U20323 ( .C1(n17307), .C2(n17102), .A(n17098), .B(n17237), .ZN(
        n17099) );
  INV_X1 U20324 ( .A(n17099), .ZN(n17100) );
  OAI211_X1 U20325 ( .C1(n17131), .C2(n19161), .A(n17101), .B(n17100), .ZN(
        P3_U2707) );
  AOI22_X1 U20326 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17157), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17156), .ZN(n17104) );
  OAI211_X1 U20327 ( .C1(n17107), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17215), .B(
        n17102), .ZN(n17103) );
  OAI211_X1 U20328 ( .C1(n17105), .C2(n17226), .A(n17104), .B(n17103), .ZN(
        P3_U2708) );
  INV_X1 U20329 ( .A(n17157), .ZN(n17149) );
  AOI22_X1 U20330 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17156), .B1(n17233), .B2(
        n17106), .ZN(n17110) );
  AOI211_X1 U20331 ( .C1(n17302), .C2(n17111), .A(n17107), .B(n17237), .ZN(
        n17108) );
  INV_X1 U20332 ( .A(n17108), .ZN(n17109) );
  OAI211_X1 U20333 ( .C1(n17149), .C2(n17193), .A(n17110), .B(n17109), .ZN(
        P3_U2709) );
  AOI22_X1 U20334 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17157), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17156), .ZN(n17114) );
  OAI211_X1 U20335 ( .C1(n17112), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17215), .B(
        n17111), .ZN(n17113) );
  OAI211_X1 U20336 ( .C1(n17115), .C2(n17226), .A(n17114), .B(n17113), .ZN(
        P3_U2710) );
  AOI22_X1 U20337 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17156), .B1(n17233), .B2(
        n17116), .ZN(n17120) );
  OAI211_X1 U20338 ( .C1(n17118), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17215), .B(
        n17117), .ZN(n17119) );
  OAI211_X1 U20339 ( .C1(n17149), .C2(n17203), .A(n17120), .B(n17119), .ZN(
        P3_U2711) );
  AOI22_X1 U20340 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17157), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17156), .ZN(n17124) );
  OAI211_X1 U20341 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17122), .A(n17225), .B(
        n17121), .ZN(n17123) );
  OAI211_X1 U20342 ( .C1(n17125), .C2(n17226), .A(n17124), .B(n17123), .ZN(
        P3_U2712) );
  INV_X1 U20343 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17285) );
  NAND2_X1 U20344 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17150), .ZN(n17146) );
  NAND2_X1 U20345 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17140), .ZN(n17137) );
  NAND2_X1 U20346 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17294), .ZN(n17130) );
  AOI22_X1 U20347 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17156), .B1(n17233), .B2(
        n17126), .ZN(n17129) );
  NAND2_X1 U20348 ( .A1(n17215), .A2(n17137), .ZN(n17135) );
  OAI21_X1 U20349 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17222), .A(n17135), .ZN(
        n17127) );
  AOI22_X1 U20350 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17157), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17127), .ZN(n17128) );
  OAI211_X1 U20351 ( .C1(n17137), .C2(n17130), .A(n17129), .B(n17128), .ZN(
        P3_U2713) );
  INV_X1 U20352 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17292) );
  INV_X1 U20353 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18086) );
  OAI22_X1 U20354 ( .A1(n17132), .A2(n17226), .B1(n18086), .B2(n17131), .ZN(
        n17133) );
  AOI21_X1 U20355 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17157), .A(n17133), .ZN(
        n17134) );
  OAI221_X1 U20356 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17137), .C1(n17292), 
        .C2(n17135), .A(n17134), .ZN(P3_U2714) );
  AOI22_X1 U20357 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17156), .B1(n17233), .B2(
        n17136), .ZN(n17139) );
  OAI211_X1 U20358 ( .C1(n17140), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17215), .B(
        n17137), .ZN(n17138) );
  OAI211_X1 U20359 ( .C1(n17149), .C2(n18079), .A(n17139), .B(n17138), .ZN(
        P3_U2715) );
  AOI22_X1 U20360 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17157), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17156), .ZN(n17143) );
  AOI211_X1 U20361 ( .C1(n20845), .C2(n17146), .A(n17140), .B(n17237), .ZN(
        n17141) );
  INV_X1 U20362 ( .A(n17141), .ZN(n17142) );
  OAI211_X1 U20363 ( .C1(n17144), .C2(n17226), .A(n17143), .B(n17142), .ZN(
        P3_U2716) );
  AOI22_X1 U20364 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17156), .B1(n17233), .B2(
        n17145), .ZN(n17148) );
  OAI211_X1 U20365 ( .C1(n17150), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17215), .B(
        n17146), .ZN(n17147) );
  OAI211_X1 U20366 ( .C1(n17149), .C2(n18068), .A(n17148), .B(n17147), .ZN(
        P3_U2717) );
  AOI22_X1 U20367 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17157), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17156), .ZN(n17154) );
  INV_X1 U20368 ( .A(n17158), .ZN(n17152) );
  INV_X1 U20369 ( .A(n17150), .ZN(n17151) );
  OAI211_X1 U20370 ( .C1(n17152), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17215), .B(
        n17151), .ZN(n17153) );
  OAI211_X1 U20371 ( .C1(n17155), .C2(n17226), .A(n17154), .B(n17153), .ZN(
        P3_U2718) );
  AOI22_X1 U20372 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17157), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17156), .ZN(n17161) );
  OAI211_X1 U20373 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17159), .A(n17225), .B(
        n17158), .ZN(n17160) );
  OAI211_X1 U20374 ( .C1(n17162), .C2(n17226), .A(n17161), .B(n17160), .ZN(
        P3_U2719) );
  OR2_X1 U20375 ( .A1(n17163), .A2(n17164), .ZN(n17167) );
  NAND2_X1 U20376 ( .A1(n17225), .A2(n17164), .ZN(n17173) );
  AOI22_X1 U20377 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17234), .B1(n17233), .B2(
        n17165), .ZN(n17166) );
  OAI221_X1 U20378 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17167), .C1(n20940), 
        .C2(n17173), .A(n17166), .ZN(P3_U2720) );
  INV_X1 U20379 ( .A(n17168), .ZN(n17169) );
  NOR2_X1 U20380 ( .A1(n17169), .A2(n17222), .ZN(n17205) );
  NAND3_X1 U20381 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(n17205), .ZN(n17195) );
  NAND2_X1 U20382 ( .A1(n17170), .A2(n17189), .ZN(n17174) );
  INV_X1 U20383 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20384 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17234), .B1(n17233), .B2(
        n17171), .ZN(n17172) );
  OAI221_X1 U20385 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17174), .C1(n17342), 
        .C2(n17173), .A(n17172), .ZN(P3_U2721) );
  INV_X1 U20386 ( .A(n17174), .ZN(n17178) );
  NAND2_X1 U20387 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17175) );
  NAND2_X1 U20388 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17189), .ZN(n17188) );
  NOR2_X1 U20389 ( .A1(n17175), .A2(n17188), .ZN(n17183) );
  AOI21_X1 U20390 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17225), .A(n17183), .ZN(
        n17177) );
  OAI222_X1 U20391 ( .A1(n17229), .A2(n17179), .B1(n17178), .B2(n17177), .C1(
        n17226), .C2(n17176), .ZN(P3_U2722) );
  INV_X1 U20392 ( .A(n17188), .ZN(n17180) );
  AOI22_X1 U20393 ( .A1(n17180), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17215), .ZN(n17182) );
  OAI222_X1 U20394 ( .A1(n17229), .A2(n17184), .B1(n17183), .B2(n17182), .C1(
        n17226), .C2(n17181), .ZN(P3_U2723) );
  NAND2_X1 U20395 ( .A1(n17225), .A2(n17188), .ZN(n17192) );
  INV_X1 U20396 ( .A(n17185), .ZN(n17186) );
  AOI22_X1 U20397 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17234), .B1(n17233), .B2(
        n17186), .ZN(n17187) );
  OAI221_X1 U20398 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17188), .C1(n17336), 
        .C2(n17192), .A(n17187), .ZN(P3_U2724) );
  NOR2_X1 U20399 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17189), .ZN(n17191) );
  OAI222_X1 U20400 ( .A1(n17229), .A2(n17193), .B1(n17192), .B2(n17191), .C1(
        n17226), .C2(n17190), .ZN(P3_U2725) );
  AOI22_X1 U20401 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17234), .B1(n17233), .B2(
        n17194), .ZN(n17197) );
  OAI211_X1 U20402 ( .C1(P3_EAX_REG_9__SCAN_IN), .C2(n17198), .A(n17225), .B(
        n17195), .ZN(n17196) );
  NAND2_X1 U20403 ( .A1(n17197), .A2(n17196), .ZN(P3_U2726) );
  AOI211_X1 U20404 ( .C1(n17329), .C2(n17199), .A(n17237), .B(n17198), .ZN(
        n17200) );
  AOI21_X1 U20405 ( .B1(n17233), .B2(n17201), .A(n17200), .ZN(n17202) );
  OAI21_X1 U20406 ( .B1(n17203), .B2(n17229), .A(n17202), .ZN(P3_U2727) );
  INV_X1 U20407 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17325) );
  INV_X1 U20408 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17321) );
  INV_X1 U20409 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17317) );
  NOR3_X1 U20410 ( .A1(n17223), .A2(n17317), .A3(n17222), .ZN(n17228) );
  NAND2_X1 U20411 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17228), .ZN(n17214) );
  NOR2_X1 U20412 ( .A1(n17321), .A2(n17214), .ZN(n17218) );
  NAND2_X1 U20413 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17218), .ZN(n17207) );
  NOR2_X1 U20414 ( .A1(n17325), .A2(n17207), .ZN(n17210) );
  AOI21_X1 U20415 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17225), .A(n17210), .ZN(
        n17206) );
  OAI222_X1 U20416 ( .A1(n17229), .A2(n20841), .B1(n17206), .B2(n17205), .C1(
        n17226), .C2(n17204), .ZN(P3_U2728) );
  INV_X1 U20417 ( .A(n17207), .ZN(n17213) );
  AOI21_X1 U20418 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17225), .A(n17213), .ZN(
        n17209) );
  OAI222_X1 U20419 ( .A1(n18090), .A2(n17229), .B1(n17210), .B2(n17209), .C1(
        n17226), .C2(n17208), .ZN(P3_U2729) );
  AOI21_X1 U20420 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17225), .A(n17218), .ZN(
        n17212) );
  OAI222_X1 U20421 ( .A1(n18084), .A2(n17229), .B1(n17213), .B2(n17212), .C1(
        n17226), .C2(n17211), .ZN(P3_U2730) );
  INV_X1 U20422 ( .A(n17214), .ZN(n17221) );
  AOI21_X1 U20423 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17215), .A(n17221), .ZN(
        n17217) );
  OAI222_X1 U20424 ( .A1(n18079), .A2(n17229), .B1(n17218), .B2(n17217), .C1(
        n17226), .C2(n17216), .ZN(P3_U2731) );
  AOI21_X1 U20425 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17225), .A(n17228), .ZN(
        n17220) );
  OAI222_X1 U20426 ( .A1(n18074), .A2(n17229), .B1(n17221), .B2(n17220), .C1(
        n17226), .C2(n17219), .ZN(P3_U2732) );
  NOR2_X1 U20427 ( .A1(n17223), .A2(n17222), .ZN(n17224) );
  AOI21_X1 U20428 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17225), .A(n17224), .ZN(
        n17227) );
  OAI222_X1 U20429 ( .A1(n18068), .A2(n17229), .B1(n17228), .B2(n17227), .C1(
        n17226), .C2(n10128), .ZN(P3_U2733) );
  NAND2_X1 U20430 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17230), .ZN(n17231) );
  XOR2_X1 U20431 ( .A(P3_EAX_REG_1__SCAN_IN), .B(n17231), .Z(n17236) );
  AOI22_X1 U20432 ( .A1(n17234), .A2(BUF2_REG_1__SCAN_IN), .B1(n17233), .B2(
        n17232), .ZN(n17235) );
  OAI21_X1 U20433 ( .B1(n17237), .B2(n17236), .A(n17235), .ZN(P3_U2734) );
  INV_X1 U20434 ( .A(n17546), .ZN(n17707) );
  NOR2_X1 U20435 ( .A1(n17709), .A2(n17707), .ZN(n17266) );
  AND2_X1 U20436 ( .A1(n17268), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20437 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17311) );
  NAND2_X1 U20438 ( .A1(n17256), .A2(n17239), .ZN(n17255) );
  AOI22_X1 U20439 ( .A1(n18703), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17240) );
  OAI21_X1 U20440 ( .B1(n17311), .B2(n17255), .A(n17240), .ZN(P3_U2737) );
  INV_X1 U20441 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20442 ( .A1(n18703), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17241) );
  OAI21_X1 U20443 ( .B1(n17309), .B2(n17255), .A(n17241), .ZN(P3_U2738) );
  AOI22_X1 U20444 ( .A1(n18703), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17242) );
  OAI21_X1 U20445 ( .B1(n17307), .B2(n17255), .A(n17242), .ZN(P3_U2739) );
  INV_X1 U20446 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U20447 ( .A1(n18703), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17243) );
  OAI21_X1 U20448 ( .B1(n17304), .B2(n17255), .A(n17243), .ZN(P3_U2740) );
  AOI22_X1 U20449 ( .A1(n18703), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17244) );
  OAI21_X1 U20450 ( .B1(n17302), .B2(n17255), .A(n17244), .ZN(P3_U2741) );
  INV_X1 U20451 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20452 ( .A1(n18703), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17245) );
  OAI21_X1 U20453 ( .B1(n17300), .B2(n17255), .A(n17245), .ZN(P3_U2742) );
  INV_X1 U20454 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U20455 ( .A1(n18703), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17246) );
  OAI21_X1 U20456 ( .B1(n17298), .B2(n17255), .A(n17246), .ZN(P3_U2743) );
  INV_X1 U20457 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20458 ( .A1(n18703), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17247) );
  OAI21_X1 U20459 ( .B1(n17296), .B2(n17255), .A(n17247), .ZN(P3_U2744) );
  AOI22_X1 U20460 ( .A1(n18703), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17248) );
  OAI21_X1 U20461 ( .B1(n17294), .B2(n17255), .A(n17248), .ZN(P3_U2745) );
  AOI22_X1 U20462 ( .A1(n17266), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17249) );
  OAI21_X1 U20463 ( .B1(n17292), .B2(n17255), .A(n17249), .ZN(P3_U2746) );
  INV_X1 U20464 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17290) );
  AOI22_X1 U20465 ( .A1(n17266), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17250) );
  OAI21_X1 U20466 ( .B1(n17290), .B2(n17255), .A(n17250), .ZN(P3_U2747) );
  AOI22_X1 U20467 ( .A1(n17266), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17251) );
  OAI21_X1 U20468 ( .B1(n20845), .B2(n17255), .A(n17251), .ZN(P3_U2748) );
  INV_X1 U20469 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20470 ( .A1(n17266), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17252) );
  OAI21_X1 U20471 ( .B1(n17287), .B2(n17255), .A(n17252), .ZN(P3_U2749) );
  AOI22_X1 U20472 ( .A1(n17266), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17253) );
  OAI21_X1 U20473 ( .B1(n17285), .B2(n17255), .A(n17253), .ZN(P3_U2750) );
  INV_X1 U20474 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20475 ( .A1(n17266), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17254) );
  OAI21_X1 U20476 ( .B1(n17283), .B2(n17255), .A(n17254), .ZN(P3_U2751) );
  AOI22_X1 U20477 ( .A1(n17266), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17257) );
  OAI21_X1 U20478 ( .B1(n20940), .B2(n17276), .A(n17257), .ZN(P3_U2752) );
  AOI22_X1 U20479 ( .A1(n17266), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17258) );
  OAI21_X1 U20480 ( .B1(n17342), .B2(n17276), .A(n17258), .ZN(P3_U2753) );
  AOI22_X1 U20481 ( .A1(n17266), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17259) );
  OAI21_X1 U20482 ( .B1(n17340), .B2(n17276), .A(n17259), .ZN(P3_U2754) );
  AOI22_X1 U20483 ( .A1(n17266), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17260) );
  OAI21_X1 U20484 ( .B1(n17338), .B2(n17276), .A(n17260), .ZN(P3_U2755) );
  AOI22_X1 U20485 ( .A1(n18703), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17261) );
  OAI21_X1 U20486 ( .B1(n17336), .B2(n17276), .A(n17261), .ZN(P3_U2756) );
  AOI22_X1 U20487 ( .A1(n18703), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17262) );
  OAI21_X1 U20488 ( .B1(n17333), .B2(n17276), .A(n17262), .ZN(P3_U2757) );
  INV_X1 U20489 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U20490 ( .A1(n18703), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17263) );
  OAI21_X1 U20491 ( .B1(n17331), .B2(n17276), .A(n17263), .ZN(P3_U2758) );
  AOI22_X1 U20492 ( .A1(n18703), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17264) );
  OAI21_X1 U20493 ( .B1(n17329), .B2(n17276), .A(n17264), .ZN(P3_U2759) );
  AOI22_X1 U20494 ( .A1(n18703), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17265) );
  OAI21_X1 U20495 ( .B1(n17327), .B2(n17276), .A(n17265), .ZN(P3_U2760) );
  AOI22_X1 U20496 ( .A1(n17266), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17267) );
  OAI21_X1 U20497 ( .B1(n17325), .B2(n17276), .A(n17267), .ZN(P3_U2761) );
  INV_X1 U20498 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20499 ( .A1(n18703), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17268), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17269) );
  OAI21_X1 U20500 ( .B1(n17323), .B2(n17276), .A(n17269), .ZN(P3_U2762) );
  AOI22_X1 U20501 ( .A1(n18703), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17270) );
  OAI21_X1 U20502 ( .B1(n17321), .B2(n17276), .A(n17270), .ZN(P3_U2763) );
  AOI22_X1 U20503 ( .A1(n18703), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17271) );
  OAI21_X1 U20504 ( .B1(n17319), .B2(n17276), .A(n17271), .ZN(P3_U2764) );
  AOI22_X1 U20505 ( .A1(n18703), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20506 ( .B1(n17317), .B2(n17276), .A(n17272), .ZN(P3_U2765) );
  INV_X1 U20507 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20508 ( .A1(n18703), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17273) );
  OAI21_X1 U20509 ( .B1(n17315), .B2(n17276), .A(n17273), .ZN(P3_U2766) );
  AOI22_X1 U20510 ( .A1(n18703), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17274), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17275) );
  OAI21_X1 U20511 ( .B1(n17313), .B2(n17276), .A(n17275), .ZN(P3_U2767) );
  INV_X1 U20512 ( .A(n17277), .ZN(n17280) );
  NOR3_X1 U20513 ( .A1(n18062), .A2(n17279), .A3(n17278), .ZN(n17305) );
  OAI211_X1 U20514 ( .C1(n18062), .C2(n18702), .A(n17281), .B(n17280), .ZN(
        n17334) );
  AOI22_X1 U20515 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17343), .ZN(n17282) );
  OAI21_X1 U20516 ( .B1(n17283), .B2(n17345), .A(n17282), .ZN(P3_U2768) );
  AOI22_X1 U20517 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17343), .ZN(n17284) );
  OAI21_X1 U20518 ( .B1(n17285), .B2(n17345), .A(n17284), .ZN(P3_U2769) );
  AOI22_X1 U20519 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17343), .ZN(n17286) );
  OAI21_X1 U20520 ( .B1(n17287), .B2(n17345), .A(n17286), .ZN(P3_U2770) );
  AOI22_X1 U20521 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17343), .ZN(n17288) );
  OAI21_X1 U20522 ( .B1(n20845), .B2(n17345), .A(n17288), .ZN(P3_U2771) );
  AOI22_X1 U20523 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17343), .ZN(n17289) );
  OAI21_X1 U20524 ( .B1(n17290), .B2(n17345), .A(n17289), .ZN(P3_U2772) );
  AOI22_X1 U20525 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17334), .ZN(n17291) );
  OAI21_X1 U20526 ( .B1(n17292), .B2(n17345), .A(n17291), .ZN(P3_U2773) );
  AOI22_X1 U20527 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17334), .ZN(n17293) );
  OAI21_X1 U20528 ( .B1(n17294), .B2(n17345), .A(n17293), .ZN(P3_U2774) );
  AOI22_X1 U20529 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17334), .ZN(n17295) );
  OAI21_X1 U20530 ( .B1(n17296), .B2(n17345), .A(n17295), .ZN(P3_U2775) );
  AOI22_X1 U20531 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17334), .ZN(n17297) );
  OAI21_X1 U20532 ( .B1(n17298), .B2(n17345), .A(n17297), .ZN(P3_U2776) );
  AOI22_X1 U20533 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17334), .ZN(n17299) );
  OAI21_X1 U20534 ( .B1(n17300), .B2(n17345), .A(n17299), .ZN(P3_U2777) );
  AOI22_X1 U20535 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17334), .ZN(n17301) );
  OAI21_X1 U20536 ( .B1(n17302), .B2(n17345), .A(n17301), .ZN(P3_U2778) );
  AOI22_X1 U20537 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17334), .ZN(n17303) );
  OAI21_X1 U20538 ( .B1(n17304), .B2(n17345), .A(n17303), .ZN(P3_U2779) );
  AOI22_X1 U20539 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17343), .ZN(n17306) );
  OAI21_X1 U20540 ( .B1(n17307), .B2(n17345), .A(n17306), .ZN(P3_U2780) );
  AOI22_X1 U20541 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17343), .ZN(n17308) );
  OAI21_X1 U20542 ( .B1(n17309), .B2(n17345), .A(n17308), .ZN(P3_U2781) );
  AOI22_X1 U20543 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n9796), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17343), .ZN(n17310) );
  OAI21_X1 U20544 ( .B1(n17311), .B2(n17345), .A(n17310), .ZN(P3_U2782) );
  AOI22_X1 U20545 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17343), .ZN(n17312) );
  OAI21_X1 U20546 ( .B1(n17313), .B2(n17345), .A(n17312), .ZN(P3_U2783) );
  AOI22_X1 U20547 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17343), .ZN(n17314) );
  OAI21_X1 U20548 ( .B1(n17315), .B2(n17345), .A(n17314), .ZN(P3_U2784) );
  AOI22_X1 U20549 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17343), .ZN(n17316) );
  OAI21_X1 U20550 ( .B1(n17317), .B2(n17345), .A(n17316), .ZN(P3_U2785) );
  AOI22_X1 U20551 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17343), .ZN(n17318) );
  OAI21_X1 U20552 ( .B1(n17319), .B2(n17345), .A(n17318), .ZN(P3_U2786) );
  AOI22_X1 U20553 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17343), .ZN(n17320) );
  OAI21_X1 U20554 ( .B1(n17321), .B2(n17345), .A(n17320), .ZN(P3_U2787) );
  AOI22_X1 U20555 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17343), .ZN(n17322) );
  OAI21_X1 U20556 ( .B1(n17323), .B2(n17345), .A(n17322), .ZN(P3_U2788) );
  AOI22_X1 U20557 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17343), .ZN(n17324) );
  OAI21_X1 U20558 ( .B1(n17325), .B2(n17345), .A(n17324), .ZN(P3_U2789) );
  AOI22_X1 U20559 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17343), .ZN(n17326) );
  OAI21_X1 U20560 ( .B1(n17327), .B2(n17345), .A(n17326), .ZN(P3_U2790) );
  AOI22_X1 U20561 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17343), .ZN(n17328) );
  OAI21_X1 U20562 ( .B1(n17329), .B2(n17345), .A(n17328), .ZN(P3_U2791) );
  AOI22_X1 U20563 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17334), .ZN(n17330) );
  OAI21_X1 U20564 ( .B1(n17331), .B2(n17345), .A(n17330), .ZN(P3_U2792) );
  AOI22_X1 U20565 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17334), .ZN(n17332) );
  OAI21_X1 U20566 ( .B1(n17333), .B2(n17345), .A(n17332), .ZN(P3_U2793) );
  AOI22_X1 U20567 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17334), .ZN(n17335) );
  OAI21_X1 U20568 ( .B1(n17336), .B2(n17345), .A(n17335), .ZN(P3_U2794) );
  AOI22_X1 U20569 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17343), .ZN(n17337) );
  OAI21_X1 U20570 ( .B1(n17338), .B2(n17345), .A(n17337), .ZN(P3_U2795) );
  AOI22_X1 U20571 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17343), .ZN(n17339) );
  OAI21_X1 U20572 ( .B1(n17340), .B2(n17345), .A(n17339), .ZN(P3_U2796) );
  AOI22_X1 U20573 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17343), .ZN(n17341) );
  OAI21_X1 U20574 ( .B1(n17342), .B2(n17345), .A(n17341), .ZN(P3_U2797) );
  AOI22_X1 U20575 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n9796), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17343), .ZN(n17344) );
  OAI21_X1 U20576 ( .B1(n20940), .B2(n17345), .A(n17344), .ZN(P3_U2798) );
  OAI21_X1 U20577 ( .B1(n17348), .B2(n17347), .A(n17346), .ZN(n17362) );
  OAI21_X1 U20578 ( .B1(n17349), .B2(n17707), .A(n17708), .ZN(n17350) );
  AOI21_X1 U20579 ( .B1(n17667), .B2(n17352), .A(n17350), .ZN(n17386) );
  OAI21_X1 U20580 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17457), .A(
        n17386), .ZN(n17363) );
  NOR3_X1 U20581 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17351), .A3(
        n17430), .ZN(n17358) );
  NOR2_X1 U20582 ( .A1(n17472), .A2(n17352), .ZN(n17368) );
  OAI211_X1 U20583 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17368), .B(n17353), .ZN(n17354) );
  OAI211_X1 U20584 ( .C1(n17549), .C2(n17356), .A(n17355), .B(n17354), .ZN(
        n17357) );
  AOI211_X1 U20585 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17363), .A(
        n17358), .B(n17357), .ZN(n17361) );
  AOI22_X1 U20586 ( .A1(n9792), .A2(n17359), .B1(n17543), .B2(n17723), .ZN(
        n17381) );
  NAND2_X1 U20587 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17381), .ZN(
        n17369) );
  OAI211_X1 U20588 ( .C1(n17698), .C2(n17543), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17369), .ZN(n17360) );
  OAI211_X1 U20589 ( .C1(n17606), .C2(n17362), .A(n17361), .B(n17360), .ZN(
        P3_U2802) );
  AOI22_X1 U20590 ( .A1(n17565), .A2(n17364), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17363), .ZN(n17373) );
  OAI21_X1 U20591 ( .B1(n17617), .B2(n17366), .A(n17365), .ZN(n17726) );
  AOI22_X1 U20592 ( .A1(n17618), .A2(n17726), .B1(n17368), .B2(n17367), .ZN(
        n17372) );
  NOR2_X1 U20593 ( .A1(n17715), .A2(n17430), .ZN(n17370) );
  OAI21_X1 U20594 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17370), .A(
        n17369), .ZN(n17371) );
  NAND2_X1 U20595 ( .A1(n18035), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17728) );
  NAND4_X1 U20596 ( .A1(n17373), .A2(n17372), .A3(n17371), .A4(n17728), .ZN(
        P3_U2803) );
  AOI21_X1 U20597 ( .B1(n17374), .B2(n18442), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17385) );
  INV_X1 U20598 ( .A(n17457), .ZN(n17375) );
  INV_X1 U20599 ( .A(n17693), .ZN(n17376) );
  AOI22_X1 U20600 ( .A1(n18035), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17377), 
        .B2(n17376), .ZN(n17384) );
  NOR3_X1 U20601 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17765), .A3(
        n17753), .ZN(n17731) );
  INV_X1 U20602 ( .A(n17378), .ZN(n17443) );
  NOR2_X1 U20603 ( .A1(n17732), .A2(n17443), .ZN(n17411) );
  AOI21_X1 U20604 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17380), .A(
        n17379), .ZN(n17740) );
  OAI22_X1 U20605 ( .A1(n17381), .A2(n17735), .B1(n17740), .B2(n17606), .ZN(
        n17382) );
  AOI21_X1 U20606 ( .B1(n17731), .B2(n17411), .A(n17382), .ZN(n17383) );
  OAI211_X1 U20607 ( .C1(n17386), .C2(n17385), .A(n17384), .B(n17383), .ZN(
        P3_U2804) );
  OAI21_X1 U20608 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17388), .A(
        n17387), .ZN(n17741) );
  INV_X1 U20609 ( .A(n17389), .ZN(n17423) );
  OAI21_X1 U20610 ( .B1(n17390), .B2(n18132), .A(n17708), .ZN(n17391) );
  AOI21_X1 U20611 ( .B1(n17546), .B2(n17423), .A(n17391), .ZN(n17422) );
  OAI21_X1 U20612 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17457), .A(
        n17422), .ZN(n17405) );
  NOR2_X1 U20613 ( .A1(n17472), .A2(n17392), .ZN(n17407) );
  OAI211_X1 U20614 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17407), .B(n17393), .ZN(n17394) );
  NAND2_X1 U20615 ( .A1(n18035), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17752) );
  OAI211_X1 U20616 ( .C1(n17549), .C2(n17395), .A(n17394), .B(n17752), .ZN(
        n17402) );
  OAI21_X1 U20617 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17397), .A(
        n17396), .ZN(n17757) );
  OAI21_X1 U20618 ( .B1(n15647), .B2(n17399), .A(n17398), .ZN(n17400) );
  XNOR2_X1 U20619 ( .A(n17400), .B(n17753), .ZN(n17742) );
  OAI22_X1 U20620 ( .A1(n17713), .A2(n17757), .B1(n17606), .B2(n17742), .ZN(
        n17401) );
  AOI211_X1 U20621 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17405), .A(
        n17402), .B(n17401), .ZN(n17403) );
  OAI21_X1 U20622 ( .B1(n17621), .B2(n17741), .A(n17403), .ZN(P3_U2805) );
  INV_X1 U20623 ( .A(n17404), .ZN(n17414) );
  NOR2_X1 U20624 ( .A1(n9800), .A2(n18630), .ZN(n17770) );
  AOI221_X1 U20625 ( .B1(n17407), .B2(n17406), .C1(n17405), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17770), .ZN(n17413) );
  AOI22_X1 U20626 ( .A1(n17698), .A2(n17758), .B1(n17543), .B2(n17762), .ZN(
        n17428) );
  AOI21_X1 U20627 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17409), .A(
        n17408), .ZN(n17772) );
  OAI22_X1 U20628 ( .A1(n17428), .A2(n17765), .B1(n17772), .B2(n17606), .ZN(
        n17410) );
  AOI21_X1 U20629 ( .B1(n17411), .B2(n17765), .A(n17410), .ZN(n17412) );
  OAI211_X1 U20630 ( .C1(n17549), .C2(n17414), .A(n17413), .B(n17412), .ZN(
        P3_U2806) );
  AOI22_X1 U20631 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15647), .B1(
        n17416), .B2(n17432), .ZN(n17417) );
  NAND2_X1 U20632 ( .A1(n17415), .A2(n17417), .ZN(n17418) );
  XNOR2_X1 U20633 ( .A(n17418), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17774) );
  AOI21_X1 U20634 ( .B1(n17419), .B2(n18442), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17421) );
  OAI22_X1 U20635 ( .A1(n17422), .A2(n17421), .B1(n17549), .B2(n17420), .ZN(
        n17426) );
  OR2_X1 U20636 ( .A1(n17457), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17424) );
  OAI22_X1 U20637 ( .A1(n9800), .A2(n18629), .B1(n17424), .B2(n17423), .ZN(
        n17425) );
  AOI211_X1 U20638 ( .C1(n17618), .C2(n17774), .A(n17426), .B(n17425), .ZN(
        n17427) );
  OAI221_X1 U20639 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17430), 
        .C1(n17429), .C2(n17428), .A(n17427), .ZN(P3_U2807) );
  INV_X1 U20640 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17793) );
  NAND2_X1 U20641 ( .A1(n17713), .A2(n17621), .ZN(n17462) );
  OAI22_X1 U20642 ( .A1(n17867), .A2(n17713), .B1(n17856), .B2(n17621), .ZN(
        n17463) );
  AOI21_X1 U20643 ( .B1(n17779), .B2(n17462), .A(n17463), .ZN(n17455) );
  INV_X1 U20644 ( .A(n17415), .ZN(n17431) );
  AOI221_X1 U20645 ( .B1(n17502), .B2(n17432), .C1(n17779), .C2(n17432), .A(
        n17431), .ZN(n17433) );
  XOR2_X1 U20646 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17433), .Z(
        n17789) );
  OAI21_X1 U20647 ( .B1(n17434), .B2(n17707), .A(n17708), .ZN(n17435) );
  AOI21_X1 U20648 ( .B1(n17667), .B2(n17437), .A(n17435), .ZN(n17459) );
  OAI21_X1 U20649 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17457), .A(
        n17459), .ZN(n17446) );
  AOI22_X1 U20650 ( .A1(n17565), .A2(n17436), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17446), .ZN(n17440) );
  NOR2_X1 U20651 ( .A1(n17472), .A2(n17437), .ZN(n17448) );
  OAI211_X1 U20652 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17448), .B(n17438), .ZN(n17439) );
  OAI211_X1 U20653 ( .C1(n20836), .C2(n9800), .A(n17440), .B(n17439), .ZN(
        n17441) );
  AOI21_X1 U20654 ( .B1(n17618), .B2(n17789), .A(n17441), .ZN(n17442) );
  OAI221_X1 U20655 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17443), 
        .C1(n17793), .C2(n17455), .A(n17442), .ZN(P3_U2808) );
  OAI22_X1 U20656 ( .A1(n9800), .A2(n18626), .B1(n17549), .B2(n17444), .ZN(
        n17445) );
  AOI221_X1 U20657 ( .B1(n17448), .B2(n17447), .C1(n17446), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17445), .ZN(n17454) );
  INV_X1 U20658 ( .A(n17452), .ZN(n17799) );
  NOR3_X1 U20659 ( .A1(n15647), .A2(n17830), .A3(n17449), .ZN(n17467) );
  INV_X1 U20660 ( .A(n17487), .ZN(n17468) );
  AOI22_X1 U20661 ( .A1(n17799), .A2(n17467), .B1(n17468), .B2(n17450), .ZN(
        n17451) );
  XNOR2_X1 U20662 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17451), .ZN(
        n17803) );
  NOR2_X1 U20663 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17452), .ZN(
        n17802) );
  NAND2_X1 U20664 ( .A1(n17827), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17794) );
  NOR2_X1 U20665 ( .A1(n17514), .A2(n17794), .ZN(n17479) );
  AOI22_X1 U20666 ( .A1(n17618), .A2(n17803), .B1(n17802), .B2(n17479), .ZN(
        n17453) );
  OAI211_X1 U20667 ( .C1(n17455), .C2(n17783), .A(n17454), .B(n17453), .ZN(
        P3_U2809) );
  INV_X1 U20668 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17780) );
  OAI221_X1 U20669 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17486), 
        .C1(n17814), .C2(n17467), .A(n17415), .ZN(n17456) );
  XNOR2_X1 U20670 ( .A(n17780), .B(n17456), .ZN(n17813) );
  AOI21_X1 U20671 ( .B1(n9869), .B2(n18442), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17458) );
  OAI22_X1 U20672 ( .A1(n17459), .A2(n17458), .B1(n9800), .B2(n18623), .ZN(
        n17460) );
  AOI221_X1 U20673 ( .B1(n17565), .B2(n17461), .C1(n17375), .C2(n17461), .A(
        n17460), .ZN(n17466) );
  INV_X1 U20674 ( .A(n17462), .ZN(n17464) );
  NOR2_X1 U20675 ( .A1(n17814), .A2(n17794), .ZN(n17809) );
  INV_X1 U20676 ( .A(n17463), .ZN(n17513) );
  OAI21_X1 U20677 ( .B1(n17464), .B2(n17809), .A(n17513), .ZN(n17478) );
  NOR2_X1 U20678 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17814), .ZN(
        n17806) );
  AOI22_X1 U20679 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17478), .B1(
        n17479), .B2(n17806), .ZN(n17465) );
  OAI211_X1 U20680 ( .C1(n17606), .C2(n17813), .A(n17466), .B(n17465), .ZN(
        P3_U2810) );
  AOI21_X1 U20681 ( .B1(n17468), .B2(n17486), .A(n17467), .ZN(n17469) );
  XNOR2_X1 U20682 ( .A(n17469), .B(n17814), .ZN(n17819) );
  INV_X1 U20683 ( .A(n17708), .ZN(n17682) );
  AOI21_X1 U20684 ( .B1(n17667), .B2(n17471), .A(n17682), .ZN(n17493) );
  OAI21_X1 U20685 ( .B1(n17470), .B2(n17707), .A(n17493), .ZN(n17483) );
  AOI22_X1 U20686 ( .A1(n18035), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17483), .ZN(n17475) );
  NOR2_X1 U20687 ( .A1(n17472), .A2(n17471), .ZN(n17485) );
  OAI211_X1 U20688 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17485), .B(n17473), .ZN(n17474) );
  OAI211_X1 U20689 ( .C1(n17549), .C2(n17476), .A(n17475), .B(n17474), .ZN(
        n17477) );
  AOI221_X1 U20690 ( .B1(n17479), .B2(n17814), .C1(n17478), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17477), .ZN(n17480) );
  OAI21_X1 U20691 ( .B1(n17819), .B2(n17606), .A(n17480), .ZN(P3_U2811) );
  NAND2_X1 U20692 ( .A1(n17827), .A2(n17830), .ZN(n17836) );
  INV_X1 U20693 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17484) );
  INV_X1 U20694 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18619) );
  OAI22_X1 U20695 ( .A1(n9800), .A2(n18619), .B1(n17549), .B2(n17481), .ZN(
        n17482) );
  AOI221_X1 U20696 ( .B1(n17485), .B2(n17484), .C1(n17483), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17482), .ZN(n17490) );
  OAI21_X1 U20697 ( .B1(n17827), .B2(n17514), .A(n17513), .ZN(n17498) );
  AOI21_X1 U20698 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17617), .A(
        n17486), .ZN(n17488) );
  XNOR2_X1 U20699 ( .A(n17488), .B(n17487), .ZN(n17833) );
  AOI22_X1 U20700 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17498), .B1(
        n17618), .B2(n17833), .ZN(n17489) );
  OAI211_X1 U20701 ( .C1(n17514), .C2(n17836), .A(n17490), .B(n17489), .ZN(
        P3_U2812) );
  NAND2_X1 U20702 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17837), .ZN(
        n17843) );
  AOI21_X1 U20703 ( .B1(n17491), .B2(n18442), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17494) );
  OAI22_X1 U20704 ( .A1(n17494), .A2(n17493), .B1(n17693), .B2(n17492), .ZN(
        n17495) );
  AOI21_X1 U20705 ( .B1(n18035), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17495), 
        .ZN(n17500) );
  OAI21_X1 U20706 ( .B1(n17497), .B2(n17837), .A(n17496), .ZN(n17840) );
  AOI22_X1 U20707 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17498), .B1(
        n17618), .B2(n17840), .ZN(n17499) );
  OAI211_X1 U20708 ( .C1(n17514), .C2(n17843), .A(n17500), .B(n17499), .ZN(
        P3_U2813) );
  AOI21_X1 U20709 ( .B1(n17617), .B2(n17502), .A(n17501), .ZN(n17503) );
  XNOR2_X1 U20710 ( .A(n17503), .B(n17848), .ZN(n17852) );
  NAND3_X1 U20711 ( .A1(n17504), .A2(n17562), .A3(n17561), .ZN(n17516) );
  OAI21_X1 U20712 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17505), .ZN(n17510) );
  AOI21_X1 U20713 ( .B1(n17667), .B2(n17506), .A(n17682), .ZN(n17532) );
  OAI21_X1 U20714 ( .B1(n17507), .B2(n17707), .A(n17532), .ZN(n17518) );
  AOI22_X1 U20715 ( .A1(n17565), .A2(n17508), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17518), .ZN(n17509) );
  NAND2_X1 U20716 ( .A1(n18035), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17853) );
  OAI211_X1 U20717 ( .C1(n17516), .C2(n17510), .A(n17509), .B(n17853), .ZN(
        n17511) );
  AOI21_X1 U20718 ( .B1(n17618), .B2(n17852), .A(n17511), .ZN(n17512) );
  OAI221_X1 U20719 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17514), 
        .C1(n17848), .C2(n17513), .A(n17512), .ZN(P3_U2814) );
  INV_X1 U20720 ( .A(n17524), .ZN(n17846) );
  NOR2_X1 U20721 ( .A1(n9952), .A2(n17846), .ZN(n17537) );
  NOR2_X1 U20722 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17537), .ZN(
        n17857) );
  OR2_X1 U20723 ( .A1(n17621), .A2(n17856), .ZN(n17528) );
  NOR2_X1 U20724 ( .A1(n9800), .A2(n18613), .ZN(n17866) );
  OAI22_X1 U20725 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17516), .B1(
        n17549), .B2(n17515), .ZN(n17517) );
  AOI211_X1 U20726 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17518), .A(
        n17866), .B(n17517), .ZN(n17527) );
  INV_X1 U20727 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17884) );
  OAI21_X1 U20728 ( .B1(n17521), .B2(n17519), .A(n17520), .ZN(n17522) );
  OAI221_X1 U20729 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17884), 
        .C1(n17903), .C2(n17617), .A(n17522), .ZN(n17523) );
  XNOR2_X1 U20730 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17523), .ZN(
        n17870) );
  NOR2_X1 U20731 ( .A1(n17867), .A2(n17713), .ZN(n17525) );
  INV_X1 U20732 ( .A(n17529), .ZN(n17913) );
  NAND2_X1 U20733 ( .A1(n17524), .A2(n17913), .ZN(n17530) );
  NAND2_X1 U20734 ( .A1(n17862), .A2(n17530), .ZN(n17868) );
  AOI22_X1 U20735 ( .A1(n17618), .A2(n17870), .B1(n17525), .B2(n17868), .ZN(
        n17526) );
  OAI211_X1 U20736 ( .C1(n17857), .C2(n17528), .A(n17527), .B(n17526), .ZN(
        P3_U2815) );
  NAND2_X1 U20737 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17906), .ZN(
        n17881) );
  NOR2_X1 U20738 ( .A1(n17529), .A2(n17881), .ZN(n17896) );
  OAI221_X1 U20739 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17896), .A(n17530), .ZN(
        n17892) );
  NOR2_X1 U20740 ( .A1(n17531), .A2(n18132), .ZN(n17612) );
  NAND2_X1 U20741 ( .A1(n9912), .A2(n17612), .ZN(n17576) );
  AOI221_X1 U20742 ( .B1(n17534), .B2(n17533), .C1(n17576), .C2(n17533), .A(
        n17532), .ZN(n17535) );
  NOR2_X1 U20743 ( .A1(n9800), .A2(n18612), .ZN(n17886) );
  AOI211_X1 U20744 ( .C1(n17536), .C2(n17376), .A(n17535), .B(n17886), .ZN(
        n17542) );
  INV_X1 U20745 ( .A(n17881), .ZN(n17877) );
  NAND2_X1 U20746 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17877), .ZN(
        n17858) );
  NOR2_X1 U20747 ( .A1(n15647), .A2(n9952), .ZN(n17596) );
  INV_X1 U20748 ( .A(n17858), .ZN(n17539) );
  AOI21_X1 U20749 ( .B1(n17596), .B2(n17539), .A(n17538), .ZN(n17540) );
  XNOR2_X1 U20750 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17540), .ZN(
        n17889) );
  AOI22_X1 U20751 ( .A1(n17543), .A2(n17887), .B1(n17618), .B2(n17889), .ZN(
        n17541) );
  OAI211_X1 U20752 ( .C1(n17713), .C2(n17892), .A(n17542), .B(n17541), .ZN(
        P3_U2816) );
  INV_X1 U20753 ( .A(n17896), .ZN(n17544) );
  NAND2_X1 U20754 ( .A1(n17916), .A2(n17877), .ZN(n17893) );
  AOI22_X1 U20755 ( .A1(n9792), .A2(n17544), .B1(n17543), .B2(n17893), .ZN(
        n17570) );
  AOI21_X1 U20756 ( .B1(n17546), .B2(n17545), .A(n17682), .ZN(n17547) );
  OAI21_X1 U20757 ( .B1(n17562), .B2(n17681), .A(n17547), .ZN(n17563) );
  NOR2_X1 U20758 ( .A1(n9800), .A2(n18609), .ZN(n17553) );
  OAI211_X1 U20759 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17562), .B(n17561), .ZN(n17550) );
  OAI22_X1 U20760 ( .A1(n17551), .A2(n17550), .B1(n17549), .B2(n17548), .ZN(
        n17552) );
  AOI211_X1 U20761 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17563), .A(
        n17553), .B(n17552), .ZN(n17557) );
  OAI22_X1 U20762 ( .A1(n17617), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n17881), .B2(n17519), .ZN(n17554) );
  OAI21_X1 U20763 ( .B1(n17617), .B2(n17559), .A(n17554), .ZN(n17555) );
  XNOR2_X1 U20764 ( .A(n17555), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17900) );
  NOR2_X1 U20765 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17881), .ZN(
        n17899) );
  AOI22_X1 U20766 ( .A1(n17618), .A2(n17900), .B1(n17899), .B2(n17603), .ZN(
        n17556) );
  OAI211_X1 U20767 ( .C1(n17570), .C2(n17558), .A(n17557), .B(n17556), .ZN(
        P3_U2817) );
  NAND2_X1 U20768 ( .A1(n17906), .A2(n17603), .ZN(n17571) );
  AOI21_X1 U20769 ( .B1(n17906), .B2(n17596), .A(n17559), .ZN(n17560) );
  XNOR2_X1 U20770 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17560), .ZN(
        n17907) );
  NAND2_X1 U20771 ( .A1(n17562), .A2(n17561), .ZN(n17567) );
  AOI22_X1 U20772 ( .A1(n17565), .A2(n17564), .B1(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17563), .ZN(n17566) );
  NAND2_X1 U20773 ( .A1(n18035), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17908) );
  OAI211_X1 U20774 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17567), .A(
        n17566), .B(n17908), .ZN(n17568) );
  AOI21_X1 U20775 ( .B1(n17618), .B2(n17907), .A(n17568), .ZN(n17569) );
  OAI221_X1 U20776 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17571), 
        .C1(n17903), .C2(n17570), .A(n17569), .ZN(P3_U2818) );
  AOI22_X1 U20777 ( .A1(n18035), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17572), 
        .B2(n17376), .ZN(n17580) );
  INV_X1 U20778 ( .A(n17596), .ZN(n17583) );
  OAI21_X1 U20779 ( .B1(n17922), .B2(n17583), .A(n17573), .ZN(n17575) );
  XNOR2_X1 U20780 ( .A(n17575), .B(n17574), .ZN(n17926) );
  NOR2_X1 U20781 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17922), .ZN(
        n17925) );
  AOI22_X1 U20782 ( .A1(n17618), .A2(n17926), .B1(n17925), .B2(n17603), .ZN(
        n17579) );
  AND2_X1 U20783 ( .A1(n17922), .A2(n17603), .ZN(n17592) );
  OAI22_X1 U20784 ( .A1(n17916), .A2(n17621), .B1(n17713), .B2(n17913), .ZN(
        n17604) );
  OAI21_X1 U20785 ( .B1(n17592), .B2(n17604), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17578) );
  NAND3_X1 U20786 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(n17612), .ZN(n17598) );
  NOR2_X1 U20787 ( .A1(n17587), .A2(n17598), .ZN(n17586) );
  OAI211_X1 U20788 ( .C1(n17586), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17634), .B(n17576), .ZN(n17577) );
  NAND4_X1 U20789 ( .A1(n17580), .A2(n17579), .A3(n17578), .A4(n17577), .ZN(
        P3_U2819) );
  INV_X1 U20790 ( .A(n17581), .ZN(n17591) );
  INV_X1 U20791 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17582) );
  OAI221_X1 U20792 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17583), 
        .C1(n17582), .C2(n17596), .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17585) );
  INV_X1 U20793 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17931) );
  NAND4_X1 U20794 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15647), .A3(
        n17931), .A4(n17519), .ZN(n17584) );
  OAI211_X1 U20795 ( .C1(n17595), .C2(n17591), .A(n17585), .B(n17584), .ZN(
        n17936) );
  INV_X1 U20796 ( .A(n17634), .ZN(n17704) );
  AOI211_X1 U20797 ( .C1(n17598), .C2(n17587), .A(n17704), .B(n17586), .ZN(
        n17589) );
  NAND2_X1 U20798 ( .A1(n18035), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n17934) );
  INV_X1 U20799 ( .A(n17934), .ZN(n17588) );
  AOI211_X1 U20800 ( .C1(n17590), .C2(n17376), .A(n17589), .B(n17588), .ZN(
        n17594) );
  AOI22_X1 U20801 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17604), .B1(
        n17592), .B2(n17591), .ZN(n17593) );
  OAI211_X1 U20802 ( .C1(n17606), .C2(n17936), .A(n17594), .B(n17593), .ZN(
        P3_U2820) );
  NOR2_X1 U20803 ( .A1(n17596), .A2(n17595), .ZN(n17597) );
  XNOR2_X1 U20804 ( .A(n17597), .B(n17931), .ZN(n17943) );
  AND2_X1 U20805 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17612), .ZN(
        n17599) );
  OAI211_X1 U20806 ( .C1(n17599), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17634), .B(n17598), .ZN(n17600) );
  NAND2_X1 U20807 ( .A1(n18035), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17940) );
  OAI211_X1 U20808 ( .C1(n17693), .C2(n17601), .A(n17600), .B(n17940), .ZN(
        n17602) );
  AOI221_X1 U20809 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17604), .C1(
        n17931), .C2(n17603), .A(n17602), .ZN(n17605) );
  OAI21_X1 U20810 ( .B1(n17943), .B2(n17606), .A(n17605), .ZN(P3_U2821) );
  AOI21_X1 U20811 ( .B1(n17667), .B2(n17607), .A(n17682), .ZN(n17633) );
  OAI21_X1 U20812 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18132), .A(
        n17633), .ZN(n17610) );
  OAI22_X1 U20813 ( .A1(n17693), .A2(n17608), .B1(n9800), .B2(n18601), .ZN(
        n17609) );
  AOI221_X1 U20814 ( .B1(n17612), .B2(n17611), .C1(n17610), .C2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(n17609), .ZN(n17620) );
  AOI21_X1 U20815 ( .B1(n17614), .B2(n17948), .A(n17613), .ZN(n17953) );
  OAI21_X1 U20816 ( .B1(n17617), .B2(n17616), .A(n17615), .ZN(n17954) );
  AOI22_X1 U20817 ( .A1(n9792), .A2(n17953), .B1(n17618), .B2(n17954), .ZN(
        n17619) );
  OAI211_X1 U20818 ( .C1(n17959), .C2(n17621), .A(n17620), .B(n17619), .ZN(
        P3_U2822) );
  NOR2_X1 U20819 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18132), .ZN(
        n17622) );
  AOI22_X1 U20820 ( .A1(n18035), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n17623), 
        .B2(n17622), .ZN(n17632) );
  AOI21_X1 U20821 ( .B1(n17625), .B2(n17962), .A(n17624), .ZN(n17965) );
  NAND2_X1 U20822 ( .A1(n17627), .A2(n17626), .ZN(n17628) );
  XNOR2_X1 U20823 ( .A(n17628), .B(n17962), .ZN(n17968) );
  OAI22_X1 U20824 ( .A1(n17693), .A2(n17629), .B1(n17713), .B2(n17968), .ZN(
        n17630) );
  AOI21_X1 U20825 ( .B1(n17701), .B2(n17965), .A(n17630), .ZN(n17631) );
  OAI211_X1 U20826 ( .C1(n17633), .C2(n10100), .A(n17632), .B(n17631), .ZN(
        P3_U2823) );
  OAI21_X1 U20827 ( .B1(n17637), .B2(n18132), .A(n17634), .ZN(n17657) );
  AOI21_X1 U20828 ( .B1(n17636), .B2(n17635), .A(n9903), .ZN(n17972) );
  NOR2_X1 U20829 ( .A1(n9800), .A2(n18596), .ZN(n17971) );
  NOR3_X1 U20830 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17637), .A3(
        n18132), .ZN(n17638) );
  AOI211_X1 U20831 ( .C1(n17701), .C2(n17972), .A(n17971), .B(n17638), .ZN(
        n17644) );
  AOI21_X1 U20832 ( .B1(n17641), .B2(n17640), .A(n17639), .ZN(n17976) );
  AOI22_X1 U20833 ( .A1(n17698), .A2(n17976), .B1(n17642), .B2(n17376), .ZN(
        n17643) );
  OAI211_X1 U20834 ( .C1(n17645), .C2(n17657), .A(n17644), .B(n17643), .ZN(
        P3_U2824) );
  AOI21_X1 U20835 ( .B1(n17646), .B2(n17708), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17658) );
  OAI21_X1 U20836 ( .B1(n17649), .B2(n17648), .A(n17647), .ZN(n17650) );
  XNOR2_X1 U20837 ( .A(n17650), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17980) );
  AOI22_X1 U20838 ( .A1(n18035), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17701), 
        .B2(n17980), .ZN(n17656) );
  AOI21_X1 U20839 ( .B1(n17653), .B2(n17652), .A(n17651), .ZN(n17979) );
  AOI22_X1 U20840 ( .A1(n9792), .A2(n17979), .B1(n17654), .B2(n17376), .ZN(
        n17655) );
  OAI211_X1 U20841 ( .C1(n17658), .C2(n17657), .A(n17656), .B(n17655), .ZN(
        P3_U2825) );
  OAI21_X1 U20842 ( .B1(n17661), .B2(n17660), .A(n17659), .ZN(n17662) );
  INV_X1 U20843 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17993) );
  XNOR2_X1 U20844 ( .A(n17662), .B(n17993), .ZN(n17988) );
  AOI22_X1 U20845 ( .A1(n18035), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18442), 
        .B2(n17663), .ZN(n17672) );
  AOI21_X1 U20846 ( .B1(n9911), .B2(n17665), .A(n17664), .ZN(n17990) );
  AOI21_X1 U20847 ( .B1(n17667), .B2(n17666), .A(n17682), .ZN(n17676) );
  OAI22_X1 U20848 ( .A1(n17693), .A2(n17669), .B1(n17676), .B2(n17668), .ZN(
        n17670) );
  AOI21_X1 U20849 ( .B1(n17701), .B2(n17990), .A(n17670), .ZN(n17671) );
  OAI211_X1 U20850 ( .C1(n17713), .C2(n17988), .A(n17672), .B(n17671), .ZN(
        P3_U2826) );
  AOI21_X1 U20851 ( .B1(n17675), .B2(n17674), .A(n17673), .ZN(n17997) );
  INV_X1 U20852 ( .A(n17676), .ZN(n17677) );
  AOI22_X1 U20853 ( .A1(n17701), .A2(n17997), .B1(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17677), .ZN(n17685) );
  AOI21_X1 U20854 ( .B1(n17680), .B2(n17679), .A(n17678), .ZN(n17996) );
  NOR2_X1 U20855 ( .A1(n9800), .A2(n18591), .ZN(n17995) );
  NOR4_X1 U20856 ( .A1(n17682), .A2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17681), .A4(n17696), .ZN(n17683) );
  AOI211_X1 U20857 ( .C1(n9792), .C2(n17996), .A(n17995), .B(n17683), .ZN(
        n17684) );
  OAI211_X1 U20858 ( .C1(n17693), .C2(n17686), .A(n17685), .B(n17684), .ZN(
        P3_U2827) );
  AOI21_X1 U20859 ( .B1(n17689), .B2(n17688), .A(n17687), .ZN(n18011) );
  NOR2_X1 U20860 ( .A1(n9800), .A2(n20808), .ZN(n18015) );
  XNOR2_X1 U20861 ( .A(n17691), .B(n17690), .ZN(n18017) );
  OAI22_X1 U20862 ( .A1(n17693), .A2(n17692), .B1(n17712), .B2(n18017), .ZN(
        n17694) );
  AOI211_X1 U20863 ( .C1(n17698), .C2(n18011), .A(n18015), .B(n17694), .ZN(
        n17695) );
  OAI221_X1 U20864 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18132), .C1(
        n17696), .C2(n17708), .A(n17695), .ZN(P3_U2828) );
  NOR2_X1 U20865 ( .A1(n17706), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17697) );
  XNOR2_X1 U20866 ( .A(n17697), .B(n17700), .ZN(n18018) );
  AOI22_X1 U20867 ( .A1(n18035), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17698), 
        .B2(n18018), .ZN(n17703) );
  AOI21_X1 U20868 ( .B1(n17705), .B2(n17700), .A(n17699), .ZN(n18020) );
  AOI22_X1 U20869 ( .A1(n17701), .A2(n18020), .B1(n21011), .B2(n17376), .ZN(
        n17702) );
  OAI211_X1 U20870 ( .C1(n17704), .C2(n21011), .A(n17703), .B(n17702), .ZN(
        P3_U2829) );
  OAI21_X1 U20871 ( .B1(n17706), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17705), .ZN(n18038) );
  INV_X1 U20872 ( .A(n18038), .ZN(n18040) );
  NAND3_X1 U20873 ( .A1(n17709), .A2(n17708), .A3(n17707), .ZN(n17710) );
  AOI22_X1 U20874 ( .A1(n18035), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17710), .ZN(n17711) );
  OAI221_X1 U20875 ( .B1(n18040), .B2(n17713), .C1(n18038), .C2(n17712), .A(
        n17711), .ZN(P3_U2830) );
  NAND2_X1 U20876 ( .A1(n9800), .A2(n18022), .ZN(n17973) );
  INV_X1 U20877 ( .A(n17773), .ZN(n17714) );
  NOR2_X1 U20878 ( .A1(n17715), .A2(n17714), .ZN(n17725) );
  AOI21_X1 U20879 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18516), .A(
        n17716), .ZN(n17782) );
  NOR2_X1 U20880 ( .A1(n17779), .A2(n17782), .ZN(n17717) );
  INV_X1 U20881 ( .A(n18003), .ZN(n17831) );
  AOI21_X1 U20882 ( .B1(n17717), .B2(n17844), .A(n17831), .ZN(n17761) );
  AOI21_X1 U20883 ( .B1(n17746), .B2(n18003), .A(n17761), .ZN(n17747) );
  AOI21_X1 U20884 ( .B1(n17719), .B2(n18003), .A(n17718), .ZN(n17720) );
  OAI211_X1 U20885 ( .C1(n17721), .C2(n17914), .A(n17747), .B(n17720), .ZN(
        n17722) );
  AOI21_X1 U20886 ( .B1(n17894), .B2(n17723), .A(n17722), .ZN(n17736) );
  INV_X1 U20887 ( .A(n17736), .ZN(n17724) );
  MUX2_X1 U20888 ( .A(n17725), .B(n17724), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17727) );
  AOI22_X1 U20889 ( .A1(n18032), .A2(n17727), .B1(n17955), .B2(n17726), .ZN(
        n17729) );
  OAI211_X1 U20890 ( .C1(n17730), .C2(n17973), .A(n17729), .B(n17728), .ZN(
        P3_U2835) );
  INV_X1 U20891 ( .A(n17731), .ZN(n17734) );
  INV_X1 U20892 ( .A(n17732), .ZN(n17733) );
  INV_X1 U20893 ( .A(n17801), .ZN(n17784) );
  NAND3_X1 U20894 ( .A1(n17733), .A2(n17785), .A3(n17784), .ZN(n17767) );
  OAI22_X1 U20895 ( .A1(n17736), .A2(n17735), .B1(n17734), .B2(n17767), .ZN(
        n17737) );
  AOI22_X1 U20896 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18024), .B1(
        n18032), .B2(n17737), .ZN(n17739) );
  NAND2_X1 U20897 ( .A1(n18035), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17738) );
  OAI211_X1 U20898 ( .C1(n17740), .C2(n17942), .A(n17739), .B(n17738), .ZN(
        P3_U2836) );
  INV_X1 U20899 ( .A(n17888), .ZN(n17958) );
  OAI22_X1 U20900 ( .A1(n17942), .A2(n17742), .B1(n17958), .B2(n17741), .ZN(
        n17755) );
  NAND2_X1 U20901 ( .A1(n17744), .A2(n17743), .ZN(n17745) );
  NOR2_X1 U20902 ( .A1(n17746), .A2(n17745), .ZN(n17750) );
  INV_X1 U20903 ( .A(n17746), .ZN(n17748) );
  OAI221_X1 U20904 ( .B1(n18524), .B2(n17763), .C1(n18524), .C2(n17748), .A(
        n17747), .ZN(n17749) );
  OAI221_X1 U20905 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17750), 
        .C1(n17753), .C2(n17749), .A(n18032), .ZN(n17751) );
  OAI211_X1 U20906 ( .C1(n17973), .C2(n17753), .A(n17752), .B(n17751), .ZN(
        n17754) );
  NOR2_X1 U20907 ( .A1(n17755), .A2(n17754), .ZN(n17756) );
  OAI21_X1 U20908 ( .B1(n17757), .B2(n18039), .A(n17756), .ZN(P3_U2837) );
  INV_X1 U20909 ( .A(n17758), .ZN(n17759) );
  OAI21_X1 U20910 ( .B1(n17759), .B2(n17914), .A(n17973), .ZN(n17760) );
  AOI211_X1 U20911 ( .C1(n17894), .C2(n17762), .A(n17761), .B(n17760), .ZN(
        n17766) );
  OAI211_X1 U20912 ( .C1(n17763), .C2(n18524), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17766), .ZN(n17764) );
  NAND2_X1 U20913 ( .A1(n9800), .A2(n17764), .ZN(n17776) );
  AOI211_X1 U20914 ( .C1(n17850), .C2(n17766), .A(n17765), .B(n17776), .ZN(
        n17769) );
  NOR3_X1 U20915 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18022), .A3(
        n17767), .ZN(n17768) );
  NOR3_X1 U20916 ( .A1(n17770), .A2(n17769), .A3(n17768), .ZN(n17771) );
  OAI21_X1 U20917 ( .B1(n17772), .B2(n17942), .A(n17771), .ZN(P3_U2838) );
  AOI21_X1 U20918 ( .B1(n17773), .B2(n17973), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17777) );
  AOI22_X1 U20919 ( .A1(n18035), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17955), 
        .B2(n17774), .ZN(n17775) );
  OAI21_X1 U20920 ( .B1(n17777), .B2(n17776), .A(n17775), .ZN(P3_U2839) );
  AOI21_X1 U20921 ( .B1(n17844), .B2(n17809), .A(n18531), .ZN(n17778) );
  AOI221_X1 U20922 ( .B1(n17830), .B2(n18506), .C1(n17829), .C2(n18506), .A(
        n17778), .ZN(n17796) );
  NAND2_X1 U20923 ( .A1(n17915), .A2(n17914), .ZN(n17921) );
  AOI22_X1 U20924 ( .A1(n17876), .A2(n17780), .B1(n17779), .B2(n17921), .ZN(
        n17798) );
  OAI211_X1 U20925 ( .C1(n17799), .C2(n18524), .A(n17796), .B(n17798), .ZN(
        n17781) );
  AOI211_X1 U20926 ( .C1(n17847), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        n17788) );
  OAI22_X1 U20927 ( .A1(n17856), .A2(n17915), .B1(n17867), .B2(n17914), .ZN(
        n17795) );
  INV_X1 U20928 ( .A(n17795), .ZN(n17787) );
  NAND2_X1 U20929 ( .A1(n17785), .A2(n17784), .ZN(n17786) );
  AOI22_X1 U20930 ( .A1(n17788), .A2(n17787), .B1(n17793), .B2(n17786), .ZN(
        n17790) );
  AOI22_X1 U20931 ( .A1(n18032), .A2(n17790), .B1(n17955), .B2(n17789), .ZN(
        n17792) );
  NAND2_X1 U20932 ( .A1(n18035), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17791) );
  OAI211_X1 U20933 ( .C1(n17973), .C2(n17793), .A(n17792), .B(n17791), .ZN(
        P3_U2840) );
  INV_X1 U20934 ( .A(n17844), .ZN(n17824) );
  NOR3_X1 U20935 ( .A1(n18031), .A2(n17824), .A3(n17794), .ZN(n17797) );
  NOR2_X1 U20936 ( .A1(n18022), .A2(n17795), .ZN(n17849) );
  OAI211_X1 U20937 ( .C1(n18516), .C2(n17797), .A(n17849), .B(n17796), .ZN(
        n17807) );
  NOR2_X1 U20938 ( .A1(n18506), .A2(n18529), .ZN(n18023) );
  OAI21_X1 U20939 ( .B1(n17799), .B2(n18023), .A(n17798), .ZN(n17800) );
  OAI21_X1 U20940 ( .B1(n17807), .B2(n17800), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17805) );
  NOR3_X1 U20941 ( .A1(n17801), .A2(n18022), .A3(n17830), .ZN(n17815) );
  AOI22_X1 U20942 ( .A1(n17955), .A2(n17803), .B1(n17802), .B2(n17815), .ZN(
        n17804) );
  OAI221_X1 U20943 ( .B1(n18035), .B2(n17805), .C1(n9800), .C2(n18626), .A(
        n17804), .ZN(P3_U2841) );
  AOI22_X1 U20944 ( .A1(n18035), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17815), 
        .B2(n17806), .ZN(n17812) );
  INV_X1 U20945 ( .A(n17807), .ZN(n17808) );
  INV_X1 U20946 ( .A(n17921), .ZN(n17826) );
  AOI221_X1 U20947 ( .B1(n17809), .B2(n17808), .C1(n17826), .C2(n17808), .A(
        n18035), .ZN(n17816) );
  NOR3_X1 U20948 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18023), .A3(
        n18720), .ZN(n17810) );
  OAI21_X1 U20949 ( .B1(n17816), .B2(n17810), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17811) );
  OAI211_X1 U20950 ( .C1(n17813), .C2(n17942), .A(n17812), .B(n17811), .ZN(
        P3_U2842) );
  AOI22_X1 U20951 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17816), .B1(
        n17815), .B2(n17814), .ZN(n17818) );
  NAND2_X1 U20952 ( .A1(n18035), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17817) );
  OAI211_X1 U20953 ( .C1(n17819), .C2(n17942), .A(n17818), .B(n17817), .ZN(
        P3_U2843) );
  INV_X1 U20954 ( .A(n17820), .ZN(n17822) );
  OAI22_X1 U20955 ( .A1(n17945), .A2(n18524), .B1(n17944), .B2(n18008), .ZN(
        n17999) );
  INV_X1 U20956 ( .A(n17999), .ZN(n17963) );
  OR2_X1 U20957 ( .A1(n17821), .A2(n17963), .ZN(n17859) );
  NAND2_X1 U20958 ( .A1(n17823), .A2(n17939), .ZN(n17855) );
  NOR2_X1 U20959 ( .A1(n18516), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18004) );
  OAI21_X1 U20960 ( .B1(n17824), .B2(n17848), .A(n18003), .ZN(n17825) );
  OAI211_X1 U20961 ( .C1(n17827), .C2(n17826), .A(n17849), .B(n17825), .ZN(
        n17828) );
  AOI211_X1 U20962 ( .C1(n18506), .C2(n17829), .A(n18004), .B(n17828), .ZN(
        n17838) );
  AOI221_X1 U20963 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17838), 
        .C1(n17831), .C2(n17838), .A(n17830), .ZN(n17832) );
  AOI22_X1 U20964 ( .A1(n17833), .A2(n17955), .B1(n17832), .B2(n9800), .ZN(
        n17835) );
  NAND2_X1 U20965 ( .A1(n18035), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17834) );
  OAI211_X1 U20966 ( .C1(n17836), .C2(n17855), .A(n17835), .B(n17834), .ZN(
        P3_U2844) );
  NOR3_X1 U20967 ( .A1(n18035), .A2(n17838), .A3(n17837), .ZN(n17839) );
  AOI21_X1 U20968 ( .B1(n17955), .B2(n17840), .A(n17839), .ZN(n17842) );
  NAND2_X1 U20969 ( .A1(n15711), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17841) );
  OAI211_X1 U20970 ( .C1(n17843), .C2(n17855), .A(n17842), .B(n17841), .ZN(
        P3_U2845) );
  AOI22_X1 U20971 ( .A1(n18516), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17844), .ZN(n17845) );
  OAI22_X1 U20972 ( .A1(n18531), .A2(n17912), .B1(n17874), .B2(n18524), .ZN(
        n17918) );
  AOI211_X1 U20973 ( .C1(n17847), .C2(n17846), .A(n17845), .B(n17918), .ZN(
        n17861) );
  AOI221_X1 U20974 ( .B1(n17850), .B2(n17849), .C1(n17861), .C2(n17849), .A(
        n17848), .ZN(n17851) );
  AOI22_X1 U20975 ( .A1(n17852), .A2(n17955), .B1(n17851), .B2(n9800), .ZN(
        n17854) );
  OAI211_X1 U20976 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17855), .A(
        n17854), .B(n17853), .ZN(P3_U2846) );
  NOR2_X1 U20977 ( .A1(n17856), .A2(n17915), .ZN(n17865) );
  INV_X1 U20978 ( .A(n17857), .ZN(n17864) );
  OR2_X1 U20979 ( .A1(n17859), .A2(n17858), .ZN(n17883) );
  AOI211_X1 U20980 ( .C1(n17862), .C2(n17883), .A(n17861), .B(n17860), .ZN(
        n17863) );
  AOI21_X1 U20981 ( .B1(n17865), .B2(n17864), .A(n17863), .ZN(n17873) );
  AOI21_X1 U20982 ( .B1(n18024), .B2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n17866), .ZN(n17872) );
  NOR2_X1 U20983 ( .A1(n17867), .A2(n18039), .ZN(n17869) );
  AOI22_X1 U20984 ( .A1(n17955), .A2(n17870), .B1(n17869), .B2(n17868), .ZN(
        n17871) );
  OAI211_X1 U20985 ( .C1(n17873), .C2(n18022), .A(n17872), .B(n17871), .ZN(
        P3_U2847) );
  NOR2_X1 U20986 ( .A1(n17874), .A2(n18524), .ZN(n17880) );
  OAI21_X1 U20987 ( .B1(n17884), .B2(n17876), .A(n17875), .ZN(n17878) );
  NAND3_X1 U20988 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17912), .A3(
        n17877), .ZN(n17905) );
  NAND2_X1 U20989 ( .A1(n18529), .A2(n17905), .ZN(n17897) );
  OAI211_X1 U20990 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18023), .A(
        n17878), .B(n17897), .ZN(n17879) );
  AOI211_X1 U20991 ( .C1(n18506), .C2(n17881), .A(n17880), .B(n17879), .ZN(
        n17882) );
  AOI211_X1 U20992 ( .C1(n17884), .C2(n17883), .A(n17882), .B(n18022), .ZN(
        n17885) );
  AOI211_X1 U20993 ( .C1(n18024), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17886), .B(n17885), .ZN(n17891) );
  AOI22_X1 U20994 ( .A1(n17955), .A2(n17889), .B1(n17888), .B2(n17887), .ZN(
        n17890) );
  OAI211_X1 U20995 ( .C1(n18039), .C2(n17892), .A(n17891), .B(n17890), .ZN(
        P3_U2848) );
  NOR2_X1 U20996 ( .A1(n17930), .A2(n17906), .ZN(n17924) );
  AOI211_X1 U20997 ( .C1(n17894), .C2(n17893), .A(n17924), .B(n17918), .ZN(
        n17895) );
  OAI21_X1 U20998 ( .B1(n17896), .B2(n17914), .A(n17895), .ZN(n17904) );
  OAI211_X1 U20999 ( .C1(n17930), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18032), .B(n17897), .ZN(n17898) );
  OAI21_X1 U21000 ( .B1(n17904), .B2(n17898), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17902) );
  AOI22_X1 U21001 ( .A1(n17955), .A2(n17900), .B1(n17939), .B2(n17899), .ZN(
        n17901) );
  OAI221_X1 U21002 ( .B1(n18035), .B2(n17902), .C1(n9800), .C2(n18609), .A(
        n17901), .ZN(P3_U2849) );
  AOI211_X1 U21003 ( .C1(n17905), .C2(n18529), .A(n17904), .B(n17903), .ZN(
        n17911) );
  AOI22_X1 U21004 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18032), .B1(
        n17906), .B2(n17939), .ZN(n17910) );
  AOI22_X1 U21005 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18024), .B1(
        n17955), .B2(n17907), .ZN(n17909) );
  OAI211_X1 U21006 ( .C1(n17911), .C2(n17910), .A(n17909), .B(n17908), .ZN(
        P3_U2850) );
  AOI21_X1 U21007 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n17912), .A(
        n18516), .ZN(n17919) );
  OAI22_X1 U21008 ( .A1(n17916), .A2(n17915), .B1(n17914), .B2(n17913), .ZN(
        n17917) );
  NOR4_X1 U21009 ( .A1(n17919), .A2(n17918), .A3(n18022), .A4(n17917), .ZN(
        n17937) );
  OAI21_X1 U21010 ( .B1(n18516), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17937), .ZN(n17920) );
  AOI21_X1 U21011 ( .B1(n17922), .B2(n17921), .A(n17920), .ZN(n17929) );
  OAI21_X1 U21012 ( .B1(n18516), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17929), .ZN(n17923) );
  OAI21_X1 U21013 ( .B1(n17924), .B2(n17923), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17928) );
  AOI22_X1 U21014 ( .A1(n17955), .A2(n17926), .B1(n17939), .B2(n17925), .ZN(
        n17927) );
  OAI221_X1 U21015 ( .B1(n15711), .B2(n17928), .C1(n9800), .C2(n18606), .A(
        n17927), .ZN(P3_U2851) );
  AOI221_X1 U21016 ( .B1(n17930), .B2(n17929), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17929), .A(n18035), .ZN(
        n17933) );
  NOR2_X1 U21017 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17931), .ZN(
        n17932) );
  AOI22_X1 U21018 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17933), .B1(
        n17939), .B2(n17932), .ZN(n17935) );
  OAI211_X1 U21019 ( .C1(n17936), .C2(n17942), .A(n17935), .B(n17934), .ZN(
        P3_U2852) );
  OAI21_X1 U21020 ( .B1(n18035), .B2(n17937), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17938) );
  OAI21_X1 U21021 ( .B1(n17939), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17938), .ZN(n17941) );
  OAI211_X1 U21022 ( .C1(n17943), .C2(n17942), .A(n17941), .B(n17940), .ZN(
        P3_U2853) );
  NAND2_X1 U21023 ( .A1(n18032), .A2(n17999), .ZN(n17982) );
  NOR2_X1 U21024 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17982), .ZN(
        n17951) );
  AOI211_X1 U21025 ( .C1(n17944), .C2(n18003), .A(n18004), .B(n17983), .ZN(
        n17946) );
  NAND2_X1 U21026 ( .A1(n18506), .A2(n17945), .ZN(n18012) );
  NAND2_X1 U21027 ( .A1(n17946), .A2(n18012), .ZN(n17998) );
  NOR3_X1 U21028 ( .A1(n17993), .A2(n10142), .A3(n17998), .ZN(n17975) );
  NAND3_X1 U21029 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n17975), .ZN(n17947) );
  NAND2_X1 U21030 ( .A1(n18026), .A2(n17947), .ZN(n17960) );
  AOI21_X1 U21031 ( .B1(n17973), .B2(n17960), .A(n17948), .ZN(n17950) );
  NOR2_X1 U21032 ( .A1(n9800), .A2(n18601), .ZN(n17949) );
  AOI211_X1 U21033 ( .C1(n17952), .C2(n17951), .A(n17950), .B(n17949), .ZN(
        n17957) );
  AOI22_X1 U21034 ( .A1(n17955), .A2(n17954), .B1(n18019), .B2(n17953), .ZN(
        n17956) );
  OAI211_X1 U21035 ( .C1(n17959), .C2(n17958), .A(n17957), .B(n17956), .ZN(
        P3_U2854) );
  AOI22_X1 U21036 ( .A1(n18035), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18024), .ZN(n17967) );
  INV_X1 U21037 ( .A(n18037), .ZN(n18021) );
  AOI221_X1 U21038 ( .B1(n17963), .B2(n17962), .C1(n17961), .C2(n17962), .A(
        n17960), .ZN(n17964) );
  AOI21_X1 U21039 ( .B1(n17965), .B2(n18021), .A(n17964), .ZN(n17966) );
  OAI211_X1 U21040 ( .C1(n18039), .C2(n17968), .A(n17967), .B(n17966), .ZN(
        P3_U2855) );
  NAND3_X1 U21041 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17969) );
  NOR3_X1 U21042 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17969), .A3(
        n17982), .ZN(n17970) );
  AOI211_X1 U21043 ( .C1(n18021), .C2(n17972), .A(n17971), .B(n17970), .ZN(
        n17978) );
  OAI21_X1 U21044 ( .B1(n17975), .B2(n17974), .A(n17973), .ZN(n17981) );
  AOI22_X1 U21045 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17981), .B1(
        n18019), .B2(n17976), .ZN(n17977) );
  NAND2_X1 U21046 ( .A1(n17978), .A2(n17977), .ZN(P3_U2856) );
  AOI22_X1 U21047 ( .A1(n15711), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18019), 
        .B2(n17979), .ZN(n17986) );
  AOI22_X1 U21048 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17981), .B1(
        n18021), .B2(n17980), .ZN(n17985) );
  NOR2_X1 U21049 ( .A1(n17983), .A2(n17982), .ZN(n17987) );
  NAND3_X1 U21050 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17987), .A3(
        n10142), .ZN(n17984) );
  NAND3_X1 U21051 ( .A1(n17986), .A2(n17985), .A3(n17984), .ZN(P3_U2857) );
  INV_X1 U21052 ( .A(n17987), .ZN(n17994) );
  AOI21_X1 U21053 ( .B1(n18026), .B2(n17998), .A(n18024), .ZN(n17992) );
  OAI22_X1 U21054 ( .A1(n9800), .A2(n18592), .B1(n18039), .B2(n17988), .ZN(
        n17989) );
  AOI21_X1 U21055 ( .B1(n18021), .B2(n17990), .A(n17989), .ZN(n17991) );
  OAI221_X1 U21056 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n17994), .C1(
        n17993), .C2(n17992), .A(n17991), .ZN(P3_U2858) );
  AOI21_X1 U21057 ( .B1(n18024), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n17995), .ZN(n18002) );
  AOI22_X1 U21058 ( .A1(n18021), .A2(n17997), .B1(n18019), .B2(n17996), .ZN(
        n18001) );
  OAI211_X1 U21059 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n17999), .A(
        n18032), .B(n17998), .ZN(n18000) );
  NAND3_X1 U21060 ( .A1(n18002), .A2(n18001), .A3(n18000), .ZN(P3_U2859) );
  OAI21_X1 U21061 ( .B1(n18004), .B2(n18668), .A(n18003), .ZN(n18007) );
  NAND2_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18006) );
  AOI221_X1 U21063 ( .B1(n18524), .B2(n18007), .C1(n18006), .C2(n18007), .A(
        n18005), .ZN(n18010) );
  NOR3_X1 U21064 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18668), .A3(
        n18008), .ZN(n18009) );
  AOI211_X1 U21065 ( .C1(n18011), .C2(n18494), .A(n18010), .B(n18009), .ZN(
        n18013) );
  AOI21_X1 U21066 ( .B1(n18013), .B2(n18012), .A(n18022), .ZN(n18014) );
  AOI211_X1 U21067 ( .C1(n18024), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18015), .B(n18014), .ZN(n18016) );
  OAI21_X1 U21068 ( .B1(n18037), .B2(n18017), .A(n18016), .ZN(P3_U2860) );
  AOI22_X1 U21069 ( .A1(n18021), .A2(n18020), .B1(n18019), .B2(n18018), .ZN(
        n18030) );
  NAND2_X1 U21070 ( .A1(n18035), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18029) );
  NOR3_X1 U21071 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18023), .A3(
        n18022), .ZN(n18033) );
  OAI21_X1 U21072 ( .B1(n18024), .B2(n18033), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18028) );
  NAND3_X1 U21073 ( .A1(n18026), .A2(n18668), .A3(n18025), .ZN(n18027) );
  NAND4_X1 U21074 ( .A1(n18030), .A2(n18029), .A3(n18028), .A4(n18027), .ZN(
        P3_U2861) );
  AOI21_X1 U21075 ( .B1(n18531), .B2(n18032), .A(n18031), .ZN(n18034) );
  AOI221_X1 U21076 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n18035), .C1(n18034), 
        .C2(n9800), .A(n18033), .ZN(n18036) );
  OAI221_X1 U21077 ( .B1(n18040), .B2(n18039), .C1(n18038), .C2(n18037), .A(
        n18036), .ZN(P3_U2862) );
  OAI211_X1 U21078 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18041), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18558)
         );
  INV_X1 U21079 ( .A(n18705), .ZN(n18042) );
  OAI21_X1 U21080 ( .B1(n18044), .B2(n18042), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18043) );
  OAI221_X1 U21081 ( .B1(n18044), .B2(n18558), .C1(n18044), .C2(n18104), .A(
        n18043), .ZN(P3_U2863) );
  NAND2_X1 U21082 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18047) );
  AOI221_X1 U21083 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18047), .C1(n18046), 
        .C2(n18047), .A(n18045), .ZN(n18052) );
  NOR2_X1 U21084 ( .A1(n18048), .A2(n18536), .ZN(n18049) );
  OAI21_X1 U21085 ( .B1(n18049), .B2(n18315), .A(n18053), .ZN(n18050) );
  AOI22_X1 U21086 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18052), .B1(
        n18050), .B2(n21014), .ZN(P3_U2865) );
  NOR2_X1 U21087 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21014), .ZN(
        n18243) );
  INV_X1 U21088 ( .A(n18243), .ZN(n18291) );
  NOR2_X1 U21089 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18543), .ZN(
        n18338) );
  NAND2_X1 U21090 ( .A1(n18315), .A2(n18338), .ZN(n18361) );
  AND2_X1 U21091 ( .A1(n18291), .A2(n18361), .ZN(n18051) );
  OAI22_X1 U21092 ( .A1(n18052), .A2(n18543), .B1(n18051), .B2(n18050), .ZN(
        P3_U2866) );
  NOR2_X1 U21093 ( .A1(n20939), .A2(n18053), .ZN(P3_U2867) );
  NAND2_X1 U21094 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18535) );
  NAND2_X1 U21095 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18103) );
  NOR2_X2 U21096 ( .A1(n18535), .A2(n18103), .ZN(n18436) );
  NAND2_X1 U21097 ( .A1(n18536), .A2(n18360), .ZN(n18537) );
  NAND2_X1 U21098 ( .A1(n21014), .A2(n18543), .ZN(n18201) );
  NOR2_X1 U21099 ( .A1(n18537), .A2(n18201), .ZN(n18150) );
  CLKBUF_X1 U21100 ( .A(n18150), .Z(n18173) );
  NOR2_X1 U21101 ( .A1(n18436), .A2(n18173), .ZN(n18133) );
  OAI21_X1 U21102 ( .B1(n18684), .B2(n18360), .A(n18364), .ZN(n18222) );
  NOR2_X1 U21103 ( .A1(n18536), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18314) );
  NOR2_X1 U21104 ( .A1(n18360), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18289) );
  NOR2_X1 U21105 ( .A1(n18314), .A2(n18289), .ZN(n18362) );
  OR2_X1 U21106 ( .A1(n18103), .A2(n18362), .ZN(n18411) );
  OAI22_X1 U21107 ( .A1(n18133), .A2(n18222), .B1(n18132), .B2(n18411), .ZN(
        n18101) );
  AND2_X1 U21108 ( .A1(n18442), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18438) );
  INV_X1 U21109 ( .A(n18103), .ZN(n18388) );
  NAND2_X1 U21110 ( .A1(n18388), .A2(n18314), .ZN(n18435) );
  INV_X1 U21111 ( .A(n18435), .ZN(n18127) );
  NOR2_X2 U21112 ( .A1(n18131), .A2(n18054), .ZN(n18437) );
  INV_X1 U21113 ( .A(n18560), .ZN(n18410) );
  NOR2_X1 U21114 ( .A1(n18410), .A2(n18133), .ZN(n18095) );
  AOI22_X1 U21115 ( .A1(n18438), .A2(n18127), .B1(n18437), .B2(n18095), .ZN(
        n18060) );
  NAND2_X1 U21116 ( .A1(n18056), .A2(n18055), .ZN(n18096) );
  NOR2_X1 U21117 ( .A1(n18057), .A2(n18096), .ZN(n18102) );
  NAND2_X1 U21118 ( .A1(n18388), .A2(n18536), .ZN(n18385) );
  NOR2_X2 U21119 ( .A1(n18360), .A2(n18385), .ZN(n18488) );
  NOR2_X2 U21120 ( .A1(n18058), .A2(n18132), .ZN(n18443) );
  AOI22_X1 U21121 ( .A1(n18173), .A2(n18102), .B1(n18488), .B2(n18443), .ZN(
        n18059) );
  OAI211_X1 U21122 ( .C1(n18061), .C2(n18101), .A(n18060), .B(n18059), .ZN(
        P3_U2868) );
  NOR2_X2 U21123 ( .A1(n14764), .A2(n18132), .ZN(n18448) );
  AND2_X1 U21124 ( .A1(n18364), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18447) );
  AOI22_X1 U21125 ( .A1(n18488), .A2(n18448), .B1(n18095), .B2(n18447), .ZN(
        n18065) );
  NOR2_X1 U21126 ( .A1(n18062), .A2(n18096), .ZN(n18107) );
  NOR2_X2 U21127 ( .A1(n18132), .A2(n18063), .ZN(n18449) );
  AOI22_X1 U21128 ( .A1(n18150), .A2(n18107), .B1(n18127), .B2(n18449), .ZN(
        n18064) );
  OAI211_X1 U21129 ( .C1(n18066), .C2(n18101), .A(n18065), .B(n18064), .ZN(
        P3_U2869) );
  NOR2_X2 U21130 ( .A1(n18132), .A2(n18067), .ZN(n18454) );
  NOR2_X2 U21131 ( .A1(n18131), .A2(n18068), .ZN(n18453) );
  AOI22_X1 U21132 ( .A1(n18127), .A2(n18454), .B1(n18095), .B2(n18453), .ZN(
        n18071) );
  NOR2_X1 U21133 ( .A1(n18069), .A2(n18096), .ZN(n18110) );
  AND2_X1 U21134 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18442), .ZN(n18455) );
  AOI22_X1 U21135 ( .A1(n18150), .A2(n18110), .B1(n18488), .B2(n18455), .ZN(
        n18070) );
  OAI211_X1 U21136 ( .C1(n18072), .C2(n18101), .A(n18071), .B(n18070), .ZN(
        P3_U2870) );
  NOR2_X2 U21137 ( .A1(n18132), .A2(n18073), .ZN(n18461) );
  NOR2_X2 U21138 ( .A1(n18131), .A2(n18074), .ZN(n18459) );
  AOI22_X1 U21139 ( .A1(n18127), .A2(n18461), .B1(n18095), .B2(n18459), .ZN(
        n18077) );
  NOR2_X1 U21140 ( .A1(n18075), .A2(n18096), .ZN(n18113) );
  NOR2_X2 U21141 ( .A1(n19155), .A2(n18132), .ZN(n18460) );
  AOI22_X1 U21142 ( .A1(n18150), .A2(n18113), .B1(n18488), .B2(n18460), .ZN(
        n18076) );
  OAI211_X1 U21143 ( .C1(n18078), .C2(n18101), .A(n18077), .B(n18076), .ZN(
        P3_U2871) );
  AND2_X1 U21144 ( .A1(n18442), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18466) );
  NOR2_X2 U21145 ( .A1(n18131), .A2(n18079), .ZN(n18465) );
  AOI22_X1 U21146 ( .A1(n18127), .A2(n18466), .B1(n18095), .B2(n18465), .ZN(
        n18082) );
  NOR2_X1 U21147 ( .A1(n18080), .A2(n18096), .ZN(n18116) );
  NOR2_X2 U21148 ( .A1(n19161), .A2(n18132), .ZN(n18467) );
  AOI22_X1 U21149 ( .A1(n18150), .A2(n18116), .B1(n18488), .B2(n18467), .ZN(
        n18081) );
  OAI211_X1 U21150 ( .C1(n18083), .C2(n18101), .A(n18082), .B(n18081), .ZN(
        P3_U2872) );
  AND2_X1 U21151 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18442), .ZN(n18471) );
  NOR2_X2 U21152 ( .A1(n18131), .A2(n18084), .ZN(n18472) );
  AOI22_X1 U21153 ( .A1(n18488), .A2(n18471), .B1(n18095), .B2(n18472), .ZN(
        n18088) );
  NOR2_X1 U21154 ( .A1(n18085), .A2(n18096), .ZN(n18119) );
  NOR2_X2 U21155 ( .A1(n18132), .A2(n18086), .ZN(n18473) );
  AOI22_X1 U21156 ( .A1(n18173), .A2(n18119), .B1(n18127), .B2(n18473), .ZN(
        n18087) );
  OAI211_X1 U21157 ( .C1(n18089), .C2(n18101), .A(n18088), .B(n18087), .ZN(
        P3_U2873) );
  NOR2_X2 U21158 ( .A1(n18132), .A2(n19170), .ZN(n18478) );
  NOR2_X2 U21159 ( .A1(n18131), .A2(n18090), .ZN(n18477) );
  AOI22_X1 U21160 ( .A1(n18127), .A2(n18478), .B1(n18095), .B2(n18477), .ZN(
        n18093) );
  NOR2_X1 U21161 ( .A1(n18091), .A2(n18096), .ZN(n18122) );
  NOR2_X2 U21162 ( .A1(n14052), .A2(n18132), .ZN(n18479) );
  AOI22_X1 U21163 ( .A1(n18150), .A2(n18122), .B1(n18488), .B2(n18479), .ZN(
        n18092) );
  OAI211_X1 U21164 ( .C1(n18094), .C2(n18101), .A(n18093), .B(n18092), .ZN(
        P3_U2874) );
  AND2_X1 U21165 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18442), .ZN(n18487) );
  NOR2_X2 U21166 ( .A1(n20841), .A2(n18131), .ZN(n18484) );
  AOI22_X1 U21167 ( .A1(n18127), .A2(n18487), .B1(n18095), .B2(n18484), .ZN(
        n18100) );
  NOR2_X1 U21168 ( .A1(n18097), .A2(n18096), .ZN(n18125) );
  NOR2_X2 U21169 ( .A1(n18132), .A2(n18098), .ZN(n18486) );
  AOI22_X1 U21170 ( .A1(n18150), .A2(n18125), .B1(n18488), .B2(n18486), .ZN(
        n18099) );
  OAI211_X1 U21171 ( .C1(n21017), .C2(n18101), .A(n18100), .B(n18099), .ZN(
        P3_U2875) );
  INV_X1 U21172 ( .A(n18201), .ZN(n18156) );
  NAND2_X1 U21173 ( .A1(n18156), .A2(n18289), .ZN(n18157) );
  NAND2_X1 U21174 ( .A1(n18536), .A2(n18560), .ZN(n18290) );
  NOR2_X1 U21175 ( .A1(n18201), .A2(n18290), .ZN(n18126) );
  AOI22_X1 U21176 ( .A1(n18443), .A2(n18127), .B1(n18437), .B2(n18126), .ZN(
        n18106) );
  NOR2_X1 U21177 ( .A1(n18536), .A2(n18103), .ZN(n18439) );
  NAND2_X1 U21178 ( .A1(n18364), .A2(n18104), .ZN(n18292) );
  NOR2_X1 U21179 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18292), .ZN(
        n18387) );
  AOI22_X1 U21180 ( .A1(n18442), .A2(n18439), .B1(n18156), .B2(n18387), .ZN(
        n18128) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18128), .B1(
        n18436), .B2(n18438), .ZN(n18105) );
  OAI211_X1 U21182 ( .C1(n18446), .C2(n18157), .A(n18106), .B(n18105), .ZN(
        P3_U2876) );
  INV_X1 U21183 ( .A(n18107), .ZN(n18452) );
  AOI22_X1 U21184 ( .A1(n18436), .A2(n18449), .B1(n18447), .B2(n18126), .ZN(
        n18109) );
  AOI22_X1 U21185 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18128), .B1(
        n18127), .B2(n18448), .ZN(n18108) );
  OAI211_X1 U21186 ( .C1(n18452), .C2(n18157), .A(n18109), .B(n18108), .ZN(
        P3_U2877) );
  INV_X1 U21187 ( .A(n18110), .ZN(n18458) );
  AOI22_X1 U21188 ( .A1(n18436), .A2(n18454), .B1(n18453), .B2(n18126), .ZN(
        n18112) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18128), .B1(
        n18127), .B2(n18455), .ZN(n18111) );
  OAI211_X1 U21190 ( .C1(n18458), .C2(n18157), .A(n18112), .B(n18111), .ZN(
        P3_U2878) );
  INV_X1 U21191 ( .A(n18113), .ZN(n18464) );
  AOI22_X1 U21192 ( .A1(n18127), .A2(n18460), .B1(n18459), .B2(n18126), .ZN(
        n18115) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18128), .B1(
        n18436), .B2(n18461), .ZN(n18114) );
  OAI211_X1 U21194 ( .C1(n18464), .C2(n18157), .A(n18115), .B(n18114), .ZN(
        P3_U2879) );
  AOI22_X1 U21195 ( .A1(n18127), .A2(n18467), .B1(n18465), .B2(n18126), .ZN(
        n18118) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18128), .B1(
        n18436), .B2(n18466), .ZN(n18117) );
  OAI211_X1 U21197 ( .C1(n18470), .C2(n18157), .A(n18118), .B(n18117), .ZN(
        P3_U2880) );
  INV_X1 U21198 ( .A(n18119), .ZN(n18476) );
  AOI22_X1 U21199 ( .A1(n18436), .A2(n18473), .B1(n18472), .B2(n18126), .ZN(
        n18121) );
  AOI22_X1 U21200 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18128), .B1(
        n18127), .B2(n18471), .ZN(n18120) );
  OAI211_X1 U21201 ( .C1(n18476), .C2(n18157), .A(n18121), .B(n18120), .ZN(
        P3_U2881) );
  INV_X1 U21202 ( .A(n18122), .ZN(n18482) );
  AOI22_X1 U21203 ( .A1(n18127), .A2(n18479), .B1(n18477), .B2(n18126), .ZN(
        n18124) );
  AOI22_X1 U21204 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18128), .B1(
        n18436), .B2(n18478), .ZN(n18123) );
  OAI211_X1 U21205 ( .C1(n18482), .C2(n18157), .A(n18124), .B(n18123), .ZN(
        P3_U2882) );
  INV_X1 U21206 ( .A(n18125), .ZN(n18492) );
  AOI22_X1 U21207 ( .A1(n18127), .A2(n18486), .B1(n18484), .B2(n18126), .ZN(
        n18130) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18128), .B1(
        n18436), .B2(n18487), .ZN(n18129) );
  OAI211_X1 U21209 ( .C1(n18492), .C2(n18157), .A(n18130), .B(n18129), .ZN(
        P3_U2883) );
  NAND2_X1 U21210 ( .A1(n18156), .A2(n18314), .ZN(n18154) );
  AOI21_X1 U21211 ( .B1(n18157), .B2(n18154), .A(n18410), .ZN(n18149) );
  AOI22_X1 U21212 ( .A1(n18150), .A2(n18438), .B1(n18437), .B2(n18149), .ZN(
        n18136) );
  INV_X1 U21213 ( .A(n18154), .ZN(n18218) );
  AOI21_X1 U21214 ( .B1(n18157), .B2(n18154), .A(n18131), .ZN(n18178) );
  NOR2_X1 U21215 ( .A1(n18133), .A2(n18132), .ZN(n18134) );
  OAI22_X1 U21216 ( .A1(n18218), .A2(n18684), .B1(n18178), .B2(n18134), .ZN(
        n18151) );
  AOI22_X1 U21217 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18151), .B1(
        n18436), .B2(n18443), .ZN(n18135) );
  OAI211_X1 U21218 ( .C1(n18446), .C2(n18154), .A(n18136), .B(n18135), .ZN(
        P3_U2884) );
  AOI22_X1 U21219 ( .A1(n18173), .A2(n18449), .B1(n18447), .B2(n18149), .ZN(
        n18138) );
  AOI22_X1 U21220 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18151), .B1(
        n18436), .B2(n18448), .ZN(n18137) );
  OAI211_X1 U21221 ( .C1(n18452), .C2(n18154), .A(n18138), .B(n18137), .ZN(
        P3_U2885) );
  AOI22_X1 U21222 ( .A1(n18173), .A2(n18454), .B1(n18453), .B2(n18149), .ZN(
        n18140) );
  AOI22_X1 U21223 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18151), .B1(
        n18436), .B2(n18455), .ZN(n18139) );
  OAI211_X1 U21224 ( .C1(n18458), .C2(n18154), .A(n18140), .B(n18139), .ZN(
        P3_U2886) );
  AOI22_X1 U21225 ( .A1(n18173), .A2(n18461), .B1(n18459), .B2(n18149), .ZN(
        n18142) );
  AOI22_X1 U21226 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18151), .B1(
        n18436), .B2(n18460), .ZN(n18141) );
  OAI211_X1 U21227 ( .C1(n18464), .C2(n18154), .A(n18142), .B(n18141), .ZN(
        P3_U2887) );
  AOI22_X1 U21228 ( .A1(n18173), .A2(n18466), .B1(n18465), .B2(n18149), .ZN(
        n18144) );
  AOI22_X1 U21229 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18151), .B1(
        n18436), .B2(n18467), .ZN(n18143) );
  OAI211_X1 U21230 ( .C1(n18470), .C2(n18154), .A(n18144), .B(n18143), .ZN(
        P3_U2888) );
  AOI22_X1 U21231 ( .A1(n18436), .A2(n18471), .B1(n18472), .B2(n18149), .ZN(
        n18146) );
  AOI22_X1 U21232 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18151), .B1(
        n18150), .B2(n18473), .ZN(n18145) );
  OAI211_X1 U21233 ( .C1(n18476), .C2(n18154), .A(n18146), .B(n18145), .ZN(
        P3_U2889) );
  AOI22_X1 U21234 ( .A1(n18173), .A2(n18478), .B1(n18477), .B2(n18149), .ZN(
        n18148) );
  AOI22_X1 U21235 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18151), .B1(
        n18436), .B2(n18479), .ZN(n18147) );
  OAI211_X1 U21236 ( .C1(n18482), .C2(n18154), .A(n18148), .B(n18147), .ZN(
        P3_U2890) );
  AOI22_X1 U21237 ( .A1(n18436), .A2(n18486), .B1(n18484), .B2(n18149), .ZN(
        n18153) );
  AOI22_X1 U21238 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18151), .B1(
        n18150), .B2(n18487), .ZN(n18152) );
  OAI211_X1 U21239 ( .C1(n18492), .C2(n18154), .A(n18153), .B(n18152), .ZN(
        P3_U2891) );
  NOR2_X2 U21240 ( .A1(n18535), .A2(n18201), .ZN(n18239) );
  INV_X1 U21241 ( .A(n18239), .ZN(n18177) );
  OAI21_X1 U21242 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18315), .A(
        n18364), .ZN(n18155) );
  AOI21_X1 U21243 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18535), .A(n18155), 
        .ZN(n18244) );
  NAND2_X1 U21244 ( .A1(n18156), .A2(n18244), .ZN(n18174) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18174), .B1(
        n18437), .B2(n18172), .ZN(n18159) );
  INV_X1 U21246 ( .A(n18157), .ZN(n18196) );
  AOI22_X1 U21247 ( .A1(n18173), .A2(n18443), .B1(n18438), .B2(n18196), .ZN(
        n18158) );
  OAI211_X1 U21248 ( .C1(n18446), .C2(n18177), .A(n18159), .B(n18158), .ZN(
        P3_U2892) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18174), .B1(
        n18447), .B2(n18172), .ZN(n18161) );
  AOI22_X1 U21250 ( .A1(n18173), .A2(n18448), .B1(n18449), .B2(n18196), .ZN(
        n18160) );
  OAI211_X1 U21251 ( .C1(n18452), .C2(n18177), .A(n18161), .B(n18160), .ZN(
        P3_U2893) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18174), .B1(
        n18453), .B2(n18172), .ZN(n18163) );
  AOI22_X1 U21253 ( .A1(n18173), .A2(n18455), .B1(n18454), .B2(n18196), .ZN(
        n18162) );
  OAI211_X1 U21254 ( .C1(n18458), .C2(n18177), .A(n18163), .B(n18162), .ZN(
        P3_U2894) );
  AOI22_X1 U21255 ( .A1(n18461), .A2(n18196), .B1(n18459), .B2(n18172), .ZN(
        n18165) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18174), .B1(
        n18173), .B2(n18460), .ZN(n18164) );
  OAI211_X1 U21257 ( .C1(n18464), .C2(n18177), .A(n18165), .B(n18164), .ZN(
        P3_U2895) );
  AOI22_X1 U21258 ( .A1(n18466), .A2(n18196), .B1(n18465), .B2(n18172), .ZN(
        n18167) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18174), .B1(
        n18173), .B2(n18467), .ZN(n18166) );
  OAI211_X1 U21260 ( .C1(n18470), .C2(n18177), .A(n18167), .B(n18166), .ZN(
        P3_U2896) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18174), .B1(
        n18472), .B2(n18172), .ZN(n18169) );
  AOI22_X1 U21262 ( .A1(n18173), .A2(n18471), .B1(n18473), .B2(n18196), .ZN(
        n18168) );
  OAI211_X1 U21263 ( .C1(n18476), .C2(n18177), .A(n18169), .B(n18168), .ZN(
        P3_U2897) );
  AOI22_X1 U21264 ( .A1(n18477), .A2(n18172), .B1(n18478), .B2(n18196), .ZN(
        n18171) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18174), .B1(
        n18173), .B2(n18479), .ZN(n18170) );
  OAI211_X1 U21266 ( .C1(n18482), .C2(n18177), .A(n18171), .B(n18170), .ZN(
        P3_U2898) );
  AOI22_X1 U21267 ( .A1(n18487), .A2(n18196), .B1(n18484), .B2(n18172), .ZN(
        n18176) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18174), .B1(
        n18173), .B2(n18486), .ZN(n18175) );
  OAI211_X1 U21269 ( .C1(n18492), .C2(n18177), .A(n18176), .B(n18175), .ZN(
        P3_U2899) );
  NOR2_X2 U21270 ( .A1(n18537), .A2(n18291), .ZN(n18261) );
  INV_X1 U21271 ( .A(n18261), .ZN(n18200) );
  NAND2_X1 U21272 ( .A1(n18177), .A2(n18200), .ZN(n18223) );
  AND2_X1 U21273 ( .A1(n18560), .A2(n18223), .ZN(n18195) );
  AOI22_X1 U21274 ( .A1(n18438), .A2(n18218), .B1(n18437), .B2(n18195), .ZN(
        n18182) );
  AOI22_X1 U21275 ( .A1(n18223), .A2(n18364), .B1(n18315), .B2(n18178), .ZN(
        n18179) );
  AOI21_X1 U21276 ( .B1(n18200), .B2(P3_STATE2_REG_3__SCAN_IN), .A(n18179), 
        .ZN(n18180) );
  INV_X1 U21277 ( .A(n18180), .ZN(n18197) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18197), .B1(
        n18443), .B2(n18196), .ZN(n18181) );
  OAI211_X1 U21279 ( .C1(n18446), .C2(n18200), .A(n18182), .B(n18181), .ZN(
        P3_U2900) );
  AOI22_X1 U21280 ( .A1(n18448), .A2(n18196), .B1(n18447), .B2(n18195), .ZN(
        n18184) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18197), .B1(
        n18449), .B2(n18218), .ZN(n18183) );
  OAI211_X1 U21282 ( .C1(n18452), .C2(n18200), .A(n18184), .B(n18183), .ZN(
        P3_U2901) );
  AOI22_X1 U21283 ( .A1(n18455), .A2(n18196), .B1(n18453), .B2(n18195), .ZN(
        n18186) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18197), .B1(
        n18454), .B2(n18218), .ZN(n18185) );
  OAI211_X1 U21285 ( .C1(n18458), .C2(n18200), .A(n18186), .B(n18185), .ZN(
        P3_U2902) );
  AOI22_X1 U21286 ( .A1(n18461), .A2(n18218), .B1(n18459), .B2(n18195), .ZN(
        n18188) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18197), .B1(
        n18460), .B2(n18196), .ZN(n18187) );
  OAI211_X1 U21288 ( .C1(n18464), .C2(n18200), .A(n18188), .B(n18187), .ZN(
        P3_U2903) );
  AOI22_X1 U21289 ( .A1(n18467), .A2(n18196), .B1(n18465), .B2(n18195), .ZN(
        n18190) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18197), .B1(
        n18466), .B2(n18218), .ZN(n18189) );
  OAI211_X1 U21291 ( .C1(n18470), .C2(n18200), .A(n18190), .B(n18189), .ZN(
        P3_U2904) );
  AOI22_X1 U21292 ( .A1(n18472), .A2(n18195), .B1(n18471), .B2(n18196), .ZN(
        n18192) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18197), .B1(
        n18473), .B2(n18218), .ZN(n18191) );
  OAI211_X1 U21294 ( .C1(n18476), .C2(n18200), .A(n18192), .B(n18191), .ZN(
        P3_U2905) );
  AOI22_X1 U21295 ( .A1(n18477), .A2(n18195), .B1(n18478), .B2(n18218), .ZN(
        n18194) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18197), .B1(
        n18479), .B2(n18196), .ZN(n18193) );
  OAI211_X1 U21297 ( .C1(n18482), .C2(n18200), .A(n18194), .B(n18193), .ZN(
        P3_U2906) );
  AOI22_X1 U21298 ( .A1(n18487), .A2(n18218), .B1(n18484), .B2(n18195), .ZN(
        n18199) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18197), .B1(
        n18486), .B2(n18196), .ZN(n18198) );
  OAI211_X1 U21300 ( .C1(n18492), .C2(n18200), .A(n18199), .B(n18198), .ZN(
        P3_U2907) );
  NAND2_X1 U21301 ( .A1(n18289), .A2(n18243), .ZN(n18245) );
  NOR2_X1 U21302 ( .A1(n18290), .A2(n18291), .ZN(n18217) );
  AOI22_X1 U21303 ( .A1(n18443), .A2(n18218), .B1(n18437), .B2(n18217), .ZN(
        n18204) );
  NOR2_X1 U21304 ( .A1(n18536), .A2(n18201), .ZN(n18202) );
  AOI22_X1 U21305 ( .A1(n18442), .A2(n18202), .B1(n18387), .B2(n18243), .ZN(
        n18219) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18219), .B1(
        n18438), .B2(n18239), .ZN(n18203) );
  OAI211_X1 U21307 ( .C1(n18446), .C2(n18245), .A(n18204), .B(n18203), .ZN(
        P3_U2908) );
  AOI22_X1 U21308 ( .A1(n18448), .A2(n18218), .B1(n18447), .B2(n18217), .ZN(
        n18206) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18219), .B1(
        n18449), .B2(n18239), .ZN(n18205) );
  OAI211_X1 U21310 ( .C1(n18452), .C2(n18245), .A(n18206), .B(n18205), .ZN(
        P3_U2909) );
  AOI22_X1 U21311 ( .A1(n18455), .A2(n18218), .B1(n18453), .B2(n18217), .ZN(
        n18208) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18219), .B1(
        n18454), .B2(n18239), .ZN(n18207) );
  OAI211_X1 U21313 ( .C1(n18458), .C2(n18245), .A(n18208), .B(n18207), .ZN(
        P3_U2910) );
  AOI22_X1 U21314 ( .A1(n18461), .A2(n18239), .B1(n18459), .B2(n18217), .ZN(
        n18210) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18219), .B1(
        n18460), .B2(n18218), .ZN(n18209) );
  OAI211_X1 U21316 ( .C1(n18464), .C2(n18245), .A(n18210), .B(n18209), .ZN(
        P3_U2911) );
  AOI22_X1 U21317 ( .A1(n18467), .A2(n18218), .B1(n18465), .B2(n18217), .ZN(
        n18212) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18219), .B1(
        n18466), .B2(n18239), .ZN(n18211) );
  OAI211_X1 U21319 ( .C1(n18470), .C2(n18245), .A(n18212), .B(n18211), .ZN(
        P3_U2912) );
  AOI22_X1 U21320 ( .A1(n18472), .A2(n18217), .B1(n18471), .B2(n18218), .ZN(
        n18214) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18219), .B1(
        n18473), .B2(n18239), .ZN(n18213) );
  OAI211_X1 U21322 ( .C1(n18476), .C2(n18245), .A(n18214), .B(n18213), .ZN(
        P3_U2913) );
  AOI22_X1 U21323 ( .A1(n18477), .A2(n18217), .B1(n18478), .B2(n18239), .ZN(
        n18216) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18219), .B1(
        n18479), .B2(n18218), .ZN(n18215) );
  OAI211_X1 U21325 ( .C1(n18482), .C2(n18245), .A(n18216), .B(n18215), .ZN(
        P3_U2914) );
  AOI22_X1 U21326 ( .A1(n18487), .A2(n18239), .B1(n18484), .B2(n18217), .ZN(
        n18221) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18219), .B1(
        n18486), .B2(n18218), .ZN(n18220) );
  OAI211_X1 U21328 ( .C1(n18492), .C2(n18245), .A(n18221), .B(n18220), .ZN(
        P3_U2915) );
  NAND2_X1 U21329 ( .A1(n18314), .A2(n18243), .ZN(n18266) );
  NAND2_X1 U21330 ( .A1(n18245), .A2(n18266), .ZN(n18267) );
  AND2_X1 U21331 ( .A1(n18560), .A2(n18267), .ZN(n18238) );
  AOI22_X1 U21332 ( .A1(n18438), .A2(n18261), .B1(n18437), .B2(n18238), .ZN(
        n18225) );
  INV_X1 U21333 ( .A(n18222), .ZN(n18414) );
  OAI221_X1 U21334 ( .B1(n18267), .B2(n18315), .C1(n18267), .C2(n18223), .A(
        n18414), .ZN(n18240) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18240), .B1(
        n18443), .B2(n18239), .ZN(n18224) );
  OAI211_X1 U21336 ( .C1(n18446), .C2(n18266), .A(n18225), .B(n18224), .ZN(
        P3_U2916) );
  AOI22_X1 U21337 ( .A1(n18448), .A2(n18239), .B1(n18447), .B2(n18238), .ZN(
        n18227) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18240), .B1(
        n18449), .B2(n18261), .ZN(n18226) );
  OAI211_X1 U21339 ( .C1(n18452), .C2(n18266), .A(n18227), .B(n18226), .ZN(
        P3_U2917) );
  AOI22_X1 U21340 ( .A1(n18455), .A2(n18239), .B1(n18453), .B2(n18238), .ZN(
        n18229) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18240), .B1(
        n18454), .B2(n18261), .ZN(n18228) );
  OAI211_X1 U21342 ( .C1(n18458), .C2(n18266), .A(n18229), .B(n18228), .ZN(
        P3_U2918) );
  AOI22_X1 U21343 ( .A1(n18460), .A2(n18239), .B1(n18459), .B2(n18238), .ZN(
        n18231) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18240), .B1(
        n18461), .B2(n18261), .ZN(n18230) );
  OAI211_X1 U21345 ( .C1(n18464), .C2(n18266), .A(n18231), .B(n18230), .ZN(
        P3_U2919) );
  AOI22_X1 U21346 ( .A1(n18467), .A2(n18239), .B1(n18465), .B2(n18238), .ZN(
        n18233) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18240), .B1(
        n18466), .B2(n18261), .ZN(n18232) );
  OAI211_X1 U21348 ( .C1(n18470), .C2(n18266), .A(n18233), .B(n18232), .ZN(
        P3_U2920) );
  AOI22_X1 U21349 ( .A1(n18473), .A2(n18261), .B1(n18472), .B2(n18238), .ZN(
        n18235) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18240), .B1(
        n18471), .B2(n18239), .ZN(n18234) );
  OAI211_X1 U21351 ( .C1(n18476), .C2(n18266), .A(n18235), .B(n18234), .ZN(
        P3_U2921) );
  AOI22_X1 U21352 ( .A1(n18477), .A2(n18238), .B1(n18478), .B2(n18261), .ZN(
        n18237) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18240), .B1(
        n18479), .B2(n18239), .ZN(n18236) );
  OAI211_X1 U21354 ( .C1(n18482), .C2(n18266), .A(n18237), .B(n18236), .ZN(
        P3_U2922) );
  AOI22_X1 U21355 ( .A1(n18487), .A2(n18261), .B1(n18484), .B2(n18238), .ZN(
        n18242) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18240), .B1(
        n18486), .B2(n18239), .ZN(n18241) );
  OAI211_X1 U21357 ( .C1(n18492), .C2(n18266), .A(n18242), .B(n18241), .ZN(
        P3_U2923) );
  NOR2_X2 U21358 ( .A1(n18535), .A2(n18291), .ZN(n18333) );
  INV_X1 U21359 ( .A(n18333), .ZN(n18265) );
  NAND2_X1 U21360 ( .A1(n18244), .A2(n18243), .ZN(n18262) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18262), .B1(
        n18437), .B2(n18260), .ZN(n18247) );
  INV_X1 U21362 ( .A(n18245), .ZN(n18285) );
  AOI22_X1 U21363 ( .A1(n18443), .A2(n18261), .B1(n18438), .B2(n18285), .ZN(
        n18246) );
  OAI211_X1 U21364 ( .C1(n18446), .C2(n18265), .A(n18247), .B(n18246), .ZN(
        P3_U2924) );
  AOI22_X1 U21365 ( .A1(n18449), .A2(n18285), .B1(n18447), .B2(n18260), .ZN(
        n18249) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18262), .B1(
        n18448), .B2(n18261), .ZN(n18248) );
  OAI211_X1 U21367 ( .C1(n18452), .C2(n18265), .A(n18249), .B(n18248), .ZN(
        P3_U2925) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18262), .B1(
        n18453), .B2(n18260), .ZN(n18251) );
  AOI22_X1 U21369 ( .A1(n18455), .A2(n18261), .B1(n18454), .B2(n18285), .ZN(
        n18250) );
  OAI211_X1 U21370 ( .C1(n18458), .C2(n18265), .A(n18251), .B(n18250), .ZN(
        P3_U2926) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18262), .B1(
        n18459), .B2(n18260), .ZN(n18253) );
  AOI22_X1 U21372 ( .A1(n18460), .A2(n18261), .B1(n18461), .B2(n18285), .ZN(
        n18252) );
  OAI211_X1 U21373 ( .C1(n18464), .C2(n18265), .A(n18253), .B(n18252), .ZN(
        P3_U2927) );
  AOI22_X1 U21374 ( .A1(n18466), .A2(n18285), .B1(n18465), .B2(n18260), .ZN(
        n18255) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18262), .B1(
        n18467), .B2(n18261), .ZN(n18254) );
  OAI211_X1 U21376 ( .C1(n18470), .C2(n18265), .A(n18255), .B(n18254), .ZN(
        P3_U2928) );
  AOI22_X1 U21377 ( .A1(n18472), .A2(n18260), .B1(n18471), .B2(n18261), .ZN(
        n18257) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18262), .B1(
        n18473), .B2(n18285), .ZN(n18256) );
  OAI211_X1 U21379 ( .C1(n18476), .C2(n18265), .A(n18257), .B(n18256), .ZN(
        P3_U2929) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18262), .B1(
        n18477), .B2(n18260), .ZN(n18259) );
  AOI22_X1 U21381 ( .A1(n18479), .A2(n18261), .B1(n18478), .B2(n18285), .ZN(
        n18258) );
  OAI211_X1 U21382 ( .C1(n18482), .C2(n18265), .A(n18259), .B(n18258), .ZN(
        P3_U2930) );
  AOI22_X1 U21383 ( .A1(n18486), .A2(n18261), .B1(n18484), .B2(n18260), .ZN(
        n18264) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18262), .B1(
        n18487), .B2(n18285), .ZN(n18263) );
  OAI211_X1 U21385 ( .C1(n18492), .C2(n18265), .A(n18264), .B(n18263), .ZN(
        P3_U2931) );
  INV_X1 U21386 ( .A(n18338), .ZN(n18386) );
  NOR2_X2 U21387 ( .A1(n18537), .A2(n18386), .ZN(n18355) );
  INV_X1 U21388 ( .A(n18355), .ZN(n18288) );
  INV_X1 U21389 ( .A(n18266), .ZN(n18310) );
  NOR2_X1 U21390 ( .A1(n18333), .A2(n18355), .ZN(n18316) );
  NOR2_X1 U21391 ( .A1(n18410), .A2(n18316), .ZN(n18283) );
  AOI22_X1 U21392 ( .A1(n18438), .A2(n18310), .B1(n18437), .B2(n18283), .ZN(
        n18270) );
  INV_X1 U21393 ( .A(n18316), .ZN(n18268) );
  OAI221_X1 U21394 ( .B1(n18268), .B2(n18315), .C1(n18268), .C2(n18267), .A(
        n18414), .ZN(n18284) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18284), .B1(
        n18443), .B2(n18285), .ZN(n18269) );
  OAI211_X1 U21396 ( .C1(n18446), .C2(n18288), .A(n18270), .B(n18269), .ZN(
        P3_U2932) );
  AOI22_X1 U21397 ( .A1(n18449), .A2(n18310), .B1(n18447), .B2(n18283), .ZN(
        n18272) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18284), .B1(
        n18448), .B2(n18285), .ZN(n18271) );
  OAI211_X1 U21399 ( .C1(n18452), .C2(n18288), .A(n18272), .B(n18271), .ZN(
        P3_U2933) );
  AOI22_X1 U21400 ( .A1(n18454), .A2(n18310), .B1(n18453), .B2(n18283), .ZN(
        n18274) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18284), .B1(
        n18455), .B2(n18285), .ZN(n18273) );
  OAI211_X1 U21402 ( .C1(n18458), .C2(n18288), .A(n18274), .B(n18273), .ZN(
        P3_U2934) );
  AOI22_X1 U21403 ( .A1(n18461), .A2(n18310), .B1(n18459), .B2(n18283), .ZN(
        n18276) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18284), .B1(
        n18460), .B2(n18285), .ZN(n18275) );
  OAI211_X1 U21405 ( .C1(n18464), .C2(n18288), .A(n18276), .B(n18275), .ZN(
        P3_U2935) );
  AOI22_X1 U21406 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18284), .B1(
        n18465), .B2(n18283), .ZN(n18278) );
  AOI22_X1 U21407 ( .A1(n18467), .A2(n18285), .B1(n18466), .B2(n18310), .ZN(
        n18277) );
  OAI211_X1 U21408 ( .C1(n18470), .C2(n18288), .A(n18278), .B(n18277), .ZN(
        P3_U2936) );
  AOI22_X1 U21409 ( .A1(n18473), .A2(n18310), .B1(n18472), .B2(n18283), .ZN(
        n18280) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18284), .B1(
        n18471), .B2(n18285), .ZN(n18279) );
  OAI211_X1 U21411 ( .C1(n18476), .C2(n18288), .A(n18280), .B(n18279), .ZN(
        P3_U2937) );
  AOI22_X1 U21412 ( .A1(n18479), .A2(n18285), .B1(n18477), .B2(n18283), .ZN(
        n18282) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18284), .B1(
        n18478), .B2(n18310), .ZN(n18281) );
  OAI211_X1 U21414 ( .C1(n18482), .C2(n18288), .A(n18282), .B(n18281), .ZN(
        P3_U2938) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18284), .B1(
        n18484), .B2(n18283), .ZN(n18287) );
  AOI22_X1 U21416 ( .A1(n18486), .A2(n18285), .B1(n18487), .B2(n18310), .ZN(
        n18286) );
  OAI211_X1 U21417 ( .C1(n18492), .C2(n18288), .A(n18287), .B(n18286), .ZN(
        P3_U2939) );
  NAND2_X1 U21418 ( .A1(n18289), .A2(n18338), .ZN(n18339) );
  NOR2_X1 U21419 ( .A1(n18290), .A2(n18386), .ZN(n18309) );
  AOI22_X1 U21420 ( .A1(n18443), .A2(n18310), .B1(n18437), .B2(n18309), .ZN(
        n18296) );
  NOR2_X1 U21421 ( .A1(n18536), .A2(n18291), .ZN(n18294) );
  INV_X1 U21422 ( .A(n18292), .ZN(n18440) );
  NOR2_X1 U21423 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18386), .ZN(
        n18293) );
  AOI22_X1 U21424 ( .A1(n18442), .A2(n18294), .B1(n18440), .B2(n18293), .ZN(
        n18311) );
  AOI22_X1 U21425 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18311), .B1(
        n18438), .B2(n18333), .ZN(n18295) );
  OAI211_X1 U21426 ( .C1(n18446), .C2(n18339), .A(n18296), .B(n18295), .ZN(
        P3_U2940) );
  AOI22_X1 U21427 ( .A1(n18449), .A2(n18333), .B1(n18447), .B2(n18309), .ZN(
        n18298) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18311), .B1(
        n18448), .B2(n18310), .ZN(n18297) );
  OAI211_X1 U21429 ( .C1(n18452), .C2(n18339), .A(n18298), .B(n18297), .ZN(
        P3_U2941) );
  AOI22_X1 U21430 ( .A1(n18455), .A2(n18310), .B1(n18453), .B2(n18309), .ZN(
        n18300) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18311), .B1(
        n18454), .B2(n18333), .ZN(n18299) );
  OAI211_X1 U21432 ( .C1(n18458), .C2(n18339), .A(n18300), .B(n18299), .ZN(
        P3_U2942) );
  AOI22_X1 U21433 ( .A1(n18460), .A2(n18310), .B1(n18459), .B2(n18309), .ZN(
        n18302) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18311), .B1(
        n18461), .B2(n18333), .ZN(n18301) );
  OAI211_X1 U21435 ( .C1(n18464), .C2(n18339), .A(n18302), .B(n18301), .ZN(
        P3_U2943) );
  AOI22_X1 U21436 ( .A1(n18467), .A2(n18310), .B1(n18465), .B2(n18309), .ZN(
        n18304) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18311), .B1(
        n18466), .B2(n18333), .ZN(n18303) );
  OAI211_X1 U21438 ( .C1(n18470), .C2(n18339), .A(n18304), .B(n18303), .ZN(
        P3_U2944) );
  AOI22_X1 U21439 ( .A1(n18473), .A2(n18333), .B1(n18472), .B2(n18309), .ZN(
        n18306) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18311), .B1(
        n18471), .B2(n18310), .ZN(n18305) );
  OAI211_X1 U21441 ( .C1(n18476), .C2(n18339), .A(n18306), .B(n18305), .ZN(
        P3_U2945) );
  AOI22_X1 U21442 ( .A1(n18479), .A2(n18310), .B1(n18477), .B2(n18309), .ZN(
        n18308) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18311), .B1(
        n18478), .B2(n18333), .ZN(n18307) );
  OAI211_X1 U21444 ( .C1(n18482), .C2(n18339), .A(n18308), .B(n18307), .ZN(
        P3_U2946) );
  AOI22_X1 U21445 ( .A1(n18486), .A2(n18310), .B1(n18484), .B2(n18309), .ZN(
        n18313) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18311), .B1(
        n18487), .B2(n18333), .ZN(n18312) );
  OAI211_X1 U21447 ( .C1(n18492), .C2(n18339), .A(n18313), .B(n18312), .ZN(
        P3_U2947) );
  NAND2_X1 U21448 ( .A1(n18314), .A2(n18338), .ZN(n18337) );
  AOI22_X1 U21449 ( .A1(n18443), .A2(n18333), .B1(n18437), .B2(n18332), .ZN(
        n18319) );
  INV_X1 U21450 ( .A(n18337), .ZN(n18405) );
  INV_X1 U21451 ( .A(n18315), .ZN(n18413) );
  AOI221_X1 U21452 ( .B1(n18316), .B2(n18339), .C1(n18413), .C2(n18339), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18317) );
  OAI21_X1 U21453 ( .B1(n18405), .B2(n18317), .A(n18364), .ZN(n18334) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18334), .B1(
        n18438), .B2(n18355), .ZN(n18318) );
  OAI211_X1 U21455 ( .C1(n18446), .C2(n18337), .A(n18319), .B(n18318), .ZN(
        P3_U2948) );
  AOI22_X1 U21456 ( .A1(n18449), .A2(n18355), .B1(n18447), .B2(n18332), .ZN(
        n18321) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18334), .B1(
        n18448), .B2(n18333), .ZN(n18320) );
  OAI211_X1 U21458 ( .C1(n18452), .C2(n18337), .A(n18321), .B(n18320), .ZN(
        P3_U2949) );
  AOI22_X1 U21459 ( .A1(n18454), .A2(n18355), .B1(n18453), .B2(n18332), .ZN(
        n18323) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18334), .B1(
        n18455), .B2(n18333), .ZN(n18322) );
  OAI211_X1 U21461 ( .C1(n18458), .C2(n18337), .A(n18323), .B(n18322), .ZN(
        P3_U2950) );
  AOI22_X1 U21462 ( .A1(n18461), .A2(n18355), .B1(n18459), .B2(n18332), .ZN(
        n18325) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18334), .B1(
        n18460), .B2(n18333), .ZN(n18324) );
  OAI211_X1 U21464 ( .C1(n18464), .C2(n18337), .A(n18325), .B(n18324), .ZN(
        P3_U2951) );
  AOI22_X1 U21465 ( .A1(n18466), .A2(n18355), .B1(n18465), .B2(n18332), .ZN(
        n18327) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18334), .B1(
        n18467), .B2(n18333), .ZN(n18326) );
  OAI211_X1 U21467 ( .C1(n18470), .C2(n18337), .A(n18327), .B(n18326), .ZN(
        P3_U2952) );
  AOI22_X1 U21468 ( .A1(n18472), .A2(n18332), .B1(n18471), .B2(n18333), .ZN(
        n18329) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18334), .B1(
        n18473), .B2(n18355), .ZN(n18328) );
  OAI211_X1 U21470 ( .C1(n18476), .C2(n18337), .A(n18329), .B(n18328), .ZN(
        P3_U2953) );
  AOI22_X1 U21471 ( .A1(n18477), .A2(n18332), .B1(n18478), .B2(n18355), .ZN(
        n18331) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18334), .B1(
        n18479), .B2(n18333), .ZN(n18330) );
  OAI211_X1 U21473 ( .C1(n18482), .C2(n18337), .A(n18331), .B(n18330), .ZN(
        P3_U2954) );
  AOI22_X1 U21474 ( .A1(n18486), .A2(n18333), .B1(n18484), .B2(n18332), .ZN(
        n18336) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18334), .B1(
        n18487), .B2(n18355), .ZN(n18335) );
  OAI211_X1 U21476 ( .C1(n18492), .C2(n18337), .A(n18336), .B(n18335), .ZN(
        P3_U2955) );
  NOR2_X2 U21477 ( .A1(n18535), .A2(n18386), .ZN(n18431) );
  INV_X1 U21478 ( .A(n18431), .ZN(n18359) );
  AOI22_X1 U21479 ( .A1(n18443), .A2(n18355), .B1(n18437), .B2(n18354), .ZN(
        n18341) );
  OAI211_X1 U21480 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18442), .A(
        n18440), .B(n18338), .ZN(n18356) );
  INV_X1 U21481 ( .A(n18339), .ZN(n18380) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18356), .B1(
        n18438), .B2(n18380), .ZN(n18340) );
  OAI211_X1 U21483 ( .C1(n18446), .C2(n18359), .A(n18341), .B(n18340), .ZN(
        P3_U2956) );
  AOI22_X1 U21484 ( .A1(n18448), .A2(n18355), .B1(n18447), .B2(n18354), .ZN(
        n18343) );
  AOI22_X1 U21485 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18356), .B1(
        n18449), .B2(n18380), .ZN(n18342) );
  OAI211_X1 U21486 ( .C1(n18452), .C2(n18359), .A(n18343), .B(n18342), .ZN(
        P3_U2957) );
  AOI22_X1 U21487 ( .A1(n18454), .A2(n18380), .B1(n18453), .B2(n18354), .ZN(
        n18345) );
  AOI22_X1 U21488 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18356), .B1(
        n18455), .B2(n18355), .ZN(n18344) );
  OAI211_X1 U21489 ( .C1(n18458), .C2(n18359), .A(n18345), .B(n18344), .ZN(
        P3_U2958) );
  AOI22_X1 U21490 ( .A1(n18460), .A2(n18355), .B1(n18459), .B2(n18354), .ZN(
        n18347) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18356), .B1(
        n18461), .B2(n18380), .ZN(n18346) );
  OAI211_X1 U21492 ( .C1(n18464), .C2(n18359), .A(n18347), .B(n18346), .ZN(
        P3_U2959) );
  AOI22_X1 U21493 ( .A1(n18466), .A2(n18380), .B1(n18465), .B2(n18354), .ZN(
        n18349) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18356), .B1(
        n18467), .B2(n18355), .ZN(n18348) );
  OAI211_X1 U21495 ( .C1(n18470), .C2(n18359), .A(n18349), .B(n18348), .ZN(
        P3_U2960) );
  AOI22_X1 U21496 ( .A1(n18472), .A2(n18354), .B1(n18471), .B2(n18355), .ZN(
        n18351) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18356), .B1(
        n18473), .B2(n18380), .ZN(n18350) );
  OAI211_X1 U21498 ( .C1(n18476), .C2(n18359), .A(n18351), .B(n18350), .ZN(
        P3_U2961) );
  AOI22_X1 U21499 ( .A1(n18477), .A2(n18354), .B1(n18478), .B2(n18380), .ZN(
        n18353) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18356), .B1(
        n18479), .B2(n18355), .ZN(n18352) );
  OAI211_X1 U21501 ( .C1(n18482), .C2(n18359), .A(n18353), .B(n18352), .ZN(
        P3_U2962) );
  AOI22_X1 U21502 ( .A1(n18486), .A2(n18355), .B1(n18484), .B2(n18354), .ZN(
        n18358) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18356), .B1(
        n18487), .B2(n18380), .ZN(n18357) );
  OAI211_X1 U21504 ( .C1(n18492), .C2(n18359), .A(n18358), .B(n18357), .ZN(
        P3_U2963) );
  INV_X1 U21505 ( .A(n18385), .ZN(n18441) );
  NAND2_X1 U21506 ( .A1(n18441), .A2(n18360), .ZN(n18384) );
  INV_X1 U21507 ( .A(n18384), .ZN(n18485) );
  NOR2_X1 U21508 ( .A1(n18431), .A2(n18485), .ZN(n18412) );
  OAI21_X1 U21509 ( .B1(n18362), .B2(n18361), .A(n18412), .ZN(n18363) );
  OAI211_X1 U21510 ( .C1(n18485), .C2(n18684), .A(n18364), .B(n18363), .ZN(
        n18381) );
  NOR2_X1 U21511 ( .A1(n18410), .A2(n18412), .ZN(n18379) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18381), .B1(
        n18437), .B2(n18379), .ZN(n18366) );
  AOI22_X1 U21513 ( .A1(n18443), .A2(n18380), .B1(n18438), .B2(n18405), .ZN(
        n18365) );
  OAI211_X1 U21514 ( .C1(n18446), .C2(n18384), .A(n18366), .B(n18365), .ZN(
        P3_U2964) );
  AOI22_X1 U21515 ( .A1(n18448), .A2(n18380), .B1(n18447), .B2(n18379), .ZN(
        n18368) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18381), .B1(
        n18449), .B2(n18405), .ZN(n18367) );
  OAI211_X1 U21517 ( .C1(n18452), .C2(n18384), .A(n18368), .B(n18367), .ZN(
        P3_U2965) );
  AOI22_X1 U21518 ( .A1(n18454), .A2(n18405), .B1(n18453), .B2(n18379), .ZN(
        n18370) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18381), .B1(
        n18455), .B2(n18380), .ZN(n18369) );
  OAI211_X1 U21520 ( .C1(n18458), .C2(n18384), .A(n18370), .B(n18369), .ZN(
        P3_U2966) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18381), .B1(
        n18459), .B2(n18379), .ZN(n18372) );
  AOI22_X1 U21522 ( .A1(n18460), .A2(n18380), .B1(n18461), .B2(n18405), .ZN(
        n18371) );
  OAI211_X1 U21523 ( .C1(n18464), .C2(n18384), .A(n18372), .B(n18371), .ZN(
        P3_U2967) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18381), .B1(
        n18465), .B2(n18379), .ZN(n18374) );
  AOI22_X1 U21525 ( .A1(n18467), .A2(n18380), .B1(n18466), .B2(n18405), .ZN(
        n18373) );
  OAI211_X1 U21526 ( .C1(n18470), .C2(n18384), .A(n18374), .B(n18373), .ZN(
        P3_U2968) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18381), .B1(
        n18472), .B2(n18379), .ZN(n18376) );
  AOI22_X1 U21528 ( .A1(n18473), .A2(n18405), .B1(n18471), .B2(n18380), .ZN(
        n18375) );
  OAI211_X1 U21529 ( .C1(n18476), .C2(n18384), .A(n18376), .B(n18375), .ZN(
        P3_U2969) );
  AOI22_X1 U21530 ( .A1(n18479), .A2(n18380), .B1(n18477), .B2(n18379), .ZN(
        n18378) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18381), .B1(
        n18478), .B2(n18405), .ZN(n18377) );
  OAI211_X1 U21532 ( .C1(n18482), .C2(n18384), .A(n18378), .B(n18377), .ZN(
        P3_U2970) );
  AOI22_X1 U21533 ( .A1(n18487), .A2(n18405), .B1(n18484), .B2(n18379), .ZN(
        n18383) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18381), .B1(
        n18486), .B2(n18380), .ZN(n18382) );
  OAI211_X1 U21535 ( .C1(n18492), .C2(n18384), .A(n18383), .B(n18382), .ZN(
        P3_U2971) );
  INV_X1 U21536 ( .A(n18488), .ZN(n18409) );
  NOR2_X1 U21537 ( .A1(n18410), .A2(n18385), .ZN(n18404) );
  AOI22_X1 U21538 ( .A1(n18443), .A2(n18405), .B1(n18437), .B2(n18404), .ZN(
        n18391) );
  NOR2_X1 U21539 ( .A1(n18536), .A2(n18386), .ZN(n18389) );
  AOI22_X1 U21540 ( .A1(n18442), .A2(n18389), .B1(n18388), .B2(n18387), .ZN(
        n18406) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18406), .B1(
        n18438), .B2(n18431), .ZN(n18390) );
  OAI211_X1 U21542 ( .C1(n18409), .C2(n18446), .A(n18391), .B(n18390), .ZN(
        P3_U2972) );
  AOI22_X1 U21543 ( .A1(n18449), .A2(n18431), .B1(n18447), .B2(n18404), .ZN(
        n18393) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18406), .B1(
        n18448), .B2(n18405), .ZN(n18392) );
  OAI211_X1 U21545 ( .C1(n18409), .C2(n18452), .A(n18393), .B(n18392), .ZN(
        P3_U2973) );
  AOI22_X1 U21546 ( .A1(n18454), .A2(n18431), .B1(n18453), .B2(n18404), .ZN(
        n18395) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18406), .B1(
        n18455), .B2(n18405), .ZN(n18394) );
  OAI211_X1 U21548 ( .C1(n18409), .C2(n18458), .A(n18395), .B(n18394), .ZN(
        P3_U2974) );
  AOI22_X1 U21549 ( .A1(n18460), .A2(n18405), .B1(n18459), .B2(n18404), .ZN(
        n18397) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18406), .B1(
        n18461), .B2(n18431), .ZN(n18396) );
  OAI211_X1 U21551 ( .C1(n18409), .C2(n18464), .A(n18397), .B(n18396), .ZN(
        P3_U2975) );
  AOI22_X1 U21552 ( .A1(n18466), .A2(n18431), .B1(n18465), .B2(n18404), .ZN(
        n18399) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18406), .B1(
        n18467), .B2(n18405), .ZN(n18398) );
  OAI211_X1 U21554 ( .C1(n18409), .C2(n18470), .A(n18399), .B(n18398), .ZN(
        P3_U2976) );
  AOI22_X1 U21555 ( .A1(n18473), .A2(n18431), .B1(n18472), .B2(n18404), .ZN(
        n18401) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18406), .B1(
        n18471), .B2(n18405), .ZN(n18400) );
  OAI211_X1 U21557 ( .C1(n18409), .C2(n18476), .A(n18401), .B(n18400), .ZN(
        P3_U2977) );
  AOI22_X1 U21558 ( .A1(n18477), .A2(n18404), .B1(n18478), .B2(n18431), .ZN(
        n18403) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18406), .B1(
        n18479), .B2(n18405), .ZN(n18402) );
  OAI211_X1 U21560 ( .C1(n18409), .C2(n18482), .A(n18403), .B(n18402), .ZN(
        P3_U2978) );
  AOI22_X1 U21561 ( .A1(n18486), .A2(n18405), .B1(n18484), .B2(n18404), .ZN(
        n18408) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18406), .B1(
        n18487), .B2(n18431), .ZN(n18407) );
  OAI211_X1 U21563 ( .C1(n18409), .C2(n18492), .A(n18408), .B(n18407), .ZN(
        P3_U2979) );
  NOR2_X1 U21564 ( .A1(n18410), .A2(n18411), .ZN(n18430) );
  AOI22_X1 U21565 ( .A1(n18443), .A2(n18431), .B1(n18437), .B2(n18430), .ZN(
        n18417) );
  OAI21_X1 U21566 ( .B1(n18413), .B2(n18412), .A(n18411), .ZN(n18415) );
  NAND2_X1 U21567 ( .A1(n18415), .A2(n18414), .ZN(n18432) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18432), .B1(
        n18438), .B2(n18485), .ZN(n18416) );
  OAI211_X1 U21569 ( .C1(n18446), .C2(n18435), .A(n18417), .B(n18416), .ZN(
        P3_U2980) );
  AOI22_X1 U21570 ( .A1(n18448), .A2(n18431), .B1(n18447), .B2(n18430), .ZN(
        n18419) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18432), .B1(
        n18449), .B2(n18485), .ZN(n18418) );
  OAI211_X1 U21572 ( .C1(n18435), .C2(n18452), .A(n18419), .B(n18418), .ZN(
        P3_U2981) );
  AOI22_X1 U21573 ( .A1(n18455), .A2(n18431), .B1(n18453), .B2(n18430), .ZN(
        n18421) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18432), .B1(
        n18454), .B2(n18485), .ZN(n18420) );
  OAI211_X1 U21575 ( .C1(n18435), .C2(n18458), .A(n18421), .B(n18420), .ZN(
        P3_U2982) );
  AOI22_X1 U21576 ( .A1(n18460), .A2(n18431), .B1(n18459), .B2(n18430), .ZN(
        n18423) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18432), .B1(
        n18461), .B2(n18485), .ZN(n18422) );
  OAI211_X1 U21578 ( .C1(n18435), .C2(n18464), .A(n18423), .B(n18422), .ZN(
        P3_U2983) );
  AOI22_X1 U21579 ( .A1(n18467), .A2(n18431), .B1(n18465), .B2(n18430), .ZN(
        n18425) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18432), .B1(
        n18466), .B2(n18485), .ZN(n18424) );
  OAI211_X1 U21581 ( .C1(n18435), .C2(n18470), .A(n18425), .B(n18424), .ZN(
        P3_U2984) );
  AOI22_X1 U21582 ( .A1(n18473), .A2(n18485), .B1(n18472), .B2(n18430), .ZN(
        n18427) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18432), .B1(
        n18471), .B2(n18431), .ZN(n18426) );
  OAI211_X1 U21584 ( .C1(n18435), .C2(n18476), .A(n18427), .B(n18426), .ZN(
        P3_U2985) );
  AOI22_X1 U21585 ( .A1(n18477), .A2(n18430), .B1(n18478), .B2(n18485), .ZN(
        n18429) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18432), .B1(
        n18479), .B2(n18431), .ZN(n18428) );
  OAI211_X1 U21587 ( .C1(n18435), .C2(n18482), .A(n18429), .B(n18428), .ZN(
        P3_U2986) );
  AOI22_X1 U21588 ( .A1(n18487), .A2(n18485), .B1(n18484), .B2(n18430), .ZN(
        n18434) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18432), .B1(
        n18486), .B2(n18431), .ZN(n18433) );
  OAI211_X1 U21590 ( .C1(n18435), .C2(n18492), .A(n18434), .B(n18433), .ZN(
        P3_U2987) );
  INV_X1 U21591 ( .A(n18436), .ZN(n18493) );
  AND2_X1 U21592 ( .A1(n18560), .A2(n18439), .ZN(n18483) );
  AOI22_X1 U21593 ( .A1(n18488), .A2(n18438), .B1(n18437), .B2(n18483), .ZN(
        n18445) );
  AOI22_X1 U21594 ( .A1(n18442), .A2(n18441), .B1(n18440), .B2(n18439), .ZN(
        n18489) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18489), .B1(
        n18443), .B2(n18485), .ZN(n18444) );
  OAI211_X1 U21596 ( .C1(n18493), .C2(n18446), .A(n18445), .B(n18444), .ZN(
        P3_U2988) );
  AOI22_X1 U21597 ( .A1(n18448), .A2(n18485), .B1(n18447), .B2(n18483), .ZN(
        n18451) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18489), .B1(
        n18488), .B2(n18449), .ZN(n18450) );
  OAI211_X1 U21599 ( .C1(n18493), .C2(n18452), .A(n18451), .B(n18450), .ZN(
        P3_U2989) );
  AOI22_X1 U21600 ( .A1(n18488), .A2(n18454), .B1(n18453), .B2(n18483), .ZN(
        n18457) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18489), .B1(
        n18455), .B2(n18485), .ZN(n18456) );
  OAI211_X1 U21602 ( .C1(n18493), .C2(n18458), .A(n18457), .B(n18456), .ZN(
        P3_U2990) );
  AOI22_X1 U21603 ( .A1(n18460), .A2(n18485), .B1(n18459), .B2(n18483), .ZN(
        n18463) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18489), .B1(
        n18488), .B2(n18461), .ZN(n18462) );
  OAI211_X1 U21605 ( .C1(n18493), .C2(n18464), .A(n18463), .B(n18462), .ZN(
        P3_U2991) );
  AOI22_X1 U21606 ( .A1(n18488), .A2(n18466), .B1(n18465), .B2(n18483), .ZN(
        n18469) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18489), .B1(
        n18467), .B2(n18485), .ZN(n18468) );
  OAI211_X1 U21608 ( .C1(n18493), .C2(n18470), .A(n18469), .B(n18468), .ZN(
        P3_U2992) );
  AOI22_X1 U21609 ( .A1(n18472), .A2(n18483), .B1(n18471), .B2(n18485), .ZN(
        n18475) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18489), .B1(
        n18488), .B2(n18473), .ZN(n18474) );
  OAI211_X1 U21611 ( .C1(n18493), .C2(n18476), .A(n18475), .B(n18474), .ZN(
        P3_U2993) );
  AOI22_X1 U21612 ( .A1(n18488), .A2(n18478), .B1(n18477), .B2(n18483), .ZN(
        n18481) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18489), .B1(
        n18479), .B2(n18485), .ZN(n18480) );
  OAI211_X1 U21614 ( .C1(n18493), .C2(n18482), .A(n18481), .B(n18480), .ZN(
        P3_U2994) );
  AOI22_X1 U21615 ( .A1(n18486), .A2(n18485), .B1(n18484), .B2(n18483), .ZN(
        n18491) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18489), .B1(
        n18488), .B2(n18487), .ZN(n18490) );
  OAI211_X1 U21617 ( .C1(n18493), .C2(n18492), .A(n18491), .B(n18490), .ZN(
        P3_U2995) );
  NOR2_X1 U21618 ( .A1(n18506), .A2(n18494), .ZN(n18497) );
  OAI222_X1 U21619 ( .A1(n18500), .A2(n18499), .B1(n18498), .B2(n18497), .C1(
        n18496), .C2(n18495), .ZN(n18701) );
  OAI21_X1 U21620 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18501), .ZN(n18502) );
  OAI211_X1 U21621 ( .C1(n18528), .C2(n18504), .A(n18503), .B(n18502), .ZN(
        n18548) );
  NAND2_X1 U21622 ( .A1(n18675), .A2(n18526), .ZN(n18505) );
  NAND2_X1 U21623 ( .A1(n18531), .A2(n18690), .ZN(n18532) );
  AOI22_X1 U21624 ( .A1(n18506), .A2(n18505), .B1(n18519), .B2(n18532), .ZN(
        n18660) );
  NOR2_X1 U21625 ( .A1(n18539), .A2(n18660), .ZN(n18513) );
  AOI21_X1 U21626 ( .B1(n18509), .B2(n18508), .A(n18507), .ZN(n18515) );
  OAI21_X1 U21627 ( .B1(n18531), .B2(n18519), .A(n18515), .ZN(n18510) );
  AOI22_X1 U21628 ( .A1(n18675), .A2(n18526), .B1(n18511), .B2(n18510), .ZN(
        n18663) );
  NAND2_X1 U21629 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18663), .ZN(
        n18512) );
  OAI22_X1 U21630 ( .A1(n18513), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18539), .B2(n18512), .ZN(n18546) );
  AOI221_X1 U21631 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18515), 
        .C1(n18514), .C2(n18515), .A(n18675), .ZN(n18527) );
  NOR2_X1 U21632 ( .A1(n18516), .A2(n18690), .ZN(n18518) );
  OAI211_X1 U21633 ( .C1(n18518), .C2(n18517), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18675), .ZN(n18523) );
  INV_X1 U21634 ( .A(n18519), .ZN(n18520) );
  OAI211_X1 U21635 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18521), .B(n18520), .ZN(
        n18522) );
  OAI211_X1 U21636 ( .C1(n18673), .C2(n18524), .A(n18523), .B(n18522), .ZN(
        n18525) );
  AOI21_X1 U21637 ( .B1(n18527), .B2(n18526), .A(n18525), .ZN(n18671) );
  AOI22_X1 U21638 ( .A1(n18539), .A2(n18675), .B1(n18671), .B2(n18528), .ZN(
        n18542) );
  NOR2_X1 U21639 ( .A1(n18530), .A2(n18529), .ZN(n18534) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18531), .B1(
        n18534), .B2(n18690), .ZN(n18685) );
  INV_X1 U21641 ( .A(n18532), .ZN(n18533) );
  OAI22_X1 U21642 ( .A1(n18534), .A2(n18676), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18533), .ZN(n18680) );
  AOI222_X1 U21643 ( .A1(n18685), .A2(n18680), .B1(n18685), .B2(n18536), .C1(
        n18680), .C2(n18535), .ZN(n18538) );
  OAI21_X1 U21644 ( .B1(n18539), .B2(n18538), .A(n18537), .ZN(n18541) );
  AND2_X1 U21645 ( .A1(n18542), .A2(n18541), .ZN(n18540) );
  OAI221_X1 U21646 ( .B1(n18542), .B2(n18541), .C1(n21014), .C2(n18540), .A(
        n20939), .ZN(n18545) );
  AOI21_X1 U21647 ( .B1(n20939), .B2(n18543), .A(n18542), .ZN(n18544) );
  AOI222_X1 U21648 ( .A1(n18546), .A2(n18545), .B1(n18546), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18545), .C2(n18544), .ZN(
        n18547) );
  OR4_X1 U21649 ( .A1(n18549), .A2(n18701), .A3(n18548), .A4(n18547), .ZN(
        n18556) );
  AOI211_X1 U21650 ( .C1(n18552), .C2(n18551), .A(n18550), .B(n18556), .ZN(
        n18657) );
  AOI21_X1 U21651 ( .B1(n18709), .B2(n18720), .A(n18657), .ZN(n18561) );
  NOR2_X1 U21652 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18714) );
  NAND2_X1 U21653 ( .A1(n18709), .A2(n18703), .ZN(n18564) );
  INV_X1 U21654 ( .A(n18564), .ZN(n18553) );
  AOI211_X1 U21655 ( .C1(n18686), .C2(n18714), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18553), .ZN(n18554) );
  AOI211_X1 U21656 ( .C1(n18706), .C2(n18556), .A(n18555), .B(n18554), .ZN(
        n18557) );
  OAI221_X1 U21657 ( .B1(n18711), .B2(n18561), .C1(n18711), .C2(n18558), .A(
        n18557), .ZN(P3_U2996) );
  NAND4_X1 U21658 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18709), .A4(n18720), .ZN(n18566) );
  INV_X1 U21659 ( .A(n18559), .ZN(n18562) );
  NAND3_X1 U21660 ( .A1(n18562), .A2(n18561), .A3(n18560), .ZN(n18563) );
  NAND4_X1 U21661 ( .A1(n18565), .A2(n18564), .A3(n18566), .A4(n18563), .ZN(
        P3_U2997) );
  INV_X1 U21662 ( .A(n18566), .ZN(n18568) );
  INV_X1 U21663 ( .A(n18658), .ZN(n18567) );
  NOR4_X1 U21664 ( .A1(n18714), .A2(n18569), .A3(n18568), .A4(n18567), .ZN(
        P3_U2998) );
  AND2_X1 U21665 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18570), .ZN(
        P3_U2999) );
  AND2_X1 U21666 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18570), .ZN(
        P3_U3000) );
  AND2_X1 U21667 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18570), .ZN(
        P3_U3001) );
  AND2_X1 U21668 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18570), .ZN(
        P3_U3002) );
  AND2_X1 U21669 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18570), .ZN(
        P3_U3003) );
  AND2_X1 U21670 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18570), .ZN(
        P3_U3004) );
  AND2_X1 U21671 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18570), .ZN(
        P3_U3005) );
  AND2_X1 U21672 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18570), .ZN(
        P3_U3006) );
  AND2_X1 U21673 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18570), .ZN(
        P3_U3007) );
  AND2_X1 U21674 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18570), .ZN(
        P3_U3008) );
  AND2_X1 U21675 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18570), .ZN(
        P3_U3009) );
  AND2_X1 U21676 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18570), .ZN(
        P3_U3010) );
  AND2_X1 U21677 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18570), .ZN(
        P3_U3011) );
  AND2_X1 U21678 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18570), .ZN(
        P3_U3012) );
  INV_X1 U21679 ( .A(P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n21030) );
  NOR2_X1 U21680 ( .A1(n21030), .A2(n18656), .ZN(P3_U3013) );
  AND2_X1 U21681 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18570), .ZN(
        P3_U3014) );
  INV_X1 U21682 ( .A(P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20844) );
  NOR2_X1 U21683 ( .A1(n20844), .A2(n18656), .ZN(P3_U3015) );
  AND2_X1 U21684 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18570), .ZN(
        P3_U3016) );
  AND2_X1 U21685 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18570), .ZN(
        P3_U3017) );
  AND2_X1 U21686 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18570), .ZN(
        P3_U3018) );
  AND2_X1 U21687 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18570), .ZN(
        P3_U3019) );
  AND2_X1 U21688 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18570), .ZN(
        P3_U3020) );
  AND2_X1 U21689 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18570), .ZN(P3_U3021) );
  AND2_X1 U21690 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18570), .ZN(P3_U3022) );
  AND2_X1 U21691 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18570), .ZN(P3_U3023) );
  AND2_X1 U21692 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18570), .ZN(P3_U3024) );
  AND2_X1 U21693 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18570), .ZN(P3_U3025) );
  AND2_X1 U21694 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18570), .ZN(P3_U3026) );
  AND2_X1 U21695 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18570), .ZN(P3_U3027) );
  AND2_X1 U21696 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18570), .ZN(P3_U3028) );
  INV_X1 U21697 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18716) );
  AOI21_X1 U21698 ( .B1(HOLD), .B2(n18571), .A(n18716), .ZN(n18574) );
  NAND2_X1 U21699 ( .A1(n18709), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18580) );
  INV_X1 U21700 ( .A(n18580), .ZN(n18579) );
  OAI21_X1 U21701 ( .B1(n18579), .B2(n18584), .A(n18586), .ZN(n18573) );
  INV_X1 U21702 ( .A(NA), .ZN(n20986) );
  OR3_X1 U21703 ( .A1(n20986), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18572) );
  OAI211_X1 U21704 ( .C1(n18652), .C2(n18574), .A(n18573), .B(n18572), .ZN(
        P3_U3029) );
  AOI21_X1 U21705 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18575) );
  AOI21_X1 U21706 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18575), .ZN(
        n18576) );
  AOI22_X1 U21707 ( .A1(n18709), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18576), .ZN(n18578) );
  NAND2_X1 U21708 ( .A1(n18578), .A2(n18577), .ZN(P3_U3030) );
  AOI221_X1 U21709 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18584), .C1(n20986), 
        .C2(n18584), .A(n18579), .ZN(n18585) );
  NOR2_X1 U21710 ( .A1(n18586), .A2(n20742), .ZN(n18582) );
  OAI22_X1 U21711 ( .A1(NA), .A2(n18580), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18581) );
  OAI22_X1 U21712 ( .A1(n18582), .A2(n18581), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18583) );
  OAI22_X1 U21713 ( .A1(n18585), .A2(n18586), .B1(n18584), .B2(n18583), .ZN(
        P3_U3031) );
  INV_X1 U21714 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18587) );
  OAI222_X1 U21715 ( .A1(n18639), .A2(n20808), .B1(n18588), .B2(n18652), .C1(
        n18587), .C2(n18636), .ZN(P3_U3032) );
  OAI222_X1 U21716 ( .A1(n18639), .A2(n18591), .B1(n18589), .B2(n18652), .C1(
        n20808), .C2(n18636), .ZN(P3_U3033) );
  OAI222_X1 U21717 ( .A1(n18591), .A2(n18636), .B1(n18590), .B2(n18652), .C1(
        n18592), .C2(n18639), .ZN(P3_U3034) );
  INV_X1 U21718 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18595) );
  OAI222_X1 U21719 ( .A1(n18639), .A2(n18595), .B1(n18593), .B2(n18652), .C1(
        n18592), .C2(n18636), .ZN(P3_U3035) );
  OAI222_X1 U21720 ( .A1(n18595), .A2(n18636), .B1(n18594), .B2(n18652), .C1(
        n18596), .C2(n18639), .ZN(P3_U3036) );
  INV_X1 U21721 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18598) );
  OAI222_X1 U21722 ( .A1(n18639), .A2(n18598), .B1(n18597), .B2(n18652), .C1(
        n18596), .C2(n18636), .ZN(P3_U3037) );
  OAI222_X1 U21723 ( .A1(n18639), .A2(n18601), .B1(n18599), .B2(n18652), .C1(
        n18598), .C2(n18636), .ZN(P3_U3038) );
  OAI222_X1 U21724 ( .A1(n18601), .A2(n18636), .B1(n18600), .B2(n18652), .C1(
        n18602), .C2(n18639), .ZN(P3_U3039) );
  OAI222_X1 U21725 ( .A1(n18639), .A2(n18604), .B1(n18603), .B2(n18652), .C1(
        n18602), .C2(n18636), .ZN(P3_U3040) );
  OAI222_X1 U21726 ( .A1(n18639), .A2(n18606), .B1(n18605), .B2(n18652), .C1(
        n18604), .C2(n18636), .ZN(P3_U3041) );
  OAI222_X1 U21727 ( .A1(n18639), .A2(n20904), .B1(n18607), .B2(n18652), .C1(
        n18606), .C2(n18636), .ZN(P3_U3042) );
  OAI222_X1 U21728 ( .A1(n18639), .A2(n18609), .B1(n18608), .B2(n18652), .C1(
        n20904), .C2(n18636), .ZN(P3_U3043) );
  OAI222_X1 U21729 ( .A1(n18639), .A2(n18612), .B1(n18610), .B2(n18652), .C1(
        n18609), .C2(n18642), .ZN(P3_U3044) );
  OAI222_X1 U21730 ( .A1(n18612), .A2(n18636), .B1(n18611), .B2(n18652), .C1(
        n18613), .C2(n18639), .ZN(P3_U3045) );
  OAI222_X1 U21731 ( .A1(n18639), .A2(n18615), .B1(n18614), .B2(n18652), .C1(
        n18613), .C2(n18642), .ZN(P3_U3046) );
  INV_X1 U21732 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18618) );
  OAI222_X1 U21733 ( .A1(n18639), .A2(n18618), .B1(n18616), .B2(n18652), .C1(
        n18615), .C2(n18642), .ZN(P3_U3047) );
  OAI222_X1 U21734 ( .A1(n18618), .A2(n18636), .B1(n18617), .B2(n18652), .C1(
        n18619), .C2(n18639), .ZN(P3_U3048) );
  INV_X1 U21735 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18622) );
  OAI222_X1 U21736 ( .A1(n18639), .A2(n18622), .B1(n18620), .B2(n18652), .C1(
        n18619), .C2(n18642), .ZN(P3_U3049) );
  OAI222_X1 U21737 ( .A1(n18622), .A2(n18636), .B1(n18621), .B2(n18652), .C1(
        n18623), .C2(n18639), .ZN(P3_U3050) );
  OAI222_X1 U21738 ( .A1(n18639), .A2(n18626), .B1(n18624), .B2(n18652), .C1(
        n18623), .C2(n18642), .ZN(P3_U3051) );
  OAI222_X1 U21739 ( .A1(n18626), .A2(n18636), .B1(n18625), .B2(n18652), .C1(
        n20836), .C2(n18639), .ZN(P3_U3052) );
  OAI222_X1 U21740 ( .A1(n18639), .A2(n18629), .B1(n18627), .B2(n18652), .C1(
        n20836), .C2(n18642), .ZN(P3_U3053) );
  OAI222_X1 U21741 ( .A1(n18629), .A2(n18636), .B1(n18628), .B2(n18652), .C1(
        n18630), .C2(n18639), .ZN(P3_U3054) );
  OAI222_X1 U21742 ( .A1(n18639), .A2(n20842), .B1(n18631), .B2(n18652), .C1(
        n18630), .C2(n18642), .ZN(P3_U3055) );
  INV_X1 U21743 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18633) );
  OAI222_X1 U21744 ( .A1(n18639), .A2(n18633), .B1(n18632), .B2(n18652), .C1(
        n20842), .C2(n18642), .ZN(P3_U3056) );
  OAI222_X1 U21745 ( .A1(n18639), .A2(n18635), .B1(n18634), .B2(n18652), .C1(
        n18633), .C2(n18636), .ZN(P3_U3057) );
  OAI222_X1 U21746 ( .A1(n18642), .A2(n18635), .B1(n20983), .B2(n18652), .C1(
        n18637), .C2(n18639), .ZN(P3_U3058) );
  OAI222_X1 U21747 ( .A1(n18639), .A2(n18640), .B1(n18638), .B2(n18652), .C1(
        n18637), .C2(n18636), .ZN(P3_U3059) );
  OAI222_X1 U21748 ( .A1(n18639), .A2(n18643), .B1(n18641), .B2(n18652), .C1(
        n18640), .C2(n18642), .ZN(P3_U3060) );
  OAI222_X1 U21749 ( .A1(n18639), .A2(n18645), .B1(n18644), .B2(n18652), .C1(
        n18643), .C2(n18642), .ZN(P3_U3061) );
  INV_X1 U21750 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18646) );
  AOI22_X1 U21751 ( .A1(n18652), .A2(n18647), .B1(n18646), .B2(n18718), .ZN(
        P3_U3274) );
  INV_X1 U21752 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18694) );
  INV_X1 U21753 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18648) );
  AOI22_X1 U21754 ( .A1(n18652), .A2(n18694), .B1(n18648), .B2(n18718), .ZN(
        P3_U3275) );
  INV_X1 U21755 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18649) );
  AOI22_X1 U21756 ( .A1(n18652), .A2(n18650), .B1(n18649), .B2(n18718), .ZN(
        P3_U3276) );
  INV_X1 U21757 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18697) );
  INV_X1 U21758 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18651) );
  AOI22_X1 U21759 ( .A1(n18652), .A2(n18697), .B1(n18651), .B2(n18718), .ZN(
        P3_U3277) );
  OAI21_X1 U21760 ( .B1(n18656), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18654), 
        .ZN(n18653) );
  INV_X1 U21761 ( .A(n18653), .ZN(P3_U3280) );
  INV_X1 U21762 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18655) );
  OAI21_X1 U21763 ( .B1(n18656), .B2(n18655), .A(n18654), .ZN(P3_U3281) );
  NOR2_X1 U21764 ( .A1(n18657), .A2(n18711), .ZN(n18659) );
  OAI21_X1 U21765 ( .B1(n18659), .B2(n18684), .A(n18658), .ZN(P3_U3282) );
  NOR3_X1 U21766 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18660), .A3(
        n18670), .ZN(n18661) );
  AOI21_X1 U21767 ( .B1(n18662), .B2(n18686), .A(n18661), .ZN(n18667) );
  INV_X1 U21768 ( .A(n18670), .ZN(n18721) );
  INV_X1 U21769 ( .A(n18663), .ZN(n18664) );
  AOI21_X1 U21770 ( .B1(n18721), .B2(n18664), .A(n18689), .ZN(n18666) );
  OAI22_X1 U21771 ( .A1(n18689), .A2(n18667), .B1(n18666), .B2(n18665), .ZN(
        P3_U3285) );
  NAND2_X1 U21772 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18683) );
  INV_X1 U21773 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18669) );
  AOI22_X1 U21774 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18669), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n18668), .ZN(n18678) );
  OAI22_X1 U21775 ( .A1(n18671), .A2(n18670), .B1(n18683), .B2(n18678), .ZN(
        n18672) );
  AOI21_X1 U21776 ( .B1(n18686), .B2(n18673), .A(n18672), .ZN(n18674) );
  INV_X1 U21777 ( .A(n18689), .ZN(n18681) );
  AOI22_X1 U21778 ( .A1(n18689), .A2(n18675), .B1(n18674), .B2(n18681), .ZN(
        P3_U3288) );
  INV_X1 U21779 ( .A(n18676), .ZN(n18679) );
  INV_X1 U21780 ( .A(n18683), .ZN(n18677) );
  AOI222_X1 U21781 ( .A1(n18680), .A2(n18721), .B1(n18686), .B2(n18679), .C1(
        n18678), .C2(n18677), .ZN(n18682) );
  AOI22_X1 U21782 ( .A1(n18689), .A2(n11599), .B1(n18682), .B2(n18681), .ZN(
        P3_U3289) );
  OAI221_X1 U21783 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18685), .C1(
        P3_STATE2_REG_1__SCAN_IN), .C2(n18684), .A(n18683), .ZN(n18688) );
  AOI21_X1 U21784 ( .B1(n18690), .B2(n18686), .A(n18689), .ZN(n18687) );
  AOI22_X1 U21785 ( .A1(n18690), .A2(n18689), .B1(n18688), .B2(n18687), .ZN(
        P3_U3290) );
  INV_X1 U21786 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18692) );
  NOR3_X1 U21787 ( .A1(n18692), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18691) );
  AOI221_X1 U21788 ( .B1(n18693), .B2(n18692), .C1(P3_REIP_REG_1__SCAN_IN), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18691), .ZN(n18695) );
  INV_X1 U21789 ( .A(n18699), .ZN(n18696) );
  AOI22_X1 U21790 ( .A1(n18699), .A2(n18695), .B1(n18694), .B2(n18696), .ZN(
        P3_U3292) );
  NOR2_X1 U21791 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18698) );
  AOI22_X1 U21792 ( .A1(n18699), .A2(n18698), .B1(n18697), .B2(n18696), .ZN(
        P3_U3293) );
  INV_X1 U21793 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n20988) );
  AOI22_X1 U21794 ( .A1(n18652), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n20988), 
        .B2(n18718), .ZN(P3_U3294) );
  MUX2_X1 U21795 ( .A(P3_MORE_REG_SCAN_IN), .B(n18701), .S(n18700), .Z(
        P3_U3295) );
  AOI21_X1 U21796 ( .B1(n18703), .B2(n18702), .A(n18723), .ZN(n18704) );
  OAI21_X1 U21797 ( .B1(n18706), .B2(n18705), .A(n18704), .ZN(n18717) );
  OAI21_X1 U21798 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18708), .A(n18707), 
        .ZN(n18710) );
  AOI211_X1 U21799 ( .C1(n18722), .C2(n18710), .A(n18709), .B(n18720), .ZN(
        n18712) );
  NOR2_X1 U21800 ( .A1(n18712), .A2(n18711), .ZN(n18713) );
  OAI21_X1 U21801 ( .B1(n18714), .B2(n18713), .A(n18717), .ZN(n18715) );
  OAI21_X1 U21802 ( .B1(n18717), .B2(n18716), .A(n18715), .ZN(P3_U3296) );
  INV_X1 U21803 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18726) );
  INV_X1 U21804 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18719) );
  AOI22_X1 U21805 ( .A1(n18652), .A2(n18726), .B1(n18719), .B2(n18718), .ZN(
        P3_U3297) );
  AOI21_X1 U21806 ( .B1(n18721), .B2(n18720), .A(n18723), .ZN(n18727) );
  INV_X1 U21807 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18724) );
  AOI22_X1 U21808 ( .A1(n18727), .A2(n18724), .B1(n18723), .B2(n18722), .ZN(
        P3_U3298) );
  AOI21_X1 U21809 ( .B1(n18727), .B2(n18726), .A(n18725), .ZN(P3_U3299) );
  INV_X1 U21810 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18728) );
  INV_X1 U21811 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19694) );
  NAND2_X1 U21812 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19694), .ZN(n19687) );
  OR2_X1 U21813 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19688) );
  OAI21_X1 U21814 ( .B1(n19683), .B2(n19687), .A(n19688), .ZN(n19753) );
  OAI21_X1 U21815 ( .B1(n19683), .B2(n18728), .A(n19679), .ZN(P2_U2815) );
  AOI22_X1 U21816 ( .A1(P2_CODEFETCH_REG_SCAN_IN), .A2(n18730), .B1(n18729), 
        .B2(n19390), .ZN(n18731) );
  INV_X1 U21817 ( .A(n18731), .ZN(P2_U2816) );
  AOI22_X1 U21818 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19806), .B1(n20741), .B2(
        n19683), .ZN(n18732) );
  OAI21_X1 U21819 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19806), .A(n18732), 
        .ZN(P2_U2817) );
  OAI21_X1 U21820 ( .B1(n20741), .B2(BS16), .A(n19753), .ZN(n19751) );
  OAI21_X1 U21821 ( .B1(n19753), .B2(n19574), .A(n19751), .ZN(P2_U2818) );
  INV_X1 U21822 ( .A(n18733), .ZN(n18735) );
  NOR2_X1 U21823 ( .A1(n18735), .A2(n18734), .ZN(n19805) );
  OAI21_X1 U21824 ( .B1(n19805), .B2(n12706), .A(n18736), .ZN(P2_U2819) );
  NOR4_X1 U21825 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n18746) );
  NOR4_X1 U21826 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18745) );
  AOI211_X1 U21827 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18737) );
  INV_X1 U21828 ( .A(P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20911) );
  INV_X1 U21829 ( .A(P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20910) );
  NAND3_X1 U21830 ( .A1(n18737), .A2(n20911), .A3(n20910), .ZN(n18743) );
  NOR4_X1 U21831 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_18__SCAN_IN), .A3(P2_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18741) );
  NOR4_X1 U21832 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_14__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n18740) );
  NOR4_X1 U21833 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18739) );
  NOR4_X1 U21834 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18738) );
  NAND4_X1 U21835 ( .A1(n18741), .A2(n18740), .A3(n18739), .A4(n18738), .ZN(
        n18742) );
  NOR4_X1 U21836 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_31__SCAN_IN), .A3(n18743), .A4(n18742), .ZN(n18744)
         );
  NAND3_X1 U21837 ( .A1(n18746), .A2(n18745), .A3(n18744), .ZN(n18752) );
  NOR2_X1 U21838 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18752), .ZN(n18747) );
  INV_X1 U21839 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U21840 ( .A1(n18747), .A2(n11908), .B1(n18752), .B2(n19749), .ZN(
        P2_U2820) );
  OR3_X1 U21841 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18751) );
  INV_X1 U21842 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U21843 ( .A1(n18747), .A2(n18751), .B1(n18752), .B2(n19747), .ZN(
        P2_U2821) );
  INV_X1 U21844 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19752) );
  NAND2_X1 U21845 ( .A1(n18747), .A2(n19752), .ZN(n18750) );
  INV_X1 U21846 ( .A(n18752), .ZN(n18753) );
  OAI21_X1 U21847 ( .B1(n11908), .B2(n19696), .A(n18753), .ZN(n18748) );
  OAI21_X1 U21848 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18753), .A(n18748), 
        .ZN(n18749) );
  OAI221_X1 U21849 ( .B1(n18750), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18750), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18749), .ZN(P2_U2822) );
  INV_X1 U21850 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19745) );
  OAI221_X1 U21851 ( .B1(n18753), .B2(n19745), .C1(n18752), .C2(n18751), .A(
        n18750), .ZN(P2_U2823) );
  AOI22_X1 U21852 ( .A1(n18950), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18949), .ZN(n18765) );
  AOI22_X1 U21853 ( .A1(n18754), .A2(n18954), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18928), .ZN(n18764) );
  AOI22_X1 U21854 ( .A1(n18756), .A2(n18939), .B1(n18952), .B2(n18755), .ZN(
        n18763) );
  INV_X1 U21855 ( .A(n18757), .ZN(n18761) );
  NOR2_X1 U21856 ( .A1(n18941), .A2(n18758), .ZN(n18760) );
  AOI21_X1 U21857 ( .B1(n18761), .B2(n18760), .A(n18967), .ZN(n18759) );
  OAI21_X1 U21858 ( .B1(n18761), .B2(n18760), .A(n18759), .ZN(n18762) );
  NAND4_X1 U21859 ( .A1(n18765), .A2(n18764), .A3(n18763), .A4(n18762), .ZN(
        P2_U2835) );
  NAND2_X1 U21860 ( .A1(n18912), .A2(n18766), .ZN(n18767) );
  XOR2_X1 U21861 ( .A(n18768), .B(n18767), .Z(n18778) );
  NAND2_X1 U21862 ( .A1(n18950), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n18770) );
  AOI21_X1 U21863 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18928), .A(
        n18885), .ZN(n18769) );
  OAI211_X1 U21864 ( .C1(n18926), .C2(n19719), .A(n18770), .B(n18769), .ZN(
        n18771) );
  AOI21_X1 U21865 ( .B1(n18772), .B2(n18954), .A(n18771), .ZN(n18777) );
  INV_X1 U21866 ( .A(n18773), .ZN(n18775) );
  AOI22_X1 U21867 ( .A1(n18775), .A2(n18939), .B1(n18774), .B2(n18952), .ZN(
        n18776) );
  OAI211_X1 U21868 ( .C1(n18967), .C2(n18778), .A(n18777), .B(n18776), .ZN(
        P2_U2836) );
  NOR2_X1 U21869 ( .A1(n18941), .A2(n18801), .ZN(n18780) );
  XOR2_X1 U21870 ( .A(n18780), .B(n18779), .Z(n18791) );
  NOR2_X1 U21871 ( .A1(n18926), .A2(n19717), .ZN(n18781) );
  AOI211_X1 U21872 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18928), .A(
        n18885), .B(n18781), .ZN(n18782) );
  OAI21_X1 U21873 ( .B1(n18783), .B2(n18925), .A(n18782), .ZN(n18784) );
  AOI21_X1 U21874 ( .B1(n18785), .B2(n18954), .A(n18784), .ZN(n18790) );
  OAI22_X1 U21875 ( .A1(n18787), .A2(n18957), .B1(n18786), .B2(n18920), .ZN(
        n18788) );
  INV_X1 U21876 ( .A(n18788), .ZN(n18789) );
  OAI211_X1 U21877 ( .C1(n18967), .C2(n18791), .A(n18790), .B(n18789), .ZN(
        P2_U2837) );
  NAND2_X1 U21878 ( .A1(n18803), .A2(n18840), .ZN(n18792) );
  OAI211_X1 U21879 ( .C1(n18793), .C2(n18961), .A(n18792), .B(n18905), .ZN(
        n18796) );
  NOR2_X1 U21880 ( .A1(n18925), .A2(n18794), .ZN(n18795) );
  AOI211_X1 U21881 ( .C1(n18949), .C2(P2_REIP_REG_17__SCAN_IN), .A(n18796), 
        .B(n18795), .ZN(n18797) );
  OAI21_X1 U21882 ( .B1(n18798), .B2(n18957), .A(n18797), .ZN(n18799) );
  AOI21_X1 U21883 ( .B1(n9843), .B2(n18954), .A(n18799), .ZN(n18807) );
  AOI211_X1 U21884 ( .C1(n18803), .C2(n18802), .A(n18801), .B(n18800), .ZN(
        n18804) );
  AOI21_X1 U21885 ( .B1(n18952), .B2(n18805), .A(n18804), .ZN(n18806) );
  NAND2_X1 U21886 ( .A1(n18807), .A2(n18806), .ZN(P2_U2838) );
  NAND2_X1 U21887 ( .A1(n18912), .A2(n18808), .ZN(n18809) );
  XOR2_X1 U21888 ( .A(n18810), .B(n18809), .Z(n18820) );
  OAI21_X1 U21889 ( .B1(n18925), .B2(n18811), .A(n18905), .ZN(n18815) );
  OAI22_X1 U21890 ( .A1(n18813), .A2(n18907), .B1(n18812), .B2(n18961), .ZN(
        n18814) );
  AOI211_X1 U21891 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18949), .A(n18815), 
        .B(n18814), .ZN(n18819) );
  INV_X1 U21892 ( .A(n18816), .ZN(n19013) );
  AOI22_X1 U21893 ( .A1(n18817), .A2(n18939), .B1(n18952), .B2(n19013), .ZN(
        n18818) );
  OAI211_X1 U21894 ( .C1(n18967), .C2(n18820), .A(n18819), .B(n18818), .ZN(
        P2_U2840) );
  OR2_X1 U21895 ( .A1(n18941), .A2(n18821), .ZN(n18832) );
  XNOR2_X1 U21896 ( .A(n18832), .B(n18822), .ZN(n18831) );
  AOI22_X1 U21897 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n18949), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18928), .ZN(n18823) );
  OAI211_X1 U21898 ( .C1(n18925), .C2(n18824), .A(n18823), .B(n18905), .ZN(
        n18825) );
  AOI21_X1 U21899 ( .B1(n18826), .B2(n18954), .A(n18825), .ZN(n18830) );
  OAI22_X1 U21900 ( .A1(n18976), .A2(n18957), .B1(n18827), .B2(n18920), .ZN(
        n18828) );
  INV_X1 U21901 ( .A(n18828), .ZN(n18829) );
  OAI211_X1 U21902 ( .C1(n18967), .C2(n18831), .A(n18830), .B(n18829), .ZN(
        P2_U2841) );
  AOI211_X1 U21903 ( .C1(n18841), .C2(n18833), .A(n18967), .B(n18832), .ZN(
        n18839) );
  OAI21_X1 U21904 ( .B1(n18926), .B2(n18834), .A(n18905), .ZN(n18835) );
  AOI21_X1 U21905 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(n18950), .A(n18835), .ZN(
        n18836) );
  OAI21_X1 U21906 ( .B1(n18837), .B2(n18907), .A(n18836), .ZN(n18838) );
  AOI211_X1 U21907 ( .C1(n18928), .C2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n18839), .B(n18838), .ZN(n18844) );
  AOI22_X1 U21908 ( .A1(n18842), .A2(n18939), .B1(n18841), .B2(n18840), .ZN(
        n18843) );
  OAI211_X1 U21909 ( .C1(n18845), .C2(n18920), .A(n18844), .B(n18843), .ZN(
        P2_U2842) );
  INV_X1 U21910 ( .A(n18846), .ZN(n18850) );
  INV_X1 U21911 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n18848) );
  NAND2_X1 U21912 ( .A1(n18949), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n18847) );
  OAI211_X1 U21913 ( .C1(n18925), .C2(n18848), .A(n18905), .B(n18847), .ZN(
        n18849) );
  AOI21_X1 U21914 ( .B1(n18850), .B2(n18954), .A(n18849), .ZN(n18856) );
  XOR2_X1 U21915 ( .A(n18852), .B(n18851), .Z(n18854) );
  OAI22_X1 U21916 ( .A1(n19018), .A2(n18920), .B1(n18983), .B2(n18957), .ZN(
        n18853) );
  AOI21_X1 U21917 ( .B1(n18854), .B2(n18916), .A(n18853), .ZN(n18855) );
  OAI211_X1 U21918 ( .C1(n10028), .C2(n18961), .A(n18856), .B(n18855), .ZN(
        P2_U2843) );
  NOR2_X1 U21919 ( .A1(n18941), .A2(n18857), .ZN(n18858) );
  XOR2_X1 U21920 ( .A(n18859), .B(n18858), .Z(n18866) );
  NOR2_X1 U21921 ( .A1(n18925), .A2(n12743), .ZN(n18860) );
  AOI211_X1 U21922 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18928), .A(
        n18885), .B(n18860), .ZN(n18861) );
  OAI21_X1 U21923 ( .B1(n18862), .B2(n18907), .A(n18861), .ZN(n18864) );
  OAI22_X1 U21924 ( .A1(n18985), .A2(n18957), .B1(n19022), .B2(n18920), .ZN(
        n18863) );
  AOI211_X1 U21925 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n18949), .A(n18864), 
        .B(n18863), .ZN(n18865) );
  OAI21_X1 U21926 ( .B1(n18967), .B2(n18866), .A(n18865), .ZN(P2_U2845) );
  OAI21_X1 U21927 ( .B1(n18925), .B2(n18867), .A(n18905), .ZN(n18872) );
  INV_X1 U21928 ( .A(n18868), .ZN(n18870) );
  OAI22_X1 U21929 ( .A1(n18870), .A2(n18907), .B1(n18869), .B2(n18961), .ZN(
        n18871) );
  AOI211_X1 U21930 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18949), .A(n18872), .B(
        n18871), .ZN(n18879) );
  NAND2_X1 U21931 ( .A1(n18912), .A2(n18873), .ZN(n18874) );
  XNOR2_X1 U21932 ( .A(n18875), .B(n18874), .ZN(n18877) );
  AOI22_X1 U21933 ( .A1(n18877), .A2(n18916), .B1(n18876), .B2(n18939), .ZN(
        n18878) );
  OAI211_X1 U21934 ( .C1(n18880), .C2(n18920), .A(n18879), .B(n18878), .ZN(
        P2_U2846) );
  NAND2_X1 U21935 ( .A1(n18912), .A2(n18881), .ZN(n18883) );
  XOR2_X1 U21936 ( .A(n18883), .B(n18882), .Z(n18893) );
  NOR2_X1 U21937 ( .A1(n18925), .A2(n13047), .ZN(n18884) );
  AOI211_X1 U21938 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18928), .A(
        n18885), .B(n18884), .ZN(n18886) );
  OAI21_X1 U21939 ( .B1(n18887), .B2(n18907), .A(n18886), .ZN(n18891) );
  OAI22_X1 U21940 ( .A1(n18889), .A2(n18957), .B1(n18920), .B2(n18888), .ZN(
        n18890) );
  AOI211_X1 U21941 ( .C1(P2_REIP_REG_7__SCAN_IN), .C2(n18949), .A(n18891), .B(
        n18890), .ZN(n18892) );
  OAI21_X1 U21942 ( .B1(n18893), .B2(n18967), .A(n18892), .ZN(P2_U2848) );
  OAI21_X1 U21943 ( .B1(n18925), .B2(n18894), .A(n18905), .ZN(n18897) );
  OAI22_X1 U21944 ( .A1(n18895), .A2(n18907), .B1(n19702), .B2(n18926), .ZN(
        n18896) );
  AOI211_X1 U21945 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18928), .A(
        n18897), .B(n18896), .ZN(n18903) );
  NOR2_X1 U21946 ( .A1(n18941), .A2(n18898), .ZN(n18900) );
  XNOR2_X1 U21947 ( .A(n18900), .B(n18899), .ZN(n18901) );
  AOI22_X1 U21948 ( .A1(n18901), .A2(n18916), .B1(n9894), .B2(n18939), .ZN(
        n18902) );
  OAI211_X1 U21949 ( .C1(n18920), .C2(n18904), .A(n18903), .B(n18902), .ZN(
        P2_U2849) );
  OAI21_X1 U21950 ( .B1(n18925), .B2(n12502), .A(n18905), .ZN(n18910) );
  OAI22_X1 U21951 ( .A1(n18908), .A2(n18907), .B1(n18906), .B2(n18961), .ZN(
        n18909) );
  AOI211_X1 U21952 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18949), .A(n18910), .B(
        n18909), .ZN(n18919) );
  NAND2_X1 U21953 ( .A1(n18912), .A2(n18911), .ZN(n18913) );
  XNOR2_X1 U21954 ( .A(n18914), .B(n18913), .ZN(n18917) );
  AOI22_X1 U21955 ( .A1(n18917), .A2(n18916), .B1(n18915), .B2(n18939), .ZN(
        n18918) );
  OAI211_X1 U21956 ( .C1(n18920), .C2(n19024), .A(n18919), .B(n18918), .ZN(
        P2_U2850) );
  NAND2_X1 U21957 ( .A1(n18921), .A2(n12962), .ZN(n18924) );
  INV_X1 U21958 ( .A(n18922), .ZN(n18923) );
  AND2_X1 U21959 ( .A1(n18924), .A2(n18923), .ZN(n19125) );
  OAI22_X1 U21960 ( .A1(n18926), .A2(n12179), .B1(n12497), .B2(n18925), .ZN(
        n18927) );
  AOI211_X1 U21961 ( .C1(n18952), .C2(n19125), .A(n19132), .B(n18927), .ZN(
        n18948) );
  AOI22_X1 U21962 ( .A1(n18929), .A2(n18954), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18928), .ZN(n18947) );
  INV_X1 U21963 ( .A(n18930), .ZN(n18931) );
  NAND3_X1 U21964 ( .A1(n18932), .A2(n12937), .A3(n18931), .ZN(n18933) );
  AND2_X1 U21965 ( .A1(n18934), .A2(n18933), .ZN(n19034) );
  NAND2_X1 U21966 ( .A1(n18936), .A2(n18935), .ZN(n18937) );
  AND2_X1 U21967 ( .A1(n18938), .A2(n18937), .ZN(n19122) );
  AOI22_X1 U21968 ( .A1(n19034), .A2(n18964), .B1(n18939), .B2(n19122), .ZN(
        n18946) );
  INV_X1 U21969 ( .A(n19119), .ZN(n18944) );
  NOR2_X1 U21970 ( .A1(n18941), .A2(n18940), .ZN(n18943) );
  AOI21_X1 U21971 ( .B1(n18944), .B2(n18943), .A(n18967), .ZN(n18942) );
  OAI21_X1 U21972 ( .B1(n18944), .B2(n18943), .A(n18942), .ZN(n18945) );
  NAND4_X1 U21973 ( .A1(n18948), .A2(n18947), .A3(n18946), .A4(n18945), .ZN(
        P2_U2851) );
  AOI22_X1 U21974 ( .A1(n18950), .A2(P2_EBX_REG_0__SCAN_IN), .B1(
        P2_REIP_REG_0__SCAN_IN), .B2(n18949), .ZN(n18956) );
  AOI22_X1 U21975 ( .A1(n18954), .A2(n18953), .B1(n18952), .B2(n18951), .ZN(
        n18955) );
  OAI211_X1 U21976 ( .C1(n18958), .C2(n18957), .A(n18956), .B(n18955), .ZN(
        n18963) );
  AOI21_X1 U21977 ( .B1(n18961), .B2(n18960), .A(n18959), .ZN(n18962) );
  AOI211_X1 U21978 ( .C1(n18964), .C2(n19791), .A(n18963), .B(n18962), .ZN(
        n18965) );
  OAI21_X1 U21979 ( .B1(n18967), .B2(n18966), .A(n18965), .ZN(P2_U2855) );
  INV_X1 U21980 ( .A(n18968), .ZN(n18969) );
  AOI21_X1 U21981 ( .B1(n18970), .B2(n13722), .A(n18969), .ZN(n19009) );
  AOI22_X1 U21982 ( .A1(n19009), .A2(n18998), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n18996), .ZN(n18971) );
  OAI21_X1 U21983 ( .B1(n18996), .B2(n18972), .A(n18971), .ZN(P2_U2871) );
  XOR2_X1 U21984 ( .A(n12993), .B(n18973), .Z(n18974) );
  AOI22_X1 U21985 ( .A1(n18974), .A2(n18998), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n18996), .ZN(n18975) );
  OAI21_X1 U21986 ( .B1(n18976), .B2(n18996), .A(n18975), .ZN(P2_U2873) );
  AOI21_X1 U21987 ( .B1(n18986), .B2(n18978), .A(n18977), .ZN(n18979) );
  NOR3_X1 U21988 ( .A1(n18980), .A2(n18979), .A3(n18992), .ZN(n18981) );
  AOI21_X1 U21989 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n18996), .A(n18981), .ZN(
        n18982) );
  OAI21_X1 U21990 ( .B1(n18983), .B2(n18996), .A(n18982), .ZN(P2_U2875) );
  OAI21_X1 U21991 ( .B1(n12730), .B2(n18984), .A(n18998), .ZN(n18987) );
  OAI22_X1 U21992 ( .A1(n18987), .A2(n18986), .B1(n18985), .B2(n18996), .ZN(
        n18988) );
  INV_X1 U21993 ( .A(n18988), .ZN(n18989) );
  OAI21_X1 U21994 ( .B1(n19000), .B2(n12743), .A(n18989), .ZN(P2_U2877) );
  AOI21_X1 U21995 ( .B1(n18991), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n18990), .ZN(n18993) );
  NOR3_X1 U21996 ( .A1(n18993), .A2(n9826), .A3(n18992), .ZN(n18994) );
  AOI21_X1 U21997 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n18996), .A(n18994), .ZN(
        n18995) );
  OAI21_X1 U21998 ( .B1(n18997), .B2(n18996), .A(n18995), .ZN(P2_U2879) );
  AOI22_X1 U21999 ( .A1(n19034), .A2(n18998), .B1(n19000), .B2(n19122), .ZN(
        n18999) );
  OAI21_X1 U22000 ( .B1(n19000), .B2(n12497), .A(n18999), .ZN(P2_U2883) );
  AOI22_X1 U22001 ( .A1(n19001), .A2(n19057), .B1(n19007), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19003) );
  AOI22_X1 U22002 ( .A1(n19006), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19056), .ZN(n19002) );
  NAND2_X1 U22003 ( .A1(n19003), .A2(n19002), .ZN(P2_U2888) );
  AOI22_X1 U22004 ( .A1(n19005), .A2(n19004), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19056), .ZN(n19012) );
  AOI22_X1 U22005 ( .A1(n19007), .A2(BUF1_REG_16__SCAN_IN), .B1(n19006), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19011) );
  AOI22_X1 U22006 ( .A1(n19009), .A2(n19038), .B1(n19057), .B2(n19008), .ZN(
        n19010) );
  NAND3_X1 U22007 ( .A1(n19012), .A2(n19011), .A3(n19010), .ZN(P2_U2903) );
  AOI22_X1 U22008 ( .A1(n19025), .A2(n19013), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n19056), .ZN(n19014) );
  OAI21_X1 U22009 ( .B1(n19065), .B2(n19015), .A(n19014), .ZN(P2_U2904) );
  AOI22_X1 U22010 ( .A1(n19020), .A2(n19016), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19056), .ZN(n19017) );
  OAI21_X1 U22011 ( .B1(n19023), .B2(n19018), .A(n19017), .ZN(P2_U2907) );
  AOI22_X1 U22012 ( .A1(n19020), .A2(n19019), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19056), .ZN(n19021) );
  OAI21_X1 U22013 ( .B1(n19023), .B2(n19022), .A(n19021), .ZN(P2_U2909) );
  NAND2_X1 U22014 ( .A1(n19034), .A2(n19125), .ZN(n19037) );
  OAI21_X1 U22015 ( .B1(n19037), .B2(n19061), .A(n19024), .ZN(n19026) );
  AOI22_X1 U22016 ( .A1(n19026), .A2(n19025), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19056), .ZN(n19027) );
  OAI21_X1 U22017 ( .B1(n19166), .B2(n19065), .A(n19027), .ZN(P2_U2914) );
  INV_X1 U22018 ( .A(n19028), .ZN(n19163) );
  AOI22_X1 U22019 ( .A1(n19057), .A2(n19125), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19056), .ZN(n19042) );
  INV_X1 U22020 ( .A(n19775), .ZN(n19032) );
  INV_X1 U22021 ( .A(n19785), .ZN(n19031) );
  XNOR2_X1 U22022 ( .A(n19783), .B(n19785), .ZN(n19059) );
  NOR2_X1 U22023 ( .A1(n19030), .A2(n19029), .ZN(n19060) );
  NOR2_X1 U22024 ( .A1(n19059), .A2(n19060), .ZN(n19058) );
  AOI21_X1 U22025 ( .B1(n19031), .B2(n19780), .A(n19058), .ZN(n19050) );
  XOR2_X1 U22026 ( .A(n19775), .B(n19772), .Z(n19051) );
  NOR2_X1 U22027 ( .A1(n19050), .A2(n19051), .ZN(n19049) );
  AOI21_X1 U22028 ( .B1(n19032), .B2(n19772), .A(n19049), .ZN(n19044) );
  XNOR2_X1 U22029 ( .A(n19423), .B(n19033), .ZN(n19045) );
  NOR2_X1 U22030 ( .A1(n19044), .A2(n19045), .ZN(n19043) );
  AOI21_X1 U22031 ( .B1(n19423), .B2(n19033), .A(n19043), .ZN(n19040) );
  INV_X1 U22032 ( .A(n19034), .ZN(n19036) );
  INV_X1 U22033 ( .A(n19125), .ZN(n19035) );
  NAND2_X1 U22034 ( .A1(n19036), .A2(n19035), .ZN(n19039) );
  OAI211_X1 U22035 ( .C1(n19040), .C2(n19039), .A(n19038), .B(n19037), .ZN(
        n19041) );
  OAI211_X1 U22036 ( .C1(n19163), .C2(n19065), .A(n19042), .B(n19041), .ZN(
        P2_U2915) );
  AOI22_X1 U22037 ( .A1(n19057), .A2(n19767), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19056), .ZN(n19048) );
  AOI21_X1 U22038 ( .B1(n19045), .B2(n19044), .A(n19043), .ZN(n19046) );
  OR2_X1 U22039 ( .A1(n19046), .A2(n19061), .ZN(n19047) );
  OAI211_X1 U22040 ( .C1(n19158), .C2(n19065), .A(n19048), .B(n19047), .ZN(
        P2_U2916) );
  AOI22_X1 U22041 ( .A1(n19775), .A2(n19057), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19056), .ZN(n19054) );
  AOI21_X1 U22042 ( .B1(n19051), .B2(n19050), .A(n19049), .ZN(n19052) );
  OR2_X1 U22043 ( .A1(n19052), .A2(n19061), .ZN(n19053) );
  OAI211_X1 U22044 ( .C1(n19055), .C2(n19065), .A(n19054), .B(n19053), .ZN(
        P2_U2917) );
  AOI22_X1 U22045 ( .A1(n19057), .A2(n19785), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19056), .ZN(n19064) );
  AOI21_X1 U22046 ( .B1(n19060), .B2(n19059), .A(n19058), .ZN(n19062) );
  OR2_X1 U22047 ( .A1(n19062), .A2(n19061), .ZN(n19063) );
  OAI211_X1 U22048 ( .C1(n19150), .C2(n19065), .A(n19064), .B(n19063), .ZN(
        P2_U2918) );
  NOR2_X1 U22049 ( .A1(n19091), .A2(n19066), .ZN(P2_U2920) );
  INV_X1 U22050 ( .A(n19089), .ZN(n19099) );
  AOI22_X1 U22051 ( .A1(n19097), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19067) );
  OAI21_X1 U22052 ( .B1(n11883), .B2(n19099), .A(n19067), .ZN(P2_U2936) );
  AOI22_X1 U22053 ( .A1(n19097), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19068) );
  OAI21_X1 U22054 ( .B1(n19069), .B2(n19099), .A(n19068), .ZN(P2_U2937) );
  AOI22_X1 U22055 ( .A1(n19097), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19070) );
  OAI21_X1 U22056 ( .B1(n19071), .B2(n19099), .A(n19070), .ZN(P2_U2938) );
  AOI22_X1 U22057 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19089), .B1(n19088), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19072) );
  OAI21_X1 U22058 ( .B1(n19091), .B2(n20869), .A(n19072), .ZN(P2_U2939) );
  AOI22_X1 U22059 ( .A1(n19097), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19073) );
  OAI21_X1 U22060 ( .B1(n19074), .B2(n19099), .A(n19073), .ZN(P2_U2940) );
  AOI22_X1 U22061 ( .A1(n19097), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19075) );
  OAI21_X1 U22062 ( .B1(n19076), .B2(n19099), .A(n19075), .ZN(P2_U2941) );
  AOI22_X1 U22063 ( .A1(n19097), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19077) );
  OAI21_X1 U22064 ( .B1(n20882), .B2(n19099), .A(n19077), .ZN(P2_U2942) );
  AOI22_X1 U22065 ( .A1(n19097), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19078) );
  OAI21_X1 U22066 ( .B1(n19079), .B2(n19099), .A(n19078), .ZN(P2_U2943) );
  AOI22_X1 U22067 ( .A1(n19097), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19080) );
  OAI21_X1 U22068 ( .B1(n19081), .B2(n19099), .A(n19080), .ZN(P2_U2944) );
  AOI22_X1 U22069 ( .A1(n19097), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19082) );
  OAI21_X1 U22070 ( .B1(n19083), .B2(n19099), .A(n19082), .ZN(P2_U2945) );
  INV_X1 U22071 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19085) );
  AOI22_X1 U22072 ( .A1(n19097), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19084) );
  OAI21_X1 U22073 ( .B1(n19085), .B2(n19099), .A(n19084), .ZN(P2_U2946) );
  INV_X1 U22074 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19087) );
  AOI22_X1 U22075 ( .A1(n19097), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19086) );
  OAI21_X1 U22076 ( .B1(n19087), .B2(n19099), .A(n19086), .ZN(P2_U2947) );
  AOI22_X1 U22077 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n19089), .B1(n19088), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n19090) );
  OAI21_X1 U22078 ( .B1(n19091), .B2(n20956), .A(n19090), .ZN(P2_U2948) );
  INV_X1 U22079 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19093) );
  AOI22_X1 U22080 ( .A1(n19097), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19092) );
  OAI21_X1 U22081 ( .B1(n19093), .B2(n19099), .A(n19092), .ZN(P2_U2949) );
  INV_X1 U22082 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19096) );
  AOI22_X1 U22083 ( .A1(n19097), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19095) );
  OAI21_X1 U22084 ( .B1(n19096), .B2(n19099), .A(n19095), .ZN(P2_U2950) );
  AOI22_X1 U22085 ( .A1(n19097), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19094), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19098) );
  OAI21_X1 U22086 ( .B1(n11888), .B2(n19099), .A(n19098), .ZN(P2_U2951) );
  AOI22_X1 U22087 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n19101), .B1(n19100), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n19103) );
  NAND2_X1 U22088 ( .A1(n19103), .A2(n19102), .ZN(P2_U2979) );
  AOI22_X1 U22089 ( .A1(n19104), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19132), .ZN(n19118) );
  AOI21_X1 U22090 ( .B1(n19107), .B2(n19106), .A(n19105), .ZN(n19110) );
  XNOR2_X1 U22091 ( .A(n19108), .B(n19123), .ZN(n19109) );
  XNOR2_X1 U22092 ( .A(n19110), .B(n19109), .ZN(n19131) );
  NAND2_X1 U22093 ( .A1(n19112), .A2(n19111), .ZN(n19113) );
  XNOR2_X1 U22094 ( .A(n19113), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19128) );
  AOI222_X1 U22095 ( .A1(n19131), .A2(n19116), .B1(n19115), .B2(n19128), .C1(
        n19114), .C2(n19122), .ZN(n19117) );
  OAI211_X1 U22096 ( .C1(n19120), .C2(n19119), .A(n19118), .B(n19117), .ZN(
        P2_U3010) );
  AOI22_X1 U22097 ( .A1(n19124), .A2(n19123), .B1(n19122), .B2(n19121), .ZN(
        n19136) );
  AOI22_X1 U22098 ( .A1(n19127), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19126), .B2(n19125), .ZN(n19135) );
  AOI22_X1 U22099 ( .A1(n19131), .A2(n19130), .B1(n19129), .B2(n19128), .ZN(
        n19134) );
  NAND2_X1 U22100 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19132), .ZN(n19133) );
  NAND4_X1 U22101 ( .A1(n19136), .A2(n19135), .A3(n19134), .A4(n19133), .ZN(
        P2_U3042) );
  NAND2_X1 U22102 ( .A1(n19213), .A2(n19787), .ZN(n19189) );
  NOR2_X1 U22103 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19189), .ZN(
        n19179) );
  AOI22_X1 U22104 ( .A1(n19663), .A2(n19626), .B1(n19618), .B2(n19179), .ZN(
        n19149) );
  INV_X1 U22105 ( .A(n19211), .ZN(n19138) );
  NOR2_X1 U22106 ( .A1(n19663), .A2(n19138), .ZN(n19139) );
  OAI21_X1 U22107 ( .B1(n19139), .B2(n19574), .A(n19771), .ZN(n19147) );
  NOR2_X1 U22108 ( .A1(n19669), .A2(n19179), .ZN(n19146) );
  INV_X1 U22109 ( .A(n19146), .ZN(n19143) );
  OAI21_X1 U22110 ( .B1(n19144), .B2(n19390), .A(n19616), .ZN(n19141) );
  INV_X1 U22111 ( .A(n19179), .ZN(n19140) );
  AOI21_X1 U22112 ( .B1(n19141), .B2(n19140), .A(n19281), .ZN(n19142) );
  OAI21_X1 U22113 ( .B1(n19144), .B2(n19179), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19145) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19181), .B1(
        n19619), .B2(n19180), .ZN(n19148) );
  OAI211_X1 U22115 ( .C1(n19629), .C2(n19211), .A(n19149), .B(n19148), .ZN(
        P2_U3048) );
  AOI22_X1 U22116 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19173), .ZN(n19591) );
  AOI22_X1 U22117 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19173), .ZN(n19635) );
  NOR2_X2 U22118 ( .A1(n10055), .A2(n19175), .ZN(n19630) );
  AOI22_X1 U22119 ( .A1(n19663), .A2(n19588), .B1(n19630), .B2(n19179), .ZN(
        n19152) );
  NOR2_X2 U22120 ( .A1(n19150), .A2(n19281), .ZN(n19631) );
  AOI22_X1 U22121 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19181), .B1(
        n19631), .B2(n19180), .ZN(n19151) );
  OAI211_X1 U22122 ( .C1(n19591), .C2(n19211), .A(n19152), .B(n19151), .ZN(
        P2_U3049) );
  AOI22_X1 U22123 ( .A1(n19663), .A2(n19638), .B1(n19636), .B2(n19179), .ZN(
        n19154) );
  AOI22_X1 U22124 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19181), .B1(
        n19637), .B2(n19180), .ZN(n19153) );
  OAI211_X1 U22125 ( .C1(n19641), .C2(n19211), .A(n19154), .B(n19153), .ZN(
        P2_U3050) );
  AOI22_X1 U22126 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19173), .ZN(n19559) );
  NOR2_X2 U22127 ( .A1(n19157), .A2(n19175), .ZN(n19642) );
  AOI22_X1 U22128 ( .A1(n19663), .A2(n19556), .B1(n19642), .B2(n19179), .ZN(
        n19160) );
  NOR2_X2 U22129 ( .A1(n19158), .A2(n19281), .ZN(n19643) );
  AOI22_X1 U22130 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19181), .B1(
        n19643), .B2(n19180), .ZN(n19159) );
  OAI211_X1 U22131 ( .C1(n19559), .C2(n19211), .A(n19160), .B(n19159), .ZN(
        P2_U3051) );
  AOI22_X1 U22132 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19173), .ZN(n19600) );
  OAI22_X2 U22133 ( .A1(n14746), .A2(n19171), .B1(n19161), .B2(n19169), .ZN(
        n19597) );
  NOR2_X2 U22134 ( .A1(n19162), .A2(n19175), .ZN(n19648) );
  AOI22_X1 U22135 ( .A1(n19663), .A2(n19597), .B1(n19648), .B2(n19179), .ZN(
        n19165) );
  NOR2_X2 U22136 ( .A1(n19163), .A2(n19281), .ZN(n19649) );
  AOI22_X1 U22137 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19181), .B1(
        n19649), .B2(n19180), .ZN(n19164) );
  OAI211_X1 U22138 ( .C1(n19600), .C2(n19211), .A(n19165), .B(n19164), .ZN(
        P2_U3052) );
  AOI22_X1 U22139 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19173), .ZN(n19659) );
  AOI22_X1 U22140 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19173), .ZN(n19507) );
  NOR2_X2 U22141 ( .A1(n13502), .A2(n19175), .ZN(n19654) );
  AOI22_X1 U22142 ( .A1(n19663), .A2(n19656), .B1(n19654), .B2(n19179), .ZN(
        n19168) );
  NOR2_X2 U22143 ( .A1(n19166), .A2(n19281), .ZN(n19655) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19181), .B1(
        n19655), .B2(n19180), .ZN(n19167) );
  OAI211_X1 U22145 ( .C1(n19659), .C2(n19211), .A(n19168), .B(n19167), .ZN(
        P2_U3053) );
  AOI22_X1 U22146 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19174), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19173), .ZN(n19667) );
  NOR2_X2 U22147 ( .A1(n12043), .A2(n19175), .ZN(n19660) );
  AOI22_X1 U22148 ( .A1(n19663), .A2(n19603), .B1(n19660), .B2(n19179), .ZN(
        n19178) );
  NOR2_X2 U22149 ( .A1(n19176), .A2(n19281), .ZN(n19661) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19181), .B1(
        n19661), .B2(n19180), .ZN(n19177) );
  OAI211_X1 U22151 ( .C1(n19606), .C2(n19211), .A(n19178), .B(n19177), .ZN(
        P2_U3054) );
  AOI22_X1 U22152 ( .A1(n19663), .A2(n19672), .B1(n19668), .B2(n19179), .ZN(
        n19183) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19181), .B1(
        n19670), .B2(n19180), .ZN(n19182) );
  OAI211_X1 U22154 ( .C1(n19678), .C2(n19211), .A(n19183), .B(n19182), .ZN(
        P2_U3055) );
  INV_X1 U22155 ( .A(n19184), .ZN(n19359) );
  INV_X1 U22156 ( .A(n19185), .ZN(n19186) );
  NAND2_X1 U22157 ( .A1(n19787), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19422) );
  NOR2_X1 U22158 ( .A1(n19422), .A2(n19244), .ZN(n19206) );
  NOR3_X1 U22159 ( .A1(n19186), .A2(n19206), .A3(n19390), .ZN(n19188) );
  AOI211_X2 U22160 ( .C1(n19189), .C2(n19390), .A(n19359), .B(n19188), .ZN(
        n19207) );
  AOI22_X1 U22161 ( .A1(n19207), .A2(n19619), .B1(n19618), .B2(n19206), .ZN(
        n19193) );
  INV_X1 U22162 ( .A(n19362), .ZN(n19187) );
  NAND2_X1 U22163 ( .A1(n19187), .A2(n19420), .ZN(n19190) );
  AOI21_X1 U22164 ( .B1(n19190), .B2(n19189), .A(n19188), .ZN(n19191) );
  OAI211_X1 U22165 ( .C1(n19206), .C2(n19616), .A(n19191), .B(n19624), .ZN(
        n19208) );
  NAND2_X1 U22166 ( .A1(n19420), .A2(n19367), .ZN(n19218) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19208), .B1(
        n19240), .B2(n19573), .ZN(n19192) );
  OAI211_X1 U22168 ( .C1(n19587), .C2(n19211), .A(n19193), .B(n19192), .ZN(
        P2_U3056) );
  AOI22_X1 U22169 ( .A1(n19207), .A2(n19631), .B1(n19630), .B2(n19206), .ZN(
        n19195) );
  INV_X1 U22170 ( .A(n19591), .ZN(n19632) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19208), .B1(
        n19240), .B2(n19632), .ZN(n19194) );
  OAI211_X1 U22172 ( .C1(n19635), .C2(n19211), .A(n19195), .B(n19194), .ZN(
        P2_U3057) );
  AOI22_X1 U22173 ( .A1(n19207), .A2(n19637), .B1(n19636), .B2(n19206), .ZN(
        n19197) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19208), .B1(
        n19240), .B2(n19523), .ZN(n19196) );
  OAI211_X1 U22175 ( .C1(n19500), .C2(n19211), .A(n19197), .B(n19196), .ZN(
        P2_U3058) );
  INV_X1 U22176 ( .A(n19556), .ZN(n19647) );
  AOI22_X1 U22177 ( .A1(n19207), .A2(n19643), .B1(n19642), .B2(n19206), .ZN(
        n19199) );
  INV_X1 U22178 ( .A(n19559), .ZN(n19644) );
  AOI22_X1 U22179 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19208), .B1(
        n19240), .B2(n19644), .ZN(n19198) );
  OAI211_X1 U22180 ( .C1(n19647), .C2(n19211), .A(n19199), .B(n19198), .ZN(
        P2_U3059) );
  INV_X1 U22181 ( .A(n19597), .ZN(n19653) );
  AOI22_X1 U22182 ( .A1(n19207), .A2(n19649), .B1(n19648), .B2(n19206), .ZN(
        n19201) );
  INV_X1 U22183 ( .A(n19600), .ZN(n19650) );
  AOI22_X1 U22184 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19208), .B1(
        n19240), .B2(n19650), .ZN(n19200) );
  OAI211_X1 U22185 ( .C1(n19653), .C2(n19211), .A(n19201), .B(n19200), .ZN(
        P2_U3060) );
  AOI22_X1 U22186 ( .A1(n19207), .A2(n19655), .B1(n19654), .B2(n19206), .ZN(
        n19203) );
  INV_X1 U22187 ( .A(n19659), .ZN(n19531) );
  AOI22_X1 U22188 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19208), .B1(
        n19240), .B2(n19531), .ZN(n19202) );
  OAI211_X1 U22189 ( .C1(n19507), .C2(n19211), .A(n19203), .B(n19202), .ZN(
        P2_U3061) );
  AOI22_X1 U22190 ( .A1(n19207), .A2(n19661), .B1(n19660), .B2(n19206), .ZN(
        n19205) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19208), .B1(
        n19240), .B2(n19662), .ZN(n19204) );
  OAI211_X1 U22192 ( .C1(n19667), .C2(n19211), .A(n19205), .B(n19204), .ZN(
        P2_U3062) );
  INV_X1 U22193 ( .A(n19672), .ZN(n19517) );
  AOI22_X1 U22194 ( .A1(n19207), .A2(n19670), .B1(n19668), .B2(n19206), .ZN(
        n19210) );
  AOI22_X1 U22195 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19208), .B1(
        n19240), .B2(n19512), .ZN(n19209) );
  OAI211_X1 U22196 ( .C1(n19517), .C2(n19211), .A(n19210), .B(n19209), .ZN(
        P2_U3063) );
  INV_X1 U22197 ( .A(n19212), .ZN(n19217) );
  NOR2_X1 U22198 ( .A1(n19787), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19454) );
  AND2_X1 U22199 ( .A1(n19454), .A2(n19213), .ZN(n19238) );
  OAI21_X1 U22200 ( .B1(n19217), .B2(n19238), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19216) );
  INV_X1 U22201 ( .A(n19214), .ZN(n19457) );
  NOR2_X1 U22202 ( .A1(n19457), .A2(n19244), .ZN(n19219) );
  INV_X1 U22203 ( .A(n19219), .ZN(n19215) );
  NAND2_X1 U22204 ( .A1(n19216), .A2(n19215), .ZN(n19239) );
  AOI22_X1 U22205 ( .A1(n19239), .A2(n19619), .B1(n19618), .B2(n19238), .ZN(
        n19225) );
  AOI21_X1 U22206 ( .B1(n19217), .B2(n19616), .A(n19238), .ZN(n19222) );
  AOI21_X1 U22207 ( .B1(n19263), .B2(n19218), .A(n19574), .ZN(n19220) );
  NOR2_X1 U22208 ( .A1(n19220), .A2(n19219), .ZN(n19221) );
  MUX2_X1 U22209 ( .A(n19222), .B(n19221), .S(n19771), .Z(n19223) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19626), .ZN(n19224) );
  OAI211_X1 U22211 ( .C1(n19629), .C2(n19263), .A(n19225), .B(n19224), .ZN(
        P2_U3064) );
  AOI22_X1 U22212 ( .A1(n19239), .A2(n19631), .B1(n19630), .B2(n19238), .ZN(
        n19227) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19588), .ZN(n19226) );
  OAI211_X1 U22214 ( .C1(n19591), .C2(n19263), .A(n19227), .B(n19226), .ZN(
        P2_U3065) );
  AOI22_X1 U22215 ( .A1(n19239), .A2(n19637), .B1(n19636), .B2(n19238), .ZN(
        n19229) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19638), .ZN(n19228) );
  OAI211_X1 U22217 ( .C1(n19641), .C2(n19263), .A(n19229), .B(n19228), .ZN(
        P2_U3066) );
  AOI22_X1 U22218 ( .A1(n19239), .A2(n19643), .B1(n19642), .B2(n19238), .ZN(
        n19231) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19556), .ZN(n19230) );
  OAI211_X1 U22220 ( .C1(n19559), .C2(n19263), .A(n19231), .B(n19230), .ZN(
        P2_U3067) );
  AOI22_X1 U22221 ( .A1(n19239), .A2(n19649), .B1(n19648), .B2(n19238), .ZN(
        n19233) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19597), .ZN(n19232) );
  OAI211_X1 U22223 ( .C1(n19600), .C2(n19263), .A(n19233), .B(n19232), .ZN(
        P2_U3068) );
  AOI22_X1 U22224 ( .A1(n19239), .A2(n19655), .B1(n19654), .B2(n19238), .ZN(
        n19235) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19656), .ZN(n19234) );
  OAI211_X1 U22226 ( .C1(n19659), .C2(n19263), .A(n19235), .B(n19234), .ZN(
        P2_U3069) );
  AOI22_X1 U22227 ( .A1(n19239), .A2(n19661), .B1(n19660), .B2(n19238), .ZN(
        n19237) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19603), .ZN(n19236) );
  OAI211_X1 U22229 ( .C1(n19606), .C2(n19263), .A(n19237), .B(n19236), .ZN(
        P2_U3070) );
  AOI22_X1 U22230 ( .A1(n19239), .A2(n19670), .B1(n19668), .B2(n19238), .ZN(
        n19243) );
  AOI22_X1 U22231 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19241), .B1(
        n19240), .B2(n19672), .ZN(n19242) );
  OAI211_X1 U22232 ( .C1(n19678), .C2(n19263), .A(n19243), .B(n19242), .ZN(
        P2_U3071) );
  INV_X1 U22233 ( .A(n19263), .ZN(n19269) );
  NOR2_X1 U22234 ( .A1(n19485), .A2(n19244), .ZN(n19268) );
  AOI22_X1 U22235 ( .A1(n19626), .A2(n19269), .B1(n19618), .B2(n19268), .ZN(
        n19254) );
  OAI21_X1 U22236 ( .B1(n19362), .B2(n19491), .A(n19771), .ZN(n19252) );
  NOR2_X1 U22237 ( .A1(n19787), .A2(n19244), .ZN(n19248) );
  INV_X1 U22238 ( .A(n19268), .ZN(n19245) );
  OAI211_X1 U22239 ( .C1(n19246), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19245), 
        .B(n19762), .ZN(n19247) );
  OAI211_X1 U22240 ( .C1(n19252), .C2(n19248), .A(n19624), .B(n19247), .ZN(
        n19271) );
  INV_X1 U22241 ( .A(n19248), .ZN(n19251) );
  OAI21_X1 U22242 ( .B1(n19249), .B2(n19268), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19250) );
  OAI21_X1 U22243 ( .B1(n19252), .B2(n19251), .A(n19250), .ZN(n19270) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19271), .B1(
        n19619), .B2(n19270), .ZN(n19253) );
  OAI211_X1 U22245 ( .C1(n19629), .C2(n19279), .A(n19254), .B(n19253), .ZN(
        P2_U3072) );
  AOI22_X1 U22246 ( .A1(n19632), .A2(n19302), .B1(n19268), .B2(n19630), .ZN(
        n19256) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19271), .B1(
        n19631), .B2(n19270), .ZN(n19255) );
  OAI211_X1 U22248 ( .C1(n19635), .C2(n19263), .A(n19256), .B(n19255), .ZN(
        P2_U3073) );
  AOI22_X1 U22249 ( .A1(n19269), .A2(n19638), .B1(n19636), .B2(n19268), .ZN(
        n19258) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19271), .B1(
        n19637), .B2(n19270), .ZN(n19257) );
  OAI211_X1 U22251 ( .C1(n19641), .C2(n19279), .A(n19258), .B(n19257), .ZN(
        P2_U3074) );
  AOI22_X1 U22252 ( .A1(n19644), .A2(n19302), .B1(n19268), .B2(n19642), .ZN(
        n19260) );
  AOI22_X1 U22253 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19271), .B1(
        n19643), .B2(n19270), .ZN(n19259) );
  OAI211_X1 U22254 ( .C1(n19647), .C2(n19263), .A(n19260), .B(n19259), .ZN(
        P2_U3075) );
  AOI22_X1 U22255 ( .A1(n19650), .A2(n19302), .B1(n19268), .B2(n19648), .ZN(
        n19262) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19271), .B1(
        n19649), .B2(n19270), .ZN(n19261) );
  OAI211_X1 U22257 ( .C1(n19653), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U3076) );
  AOI22_X1 U22258 ( .A1(n19269), .A2(n19656), .B1(n19268), .B2(n19654), .ZN(
        n19265) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19271), .B1(
        n19655), .B2(n19270), .ZN(n19264) );
  OAI211_X1 U22260 ( .C1(n19659), .C2(n19279), .A(n19265), .B(n19264), .ZN(
        P2_U3077) );
  AOI22_X1 U22261 ( .A1(n19269), .A2(n19603), .B1(n19268), .B2(n19660), .ZN(
        n19267) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19271), .B1(
        n19661), .B2(n19270), .ZN(n19266) );
  OAI211_X1 U22263 ( .C1(n19606), .C2(n19279), .A(n19267), .B(n19266), .ZN(
        P2_U3078) );
  AOI22_X1 U22264 ( .A1(n19672), .A2(n19269), .B1(n19668), .B2(n19268), .ZN(
        n19273) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19271), .B1(
        n19670), .B2(n19270), .ZN(n19272) );
  OAI211_X1 U22266 ( .C1(n19678), .C2(n19279), .A(n19273), .B(n19272), .ZN(
        P2_U3079) );
  NAND2_X1 U22267 ( .A1(n19274), .A2(n19770), .ZN(n19278) );
  OR2_X1 U22268 ( .A1(n19278), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19277) );
  INV_X1 U22269 ( .A(n13305), .ZN(n19276) );
  NOR2_X1 U22270 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19275), .ZN(
        n19300) );
  NOR3_X1 U22271 ( .A1(n19276), .A2(n19300), .A3(n19390), .ZN(n19280) );
  AOI21_X1 U22272 ( .B1(n19390), .B2(n19277), .A(n19280), .ZN(n19301) );
  AOI22_X1 U22273 ( .A1(n19301), .A2(n19619), .B1(n19618), .B2(n19300), .ZN(
        n19287) );
  INV_X1 U22274 ( .A(n19278), .ZN(n19285) );
  AOI21_X1 U22275 ( .B1(n19279), .B2(n19322), .A(n19574), .ZN(n19284) );
  INV_X1 U22276 ( .A(n19300), .ZN(n19282) );
  AOI211_X1 U22277 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19282), .A(n19281), 
        .B(n19280), .ZN(n19283) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19626), .ZN(n19286) );
  OAI211_X1 U22279 ( .C1(n19629), .C2(n19322), .A(n19287), .B(n19286), .ZN(
        P2_U3080) );
  AOI22_X1 U22280 ( .A1(n19301), .A2(n19631), .B1(n19630), .B2(n19300), .ZN(
        n19289) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19588), .ZN(n19288) );
  OAI211_X1 U22282 ( .C1(n19591), .C2(n19322), .A(n19289), .B(n19288), .ZN(
        P2_U3081) );
  AOI22_X1 U22283 ( .A1(n19301), .A2(n19637), .B1(n19636), .B2(n19300), .ZN(
        n19291) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19638), .ZN(n19290) );
  OAI211_X1 U22285 ( .C1(n19641), .C2(n19322), .A(n19291), .B(n19290), .ZN(
        P2_U3082) );
  AOI22_X1 U22286 ( .A1(n19301), .A2(n19643), .B1(n19642), .B2(n19300), .ZN(
        n19293) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19556), .ZN(n19292) );
  OAI211_X1 U22288 ( .C1(n19559), .C2(n19322), .A(n19293), .B(n19292), .ZN(
        P2_U3083) );
  AOI22_X1 U22289 ( .A1(n19301), .A2(n19649), .B1(n19648), .B2(n19300), .ZN(
        n19295) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19597), .ZN(n19294) );
  OAI211_X1 U22291 ( .C1(n19600), .C2(n19322), .A(n19295), .B(n19294), .ZN(
        P2_U3084) );
  AOI22_X1 U22292 ( .A1(n19301), .A2(n19655), .B1(n19654), .B2(n19300), .ZN(
        n19297) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19656), .ZN(n19296) );
  OAI211_X1 U22294 ( .C1(n19659), .C2(n19322), .A(n19297), .B(n19296), .ZN(
        P2_U3085) );
  AOI22_X1 U22295 ( .A1(n19301), .A2(n19661), .B1(n19660), .B2(n19300), .ZN(
        n19299) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19603), .ZN(n19298) );
  OAI211_X1 U22297 ( .C1(n19606), .C2(n19322), .A(n19299), .B(n19298), .ZN(
        P2_U3086) );
  AOI22_X1 U22298 ( .A1(n19301), .A2(n19670), .B1(n19668), .B2(n19300), .ZN(
        n19305) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19303), .B1(
        n19302), .B2(n19672), .ZN(n19304) );
  OAI211_X1 U22300 ( .C1(n19678), .C2(n19322), .A(n19305), .B(n19304), .ZN(
        P2_U3087) );
  INV_X1 U22301 ( .A(n19322), .ZN(n19306) );
  AOI22_X1 U22302 ( .A1(n19306), .A2(n19588), .B1(n19330), .B2(n19630), .ZN(
        n19308) );
  AOI22_X1 U22303 ( .A1(n19631), .A2(n19318), .B1(n19353), .B2(n19632), .ZN(
        n19307) );
  OAI211_X1 U22304 ( .C1(n19309), .C2(n13286), .A(n19308), .B(n19307), .ZN(
        P2_U3089) );
  AOI22_X1 U22305 ( .A1(n19644), .A2(n19353), .B1(n19330), .B2(n19642), .ZN(
        n19311) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19319), .B1(
        n19643), .B2(n19318), .ZN(n19310) );
  OAI211_X1 U22307 ( .C1(n19647), .C2(n19322), .A(n19311), .B(n19310), .ZN(
        P2_U3091) );
  AOI22_X1 U22308 ( .A1(n19650), .A2(n19353), .B1(n19330), .B2(n19648), .ZN(
        n19313) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19319), .B1(
        n19649), .B2(n19318), .ZN(n19312) );
  OAI211_X1 U22310 ( .C1(n19653), .C2(n19322), .A(n19313), .B(n19312), .ZN(
        P2_U3092) );
  AOI22_X1 U22311 ( .A1(n19531), .A2(n19353), .B1(n19330), .B2(n19654), .ZN(
        n19315) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19319), .B1(
        n19655), .B2(n19318), .ZN(n19314) );
  OAI211_X1 U22313 ( .C1(n19507), .C2(n19322), .A(n19315), .B(n19314), .ZN(
        P2_U3093) );
  AOI22_X1 U22314 ( .A1(n19662), .A2(n19353), .B1(n19330), .B2(n19660), .ZN(
        n19317) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19319), .B1(
        n19661), .B2(n19318), .ZN(n19316) );
  OAI211_X1 U22316 ( .C1(n19667), .C2(n19322), .A(n19317), .B(n19316), .ZN(
        P2_U3094) );
  AOI22_X1 U22317 ( .A1(n19512), .A2(n19353), .B1(n19668), .B2(n19330), .ZN(
        n19321) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19319), .B1(
        n19670), .B2(n19318), .ZN(n19320) );
  OAI211_X1 U22319 ( .C1(n19517), .C2(n19322), .A(n19321), .B(n19320), .ZN(
        P2_U3095) );
  INV_X1 U22320 ( .A(n19353), .ZN(n19350) );
  AOI21_X1 U22321 ( .B1(n19350), .B2(n19380), .A(n19574), .ZN(n19324) );
  NOR2_X1 U22322 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19572), .ZN(
        n19366) );
  INV_X1 U22323 ( .A(n19366), .ZN(n19360) );
  NOR2_X1 U22324 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19360), .ZN(
        n19351) );
  AOI221_X1 U22325 ( .B1(n19330), .B2(n19616), .C1(n19324), .C2(n19616), .A(
        n19351), .ZN(n19329) );
  INV_X1 U22326 ( .A(n19351), .ZN(n19325) );
  AND2_X1 U22327 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19325), .ZN(n19326) );
  NAND2_X1 U22328 ( .A1(n19327), .A2(n19326), .ZN(n19331) );
  NAND2_X1 U22329 ( .A1(n19331), .A2(n19624), .ZN(n19328) );
  INV_X1 U22330 ( .A(n19354), .ZN(n19337) );
  INV_X1 U22331 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19336) );
  NOR2_X1 U22332 ( .A1(n19330), .A2(n19351), .ZN(n19333) );
  INV_X1 U22333 ( .A(n19331), .ZN(n19332) );
  AOI211_X2 U22334 ( .C1(n19333), .C2(n19390), .A(n19359), .B(n19332), .ZN(
        n19352) );
  AOI22_X1 U22335 ( .A1(n19352), .A2(n19619), .B1(n19618), .B2(n19351), .ZN(
        n19335) );
  INV_X1 U22336 ( .A(n19380), .ZN(n19384) );
  AOI22_X1 U22337 ( .A1(n19353), .A2(n19626), .B1(n19384), .B2(n19573), .ZN(
        n19334) );
  OAI211_X1 U22338 ( .C1(n19337), .C2(n19336), .A(n19335), .B(n19334), .ZN(
        P2_U3096) );
  AOI22_X1 U22339 ( .A1(n19352), .A2(n19631), .B1(n19630), .B2(n19351), .ZN(
        n19339) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19588), .ZN(n19338) );
  OAI211_X1 U22341 ( .C1(n19591), .C2(n19380), .A(n19339), .B(n19338), .ZN(
        P2_U3097) );
  AOI22_X1 U22342 ( .A1(n19352), .A2(n19637), .B1(n19636), .B2(n19351), .ZN(
        n19341) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19638), .ZN(n19340) );
  OAI211_X1 U22344 ( .C1(n19641), .C2(n19380), .A(n19341), .B(n19340), .ZN(
        P2_U3098) );
  AOI22_X1 U22345 ( .A1(n19352), .A2(n19643), .B1(n19642), .B2(n19351), .ZN(
        n19343) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19556), .ZN(n19342) );
  OAI211_X1 U22347 ( .C1(n19559), .C2(n19380), .A(n19343), .B(n19342), .ZN(
        P2_U3099) );
  AOI22_X1 U22348 ( .A1(n19352), .A2(n19649), .B1(n19648), .B2(n19351), .ZN(
        n19345) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19597), .ZN(n19344) );
  OAI211_X1 U22350 ( .C1(n19600), .C2(n19380), .A(n19345), .B(n19344), .ZN(
        P2_U3100) );
  AOI22_X1 U22351 ( .A1(n19352), .A2(n19655), .B1(n19654), .B2(n19351), .ZN(
        n19347) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19656), .ZN(n19346) );
  OAI211_X1 U22353 ( .C1(n19659), .C2(n19380), .A(n19347), .B(n19346), .ZN(
        P2_U3101) );
  AOI22_X1 U22354 ( .A1(n19352), .A2(n19661), .B1(n19660), .B2(n19351), .ZN(
        n19349) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19354), .B1(
        n19384), .B2(n19662), .ZN(n19348) );
  OAI211_X1 U22356 ( .C1(n19667), .C2(n19350), .A(n19349), .B(n19348), .ZN(
        P2_U3102) );
  AOI22_X1 U22357 ( .A1(n19352), .A2(n19670), .B1(n19668), .B2(n19351), .ZN(
        n19356) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19354), .B1(
        n19353), .B2(n19672), .ZN(n19355) );
  OAI211_X1 U22359 ( .C1(n19678), .C2(n19380), .A(n19356), .B(n19355), .ZN(
        P2_U3103) );
  NAND2_X1 U22360 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19366), .ZN(
        n19392) );
  AND2_X1 U22361 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19392), .ZN(n19357) );
  AOI211_X2 U22362 ( .C1(n19360), .C2(n19390), .A(n19359), .B(n19364), .ZN(
        n19383) );
  INV_X1 U22363 ( .A(n19392), .ZN(n19395) );
  AOI22_X1 U22364 ( .A1(n19383), .A2(n19619), .B1(n19618), .B2(n19395), .ZN(
        n19369) );
  NOR2_X1 U22365 ( .A1(n19362), .A2(n19361), .ZN(n19766) );
  OAI21_X1 U22366 ( .B1(n19616), .B2(n19395), .A(n19624), .ZN(n19363) );
  NOR2_X1 U22367 ( .A1(n19364), .A2(n19363), .ZN(n19365) );
  OAI21_X1 U22368 ( .B1(n19366), .B2(n19766), .A(n19365), .ZN(n19385) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19385), .B1(
        n19415), .B2(n19573), .ZN(n19368) );
  OAI211_X1 U22370 ( .C1(n19587), .C2(n19380), .A(n19369), .B(n19368), .ZN(
        P2_U3104) );
  AOI22_X1 U22371 ( .A1(n19383), .A2(n19631), .B1(n19630), .B2(n19395), .ZN(
        n19371) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19385), .B1(
        n19415), .B2(n19632), .ZN(n19370) );
  OAI211_X1 U22373 ( .C1(n19635), .C2(n19380), .A(n19371), .B(n19370), .ZN(
        P2_U3105) );
  AOI22_X1 U22374 ( .A1(n19383), .A2(n19637), .B1(n19636), .B2(n19395), .ZN(
        n19373) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19385), .B1(
        n19415), .B2(n19523), .ZN(n19372) );
  OAI211_X1 U22376 ( .C1(n19500), .C2(n19380), .A(n19373), .B(n19372), .ZN(
        P2_U3106) );
  AOI22_X1 U22377 ( .A1(n19383), .A2(n19643), .B1(n19642), .B2(n19395), .ZN(
        n19375) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19385), .B1(
        n19415), .B2(n19644), .ZN(n19374) );
  OAI211_X1 U22379 ( .C1(n19647), .C2(n19380), .A(n19375), .B(n19374), .ZN(
        P2_U3107) );
  AOI22_X1 U22380 ( .A1(n19383), .A2(n19649), .B1(n19648), .B2(n19395), .ZN(
        n19377) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19597), .ZN(n19376) );
  OAI211_X1 U22382 ( .C1(n19600), .C2(n19413), .A(n19377), .B(n19376), .ZN(
        P2_U3108) );
  AOI22_X1 U22383 ( .A1(n19383), .A2(n19655), .B1(n19654), .B2(n19395), .ZN(
        n19379) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19385), .B1(
        n19415), .B2(n19531), .ZN(n19378) );
  OAI211_X1 U22385 ( .C1(n19507), .C2(n19380), .A(n19379), .B(n19378), .ZN(
        P2_U3109) );
  AOI22_X1 U22386 ( .A1(n19383), .A2(n19661), .B1(n19660), .B2(n19395), .ZN(
        n19382) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19603), .ZN(n19381) );
  OAI211_X1 U22388 ( .C1(n19606), .C2(n19413), .A(n19382), .B(n19381), .ZN(
        P2_U3110) );
  AOI22_X1 U22389 ( .A1(n19383), .A2(n19670), .B1(n19668), .B2(n19395), .ZN(
        n19387) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19385), .B1(
        n19384), .B2(n19672), .ZN(n19386) );
  OAI211_X1 U22391 ( .C1(n19678), .C2(n19413), .A(n19387), .B(n19386), .ZN(
        P2_U3111) );
  NOR2_X1 U22392 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19770), .ZN(
        n19484) );
  NAND2_X1 U22393 ( .A1(n19484), .A2(n19787), .ZN(n19431) );
  NOR2_X1 U22394 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19431), .ZN(
        n19414) );
  AOI22_X1 U22395 ( .A1(n19626), .A2(n19415), .B1(n19618), .B2(n19414), .ZN(
        n19400) );
  NAND2_X1 U22396 ( .A1(n19452), .A2(n19413), .ZN(n19388) );
  AOI21_X1 U22397 ( .B1(n19388), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19762), 
        .ZN(n19394) );
  INV_X1 U22398 ( .A(n19389), .ZN(n19396) );
  OAI21_X1 U22399 ( .B1(n19396), .B2(n19390), .A(n19616), .ZN(n19391) );
  AOI21_X1 U22400 ( .B1(n19394), .B2(n19392), .A(n19391), .ZN(n19393) );
  OAI21_X1 U22401 ( .B1(n19414), .B2(n19395), .A(n19394), .ZN(n19398) );
  OAI21_X1 U22402 ( .B1(n19396), .B2(n19414), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19397) );
  NAND2_X1 U22403 ( .A1(n19398), .A2(n19397), .ZN(n19416) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19417), .B1(
        n19619), .B2(n19416), .ZN(n19399) );
  OAI211_X1 U22405 ( .C1(n19629), .C2(n19452), .A(n19400), .B(n19399), .ZN(
        P2_U3112) );
  AOI22_X1 U22406 ( .A1(n19441), .A2(n19632), .B1(n19630), .B2(n19414), .ZN(
        n19402) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19631), .ZN(n19401) );
  OAI211_X1 U22408 ( .C1(n19635), .C2(n19413), .A(n19402), .B(n19401), .ZN(
        P2_U3113) );
  AOI22_X1 U22409 ( .A1(n19441), .A2(n19523), .B1(n19636), .B2(n19414), .ZN(
        n19404) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19637), .ZN(n19403) );
  OAI211_X1 U22411 ( .C1(n19500), .C2(n19413), .A(n19404), .B(n19403), .ZN(
        P2_U3114) );
  AOI22_X1 U22412 ( .A1(n19556), .A2(n19415), .B1(n19414), .B2(n19642), .ZN(
        n19406) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19643), .ZN(n19405) );
  OAI211_X1 U22414 ( .C1(n19559), .C2(n19452), .A(n19406), .B(n19405), .ZN(
        P2_U3115) );
  AOI22_X1 U22415 ( .A1(n19597), .A2(n19415), .B1(n19648), .B2(n19414), .ZN(
        n19408) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19649), .ZN(n19407) );
  OAI211_X1 U22417 ( .C1(n19600), .C2(n19452), .A(n19408), .B(n19407), .ZN(
        P2_U3116) );
  AOI22_X1 U22418 ( .A1(n19441), .A2(n19531), .B1(n19654), .B2(n19414), .ZN(
        n19410) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19655), .ZN(n19409) );
  OAI211_X1 U22420 ( .C1(n19507), .C2(n19413), .A(n19410), .B(n19409), .ZN(
        P2_U3117) );
  AOI22_X1 U22421 ( .A1(n19441), .A2(n19662), .B1(n19660), .B2(n19414), .ZN(
        n19412) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19661), .ZN(n19411) );
  OAI211_X1 U22423 ( .C1(n19667), .C2(n19413), .A(n19412), .B(n19411), .ZN(
        P2_U3118) );
  AOI22_X1 U22424 ( .A1(n19672), .A2(n19415), .B1(n19668), .B2(n19414), .ZN(
        n19419) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19670), .ZN(n19418) );
  OAI211_X1 U22426 ( .C1(n19678), .C2(n19452), .A(n19419), .B(n19418), .ZN(
        P2_U3119) );
  INV_X1 U22427 ( .A(n19484), .ZN(n19490) );
  NOR2_X1 U22428 ( .A1(n19422), .A2(n19490), .ZN(n19459) );
  AOI22_X1 U22429 ( .A1(n19480), .A2(n19573), .B1(n19618), .B2(n19459), .ZN(
        n19434) );
  INV_X1 U22430 ( .A(n19423), .ZN(n19768) );
  NAND2_X1 U22431 ( .A1(n19768), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19544) );
  OAI21_X1 U22432 ( .B1(n19544), .B2(n19424), .A(n19771), .ZN(n19432) );
  INV_X1 U22433 ( .A(n19431), .ZN(n19427) );
  INV_X1 U22434 ( .A(n19459), .ZN(n19425) );
  OAI211_X1 U22435 ( .C1(n19428), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19425), 
        .B(n19762), .ZN(n19426) );
  OAI211_X1 U22436 ( .C1(n19432), .C2(n19427), .A(n19624), .B(n19426), .ZN(
        n19449) );
  INV_X1 U22437 ( .A(n19428), .ZN(n19429) );
  OAI21_X1 U22438 ( .B1(n19429), .B2(n19459), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19430) );
  OAI21_X1 U22439 ( .B1(n19432), .B2(n19431), .A(n19430), .ZN(n19448) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19449), .B1(
        n19619), .B2(n19448), .ZN(n19433) );
  OAI211_X1 U22441 ( .C1(n19587), .C2(n19452), .A(n19434), .B(n19433), .ZN(
        P2_U3120) );
  AOI22_X1 U22442 ( .A1(n19441), .A2(n19588), .B1(n19630), .B2(n19459), .ZN(
        n19436) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19449), .B1(
        n19631), .B2(n19448), .ZN(n19435) );
  OAI211_X1 U22444 ( .C1(n19591), .C2(n19458), .A(n19436), .B(n19435), .ZN(
        P2_U3121) );
  AOI22_X1 U22445 ( .A1(n19523), .A2(n19480), .B1(n19636), .B2(n19459), .ZN(
        n19438) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19449), .B1(
        n19637), .B2(n19448), .ZN(n19437) );
  OAI211_X1 U22447 ( .C1(n19500), .C2(n19452), .A(n19438), .B(n19437), .ZN(
        P2_U3122) );
  AOI22_X1 U22448 ( .A1(n19441), .A2(n19556), .B1(n19459), .B2(n19642), .ZN(
        n19440) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19449), .B1(
        n19643), .B2(n19448), .ZN(n19439) );
  OAI211_X1 U22450 ( .C1(n19559), .C2(n19458), .A(n19440), .B(n19439), .ZN(
        P2_U3123) );
  AOI22_X1 U22451 ( .A1(n19441), .A2(n19597), .B1(n19648), .B2(n19459), .ZN(
        n19443) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19449), .B1(
        n19649), .B2(n19448), .ZN(n19442) );
  OAI211_X1 U22453 ( .C1(n19600), .C2(n19458), .A(n19443), .B(n19442), .ZN(
        P2_U3124) );
  AOI22_X1 U22454 ( .A1(n19480), .A2(n19531), .B1(n19654), .B2(n19459), .ZN(
        n19445) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19449), .B1(
        n19655), .B2(n19448), .ZN(n19444) );
  OAI211_X1 U22456 ( .C1(n19507), .C2(n19452), .A(n19445), .B(n19444), .ZN(
        P2_U3125) );
  AOI22_X1 U22457 ( .A1(n19662), .A2(n19480), .B1(n19660), .B2(n19459), .ZN(
        n19447) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19449), .B1(
        n19661), .B2(n19448), .ZN(n19446) );
  OAI211_X1 U22459 ( .C1(n19667), .C2(n19452), .A(n19447), .B(n19446), .ZN(
        P2_U3126) );
  AOI22_X1 U22460 ( .A1(n19512), .A2(n19480), .B1(n19668), .B2(n19459), .ZN(
        n19451) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19449), .B1(
        n19670), .B2(n19448), .ZN(n19450) );
  OAI211_X1 U22462 ( .C1(n19517), .C2(n19452), .A(n19451), .B(n19450), .ZN(
        P2_U3127) );
  INV_X1 U22463 ( .A(n19462), .ZN(n19455) );
  AND2_X1 U22464 ( .A1(n19454), .A2(n19484), .ZN(n19478) );
  OAI21_X1 U22465 ( .B1(n19455), .B2(n19478), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19456) );
  OAI21_X1 U22466 ( .B1(n19490), .B2(n19457), .A(n19456), .ZN(n19479) );
  AOI22_X1 U22467 ( .A1(n19479), .A2(n19619), .B1(n19618), .B2(n19478), .ZN(
        n19465) );
  AOI21_X1 U22468 ( .B1(n19458), .B2(n19516), .A(n19574), .ZN(n19460) );
  NOR2_X1 U22469 ( .A1(n19460), .A2(n19459), .ZN(n19461) );
  AOI211_X1 U22470 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19462), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19461), .ZN(n19463) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19481), .B1(
        n19480), .B2(n19626), .ZN(n19464) );
  OAI211_X1 U22472 ( .C1(n19629), .C2(n19516), .A(n19465), .B(n19464), .ZN(
        P2_U3128) );
  AOI22_X1 U22473 ( .A1(n19479), .A2(n19631), .B1(n19630), .B2(n19478), .ZN(
        n19467) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19481), .B1(
        n19480), .B2(n19588), .ZN(n19466) );
  OAI211_X1 U22475 ( .C1(n19591), .C2(n19516), .A(n19467), .B(n19466), .ZN(
        P2_U3129) );
  AOI22_X1 U22476 ( .A1(n19479), .A2(n19637), .B1(n19636), .B2(n19478), .ZN(
        n19469) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19481), .B1(
        n19480), .B2(n19638), .ZN(n19468) );
  OAI211_X1 U22478 ( .C1(n19641), .C2(n19516), .A(n19469), .B(n19468), .ZN(
        P2_U3130) );
  AOI22_X1 U22479 ( .A1(n19479), .A2(n19643), .B1(n19642), .B2(n19478), .ZN(
        n19471) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19481), .B1(
        n19480), .B2(n19556), .ZN(n19470) );
  OAI211_X1 U22481 ( .C1(n19559), .C2(n19516), .A(n19471), .B(n19470), .ZN(
        P2_U3131) );
  AOI22_X1 U22482 ( .A1(n19479), .A2(n19649), .B1(n19648), .B2(n19478), .ZN(
        n19473) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19481), .B1(
        n19480), .B2(n19597), .ZN(n19472) );
  OAI211_X1 U22484 ( .C1(n19600), .C2(n19516), .A(n19473), .B(n19472), .ZN(
        P2_U3132) );
  AOI22_X1 U22485 ( .A1(n19479), .A2(n19655), .B1(n19654), .B2(n19478), .ZN(
        n19475) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19481), .B1(
        n19480), .B2(n19656), .ZN(n19474) );
  OAI211_X1 U22487 ( .C1(n19659), .C2(n19516), .A(n19475), .B(n19474), .ZN(
        P2_U3133) );
  AOI22_X1 U22488 ( .A1(n19479), .A2(n19661), .B1(n19660), .B2(n19478), .ZN(
        n19477) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19481), .B1(
        n19480), .B2(n19603), .ZN(n19476) );
  OAI211_X1 U22490 ( .C1(n19606), .C2(n19516), .A(n19477), .B(n19476), .ZN(
        P2_U3134) );
  AOI22_X1 U22491 ( .A1(n19479), .A2(n19670), .B1(n19668), .B2(n19478), .ZN(
        n19483) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19481), .B1(
        n19480), .B2(n19672), .ZN(n19482) );
  OAI211_X1 U22493 ( .C1(n19678), .C2(n19516), .A(n19483), .B(n19482), .ZN(
        P2_U3135) );
  NAND2_X1 U22494 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19484), .ZN(
        n19488) );
  INV_X1 U22495 ( .A(n19489), .ZN(n19486) );
  NOR2_X1 U22496 ( .A1(n19490), .A2(n19485), .ZN(n19510) );
  OAI21_X1 U22497 ( .B1(n19486), .B2(n19510), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19487) );
  OAI21_X1 U22498 ( .B1(n19488), .B2(n19762), .A(n19487), .ZN(n19511) );
  AOI22_X1 U22499 ( .A1(n19511), .A2(n19619), .B1(n19618), .B2(n19510), .ZN(
        n19495) );
  AOI21_X1 U22500 ( .B1(n19489), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19493) );
  OAI22_X1 U22501 ( .A1(n19544), .A2(n19491), .B1(n19490), .B2(n19787), .ZN(
        n19492) );
  OAI211_X1 U22502 ( .C1(n19510), .C2(n19493), .A(n19492), .B(n19624), .ZN(
        n19513) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19513), .B1(
        n19536), .B2(n19573), .ZN(n19494) );
  OAI211_X1 U22504 ( .C1(n19587), .C2(n19516), .A(n19495), .B(n19494), .ZN(
        P2_U3136) );
  AOI22_X1 U22505 ( .A1(n19511), .A2(n19631), .B1(n19630), .B2(n19510), .ZN(
        n19497) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19513), .B1(
        n19536), .B2(n19632), .ZN(n19496) );
  OAI211_X1 U22507 ( .C1(n19635), .C2(n19516), .A(n19497), .B(n19496), .ZN(
        P2_U3137) );
  AOI22_X1 U22508 ( .A1(n19511), .A2(n19637), .B1(n19636), .B2(n19510), .ZN(
        n19499) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19513), .B1(
        n19536), .B2(n19523), .ZN(n19498) );
  OAI211_X1 U22510 ( .C1(n19500), .C2(n19516), .A(n19499), .B(n19498), .ZN(
        P2_U3138) );
  AOI22_X1 U22511 ( .A1(n19511), .A2(n19643), .B1(n19642), .B2(n19510), .ZN(
        n19502) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19513), .B1(
        n19536), .B2(n19644), .ZN(n19501) );
  OAI211_X1 U22513 ( .C1(n19647), .C2(n19516), .A(n19502), .B(n19501), .ZN(
        P2_U3139) );
  AOI22_X1 U22514 ( .A1(n19511), .A2(n19649), .B1(n19648), .B2(n19510), .ZN(
        n19504) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19513), .B1(
        n19536), .B2(n19650), .ZN(n19503) );
  OAI211_X1 U22516 ( .C1(n19653), .C2(n19516), .A(n19504), .B(n19503), .ZN(
        P2_U3140) );
  AOI22_X1 U22517 ( .A1(n19511), .A2(n19655), .B1(n19654), .B2(n19510), .ZN(
        n19506) );
  AOI22_X1 U22518 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19513), .B1(
        n19536), .B2(n19531), .ZN(n19505) );
  OAI211_X1 U22519 ( .C1(n19507), .C2(n19516), .A(n19506), .B(n19505), .ZN(
        P2_U3141) );
  AOI22_X1 U22520 ( .A1(n19511), .A2(n19661), .B1(n19660), .B2(n19510), .ZN(
        n19509) );
  AOI22_X1 U22521 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19513), .B1(
        n19536), .B2(n19662), .ZN(n19508) );
  OAI211_X1 U22522 ( .C1(n19667), .C2(n19516), .A(n19509), .B(n19508), .ZN(
        P2_U3142) );
  AOI22_X1 U22523 ( .A1(n19511), .A2(n19670), .B1(n19668), .B2(n19510), .ZN(
        n19515) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19513), .B1(
        n19536), .B2(n19512), .ZN(n19514) );
  OAI211_X1 U22525 ( .C1(n19517), .C2(n19516), .A(n19515), .B(n19514), .ZN(
        P2_U3143) );
  INV_X1 U22526 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n19520) );
  AOI22_X1 U22527 ( .A1(n19535), .A2(n19619), .B1(n19534), .B2(n19618), .ZN(
        n19519) );
  AOI22_X1 U22528 ( .A1(n19536), .A2(n19626), .B1(n19567), .B2(n19573), .ZN(
        n19518) );
  OAI211_X1 U22529 ( .C1(n19539), .C2(n19520), .A(n19519), .B(n19518), .ZN(
        P2_U3144) );
  AOI22_X1 U22530 ( .A1(n19535), .A2(n19631), .B1(n19534), .B2(n19630), .ZN(
        n19522) );
  AOI22_X1 U22531 ( .A1(n19567), .A2(n19632), .B1(n19536), .B2(n19588), .ZN(
        n19521) );
  OAI211_X1 U22532 ( .C1(n19539), .C2(n13772), .A(n19522), .B(n19521), .ZN(
        P2_U3145) );
  AOI22_X1 U22533 ( .A1(n19535), .A2(n19637), .B1(n19534), .B2(n19636), .ZN(
        n19525) );
  AOI22_X1 U22534 ( .A1(n19567), .A2(n19523), .B1(n19536), .B2(n19638), .ZN(
        n19524) );
  OAI211_X1 U22535 ( .C1(n19539), .C2(n13879), .A(n19525), .B(n19524), .ZN(
        P2_U3146) );
  AOI22_X1 U22536 ( .A1(n19535), .A2(n19643), .B1(n19534), .B2(n19642), .ZN(
        n19527) );
  AOI22_X1 U22537 ( .A1(n19536), .A2(n19556), .B1(n19567), .B2(n19644), .ZN(
        n19526) );
  OAI211_X1 U22538 ( .C1(n19539), .C2(n13912), .A(n19527), .B(n19526), .ZN(
        P2_U3147) );
  AOI22_X1 U22539 ( .A1(n19535), .A2(n19649), .B1(n19534), .B2(n19648), .ZN(
        n19529) );
  AOI22_X1 U22540 ( .A1(n19536), .A2(n19597), .B1(n19567), .B2(n19650), .ZN(
        n19528) );
  OAI211_X1 U22541 ( .C1(n19539), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P2_U3148) );
  AOI22_X1 U22542 ( .A1(n19535), .A2(n19655), .B1(n19534), .B2(n19654), .ZN(
        n19533) );
  AOI22_X1 U22543 ( .A1(n19567), .A2(n19531), .B1(n19536), .B2(n19656), .ZN(
        n19532) );
  OAI211_X1 U22544 ( .C1(n19539), .C2(n13973), .A(n19533), .B(n19532), .ZN(
        P2_U3149) );
  AOI22_X1 U22545 ( .A1(n19535), .A2(n19661), .B1(n19534), .B2(n19660), .ZN(
        n19538) );
  AOI22_X1 U22546 ( .A1(n19567), .A2(n19662), .B1(n19536), .B2(n19603), .ZN(
        n19537) );
  OAI211_X1 U22547 ( .C1(n19539), .C2(n13357), .A(n19538), .B(n19537), .ZN(
        P2_U3150) );
  INV_X1 U22548 ( .A(n13311), .ZN(n19541) );
  NOR2_X1 U22549 ( .A1(n19794), .A2(n19547), .ZN(n19576) );
  NOR3_X1 U22550 ( .A1(n19541), .A2(n19576), .A3(n19390), .ZN(n19546) );
  INV_X1 U22551 ( .A(n19547), .ZN(n19542) );
  AOI21_X1 U22552 ( .B1(n19616), .B2(n19542), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19543) );
  NOR2_X1 U22553 ( .A1(n19546), .A2(n19543), .ZN(n19566) );
  AOI22_X1 U22554 ( .A1(n19566), .A2(n19619), .B1(n19618), .B2(n19576), .ZN(
        n19551) );
  INV_X1 U22555 ( .A(n19544), .ZN(n19620) );
  NAND2_X1 U22556 ( .A1(n19620), .A2(n19545), .ZN(n19548) );
  AOI21_X1 U22557 ( .B1(n19548), .B2(n19547), .A(n19546), .ZN(n19549) );
  OAI211_X1 U22558 ( .C1(n19576), .C2(n19616), .A(n19549), .B(n19624), .ZN(
        n19568) );
  AOI22_X1 U22559 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19626), .ZN(n19550) );
  OAI211_X1 U22560 ( .C1(n19629), .C2(n19596), .A(n19551), .B(n19550), .ZN(
        P2_U3152) );
  AOI22_X1 U22561 ( .A1(n19566), .A2(n19631), .B1(n19630), .B2(n19576), .ZN(
        n19553) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19588), .ZN(n19552) );
  OAI211_X1 U22563 ( .C1(n19591), .C2(n19596), .A(n19553), .B(n19552), .ZN(
        P2_U3153) );
  AOI22_X1 U22564 ( .A1(n19566), .A2(n19637), .B1(n19636), .B2(n19576), .ZN(
        n19555) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19638), .ZN(n19554) );
  OAI211_X1 U22566 ( .C1(n19641), .C2(n19596), .A(n19555), .B(n19554), .ZN(
        P2_U3154) );
  AOI22_X1 U22567 ( .A1(n19566), .A2(n19643), .B1(n19642), .B2(n19576), .ZN(
        n19558) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19556), .ZN(n19557) );
  OAI211_X1 U22569 ( .C1(n19559), .C2(n19596), .A(n19558), .B(n19557), .ZN(
        P2_U3155) );
  AOI22_X1 U22570 ( .A1(n19566), .A2(n19649), .B1(n19648), .B2(n19576), .ZN(
        n19561) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19597), .ZN(n19560) );
  OAI211_X1 U22572 ( .C1(n19600), .C2(n19596), .A(n19561), .B(n19560), .ZN(
        P2_U3156) );
  AOI22_X1 U22573 ( .A1(n19566), .A2(n19655), .B1(n19654), .B2(n19576), .ZN(
        n19563) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19656), .ZN(n19562) );
  OAI211_X1 U22575 ( .C1(n19659), .C2(n19596), .A(n19563), .B(n19562), .ZN(
        P2_U3157) );
  AOI22_X1 U22576 ( .A1(n19566), .A2(n19661), .B1(n19660), .B2(n19576), .ZN(
        n19565) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19603), .ZN(n19564) );
  OAI211_X1 U22578 ( .C1(n19606), .C2(n19596), .A(n19565), .B(n19564), .ZN(
        P2_U3158) );
  AOI22_X1 U22579 ( .A1(n19566), .A2(n19670), .B1(n19668), .B2(n19576), .ZN(
        n19570) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19672), .ZN(n19569) );
  OAI211_X1 U22581 ( .C1(n19678), .C2(n19596), .A(n19570), .B(n19569), .ZN(
        P2_U3159) );
  OR2_X1 U22582 ( .A1(n19770), .A2(n19572), .ZN(n19622) );
  NOR2_X1 U22583 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19622), .ZN(
        n19607) );
  AOI22_X1 U22584 ( .A1(n19673), .A2(n19573), .B1(n19618), .B2(n19607), .ZN(
        n19586) );
  NOR2_X1 U22585 ( .A1(n19673), .A2(n19608), .ZN(n19575) );
  OAI21_X1 U22586 ( .B1(n19575), .B2(n19574), .A(n19771), .ZN(n19584) );
  NOR2_X1 U22587 ( .A1(n19607), .A2(n19576), .ZN(n19583) );
  INV_X1 U22588 ( .A(n19583), .ZN(n19580) );
  INV_X1 U22589 ( .A(n19607), .ZN(n19577) );
  OAI211_X1 U22590 ( .C1(n19578), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19577), 
        .B(n19762), .ZN(n19579) );
  OAI211_X1 U22591 ( .C1(n19584), .C2(n19580), .A(n19624), .B(n19579), .ZN(
        n19610) );
  OAI21_X1 U22592 ( .B1(n19581), .B2(n19607), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19582) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19610), .B1(
        n19619), .B2(n19609), .ZN(n19585) );
  OAI211_X1 U22594 ( .C1(n19587), .C2(n19596), .A(n19586), .B(n19585), .ZN(
        P2_U3160) );
  AOI22_X1 U22595 ( .A1(n19608), .A2(n19588), .B1(n19630), .B2(n19607), .ZN(
        n19590) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19610), .B1(
        n19631), .B2(n19609), .ZN(n19589) );
  OAI211_X1 U22597 ( .C1(n19591), .C2(n19666), .A(n19590), .B(n19589), .ZN(
        P2_U3161) );
  AOI22_X1 U22598 ( .A1(n19608), .A2(n19638), .B1(n19636), .B2(n19607), .ZN(
        n19593) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19610), .B1(
        n19637), .B2(n19609), .ZN(n19592) );
  OAI211_X1 U22600 ( .C1(n19641), .C2(n19666), .A(n19593), .B(n19592), .ZN(
        P2_U3162) );
  AOI22_X1 U22601 ( .A1(n19673), .A2(n19644), .B1(n19607), .B2(n19642), .ZN(
        n19595) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19610), .B1(
        n19643), .B2(n19609), .ZN(n19594) );
  OAI211_X1 U22603 ( .C1(n19647), .C2(n19596), .A(n19595), .B(n19594), .ZN(
        P2_U3163) );
  AOI22_X1 U22604 ( .A1(n19608), .A2(n19597), .B1(n19607), .B2(n19648), .ZN(
        n19599) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19610), .B1(
        n19649), .B2(n19609), .ZN(n19598) );
  OAI211_X1 U22606 ( .C1(n19600), .C2(n19666), .A(n19599), .B(n19598), .ZN(
        P2_U3164) );
  AOI22_X1 U22607 ( .A1(n19608), .A2(n19656), .B1(n19607), .B2(n19654), .ZN(
        n19602) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19610), .B1(
        n19655), .B2(n19609), .ZN(n19601) );
  OAI211_X1 U22609 ( .C1(n19659), .C2(n19666), .A(n19602), .B(n19601), .ZN(
        P2_U3165) );
  AOI22_X1 U22610 ( .A1(n19608), .A2(n19603), .B1(n19607), .B2(n19660), .ZN(
        n19605) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19610), .B1(
        n19661), .B2(n19609), .ZN(n19604) );
  OAI211_X1 U22612 ( .C1(n19606), .C2(n19666), .A(n19605), .B(n19604), .ZN(
        P2_U3166) );
  AOI22_X1 U22613 ( .A1(n19608), .A2(n19672), .B1(n19668), .B2(n19607), .ZN(
        n19612) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19610), .B1(
        n19670), .B2(n19609), .ZN(n19611) );
  OAI211_X1 U22615 ( .C1(n19678), .C2(n19666), .A(n19612), .B(n19611), .ZN(
        P2_U3167) );
  INV_X1 U22616 ( .A(n19613), .ZN(n19614) );
  NOR3_X1 U22617 ( .A1(n19614), .A2(n19669), .A3(n19390), .ZN(n19621) );
  INV_X1 U22618 ( .A(n19622), .ZN(n19615) );
  AOI21_X1 U22619 ( .B1(n19616), .B2(n19615), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19617) );
  NOR2_X1 U22620 ( .A1(n19621), .A2(n19617), .ZN(n19671) );
  AOI22_X1 U22621 ( .A1(n19671), .A2(n19619), .B1(n19669), .B2(n19618), .ZN(
        n19628) );
  NAND2_X1 U22622 ( .A1(n19620), .A2(n19763), .ZN(n19623) );
  AOI21_X1 U22623 ( .B1(n19623), .B2(n19622), .A(n19621), .ZN(n19625) );
  OAI211_X1 U22624 ( .C1(n19669), .C2(n19616), .A(n19625), .B(n19624), .ZN(
        n19674) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19674), .B1(
        n19673), .B2(n19626), .ZN(n19627) );
  OAI211_X1 U22626 ( .C1(n19629), .C2(n19677), .A(n19628), .B(n19627), .ZN(
        P2_U3168) );
  AOI22_X1 U22627 ( .A1(n19671), .A2(n19631), .B1(n19669), .B2(n19630), .ZN(
        n19634) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19674), .B1(
        n19663), .B2(n19632), .ZN(n19633) );
  OAI211_X1 U22629 ( .C1(n19635), .C2(n19666), .A(n19634), .B(n19633), .ZN(
        P2_U3169) );
  AOI22_X1 U22630 ( .A1(n19671), .A2(n19637), .B1(n19669), .B2(n19636), .ZN(
        n19640) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19674), .B1(
        n19673), .B2(n19638), .ZN(n19639) );
  OAI211_X1 U22632 ( .C1(n19641), .C2(n19677), .A(n19640), .B(n19639), .ZN(
        P2_U3170) );
  AOI22_X1 U22633 ( .A1(n19671), .A2(n19643), .B1(n19669), .B2(n19642), .ZN(
        n19646) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19674), .B1(
        n19663), .B2(n19644), .ZN(n19645) );
  OAI211_X1 U22635 ( .C1(n19647), .C2(n19666), .A(n19646), .B(n19645), .ZN(
        P2_U3171) );
  AOI22_X1 U22636 ( .A1(n19671), .A2(n19649), .B1(n19669), .B2(n19648), .ZN(
        n19652) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19674), .B1(
        n19663), .B2(n19650), .ZN(n19651) );
  OAI211_X1 U22638 ( .C1(n19653), .C2(n19666), .A(n19652), .B(n19651), .ZN(
        P2_U3172) );
  AOI22_X1 U22639 ( .A1(n19671), .A2(n19655), .B1(n19669), .B2(n19654), .ZN(
        n19658) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19674), .B1(
        n19673), .B2(n19656), .ZN(n19657) );
  OAI211_X1 U22641 ( .C1(n19659), .C2(n19677), .A(n19658), .B(n19657), .ZN(
        P2_U3173) );
  AOI22_X1 U22642 ( .A1(n19671), .A2(n19661), .B1(n19669), .B2(n19660), .ZN(
        n19665) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19674), .B1(
        n19663), .B2(n19662), .ZN(n19664) );
  OAI211_X1 U22644 ( .C1(n19667), .C2(n19666), .A(n19665), .B(n19664), .ZN(
        P2_U3174) );
  AOI22_X1 U22645 ( .A1(n19671), .A2(n19670), .B1(n19669), .B2(n19668), .ZN(
        n19676) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19674), .B1(
        n19673), .B2(n19672), .ZN(n19675) );
  OAI211_X1 U22647 ( .C1(n19678), .C2(n19677), .A(n19676), .B(n19675), .ZN(
        P2_U3175) );
  INV_X1 U22648 ( .A(P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20858) );
  NOR2_X1 U22649 ( .A1(n20858), .A2(n19753), .ZN(P2_U3179) );
  AND2_X1 U22650 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19679), .ZN(
        P2_U3180) );
  AND2_X1 U22651 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19679), .ZN(
        P2_U3181) );
  AND2_X1 U22652 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19679), .ZN(
        P2_U3182) );
  AND2_X1 U22653 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19679), .ZN(
        P2_U3183) );
  AND2_X1 U22654 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19679), .ZN(
        P2_U3184) );
  AND2_X1 U22655 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19679), .ZN(
        P2_U3185) );
  AND2_X1 U22656 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19679), .ZN(
        P2_U3186) );
  AND2_X1 U22657 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19679), .ZN(
        P2_U3187) );
  AND2_X1 U22658 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19679), .ZN(
        P2_U3188) );
  NOR2_X1 U22659 ( .A1(n20911), .A2(n19753), .ZN(P2_U3189) );
  AND2_X1 U22660 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19679), .ZN(
        P2_U3190) );
  NOR2_X1 U22661 ( .A1(n20910), .A2(n19753), .ZN(P2_U3191) );
  AND2_X1 U22662 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19679), .ZN(
        P2_U3192) );
  AND2_X1 U22663 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19679), .ZN(
        P2_U3193) );
  AND2_X1 U22664 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19679), .ZN(
        P2_U3194) );
  AND2_X1 U22665 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19679), .ZN(
        P2_U3195) );
  AND2_X1 U22666 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19679), .ZN(
        P2_U3196) );
  AND2_X1 U22667 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19679), .ZN(
        P2_U3197) );
  AND2_X1 U22668 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19679), .ZN(
        P2_U3198) );
  AND2_X1 U22669 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19679), .ZN(
        P2_U3199) );
  INV_X1 U22670 ( .A(P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21046) );
  NOR2_X1 U22671 ( .A1(n21046), .A2(n19753), .ZN(P2_U3200) );
  AND2_X1 U22672 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19679), .ZN(P2_U3201) );
  AND2_X1 U22673 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19679), .ZN(P2_U3202) );
  AND2_X1 U22674 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19679), .ZN(P2_U3203) );
  AND2_X1 U22675 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19679), .ZN(P2_U3204) );
  AND2_X1 U22676 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19679), .ZN(P2_U3205) );
  AND2_X1 U22677 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19679), .ZN(P2_U3206) );
  AND2_X1 U22678 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19679), .ZN(P2_U3207) );
  AND2_X1 U22679 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19679), .ZN(P2_U3208) );
  NAND2_X1 U22680 ( .A1(n20742), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19682) );
  NAND2_X1 U22681 ( .A1(n19680), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19689) );
  OAI211_X1 U22682 ( .C1(n19683), .C2(n19682), .A(n19689), .B(n19681), .ZN(
        n19684) );
  INV_X1 U22683 ( .A(n19684), .ZN(n19686) );
  NAND3_X1 U22684 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19694), .A3(
        n19688), .ZN(n19685) );
  OAI211_X1 U22685 ( .C1(n19687), .C2(n20742), .A(n19686), .B(n19685), .ZN(
        P2_U3210) );
  NAND2_X1 U22686 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19689), .ZN(n20744) );
  NOR2_X1 U22687 ( .A1(HOLD), .A2(n20744), .ZN(n19693) );
  OAI21_X1 U22688 ( .B1(n19688), .B2(n20986), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20745) );
  OAI22_X1 U22689 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19690), .B1(NA), 
        .B2(n19689), .ZN(n19691) );
  OAI211_X1 U22690 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19691), .ZN(n19692) );
  OAI21_X1 U22691 ( .B1(n19693), .B2(n20745), .A(n19692), .ZN(P2_U3211) );
  OAI222_X1 U22692 ( .A1(n19741), .A2(n19696), .B1(n19695), .B2(n20740), .C1(
        n19697), .C2(n19743), .ZN(P2_U3212) );
  OAI222_X1 U22693 ( .A1(n19743), .A2(n12199), .B1(n19698), .B2(n20740), .C1(
        n19697), .C2(n19741), .ZN(P2_U3213) );
  OAI222_X1 U22694 ( .A1(n19743), .A2(n12179), .B1(n19699), .B2(n20740), .C1(
        n12199), .C2(n19741), .ZN(P2_U3214) );
  OAI222_X1 U22695 ( .A1(n19743), .A2(n15380), .B1(n19700), .B2(n20740), .C1(
        n12179), .C2(n19741), .ZN(P2_U3215) );
  OAI222_X1 U22696 ( .A1(n19743), .A2(n19702), .B1(n19701), .B2(n20740), .C1(
        n15380), .C2(n19741), .ZN(P2_U3216) );
  OAI222_X1 U22697 ( .A1(n19743), .A2(n19703), .B1(n20918), .B2(n20740), .C1(
        n19702), .C2(n19741), .ZN(P2_U3217) );
  OAI222_X1 U22698 ( .A1(n19743), .A2(n12293), .B1(n19704), .B2(n20740), .C1(
        n19703), .C2(n19741), .ZN(P2_U3218) );
  OAI222_X1 U22699 ( .A1(n19743), .A2(n12364), .B1(n19705), .B2(n20740), .C1(
        n12293), .C2(n19741), .ZN(P2_U3219) );
  OAI222_X1 U22700 ( .A1(n19743), .A2(n12540), .B1(n19706), .B2(n20740), .C1(
        n12364), .C2(n19741), .ZN(P2_U3220) );
  OAI222_X1 U22701 ( .A1(n19743), .A2(n20894), .B1(n19707), .B2(n20740), .C1(
        n12540), .C2(n19741), .ZN(P2_U3221) );
  OAI222_X1 U22702 ( .A1(n19743), .A2(n12628), .B1(n19708), .B2(n20740), .C1(
        n20894), .C2(n19741), .ZN(P2_U3222) );
  OAI222_X1 U22703 ( .A1(n19743), .A2(n18834), .B1(n19709), .B2(n20740), .C1(
        n12628), .C2(n19741), .ZN(P2_U3223) );
  OAI222_X1 U22704 ( .A1(n19743), .A2(n12774), .B1(n19710), .B2(n20740), .C1(
        n18834), .C2(n19741), .ZN(P2_U3224) );
  OAI222_X1 U22705 ( .A1(n19743), .A2(n15012), .B1(n19711), .B2(n20740), .C1(
        n12774), .C2(n19741), .ZN(P2_U3225) );
  OAI222_X1 U22706 ( .A1(n19743), .A2(n19713), .B1(n19712), .B2(n20740), .C1(
        n15012), .C2(n19741), .ZN(P2_U3226) );
  OAI222_X1 U22707 ( .A1(n19743), .A2(n19715), .B1(n19714), .B2(n20740), .C1(
        n19713), .C2(n19741), .ZN(P2_U3227) );
  OAI222_X1 U22708 ( .A1(n19743), .A2(n19717), .B1(n19716), .B2(n20740), .C1(
        n19715), .C2(n19741), .ZN(P2_U3228) );
  OAI222_X1 U22709 ( .A1(n19743), .A2(n19719), .B1(n19718), .B2(n20740), .C1(
        n19717), .C2(n19741), .ZN(P2_U3229) );
  OAI222_X1 U22710 ( .A1(n19743), .A2(n19721), .B1(n19720), .B2(n20740), .C1(
        n19719), .C2(n19741), .ZN(P2_U3230) );
  OAI222_X1 U22711 ( .A1(n19743), .A2(n19723), .B1(n19722), .B2(n20740), .C1(
        n19721), .C2(n19741), .ZN(P2_U3231) );
  OAI222_X1 U22712 ( .A1(n19743), .A2(n19725), .B1(n19724), .B2(n20740), .C1(
        n19723), .C2(n19741), .ZN(P2_U3232) );
  OAI222_X1 U22713 ( .A1(n19743), .A2(n19727), .B1(n19726), .B2(n20740), .C1(
        n19725), .C2(n19741), .ZN(P2_U3233) );
  OAI222_X1 U22714 ( .A1(n19743), .A2(n19729), .B1(n19728), .B2(n20740), .C1(
        n19727), .C2(n19741), .ZN(P2_U3234) );
  OAI222_X1 U22715 ( .A1(n19743), .A2(n19731), .B1(n19730), .B2(n20740), .C1(
        n19729), .C2(n19741), .ZN(P2_U3235) );
  OAI222_X1 U22716 ( .A1(n19743), .A2(n19733), .B1(n19732), .B2(n20740), .C1(
        n19731), .C2(n19741), .ZN(P2_U3236) );
  OAI222_X1 U22717 ( .A1(n19743), .A2(n19736), .B1(n19734), .B2(n20740), .C1(
        n19733), .C2(n19741), .ZN(P2_U3237) );
  OAI222_X1 U22718 ( .A1(n19741), .A2(n19736), .B1(n19735), .B2(n20740), .C1(
        n19737), .C2(n19743), .ZN(P2_U3238) );
  OAI222_X1 U22719 ( .A1(n19743), .A2(n19739), .B1(n19738), .B2(n20740), .C1(
        n19737), .C2(n19741), .ZN(P2_U3239) );
  INV_X1 U22720 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n21028) );
  OAI222_X1 U22721 ( .A1(n19743), .A2(n21028), .B1(n19740), .B2(n20740), .C1(
        n19739), .C2(n19741), .ZN(P2_U3240) );
  INV_X1 U22722 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n21037) );
  OAI222_X1 U22723 ( .A1(n19743), .A2(n21037), .B1(n19742), .B2(n20740), .C1(
        n21028), .C2(n19741), .ZN(P2_U3241) );
  INV_X1 U22724 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U22725 ( .A1(n20740), .A2(n19745), .B1(n19744), .B2(n19806), .ZN(
        P2_U3585) );
  MUX2_X1 U22726 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20740), .Z(P2_U3586) );
  INV_X1 U22727 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U22728 ( .A1(n20740), .A2(n19747), .B1(n19746), .B2(n19806), .ZN(
        P2_U3587) );
  INV_X1 U22729 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19748) );
  AOI22_X1 U22730 ( .A1(n20740), .A2(n19749), .B1(n19748), .B2(n19806), .ZN(
        P2_U3588) );
  OAI21_X1 U22731 ( .B1(n19753), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19751), 
        .ZN(n19750) );
  INV_X1 U22732 ( .A(n19750), .ZN(P2_U3591) );
  OAI21_X1 U22733 ( .B1(n19753), .B2(n19752), .A(n19751), .ZN(P2_U3592) );
  INV_X1 U22734 ( .A(n19754), .ZN(n19755) );
  OAI222_X1 U22735 ( .A1(n19772), .A2(n19759), .B1(n19758), .B2(n19757), .C1(
        n19756), .C2(n19755), .ZN(n19761) );
  MUX2_X1 U22736 ( .A(n19761), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19760), .Z(P2_U3599) );
  AOI21_X1 U22737 ( .B1(n19763), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19762), 
        .ZN(n19765) );
  OR2_X1 U22738 ( .A1(n19765), .A2(n19764), .ZN(n19774) );
  AOI222_X1 U22739 ( .A1(n19774), .A2(n19768), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19767), .C1(n19771), .C2(n19766), .ZN(n19769) );
  AOI22_X1 U22740 ( .A1(n19795), .A2(n19770), .B1(n19769), .B2(n19792), .ZN(
        P2_U3602) );
  NAND2_X1 U22741 ( .A1(n19771), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19782) );
  OAI21_X1 U22742 ( .B1(n19780), .B2(n19782), .A(n19772), .ZN(n19773) );
  AOI22_X1 U22743 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19775), .B1(n19774), 
        .B2(n19773), .ZN(n19776) );
  AOI22_X1 U22744 ( .A1(n19795), .A2(n19777), .B1(n19776), .B2(n19792), .ZN(
        P2_U3603) );
  INV_X1 U22745 ( .A(n19790), .ZN(n19779) );
  AND2_X1 U22746 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19778) );
  OR3_X1 U22747 ( .A1(n19780), .A2(n19779), .A3(n19778), .ZN(n19781) );
  OAI21_X1 U22748 ( .B1(n19783), .B2(n19782), .A(n19781), .ZN(n19784) );
  AOI21_X1 U22749 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19785), .A(n19784), 
        .ZN(n19786) );
  AOI22_X1 U22750 ( .A1(n19795), .A2(n19787), .B1(n19786), .B2(n19792), .ZN(
        P2_U3604) );
  NOR2_X1 U22751 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19616), .ZN(
        n19789) );
  AOI211_X1 U22752 ( .C1(n19791), .C2(n19790), .A(n19789), .B(n19788), .ZN(
        n19793) );
  AOI22_X1 U22753 ( .A1(n19795), .A2(n19794), .B1(n19793), .B2(n19792), .ZN(
        P2_U3605) );
  INV_X1 U22754 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20813) );
  AOI22_X1 U22755 ( .A1(n20740), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20813), 
        .B2(n19806), .ZN(P2_U3608) );
  INV_X1 U22756 ( .A(n19796), .ZN(n19800) );
  INV_X1 U22757 ( .A(n19797), .ZN(n19799) );
  OAI22_X1 U22758 ( .A1(n19801), .A2(n19800), .B1(n19799), .B2(n19798), .ZN(
        n19803) );
  OAI21_X1 U22759 ( .B1(n19803), .B2(n19802), .A(n19805), .ZN(n19804) );
  OAI21_X1 U22760 ( .B1(n19805), .B2(n12705), .A(n19804), .ZN(P2_U3609) );
  INV_X1 U22761 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n19807) );
  AOI22_X1 U22762 ( .A1(n20740), .A2(n19808), .B1(n19807), .B2(n19806), .ZN(
        P2_U3611) );
  AND2_X1 U22763 ( .A1(n20634), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n19810) );
  INV_X1 U22764 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19809) );
  NAND2_X1 U22765 ( .A1(n20630), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20736) );
  AOI21_X1 U22766 ( .B1(n19810), .B2(n19809), .A(n20667), .ZN(P1_U2802) );
  OAI21_X1 U22767 ( .B1(n19812), .B2(n19811), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19813) );
  OAI21_X1 U22768 ( .B1(n19814), .B2(n10081), .A(n19813), .ZN(P1_U2803) );
  NOR2_X1 U22769 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19816) );
  OAI21_X1 U22770 ( .B1(n19816), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20736), .ZN(
        n19815) );
  OAI21_X1 U22771 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20736), .A(n19815), 
        .ZN(P1_U2804) );
  AOI21_X1 U22772 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20634), .A(n20739), 
        .ZN(n20703) );
  OAI21_X1 U22773 ( .B1(BS16), .B2(n19816), .A(n20703), .ZN(n20701) );
  OAI21_X1 U22774 ( .B1(n20703), .B2(n20207), .A(n20701), .ZN(P1_U2805) );
  OAI21_X1 U22775 ( .B1(n19819), .B2(n19818), .A(n19817), .ZN(P1_U2806) );
  NOR4_X1 U22776 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19829) );
  NOR4_X1 U22777 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_6__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19828) );
  INV_X1 U22778 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20702) );
  INV_X1 U22779 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20700) );
  NOR4_X1 U22780 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_2__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19820) );
  OAI21_X1 U22781 ( .B1(n20702), .B2(n20700), .A(n19820), .ZN(n19826) );
  NOR4_X1 U22782 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19824) );
  NOR4_X1 U22783 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19823) );
  NOR4_X1 U22784 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19822) );
  NOR4_X1 U22785 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19821) );
  NAND4_X1 U22786 ( .A1(n19824), .A2(n19823), .A3(n19822), .A4(n19821), .ZN(
        n19825) );
  NOR4_X1 U22787 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(n19826), .A4(n19825), .ZN(n19827)
         );
  NAND3_X1 U22788 ( .A1(n19829), .A2(n19828), .A3(n19827), .ZN(n20720) );
  NOR2_X1 U22789 ( .A1(n20720), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20722) );
  NAND3_X1 U22790 ( .A1(n20721), .A2(n20702), .A3(n20700), .ZN(n19831) );
  INV_X1 U22791 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20696) );
  AOI22_X1 U22792 ( .A1(n20722), .A2(n19831), .B1(n20696), .B2(n20720), .ZN(
        P1_U2807) );
  AOI22_X1 U22793 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(n20720), .B1(n20722), .B2(n20702), .ZN(n19830) );
  OAI21_X1 U22794 ( .B1(n20720), .B2(n19831), .A(n19830), .ZN(P1_U2808) );
  NAND2_X1 U22795 ( .A1(n19885), .A2(n19832), .ZN(n19852) );
  AOI22_X1 U22796 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(n19901), .B1(n19880), .B2(
        n19907), .ZN(n19833) );
  OAI21_X1 U22797 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n19834), .A(n19833), .ZN(
        n19835) );
  AOI211_X1 U22798 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n19895), .B(n19835), .ZN(n19840) );
  INV_X1 U22799 ( .A(n19836), .ZN(n19909) );
  AOI22_X1 U22800 ( .A1(n19909), .A2(n19873), .B1(n19838), .B2(n19837), .ZN(
        n19839) );
  OAI211_X1 U22801 ( .C1(n13104), .C2(n19852), .A(n19840), .B(n19839), .ZN(
        P1_U2831) );
  AOI21_X1 U22802 ( .B1(n19897), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n19895), .ZN(n19843) );
  NAND3_X1 U22803 ( .A1(n19878), .A2(n19841), .A3(n21024), .ZN(n19842) );
  OAI211_X1 U22804 ( .C1(n19844), .C2(n19892), .A(n19843), .B(n19842), .ZN(
        n19845) );
  AOI21_X1 U22805 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n19901), .A(n19845), .ZN(
        n19851) );
  OAI22_X1 U22806 ( .A1(n19848), .A2(n19847), .B1(n19846), .B2(n19906), .ZN(
        n19849) );
  INV_X1 U22807 ( .A(n19849), .ZN(n19850) );
  OAI211_X1 U22808 ( .C1(n21024), .C2(n19852), .A(n19851), .B(n19850), .ZN(
        P1_U2832) );
  NAND2_X1 U22809 ( .A1(n19878), .A2(n20654), .ZN(n19853) );
  OAI22_X1 U22810 ( .A1(n19892), .A2(n19855), .B1(n19854), .B2(n19853), .ZN(
        n19856) );
  AOI211_X1 U22811 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19895), .B(n19856), .ZN(n19863) );
  NAND2_X1 U22812 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19858) );
  NAND2_X1 U22813 ( .A1(n19877), .A2(n19857), .ZN(n19886) );
  OAI21_X1 U22814 ( .B1(n19858), .B2(n19886), .A(n19885), .ZN(n19870) );
  OAI22_X1 U22815 ( .A1(n19906), .A2(n19859), .B1(n19870), .B2(n20654), .ZN(
        n19860) );
  AOI21_X1 U22816 ( .B1(n19873), .B2(n19861), .A(n19860), .ZN(n19862) );
  OAI211_X1 U22817 ( .C1(n19864), .C2(n19866), .A(n19863), .B(n19862), .ZN(
        P1_U2833) );
  NAND3_X1 U22818 ( .A1(n19878), .A2(n19877), .A3(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19871) );
  OAI22_X1 U22819 ( .A1(n19867), .A2(n19866), .B1(n19892), .B2(n19865), .ZN(
        n19868) );
  AOI211_X1 U22820 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19895), .B(n19868), .ZN(n19869) );
  OAI221_X1 U22821 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n19871), .C1(n13022), 
        .C2(n19870), .A(n19869), .ZN(n19872) );
  AOI21_X1 U22822 ( .B1(n19874), .B2(n19873), .A(n19872), .ZN(n19875) );
  OAI21_X1 U22823 ( .B1(n19876), .B2(n19906), .A(n19875), .ZN(P1_U2834) );
  NAND2_X1 U22824 ( .A1(n19878), .A2(n19877), .ZN(n19882) );
  AOI22_X1 U22825 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(n19901), .B1(n19880), .B2(
        n19879), .ZN(n19881) );
  OAI21_X1 U22826 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n19882), .A(n19881), .ZN(
        n19883) );
  AOI211_X1 U22827 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n19895), .B(n19883), .ZN(n19888) );
  INV_X1 U22828 ( .A(n19884), .ZN(n19903) );
  AND2_X1 U22829 ( .A1(n19886), .A2(n19885), .ZN(n19902) );
  AOI22_X1 U22830 ( .A1(n19903), .A2(n19916), .B1(n19902), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n19887) );
  OAI211_X1 U22831 ( .C1(n19889), .C2(n19906), .A(n19888), .B(n19887), .ZN(
        P1_U2835) );
  NOR3_X1 U22832 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19891), .A3(n19890), .ZN(
        n19900) );
  OAI22_X1 U22833 ( .A1(n19894), .A2(n19893), .B1(n19892), .B2(n20004), .ZN(
        n19896) );
  AOI211_X1 U22834 ( .C1(n19897), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19896), .B(n19895), .ZN(n19898) );
  INV_X1 U22835 ( .A(n19898), .ZN(n19899) );
  AOI211_X1 U22836 ( .C1(n19901), .C2(P1_EBX_REG_4__SCAN_IN), .A(n19900), .B(
        n19899), .ZN(n19905) );
  AOI22_X1 U22837 ( .A1(n19903), .A2(n19992), .B1(P1_REIP_REG_4__SCAN_IN), 
        .B2(n19902), .ZN(n19904) );
  OAI211_X1 U22838 ( .C1(n19997), .C2(n19906), .A(n19905), .B(n19904), .ZN(
        P1_U2836) );
  AOI22_X1 U22839 ( .A1(n19909), .A2(n19915), .B1(n19908), .B2(n19907), .ZN(
        n19910) );
  OAI21_X1 U22840 ( .B1(n19919), .B2(n19911), .A(n19910), .ZN(P1_U2863) );
  NOR2_X1 U22841 ( .A1(n19913), .A2(n19912), .ZN(n19914) );
  AOI21_X1 U22842 ( .B1(n19916), .B2(n19915), .A(n19914), .ZN(n19917) );
  OAI21_X1 U22843 ( .B1(n19919), .B2(n19918), .A(n19917), .ZN(P1_U2867) );
  INV_X1 U22844 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n19923) );
  INV_X1 U22845 ( .A(n19920), .ZN(n19921) );
  AOI22_X1 U22846 ( .A1(n19921), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20727), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n19922) );
  OAI21_X1 U22847 ( .B1(n19923), .B2(n19925), .A(n19922), .ZN(P1_U2906) );
  OAI222_X1 U22848 ( .A1(n19928), .A2(n19927), .B1(n19952), .B2(n19926), .C1(
        n19925), .C2(n19924), .ZN(P1_U2921) );
  AOI22_X1 U22849 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19929) );
  OAI21_X1 U22850 ( .B1(n14272), .B2(n19952), .A(n19929), .ZN(P1_U2922) );
  AOI22_X1 U22851 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19930) );
  OAI21_X1 U22852 ( .B1(n13142), .B2(n19952), .A(n19930), .ZN(P1_U2923) );
  INV_X1 U22853 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n19932) );
  AOI22_X1 U22854 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19931) );
  OAI21_X1 U22855 ( .B1(n19932), .B2(n19952), .A(n19931), .ZN(P1_U2924) );
  AOI22_X1 U22856 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19933) );
  OAI21_X1 U22857 ( .B1(n13117), .B2(n19952), .A(n19933), .ZN(P1_U2925) );
  AOI22_X1 U22858 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19934) );
  OAI21_X1 U22859 ( .B1(n13101), .B2(n19952), .A(n19934), .ZN(P1_U2926) );
  INV_X1 U22860 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n19936) );
  AOI22_X1 U22861 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19935) );
  OAI21_X1 U22862 ( .B1(n19936), .B2(n19952), .A(n19935), .ZN(P1_U2927) );
  AOI22_X1 U22863 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19937) );
  OAI21_X1 U22864 ( .B1(n13079), .B2(n19952), .A(n19937), .ZN(P1_U2928) );
  AOI22_X1 U22865 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19938) );
  OAI21_X1 U22866 ( .B1(n10615), .B2(n19952), .A(n19938), .ZN(P1_U2929) );
  AOI22_X1 U22867 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19939) );
  OAI21_X1 U22868 ( .B1(n10679), .B2(n19952), .A(n19939), .ZN(P1_U2930) );
  AOI22_X1 U22869 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19940) );
  OAI21_X1 U22870 ( .B1(n19941), .B2(n19952), .A(n19940), .ZN(P1_U2931) );
  AOI22_X1 U22871 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19942) );
  OAI21_X1 U22872 ( .B1(n19943), .B2(n19952), .A(n19942), .ZN(P1_U2932) );
  AOI22_X1 U22873 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19944) );
  OAI21_X1 U22874 ( .B1(n19945), .B2(n19952), .A(n19944), .ZN(P1_U2933) );
  AOI22_X1 U22875 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19946) );
  OAI21_X1 U22876 ( .B1(n19947), .B2(n19952), .A(n19946), .ZN(P1_U2934) );
  AOI22_X1 U22877 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19948) );
  OAI21_X1 U22878 ( .B1(n19949), .B2(n19952), .A(n19948), .ZN(P1_U2935) );
  AOI22_X1 U22879 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20727), .B1(n19950), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19951) );
  OAI21_X1 U22880 ( .B1(n19953), .B2(n19952), .A(n19951), .ZN(P1_U2936) );
  AOI22_X1 U22881 ( .A1(n19983), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n9795), .ZN(n19956) );
  INV_X1 U22882 ( .A(n19954), .ZN(n19955) );
  NAND2_X1 U22883 ( .A1(n19969), .A2(n19955), .ZN(n19971) );
  NAND2_X1 U22884 ( .A1(n19956), .A2(n19971), .ZN(P1_U2945) );
  AOI22_X1 U22885 ( .A1(n19983), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n9795), .ZN(n19958) );
  NAND2_X1 U22886 ( .A1(n19969), .A2(n19957), .ZN(n19973) );
  NAND2_X1 U22887 ( .A1(n19958), .A2(n19973), .ZN(P1_U2946) );
  AOI22_X1 U22888 ( .A1(n19959), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n9795), .ZN(n19962) );
  INV_X1 U22889 ( .A(n19960), .ZN(n19961) );
  NAND2_X1 U22890 ( .A1(n19969), .A2(n19961), .ZN(n19975) );
  NAND2_X1 U22891 ( .A1(n19962), .A2(n19975), .ZN(P1_U2947) );
  AOI22_X1 U22892 ( .A1(n19983), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n9795), .ZN(n19964) );
  NAND2_X1 U22893 ( .A1(n19969), .A2(n19963), .ZN(n19977) );
  NAND2_X1 U22894 ( .A1(n19964), .A2(n19977), .ZN(P1_U2948) );
  AOI22_X1 U22895 ( .A1(n19983), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n9795), .ZN(n19966) );
  NAND2_X1 U22896 ( .A1(n19969), .A2(n19965), .ZN(n19979) );
  NAND2_X1 U22897 ( .A1(n19966), .A2(n19979), .ZN(P1_U2949) );
  AOI22_X1 U22898 ( .A1(n19983), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n9795), .ZN(n19970) );
  INV_X1 U22899 ( .A(n19967), .ZN(n19968) );
  NAND2_X1 U22900 ( .A1(n19969), .A2(n19968), .ZN(n19984) );
  NAND2_X1 U22901 ( .A1(n19970), .A2(n19984), .ZN(P1_U2951) );
  AOI22_X1 U22902 ( .A1(n19983), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n9795), .ZN(n19972) );
  NAND2_X1 U22903 ( .A1(n19972), .A2(n19971), .ZN(P1_U2960) );
  AOI22_X1 U22904 ( .A1(n19983), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n9795), .ZN(n19974) );
  NAND2_X1 U22905 ( .A1(n19974), .A2(n19973), .ZN(P1_U2961) );
  AOI22_X1 U22906 ( .A1(n19983), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n9795), .ZN(n19976) );
  NAND2_X1 U22907 ( .A1(n19976), .A2(n19975), .ZN(P1_U2962) );
  AOI22_X1 U22908 ( .A1(n19983), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n9795), .ZN(n19978) );
  NAND2_X1 U22909 ( .A1(n19978), .A2(n19977), .ZN(P1_U2963) );
  AOI22_X1 U22910 ( .A1(n19983), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n9795), .ZN(n19980) );
  NAND2_X1 U22911 ( .A1(n19980), .A2(n19979), .ZN(P1_U2964) );
  AOI22_X1 U22912 ( .A1(n19983), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n9795), .ZN(n19982) );
  NAND2_X1 U22913 ( .A1(n19982), .A2(n19981), .ZN(P1_U2965) );
  AOI22_X1 U22914 ( .A1(n19983), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n9795), .ZN(n19985) );
  NAND2_X1 U22915 ( .A1(n19985), .A2(n19984), .ZN(P1_U2966) );
  AOI22_X1 U22916 ( .A1(n19987), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19986), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19996) );
  OAI21_X1 U22917 ( .B1(n19990), .B2(n19989), .A(n19988), .ZN(n19991) );
  INV_X1 U22918 ( .A(n19991), .ZN(n20008) );
  AOI22_X1 U22919 ( .A1(n20008), .A2(n19994), .B1(n19993), .B2(n19992), .ZN(
        n19995) );
  OAI211_X1 U22920 ( .C1(n19998), .C2(n19997), .A(n19996), .B(n19995), .ZN(
        P1_U2995) );
  NOR2_X1 U22921 ( .A1(n20024), .A2(n19999), .ZN(n20026) );
  OAI21_X1 U22922 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20001), .A(
        n20000), .ZN(n20032) );
  AOI211_X1 U22923 ( .C1(n20036), .C2(n20035), .A(n20026), .B(n20032), .ZN(
        n20020) );
  OAI22_X1 U22924 ( .A1(n20004), .A2(n20003), .B1(n20647), .B2(n20002), .ZN(
        n20007) );
  AOI211_X1 U22925 ( .C1(n20010), .C2(n20019), .A(n20014), .B(n20005), .ZN(
        n20006) );
  AOI211_X1 U22926 ( .C1(n20008), .C2(n20031), .A(n20007), .B(n20006), .ZN(
        n20009) );
  OAI21_X1 U22927 ( .B1(n20020), .B2(n20010), .A(n20009), .ZN(P1_U3027) );
  INV_X1 U22928 ( .A(n20011), .ZN(n20013) );
  AOI21_X1 U22929 ( .B1(n20013), .B2(n20027), .A(n20012), .ZN(n20018) );
  INV_X1 U22930 ( .A(n20014), .ZN(n20015) );
  AOI22_X1 U22931 ( .A1(n20016), .A2(n20031), .B1(n20019), .B2(n20015), .ZN(
        n20017) );
  OAI211_X1 U22932 ( .C1(n20020), .C2(n20019), .A(n20018), .B(n20017), .ZN(
        P1_U3028) );
  INV_X1 U22933 ( .A(n20021), .ZN(n20028) );
  NOR4_X1 U22934 ( .A1(n20024), .A2(n20023), .A3(n20036), .A4(n20022), .ZN(
        n20025) );
  AOI211_X1 U22935 ( .C1(n20028), .C2(n20027), .A(n20026), .B(n20025), .ZN(
        n20040) );
  INV_X1 U22936 ( .A(n20029), .ZN(n20030) );
  AOI22_X1 U22937 ( .A1(n20032), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20031), .B2(n20030), .ZN(n20039) );
  NAND2_X1 U22938 ( .A1(n20033), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20038) );
  NAND4_X1 U22939 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20036), .A3(
        n20035), .A4(n20034), .ZN(n20037) );
  NAND4_X1 U22940 ( .A1(n20040), .A2(n20039), .A3(n20038), .A4(n20037), .ZN(
        P1_U3029) );
  NOR2_X1 U22941 ( .A1(n20042), .A2(n20041), .ZN(P1_U3032) );
  NOR2_X2 U22942 ( .A1(n20044), .A2(n20043), .ZN(n20090) );
  AOI22_X1 U22943 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20090), .B1(DATAI_16_), 
        .B2(n20046), .ZN(n20579) );
  INV_X1 U22944 ( .A(n11114), .ZN(n20049) );
  INV_X1 U22945 ( .A(n20456), .ZN(n20322) );
  INV_X1 U22946 ( .A(n20424), .ZN(n20298) );
  AOI22_X1 U22947 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20090), .B1(DATAI_24_), 
        .B2(n20046), .ZN(n20531) );
  INV_X1 U22948 ( .A(n20531), .ZN(n20576) );
  NOR2_X2 U22949 ( .A1(n20092), .A2(n20051), .ZN(n20568) );
  NAND3_X1 U22950 ( .A1(n20380), .A2(n20375), .A3(n20457), .ZN(n20102) );
  NOR2_X1 U22951 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20102), .ZN(
        n20093) );
  AOI22_X1 U22952 ( .A1(n20094), .A2(n20576), .B1(n20568), .B2(n20093), .ZN(
        n20065) );
  INV_X1 U22953 ( .A(n20381), .ZN(n20052) );
  NOR2_X1 U22954 ( .A1(n20052), .A2(n20324), .ZN(n20061) );
  NAND2_X1 U22955 ( .A1(n20060), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20519) );
  AND2_X1 U22956 ( .A1(n20519), .A2(n20053), .ZN(n20384) );
  NAND3_X1 U22957 ( .A1(n20128), .A2(n20496), .A3(n20625), .ZN(n20054) );
  NAND2_X1 U22958 ( .A1(n20496), .A2(n20207), .ZN(n20459) );
  NAND2_X1 U22959 ( .A1(n20054), .A2(n20459), .ZN(n20059) );
  OR2_X1 U22960 ( .A1(n20323), .A2(n20055), .ZN(n20167) );
  OR2_X1 U22961 ( .A1(n20167), .A2(n20517), .ZN(n20062) );
  INV_X1 U22962 ( .A(n20093), .ZN(n20056) );
  AOI22_X1 U22963 ( .A1(n20059), .A2(n20062), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20056), .ZN(n20057) );
  OAI211_X1 U22964 ( .C1(n20061), .C2(n10613), .A(n20384), .B(n20057), .ZN(
        n20097) );
  NOR2_X2 U22965 ( .A1(n20058), .A2(n20210), .ZN(n20569) );
  INV_X1 U22966 ( .A(n20059), .ZN(n20063) );
  NOR2_X1 U22967 ( .A1(n20060), .A2(n10613), .ZN(n20211) );
  INV_X1 U22968 ( .A(n20211), .ZN(n20387) );
  INV_X1 U22969 ( .A(n20061), .ZN(n20206) );
  AOI22_X1 U22970 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20097), .B1(
        n20569), .B2(n20096), .ZN(n20064) );
  OAI211_X1 U22971 ( .C1(n20579), .C2(n20128), .A(n20065), .B(n20064), .ZN(
        P1_U3033) );
  AOI22_X1 U22972 ( .A1(DATAI_17_), .A2(n20046), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20090), .ZN(n20585) );
  AOI22_X1 U22973 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20090), .B1(DATAI_25_), 
        .B2(n20046), .ZN(n20535) );
  INV_X1 U22974 ( .A(n20535), .ZN(n20582) );
  NOR2_X2 U22975 ( .A1(n20092), .A2(n20066), .ZN(n20580) );
  AOI22_X1 U22976 ( .A1(n20094), .A2(n20582), .B1(n20580), .B2(n20093), .ZN(
        n20069) );
  NOR2_X2 U22977 ( .A1(n20067), .A2(n20210), .ZN(n20581) );
  AOI22_X1 U22978 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20097), .B1(
        n20581), .B2(n20096), .ZN(n20068) );
  OAI211_X1 U22979 ( .C1(n20585), .C2(n20128), .A(n20069), .B(n20068), .ZN(
        P1_U3034) );
  AOI22_X1 U22980 ( .A1(DATAI_18_), .A2(n20046), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20090), .ZN(n20591) );
  AOI22_X1 U22981 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20090), .B1(DATAI_26_), 
        .B2(n20046), .ZN(n20539) );
  INV_X1 U22982 ( .A(n20539), .ZN(n20588) );
  NOR2_X2 U22983 ( .A1(n20092), .A2(n20070), .ZN(n20586) );
  AOI22_X1 U22984 ( .A1(n20094), .A2(n20588), .B1(n20586), .B2(n20093), .ZN(
        n20073) );
  NOR2_X2 U22985 ( .A1(n20071), .A2(n20210), .ZN(n20587) );
  AOI22_X1 U22986 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20097), .B1(
        n20587), .B2(n20096), .ZN(n20072) );
  OAI211_X1 U22987 ( .C1(n20591), .C2(n20128), .A(n20073), .B(n20072), .ZN(
        P1_U3035) );
  AOI22_X1 U22988 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20090), .B1(DATAI_27_), 
        .B2(n20046), .ZN(n20543) );
  INV_X1 U22989 ( .A(n20543), .ZN(n20594) );
  INV_X1 U22990 ( .A(n20074), .ZN(n20075) );
  NOR2_X2 U22991 ( .A1(n20092), .A2(n20075), .ZN(n20592) );
  AOI22_X1 U22992 ( .A1(n20094), .A2(n20594), .B1(n20592), .B2(n20093), .ZN(
        n20078) );
  NOR2_X2 U22993 ( .A1(n20076), .A2(n20210), .ZN(n20593) );
  AOI22_X1 U22994 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20097), .B1(
        n20593), .B2(n20096), .ZN(n20077) );
  OAI211_X1 U22995 ( .C1(n20597), .C2(n20128), .A(n20078), .B(n20077), .ZN(
        P1_U3036) );
  AOI22_X1 U22996 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20090), .B1(DATAI_28_), 
        .B2(n20046), .ZN(n20547) );
  INV_X1 U22997 ( .A(n20547), .ZN(n20600) );
  NOR2_X2 U22998 ( .A1(n20092), .A2(n20079), .ZN(n20598) );
  AOI22_X1 U22999 ( .A1(n20094), .A2(n20600), .B1(n20598), .B2(n20093), .ZN(
        n20082) );
  NOR2_X2 U23000 ( .A1(n20080), .A2(n20210), .ZN(n20599) );
  AOI22_X1 U23001 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20097), .B1(
        n20599), .B2(n20096), .ZN(n20081) );
  OAI211_X1 U23002 ( .C1(n20603), .C2(n20128), .A(n20082), .B(n20081), .ZN(
        P1_U3037) );
  AOI22_X1 U23003 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20090), .B1(DATAI_29_), 
        .B2(n20046), .ZN(n20551) );
  INV_X1 U23004 ( .A(n20551), .ZN(n20606) );
  NOR2_X2 U23005 ( .A1(n20092), .A2(n20083), .ZN(n20604) );
  AOI22_X1 U23006 ( .A1(n20094), .A2(n20606), .B1(n20604), .B2(n20093), .ZN(
        n20086) );
  NOR2_X2 U23007 ( .A1(n20084), .A2(n20210), .ZN(n20605) );
  AOI22_X1 U23008 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20097), .B1(
        n20605), .B2(n20096), .ZN(n20085) );
  OAI211_X1 U23009 ( .C1(n20609), .C2(n20128), .A(n20086), .B(n20085), .ZN(
        P1_U3038) );
  AOI22_X1 U23010 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20090), .B1(DATAI_22_), 
        .B2(n20046), .ZN(n20615) );
  INV_X1 U23011 ( .A(n20555), .ZN(n20612) );
  AOI22_X1 U23012 ( .A1(n20094), .A2(n20612), .B1(n20610), .B2(n20093), .ZN(
        n20089) );
  NOR2_X2 U23013 ( .A1(n20087), .A2(n20210), .ZN(n20611) );
  AOI22_X1 U23014 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20097), .B1(
        n20611), .B2(n20096), .ZN(n20088) );
  OAI211_X1 U23015 ( .C1(n20615), .C2(n20128), .A(n20089), .B(n20088), .ZN(
        P1_U3039) );
  AOI22_X1 U23016 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20090), .B1(DATAI_23_), 
        .B2(n20046), .ZN(n20626) );
  AOI22_X1 U23017 ( .A1(DATAI_31_), .A2(n20046), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20090), .ZN(n20563) );
  INV_X1 U23018 ( .A(n20563), .ZN(n20620) );
  NOR2_X2 U23019 ( .A1(n20092), .A2(n20091), .ZN(n20617) );
  AOI22_X1 U23020 ( .A1(n20094), .A2(n20620), .B1(n20617), .B2(n20093), .ZN(
        n20099) );
  NOR2_X2 U23021 ( .A1(n20095), .A2(n20210), .ZN(n20619) );
  AOI22_X1 U23022 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20097), .B1(
        n20619), .B2(n20096), .ZN(n20098) );
  OAI211_X1 U23023 ( .C1(n20626), .C2(n20128), .A(n20099), .B(n20098), .ZN(
        P1_U3040) );
  INV_X1 U23024 ( .A(n20167), .ZN(n20101) );
  INV_X1 U23025 ( .A(n20100), .ZN(n20490) );
  NOR2_X1 U23026 ( .A1(n20489), .A2(n20102), .ZN(n20122) );
  AOI21_X1 U23027 ( .B1(n20101), .B2(n20490), .A(n20122), .ZN(n20103) );
  OAI22_X1 U23028 ( .A1(n20103), .A2(n20565), .B1(n20102), .B2(n10613), .ZN(
        n20123) );
  AOI22_X1 U23029 ( .A1(n20569), .A2(n20123), .B1(n20568), .B2(n20122), .ZN(
        n20108) );
  INV_X1 U23030 ( .A(n20102), .ZN(n20106) );
  INV_X1 U23031 ( .A(n20171), .ZN(n20104) );
  OAI21_X1 U23032 ( .B1(n20104), .B2(n20351), .A(n20103), .ZN(n20105) );
  OAI221_X1 U23033 ( .B1(n20496), .B2(n20106), .C1(n20565), .C2(n20105), .A(
        n20573), .ZN(n20125) );
  INV_X1 U23034 ( .A(n20579), .ZN(n20528) );
  AOI22_X1 U23035 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20125), .B1(
        n20124), .B2(n20528), .ZN(n20107) );
  OAI211_X1 U23036 ( .C1(n20531), .C2(n20128), .A(n20108), .B(n20107), .ZN(
        P1_U3041) );
  AOI22_X1 U23037 ( .A1(n20581), .A2(n20123), .B1(n20580), .B2(n20122), .ZN(
        n20110) );
  INV_X1 U23038 ( .A(n20585), .ZN(n20532) );
  AOI22_X1 U23039 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20125), .B1(
        n20124), .B2(n20532), .ZN(n20109) );
  OAI211_X1 U23040 ( .C1(n20535), .C2(n20128), .A(n20110), .B(n20109), .ZN(
        P1_U3042) );
  AOI22_X1 U23041 ( .A1(n20587), .A2(n20123), .B1(n20586), .B2(n20122), .ZN(
        n20112) );
  INV_X1 U23042 ( .A(n20591), .ZN(n20536) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20125), .B1(
        n20124), .B2(n20536), .ZN(n20111) );
  OAI211_X1 U23044 ( .C1(n20539), .C2(n20128), .A(n20112), .B(n20111), .ZN(
        P1_U3043) );
  AOI22_X1 U23045 ( .A1(n20593), .A2(n20123), .B1(n20592), .B2(n20122), .ZN(
        n20114) );
  INV_X1 U23046 ( .A(n20597), .ZN(n20540) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20125), .B1(
        n20124), .B2(n20540), .ZN(n20113) );
  OAI211_X1 U23048 ( .C1(n20543), .C2(n20128), .A(n20114), .B(n20113), .ZN(
        P1_U3044) );
  AOI22_X1 U23049 ( .A1(n20599), .A2(n20123), .B1(n20598), .B2(n20122), .ZN(
        n20117) );
  INV_X1 U23050 ( .A(n20128), .ZN(n20115) );
  AOI22_X1 U23051 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20125), .B1(
        n20115), .B2(n20600), .ZN(n20116) );
  OAI211_X1 U23052 ( .C1(n20603), .C2(n20157), .A(n20117), .B(n20116), .ZN(
        P1_U3045) );
  AOI22_X1 U23053 ( .A1(n20605), .A2(n20123), .B1(n20604), .B2(n20122), .ZN(
        n20119) );
  INV_X1 U23054 ( .A(n20609), .ZN(n20548) );
  AOI22_X1 U23055 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20125), .B1(
        n20124), .B2(n20548), .ZN(n20118) );
  OAI211_X1 U23056 ( .C1(n20551), .C2(n20128), .A(n20119), .B(n20118), .ZN(
        P1_U3046) );
  AOI22_X1 U23057 ( .A1(n20611), .A2(n20123), .B1(n20610), .B2(n20122), .ZN(
        n20121) );
  INV_X1 U23058 ( .A(n20615), .ZN(n20552) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20125), .B1(
        n20124), .B2(n20552), .ZN(n20120) );
  OAI211_X1 U23060 ( .C1(n20555), .C2(n20128), .A(n20121), .B(n20120), .ZN(
        P1_U3047) );
  AOI22_X1 U23061 ( .A1(n20619), .A2(n20123), .B1(n20617), .B2(n20122), .ZN(
        n20127) );
  INV_X1 U23062 ( .A(n20626), .ZN(n20558) );
  AOI22_X1 U23063 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20125), .B1(
        n20124), .B2(n20558), .ZN(n20126) );
  OAI211_X1 U23064 ( .C1(n20563), .C2(n20128), .A(n20127), .B(n20126), .ZN(
        P1_U3048) );
  INV_X1 U23065 ( .A(n20568), .ZN(n20376) );
  NAND3_X1 U23066 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20380), .A3(
        n20375), .ZN(n20174) );
  OR2_X1 U23067 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20174), .ZN(
        n20156) );
  OAI22_X1 U23068 ( .A1(n20198), .A2(n20579), .B1(n20376), .B2(n20156), .ZN(
        n20130) );
  INV_X1 U23069 ( .A(n20130), .ZN(n20137) );
  NAND3_X1 U23070 ( .A1(n20198), .A2(n20157), .A3(n20496), .ZN(n20131) );
  NAND2_X1 U23071 ( .A1(n20131), .A2(n20459), .ZN(n20133) );
  OR2_X1 U23072 ( .A1(n20167), .A2(n12799), .ZN(n20134) );
  AOI22_X1 U23073 ( .A1(n20133), .A2(n20134), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20156), .ZN(n20132) );
  OR2_X1 U23074 ( .A1(n20381), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20265) );
  NAND2_X1 U23075 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20265), .ZN(n20262) );
  NAND3_X1 U23076 ( .A1(n20384), .A2(n20132), .A3(n20262), .ZN(n20160) );
  INV_X1 U23077 ( .A(n20133), .ZN(n20135) );
  AOI22_X1 U23078 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20160), .B1(
        n20569), .B2(n20159), .ZN(n20136) );
  OAI211_X1 U23079 ( .C1(n20531), .C2(n20157), .A(n20137), .B(n20136), .ZN(
        P1_U3049) );
  INV_X1 U23080 ( .A(n20580), .ZN(n20392) );
  OAI22_X1 U23081 ( .A1(n20198), .A2(n20585), .B1(n20156), .B2(n20392), .ZN(
        n20138) );
  INV_X1 U23082 ( .A(n20138), .ZN(n20140) );
  AOI22_X1 U23083 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20160), .B1(
        n20581), .B2(n20159), .ZN(n20139) );
  OAI211_X1 U23084 ( .C1(n20535), .C2(n20157), .A(n20140), .B(n20139), .ZN(
        P1_U3050) );
  INV_X1 U23085 ( .A(n20586), .ZN(n20396) );
  OAI22_X1 U23086 ( .A1(n20198), .A2(n20591), .B1(n20396), .B2(n20156), .ZN(
        n20141) );
  INV_X1 U23087 ( .A(n20141), .ZN(n20143) );
  AOI22_X1 U23088 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20160), .B1(
        n20587), .B2(n20159), .ZN(n20142) );
  OAI211_X1 U23089 ( .C1(n20539), .C2(n20157), .A(n20143), .B(n20142), .ZN(
        P1_U3051) );
  INV_X1 U23090 ( .A(n20592), .ZN(n20400) );
  OAI22_X1 U23091 ( .A1(n20198), .A2(n20597), .B1(n20156), .B2(n20400), .ZN(
        n20144) );
  INV_X1 U23092 ( .A(n20144), .ZN(n20146) );
  AOI22_X1 U23093 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20160), .B1(
        n20593), .B2(n20159), .ZN(n20145) );
  OAI211_X1 U23094 ( .C1(n20543), .C2(n20157), .A(n20146), .B(n20145), .ZN(
        P1_U3052) );
  INV_X1 U23095 ( .A(n20598), .ZN(n20404) );
  OAI22_X1 U23096 ( .A1(n20157), .A2(n20547), .B1(n20156), .B2(n20404), .ZN(
        n20147) );
  INV_X1 U23097 ( .A(n20147), .ZN(n20149) );
  AOI22_X1 U23098 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20160), .B1(
        n20599), .B2(n20159), .ZN(n20148) );
  OAI211_X1 U23099 ( .C1(n20603), .C2(n20198), .A(n20149), .B(n20148), .ZN(
        P1_U3053) );
  INV_X1 U23100 ( .A(n20604), .ZN(n20408) );
  OAI22_X1 U23101 ( .A1(n20157), .A2(n20551), .B1(n20156), .B2(n20408), .ZN(
        n20150) );
  INV_X1 U23102 ( .A(n20150), .ZN(n20152) );
  AOI22_X1 U23103 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20160), .B1(
        n20605), .B2(n20159), .ZN(n20151) );
  OAI211_X1 U23104 ( .C1(n20609), .C2(n20198), .A(n20152), .B(n20151), .ZN(
        P1_U3054) );
  INV_X1 U23105 ( .A(n20610), .ZN(n20412) );
  OAI22_X1 U23106 ( .A1(n20157), .A2(n20555), .B1(n20156), .B2(n20412), .ZN(
        n20153) );
  INV_X1 U23107 ( .A(n20153), .ZN(n20155) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20160), .B1(
        n20611), .B2(n20159), .ZN(n20154) );
  OAI211_X1 U23109 ( .C1(n20615), .C2(n20198), .A(n20155), .B(n20154), .ZN(
        P1_U3055) );
  INV_X1 U23110 ( .A(n20617), .ZN(n20416) );
  OAI22_X1 U23111 ( .A1(n20157), .A2(n20563), .B1(n20416), .B2(n20156), .ZN(
        n20158) );
  INV_X1 U23112 ( .A(n20158), .ZN(n20162) );
  AOI22_X1 U23113 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20160), .B1(
        n20619), .B2(n20159), .ZN(n20161) );
  OAI211_X1 U23114 ( .C1(n20626), .C2(n20198), .A(n20162), .B(n20161), .ZN(
        P1_U3056) );
  NAND2_X1 U23115 ( .A1(n20171), .A2(n20424), .ZN(n20213) );
  INV_X1 U23116 ( .A(n20163), .ZN(n20427) );
  NAND2_X1 U23117 ( .A1(n20427), .A2(n20380), .ZN(n20197) );
  OAI22_X1 U23118 ( .A1(n20198), .A2(n20531), .B1(n20376), .B2(n20197), .ZN(
        n20164) );
  INV_X1 U23119 ( .A(n20164), .ZN(n20178) );
  NOR3_X1 U23120 ( .A1(n20167), .A2(n20165), .A3(n20166), .ZN(n20169) );
  INV_X1 U23121 ( .A(n20197), .ZN(n20168) );
  NOR2_X1 U23122 ( .A1(n20169), .A2(n20168), .ZN(n20176) );
  INV_X1 U23123 ( .A(n20295), .ZN(n20170) );
  AOI21_X1 U23124 ( .B1(n20171), .B2(n20170), .A(n20565), .ZN(n20173) );
  AOI22_X1 U23125 ( .A1(n20176), .A2(n20173), .B1(n20565), .B2(n20174), .ZN(
        n20172) );
  NAND2_X1 U23126 ( .A1(n20573), .A2(n20172), .ZN(n20201) );
  INV_X1 U23127 ( .A(n20173), .ZN(n20175) );
  OAI22_X1 U23128 ( .A1(n20176), .A2(n20175), .B1(n10613), .B2(n20174), .ZN(
        n20200) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20201), .B1(
        n20569), .B2(n20200), .ZN(n20177) );
  OAI211_X1 U23130 ( .C1(n20579), .C2(n20213), .A(n20178), .B(n20177), .ZN(
        P1_U3057) );
  OAI22_X1 U23131 ( .A1(n20198), .A2(n20535), .B1(n20392), .B2(n20197), .ZN(
        n20179) );
  INV_X1 U23132 ( .A(n20179), .ZN(n20181) );
  AOI22_X1 U23133 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20201), .B1(
        n20581), .B2(n20200), .ZN(n20180) );
  OAI211_X1 U23134 ( .C1(n20585), .C2(n20213), .A(n20181), .B(n20180), .ZN(
        P1_U3058) );
  OAI22_X1 U23135 ( .A1(n20213), .A2(n20591), .B1(n20396), .B2(n20197), .ZN(
        n20182) );
  INV_X1 U23136 ( .A(n20182), .ZN(n20184) );
  AOI22_X1 U23137 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20201), .B1(
        n20587), .B2(n20200), .ZN(n20183) );
  OAI211_X1 U23138 ( .C1(n20539), .C2(n20198), .A(n20184), .B(n20183), .ZN(
        P1_U3059) );
  OAI22_X1 U23139 ( .A1(n20213), .A2(n20597), .B1(n20400), .B2(n20197), .ZN(
        n20185) );
  INV_X1 U23140 ( .A(n20185), .ZN(n20187) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20201), .B1(
        n20593), .B2(n20200), .ZN(n20186) );
  OAI211_X1 U23142 ( .C1(n20543), .C2(n20198), .A(n20187), .B(n20186), .ZN(
        P1_U3060) );
  OAI22_X1 U23143 ( .A1(n20198), .A2(n20547), .B1(n20197), .B2(n20404), .ZN(
        n20188) );
  INV_X1 U23144 ( .A(n20188), .ZN(n20190) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20201), .B1(
        n20599), .B2(n20200), .ZN(n20189) );
  OAI211_X1 U23146 ( .C1(n20603), .C2(n20213), .A(n20190), .B(n20189), .ZN(
        P1_U3061) );
  OAI22_X1 U23147 ( .A1(n20198), .A2(n20551), .B1(n20197), .B2(n20408), .ZN(
        n20191) );
  INV_X1 U23148 ( .A(n20191), .ZN(n20193) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20201), .B1(
        n20605), .B2(n20200), .ZN(n20192) );
  OAI211_X1 U23150 ( .C1(n20609), .C2(n20213), .A(n20193), .B(n20192), .ZN(
        P1_U3062) );
  OAI22_X1 U23151 ( .A1(n20213), .A2(n20615), .B1(n20197), .B2(n20412), .ZN(
        n20194) );
  INV_X1 U23152 ( .A(n20194), .ZN(n20196) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20201), .B1(
        n20611), .B2(n20200), .ZN(n20195) );
  OAI211_X1 U23154 ( .C1(n20555), .C2(n20198), .A(n20196), .B(n20195), .ZN(
        P1_U3063) );
  OAI22_X1 U23155 ( .A1(n20198), .A2(n20563), .B1(n20416), .B2(n20197), .ZN(
        n20199) );
  INV_X1 U23156 ( .A(n20199), .ZN(n20203) );
  AOI22_X1 U23157 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20201), .B1(
        n20619), .B2(n20200), .ZN(n20202) );
  OAI211_X1 U23158 ( .C1(n20626), .C2(n20213), .A(n20203), .B(n20202), .ZN(
        P1_U3064) );
  NOR2_X1 U23159 ( .A1(n12324), .A2(n20204), .ZN(n20291) );
  NAND3_X1 U23160 ( .A1(n20291), .A2(n20496), .A3(n12799), .ZN(n20205) );
  OAI21_X1 U23161 ( .B1(n20519), .B2(n20206), .A(n20205), .ZN(n20229) );
  NAND3_X1 U23162 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20380), .A3(
        n20457), .ZN(n20234) );
  NOR2_X1 U23163 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20234), .ZN(
        n20228) );
  AOI22_X1 U23164 ( .A1(n20569), .A2(n20229), .B1(n20568), .B2(n20228), .ZN(
        n20215) );
  AOI21_X1 U23165 ( .B1(n20213), .B2(n20259), .A(n20207), .ZN(n20208) );
  AOI21_X1 U23166 ( .B1(n20291), .B2(n12799), .A(n20208), .ZN(n20209) );
  NOR2_X1 U23167 ( .A1(n20209), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20212) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20231), .B1(
        n20230), .B2(n20576), .ZN(n20214) );
  OAI211_X1 U23169 ( .C1(n20579), .C2(n20259), .A(n20215), .B(n20214), .ZN(
        P1_U3065) );
  AOI22_X1 U23170 ( .A1(n20581), .A2(n20229), .B1(n20580), .B2(n20228), .ZN(
        n20217) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20231), .B1(
        n20230), .B2(n20582), .ZN(n20216) );
  OAI211_X1 U23172 ( .C1(n20585), .C2(n20259), .A(n20217), .B(n20216), .ZN(
        P1_U3066) );
  AOI22_X1 U23173 ( .A1(n20587), .A2(n20229), .B1(n20586), .B2(n20228), .ZN(
        n20219) );
  AOI22_X1 U23174 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20231), .B1(
        n20230), .B2(n20588), .ZN(n20218) );
  OAI211_X1 U23175 ( .C1(n20591), .C2(n20259), .A(n20219), .B(n20218), .ZN(
        P1_U3067) );
  AOI22_X1 U23176 ( .A1(n20593), .A2(n20229), .B1(n20592), .B2(n20228), .ZN(
        n20221) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20231), .B1(
        n20230), .B2(n20594), .ZN(n20220) );
  OAI211_X1 U23178 ( .C1(n20597), .C2(n20259), .A(n20221), .B(n20220), .ZN(
        P1_U3068) );
  AOI22_X1 U23179 ( .A1(n20599), .A2(n20229), .B1(n20598), .B2(n20228), .ZN(
        n20223) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20231), .B1(
        n20230), .B2(n20600), .ZN(n20222) );
  OAI211_X1 U23181 ( .C1(n20603), .C2(n20259), .A(n20223), .B(n20222), .ZN(
        P1_U3069) );
  AOI22_X1 U23182 ( .A1(n20605), .A2(n20229), .B1(n20604), .B2(n20228), .ZN(
        n20225) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20231), .B1(
        n20230), .B2(n20606), .ZN(n20224) );
  OAI211_X1 U23184 ( .C1(n20609), .C2(n20259), .A(n20225), .B(n20224), .ZN(
        P1_U3070) );
  AOI22_X1 U23185 ( .A1(n20611), .A2(n20229), .B1(n20610), .B2(n20228), .ZN(
        n20227) );
  AOI22_X1 U23186 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20231), .B1(
        n20230), .B2(n20612), .ZN(n20226) );
  OAI211_X1 U23187 ( .C1(n20615), .C2(n20259), .A(n20227), .B(n20226), .ZN(
        P1_U3071) );
  AOI22_X1 U23188 ( .A1(n20619), .A2(n20229), .B1(n20617), .B2(n20228), .ZN(
        n20233) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20231), .B1(
        n20230), .B2(n20620), .ZN(n20232) );
  OAI211_X1 U23190 ( .C1(n20626), .C2(n20259), .A(n20233), .B(n20232), .ZN(
        P1_U3072) );
  NOR2_X1 U23191 ( .A1(n20489), .A2(n20234), .ZN(n20254) );
  AOI21_X1 U23192 ( .B1(n20291), .B2(n20490), .A(n20254), .ZN(n20235) );
  OAI22_X1 U23193 ( .A1(n20235), .A2(n20565), .B1(n20234), .B2(n10613), .ZN(
        n20255) );
  AOI22_X1 U23194 ( .A1(n20569), .A2(n20255), .B1(n20568), .B2(n20254), .ZN(
        n20240) );
  INV_X1 U23195 ( .A(n20234), .ZN(n20237) );
  OAI21_X1 U23196 ( .B1(n20299), .B2(n20351), .A(n20235), .ZN(n20236) );
  OAI221_X1 U23197 ( .B1(n20496), .B2(n20237), .C1(n20565), .C2(n20236), .A(
        n20573), .ZN(n20256) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20256), .B1(
        n20278), .B2(n20528), .ZN(n20239) );
  OAI211_X1 U23199 ( .C1(n20531), .C2(n20259), .A(n20240), .B(n20239), .ZN(
        P1_U3073) );
  AOI22_X1 U23200 ( .A1(n20581), .A2(n20255), .B1(n20580), .B2(n20254), .ZN(
        n20242) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20256), .B1(
        n20278), .B2(n20532), .ZN(n20241) );
  OAI211_X1 U23202 ( .C1(n20535), .C2(n20259), .A(n20242), .B(n20241), .ZN(
        P1_U3074) );
  AOI22_X1 U23203 ( .A1(n20587), .A2(n20255), .B1(n20586), .B2(n20254), .ZN(
        n20244) );
  INV_X1 U23204 ( .A(n20259), .ZN(n20247) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20256), .B1(
        n20247), .B2(n20588), .ZN(n20243) );
  OAI211_X1 U23206 ( .C1(n20591), .C2(n20288), .A(n20244), .B(n20243), .ZN(
        P1_U3075) );
  AOI22_X1 U23207 ( .A1(n20593), .A2(n20255), .B1(n20592), .B2(n20254), .ZN(
        n20246) );
  AOI22_X1 U23208 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20256), .B1(
        n20247), .B2(n20594), .ZN(n20245) );
  OAI211_X1 U23209 ( .C1(n20597), .C2(n20288), .A(n20246), .B(n20245), .ZN(
        P1_U3076) );
  AOI22_X1 U23210 ( .A1(n20599), .A2(n20255), .B1(n20598), .B2(n20254), .ZN(
        n20249) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20256), .B1(
        n20247), .B2(n20600), .ZN(n20248) );
  OAI211_X1 U23212 ( .C1(n20603), .C2(n20288), .A(n20249), .B(n20248), .ZN(
        P1_U3077) );
  AOI22_X1 U23213 ( .A1(n20605), .A2(n20255), .B1(n20604), .B2(n20254), .ZN(
        n20251) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20256), .B1(
        n20278), .B2(n20548), .ZN(n20250) );
  OAI211_X1 U23215 ( .C1(n20551), .C2(n20259), .A(n20251), .B(n20250), .ZN(
        P1_U3078) );
  AOI22_X1 U23216 ( .A1(n20611), .A2(n20255), .B1(n20610), .B2(n20254), .ZN(
        n20253) );
  AOI22_X1 U23217 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20256), .B1(
        n20278), .B2(n20552), .ZN(n20252) );
  OAI211_X1 U23218 ( .C1(n20555), .C2(n20259), .A(n20253), .B(n20252), .ZN(
        P1_U3079) );
  AOI22_X1 U23219 ( .A1(n20619), .A2(n20255), .B1(n20617), .B2(n20254), .ZN(
        n20258) );
  AOI22_X1 U23220 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20256), .B1(
        n20278), .B2(n20558), .ZN(n20257) );
  OAI211_X1 U23221 ( .C1(n20563), .C2(n20259), .A(n20258), .B(n20257), .ZN(
        P1_U3080) );
  INV_X1 U23222 ( .A(n20314), .ZN(n20317) );
  INV_X1 U23223 ( .A(n20297), .ZN(n20293) );
  NOR2_X1 U23224 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20293), .ZN(
        n20283) );
  AOI22_X1 U23225 ( .A1(n20317), .A2(n20528), .B1(n20283), .B2(n20568), .ZN(
        n20269) );
  NAND3_X1 U23226 ( .A1(n20314), .A2(n20288), .A3(n20496), .ZN(n20260) );
  NAND2_X1 U23227 ( .A1(n20260), .A2(n20459), .ZN(n20264) );
  NAND2_X1 U23228 ( .A1(n20291), .A2(n20517), .ZN(n20266) );
  INV_X1 U23229 ( .A(n20283), .ZN(n20261) );
  AOI22_X1 U23230 ( .A1(n20264), .A2(n20266), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20261), .ZN(n20263) );
  NAND3_X1 U23231 ( .A1(n20526), .A2(n20263), .A3(n20262), .ZN(n20285) );
  INV_X1 U23232 ( .A(n20264), .ZN(n20267) );
  OAI22_X1 U23233 ( .A1(n20267), .A2(n20266), .B1(n20265), .B2(n20519), .ZN(
        n20284) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20285), .B1(
        n20569), .B2(n20284), .ZN(n20268) );
  OAI211_X1 U23235 ( .C1(n20531), .C2(n20288), .A(n20269), .B(n20268), .ZN(
        P1_U3081) );
  AOI22_X1 U23236 ( .A1(n20278), .A2(n20582), .B1(n20580), .B2(n20283), .ZN(
        n20271) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20285), .B1(
        n20581), .B2(n20284), .ZN(n20270) );
  OAI211_X1 U23238 ( .C1(n20585), .C2(n20314), .A(n20271), .B(n20270), .ZN(
        P1_U3082) );
  AOI22_X1 U23239 ( .A1(n20317), .A2(n20536), .B1(n20283), .B2(n20586), .ZN(
        n20273) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20285), .B1(
        n20587), .B2(n20284), .ZN(n20272) );
  OAI211_X1 U23241 ( .C1(n20539), .C2(n20288), .A(n20273), .B(n20272), .ZN(
        P1_U3083) );
  AOI22_X1 U23242 ( .A1(n20278), .A2(n20594), .B1(n20592), .B2(n20283), .ZN(
        n20275) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20285), .B1(
        n20593), .B2(n20284), .ZN(n20274) );
  OAI211_X1 U23244 ( .C1(n20597), .C2(n20314), .A(n20275), .B(n20274), .ZN(
        P1_U3084) );
  AOI22_X1 U23245 ( .A1(n20278), .A2(n20600), .B1(n20598), .B2(n20283), .ZN(
        n20277) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20285), .B1(
        n20599), .B2(n20284), .ZN(n20276) );
  OAI211_X1 U23247 ( .C1(n20603), .C2(n20314), .A(n20277), .B(n20276), .ZN(
        P1_U3085) );
  AOI22_X1 U23248 ( .A1(n20278), .A2(n20606), .B1(n20283), .B2(n20604), .ZN(
        n20280) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20285), .B1(
        n20605), .B2(n20284), .ZN(n20279) );
  OAI211_X1 U23250 ( .C1(n20609), .C2(n20314), .A(n20280), .B(n20279), .ZN(
        P1_U3086) );
  AOI22_X1 U23251 ( .A1(n20317), .A2(n20552), .B1(n20283), .B2(n20610), .ZN(
        n20282) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20285), .B1(
        n20611), .B2(n20284), .ZN(n20281) );
  OAI211_X1 U23253 ( .C1(n20555), .C2(n20288), .A(n20282), .B(n20281), .ZN(
        P1_U3087) );
  AOI22_X1 U23254 ( .A1(n20317), .A2(n20558), .B1(n20283), .B2(n20617), .ZN(
        n20287) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20285), .B1(
        n20619), .B2(n20284), .ZN(n20286) );
  OAI211_X1 U23256 ( .C1(n20563), .C2(n20288), .A(n20287), .B(n20286), .ZN(
        P1_U3088) );
  INV_X1 U23257 ( .A(n20165), .ZN(n20290) );
  NAND3_X1 U23258 ( .A1(n20290), .A2(n20289), .A3(n20496), .ZN(n20567) );
  INV_X1 U23259 ( .A(n20291), .ZN(n20294) );
  INV_X1 U23260 ( .A(n20292), .ZN(n20315) );
  OAI222_X1 U23261 ( .A1(n20567), .A2(n20294), .B1(n10613), .B2(n20293), .C1(
        n20565), .C2(n20292), .ZN(n20316) );
  AOI22_X1 U23262 ( .A1(n20569), .A2(n20316), .B1(n20568), .B2(n20315), .ZN(
        n20301) );
  OR2_X1 U23263 ( .A1(n20295), .A2(n20565), .ZN(n20571) );
  NOR2_X1 U23264 ( .A1(n20299), .A2(n20571), .ZN(n20296) );
  OAI21_X1 U23265 ( .B1(n20297), .B2(n20296), .A(n20573), .ZN(n20318) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20318), .B1(
        n20345), .B2(n20528), .ZN(n20300) );
  OAI211_X1 U23267 ( .C1(n20531), .C2(n20314), .A(n20301), .B(n20300), .ZN(
        P1_U3089) );
  AOI22_X1 U23268 ( .A1(n20581), .A2(n20316), .B1(n20580), .B2(n20315), .ZN(
        n20303) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20318), .B1(
        n20345), .B2(n20532), .ZN(n20302) );
  OAI211_X1 U23270 ( .C1(n20535), .C2(n20314), .A(n20303), .B(n20302), .ZN(
        P1_U3090) );
  AOI22_X1 U23271 ( .A1(n20587), .A2(n20316), .B1(n20586), .B2(n20315), .ZN(
        n20305) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20318), .B1(
        n20345), .B2(n20536), .ZN(n20304) );
  OAI211_X1 U23273 ( .C1(n20539), .C2(n20314), .A(n20305), .B(n20304), .ZN(
        P1_U3091) );
  AOI22_X1 U23274 ( .A1(n20593), .A2(n20316), .B1(n20592), .B2(n20315), .ZN(
        n20307) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20594), .ZN(n20306) );
  OAI211_X1 U23276 ( .C1(n20597), .C2(n20321), .A(n20307), .B(n20306), .ZN(
        P1_U3092) );
  AOI22_X1 U23277 ( .A1(n20599), .A2(n20316), .B1(n20598), .B2(n20315), .ZN(
        n20309) );
  INV_X1 U23278 ( .A(n20603), .ZN(n20544) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20318), .B1(
        n20345), .B2(n20544), .ZN(n20308) );
  OAI211_X1 U23280 ( .C1(n20547), .C2(n20314), .A(n20309), .B(n20308), .ZN(
        P1_U3093) );
  AOI22_X1 U23281 ( .A1(n20605), .A2(n20316), .B1(n20604), .B2(n20315), .ZN(
        n20311) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20606), .ZN(n20310) );
  OAI211_X1 U23283 ( .C1(n20609), .C2(n20321), .A(n20311), .B(n20310), .ZN(
        P1_U3094) );
  AOI22_X1 U23284 ( .A1(n20611), .A2(n20316), .B1(n20610), .B2(n20315), .ZN(
        n20313) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20318), .B1(
        n20345), .B2(n20552), .ZN(n20312) );
  OAI211_X1 U23286 ( .C1(n20555), .C2(n20314), .A(n20313), .B(n20312), .ZN(
        P1_U3095) );
  AOI22_X1 U23287 ( .A1(n20619), .A2(n20316), .B1(n20617), .B2(n20315), .ZN(
        n20320) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20318), .B1(
        n20317), .B2(n20620), .ZN(n20319) );
  OAI211_X1 U23289 ( .C1(n20626), .C2(n20321), .A(n20320), .B(n20319), .ZN(
        P1_U3096) );
  AND2_X1 U23290 ( .A1(n20323), .A2(n12324), .ZN(n20426) );
  NAND3_X1 U23291 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20375), .A3(
        n20457), .ZN(n20349) );
  NOR2_X1 U23292 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20349), .ZN(
        n20343) );
  AOI21_X1 U23293 ( .B1(n20426), .B2(n12799), .A(n20343), .ZN(n20326) );
  NAND2_X1 U23294 ( .A1(n20324), .A2(n20381), .ZN(n20464) );
  OAI22_X1 U23295 ( .A1(n20326), .A2(n20565), .B1(n20387), .B2(n20464), .ZN(
        n20344) );
  AOI22_X1 U23296 ( .A1(n20569), .A2(n20344), .B1(n20568), .B2(n20343), .ZN(
        n20330) );
  INV_X1 U23297 ( .A(n20373), .ZN(n20325) );
  OAI21_X1 U23298 ( .B1(n20325), .B2(n20345), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20327) );
  NAND2_X1 U23299 ( .A1(n20327), .A2(n20326), .ZN(n20328) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20576), .ZN(n20329) );
  OAI211_X1 U23301 ( .C1(n20579), .C2(n20373), .A(n20330), .B(n20329), .ZN(
        P1_U3097) );
  AOI22_X1 U23302 ( .A1(n20581), .A2(n20344), .B1(n20580), .B2(n20343), .ZN(
        n20332) );
  AOI22_X1 U23303 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20582), .ZN(n20331) );
  OAI211_X1 U23304 ( .C1(n20585), .C2(n20373), .A(n20332), .B(n20331), .ZN(
        P1_U3098) );
  AOI22_X1 U23305 ( .A1(n20587), .A2(n20344), .B1(n20586), .B2(n20343), .ZN(
        n20334) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20588), .ZN(n20333) );
  OAI211_X1 U23307 ( .C1(n20591), .C2(n20373), .A(n20334), .B(n20333), .ZN(
        P1_U3099) );
  AOI22_X1 U23308 ( .A1(n20593), .A2(n20344), .B1(n20592), .B2(n20343), .ZN(
        n20336) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20594), .ZN(n20335) );
  OAI211_X1 U23310 ( .C1(n20597), .C2(n20373), .A(n20336), .B(n20335), .ZN(
        P1_U3100) );
  AOI22_X1 U23311 ( .A1(n20599), .A2(n20344), .B1(n20598), .B2(n20343), .ZN(
        n20338) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20600), .ZN(n20337) );
  OAI211_X1 U23313 ( .C1(n20603), .C2(n20373), .A(n20338), .B(n20337), .ZN(
        P1_U3101) );
  AOI22_X1 U23314 ( .A1(n20605), .A2(n20344), .B1(n20604), .B2(n20343), .ZN(
        n20340) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20606), .ZN(n20339) );
  OAI211_X1 U23316 ( .C1(n20609), .C2(n20373), .A(n20340), .B(n20339), .ZN(
        P1_U3102) );
  AOI22_X1 U23317 ( .A1(n20611), .A2(n20344), .B1(n20610), .B2(n20343), .ZN(
        n20342) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20612), .ZN(n20341) );
  OAI211_X1 U23319 ( .C1(n20615), .C2(n20373), .A(n20342), .B(n20341), .ZN(
        P1_U3103) );
  AOI22_X1 U23320 ( .A1(n20619), .A2(n20344), .B1(n20617), .B2(n20343), .ZN(
        n20348) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20620), .ZN(n20347) );
  OAI211_X1 U23322 ( .C1(n20626), .C2(n20373), .A(n20348), .B(n20347), .ZN(
        P1_U3104) );
  NOR2_X1 U23323 ( .A1(n20489), .A2(n20349), .ZN(n20368) );
  AOI21_X1 U23324 ( .B1(n20426), .B2(n20490), .A(n20368), .ZN(n20350) );
  OAI22_X1 U23325 ( .A1(n20350), .A2(n20565), .B1(n20349), .B2(n10613), .ZN(
        n20369) );
  AOI22_X1 U23326 ( .A1(n20569), .A2(n20369), .B1(n20568), .B2(n20368), .ZN(
        n20355) );
  INV_X1 U23327 ( .A(n20349), .ZN(n20353) );
  INV_X1 U23328 ( .A(n20425), .ZN(n20430) );
  OAI21_X1 U23329 ( .B1(n20430), .B2(n20351), .A(n20350), .ZN(n20352) );
  OAI221_X1 U23330 ( .B1(n20496), .B2(n20353), .C1(n20565), .C2(n20352), .A(
        n20573), .ZN(n20370) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20370), .B1(
        n20378), .B2(n20528), .ZN(n20354) );
  OAI211_X1 U23332 ( .C1(n20531), .C2(n20373), .A(n20355), .B(n20354), .ZN(
        P1_U3105) );
  AOI22_X1 U23333 ( .A1(n20581), .A2(n20369), .B1(n20580), .B2(n20368), .ZN(
        n20357) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20370), .B1(
        n20378), .B2(n20532), .ZN(n20356) );
  OAI211_X1 U23335 ( .C1(n20535), .C2(n20373), .A(n20357), .B(n20356), .ZN(
        P1_U3106) );
  AOI22_X1 U23336 ( .A1(n20587), .A2(n20369), .B1(n20586), .B2(n20368), .ZN(
        n20359) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20370), .B1(
        n20378), .B2(n20536), .ZN(n20358) );
  OAI211_X1 U23338 ( .C1(n20539), .C2(n20373), .A(n20359), .B(n20358), .ZN(
        P1_U3107) );
  AOI22_X1 U23339 ( .A1(n20593), .A2(n20369), .B1(n20592), .B2(n20368), .ZN(
        n20361) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20370), .B1(
        n20378), .B2(n20540), .ZN(n20360) );
  OAI211_X1 U23341 ( .C1(n20543), .C2(n20373), .A(n20361), .B(n20360), .ZN(
        P1_U3108) );
  AOI22_X1 U23342 ( .A1(n20599), .A2(n20369), .B1(n20598), .B2(n20368), .ZN(
        n20363) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20370), .B1(
        n20378), .B2(n20544), .ZN(n20362) );
  OAI211_X1 U23344 ( .C1(n20547), .C2(n20373), .A(n20363), .B(n20362), .ZN(
        P1_U3109) );
  AOI22_X1 U23345 ( .A1(n20605), .A2(n20369), .B1(n20604), .B2(n20368), .ZN(
        n20365) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20370), .B1(
        n20378), .B2(n20548), .ZN(n20364) );
  OAI211_X1 U23347 ( .C1(n20551), .C2(n20373), .A(n20365), .B(n20364), .ZN(
        P1_U3110) );
  AOI22_X1 U23348 ( .A1(n20611), .A2(n20369), .B1(n20610), .B2(n20368), .ZN(
        n20367) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20370), .B1(
        n20378), .B2(n20552), .ZN(n20366) );
  OAI211_X1 U23350 ( .C1(n20555), .C2(n20373), .A(n20367), .B(n20366), .ZN(
        P1_U3111) );
  AOI22_X1 U23351 ( .A1(n20619), .A2(n20369), .B1(n20617), .B2(n20368), .ZN(
        n20372) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20370), .B1(
        n20378), .B2(n20558), .ZN(n20371) );
  OAI211_X1 U23353 ( .C1(n20563), .C2(n20373), .A(n20372), .B(n20371), .ZN(
        P1_U3112) );
  NAND3_X1 U23354 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20375), .ZN(n20431) );
  NOR2_X1 U23355 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20431), .ZN(
        n20382) );
  INV_X1 U23356 ( .A(n20382), .ZN(n20417) );
  OAI22_X1 U23357 ( .A1(n20449), .A2(n20579), .B1(n20376), .B2(n20417), .ZN(
        n20377) );
  INV_X1 U23358 ( .A(n20377), .ZN(n20391) );
  OAI21_X1 U23359 ( .B1(n20452), .B2(n20378), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20379) );
  NAND2_X1 U23360 ( .A1(n20379), .A2(n20496), .ZN(n20389) );
  AND2_X1 U23361 ( .A1(n20426), .A2(n20517), .ZN(n20386) );
  OR2_X1 U23362 ( .A1(n20381), .A2(n20380), .ZN(n20520) );
  NAND2_X1 U23363 ( .A1(n20520), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20525) );
  OAI21_X1 U23364 ( .B1(n20704), .B2(n20382), .A(n20525), .ZN(n20383) );
  INV_X1 U23365 ( .A(n20383), .ZN(n20385) );
  OAI211_X1 U23366 ( .C1(n20389), .C2(n20386), .A(n20385), .B(n20384), .ZN(
        n20420) );
  INV_X1 U23367 ( .A(n20386), .ZN(n20388) );
  OAI22_X1 U23368 ( .A1(n20389), .A2(n20388), .B1(n20387), .B2(n20520), .ZN(
        n20419) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20420), .B1(
        n20569), .B2(n20419), .ZN(n20390) );
  OAI211_X1 U23370 ( .C1(n20531), .C2(n20423), .A(n20391), .B(n20390), .ZN(
        P1_U3113) );
  OAI22_X1 U23371 ( .A1(n20423), .A2(n20535), .B1(n20417), .B2(n20392), .ZN(
        n20393) );
  INV_X1 U23372 ( .A(n20393), .ZN(n20395) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20420), .B1(
        n20581), .B2(n20419), .ZN(n20394) );
  OAI211_X1 U23374 ( .C1(n20585), .C2(n20449), .A(n20395), .B(n20394), .ZN(
        P1_U3114) );
  OAI22_X1 U23375 ( .A1(n20449), .A2(n20591), .B1(n20417), .B2(n20396), .ZN(
        n20397) );
  INV_X1 U23376 ( .A(n20397), .ZN(n20399) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20420), .B1(
        n20587), .B2(n20419), .ZN(n20398) );
  OAI211_X1 U23378 ( .C1(n20539), .C2(n20423), .A(n20399), .B(n20398), .ZN(
        P1_U3115) );
  OAI22_X1 U23379 ( .A1(n20423), .A2(n20543), .B1(n20417), .B2(n20400), .ZN(
        n20401) );
  INV_X1 U23380 ( .A(n20401), .ZN(n20403) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20420), .B1(
        n20593), .B2(n20419), .ZN(n20402) );
  OAI211_X1 U23382 ( .C1(n20597), .C2(n20449), .A(n20403), .B(n20402), .ZN(
        P1_U3116) );
  OAI22_X1 U23383 ( .A1(n20423), .A2(n20547), .B1(n20417), .B2(n20404), .ZN(
        n20405) );
  INV_X1 U23384 ( .A(n20405), .ZN(n20407) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20420), .B1(
        n20599), .B2(n20419), .ZN(n20406) );
  OAI211_X1 U23386 ( .C1(n20603), .C2(n20449), .A(n20407), .B(n20406), .ZN(
        P1_U3117) );
  OAI22_X1 U23387 ( .A1(n20423), .A2(n20551), .B1(n20417), .B2(n20408), .ZN(
        n20409) );
  INV_X1 U23388 ( .A(n20409), .ZN(n20411) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20420), .B1(
        n20605), .B2(n20419), .ZN(n20410) );
  OAI211_X1 U23390 ( .C1(n20609), .C2(n20449), .A(n20411), .B(n20410), .ZN(
        P1_U3118) );
  OAI22_X1 U23391 ( .A1(n20423), .A2(n20555), .B1(n20417), .B2(n20412), .ZN(
        n20413) );
  INV_X1 U23392 ( .A(n20413), .ZN(n20415) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20420), .B1(
        n20611), .B2(n20419), .ZN(n20414) );
  OAI211_X1 U23394 ( .C1(n20615), .C2(n20449), .A(n20415), .B(n20414), .ZN(
        P1_U3119) );
  OAI22_X1 U23395 ( .A1(n20449), .A2(n20626), .B1(n20417), .B2(n20416), .ZN(
        n20418) );
  INV_X1 U23396 ( .A(n20418), .ZN(n20422) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20420), .B1(
        n20619), .B2(n20419), .ZN(n20421) );
  OAI211_X1 U23398 ( .C1(n20563), .C2(n20423), .A(n20422), .B(n20421), .ZN(
        P1_U3120) );
  INV_X1 U23399 ( .A(n20426), .ZN(n20428) );
  NAND2_X1 U23400 ( .A1(n20427), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20429) );
  OAI222_X1 U23401 ( .A1(n20567), .A2(n20428), .B1(n10613), .B2(n20431), .C1(
        n20565), .C2(n20429), .ZN(n20451) );
  INV_X1 U23402 ( .A(n20429), .ZN(n20450) );
  AOI22_X1 U23403 ( .A1(n20569), .A2(n20451), .B1(n20568), .B2(n20450), .ZN(
        n20435) );
  NOR2_X1 U23404 ( .A1(n20430), .A2(n20571), .ZN(n20433) );
  INV_X1 U23405 ( .A(n20431), .ZN(n20432) );
  OAI21_X1 U23406 ( .B1(n20433), .B2(n20432), .A(n20573), .ZN(n20453) );
  AOI22_X1 U23407 ( .A1(n20453), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n20452), .B2(n20576), .ZN(n20434) );
  OAI211_X1 U23408 ( .C1(n20579), .C2(n20486), .A(n20435), .B(n20434), .ZN(
        P1_U3121) );
  AOI22_X1 U23409 ( .A1(n20581), .A2(n20451), .B1(n20580), .B2(n20450), .ZN(
        n20437) );
  INV_X1 U23410 ( .A(n20486), .ZN(n20446) );
  AOI22_X1 U23411 ( .A1(n20453), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n20446), .B2(n20532), .ZN(n20436) );
  OAI211_X1 U23412 ( .C1(n20535), .C2(n20449), .A(n20437), .B(n20436), .ZN(
        P1_U3122) );
  AOI22_X1 U23413 ( .A1(n20587), .A2(n20451), .B1(n20586), .B2(n20450), .ZN(
        n20439) );
  AOI22_X1 U23414 ( .A1(n20453), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n20446), .B2(n20536), .ZN(n20438) );
  OAI211_X1 U23415 ( .C1(n20539), .C2(n20449), .A(n20439), .B(n20438), .ZN(
        P1_U3123) );
  AOI22_X1 U23416 ( .A1(n20593), .A2(n20451), .B1(n20592), .B2(n20450), .ZN(
        n20441) );
  AOI22_X1 U23417 ( .A1(n20453), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n20446), .B2(n20540), .ZN(n20440) );
  OAI211_X1 U23418 ( .C1(n20543), .C2(n20449), .A(n20441), .B(n20440), .ZN(
        P1_U3124) );
  AOI22_X1 U23419 ( .A1(n20599), .A2(n20451), .B1(n20598), .B2(n20450), .ZN(
        n20443) );
  AOI22_X1 U23420 ( .A1(n20453), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n20446), .B2(n20544), .ZN(n20442) );
  OAI211_X1 U23421 ( .C1(n20547), .C2(n20449), .A(n20443), .B(n20442), .ZN(
        P1_U3125) );
  AOI22_X1 U23422 ( .A1(n20605), .A2(n20451), .B1(n20604), .B2(n20450), .ZN(
        n20445) );
  AOI22_X1 U23423 ( .A1(n20453), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n20452), .B2(n20606), .ZN(n20444) );
  OAI211_X1 U23424 ( .C1(n20609), .C2(n20486), .A(n20445), .B(n20444), .ZN(
        P1_U3126) );
  AOI22_X1 U23425 ( .A1(n20611), .A2(n20451), .B1(n20610), .B2(n20450), .ZN(
        n20448) );
  AOI22_X1 U23426 ( .A1(n20453), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n20446), .B2(n20552), .ZN(n20447) );
  OAI211_X1 U23427 ( .C1(n20555), .C2(n20449), .A(n20448), .B(n20447), .ZN(
        P1_U3127) );
  AOI22_X1 U23428 ( .A1(n20619), .A2(n20451), .B1(n20617), .B2(n20450), .ZN(
        n20455) );
  AOI22_X1 U23429 ( .A1(n20453), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n20452), .B2(n20620), .ZN(n20454) );
  OAI211_X1 U23430 ( .C1(n20626), .C2(n20486), .A(n20455), .B(n20454), .ZN(
        P1_U3128) );
  NAND3_X1 U23431 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20457), .ZN(n20491) );
  NOR2_X1 U23432 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20491), .ZN(
        n20481) );
  AOI22_X1 U23433 ( .A1(n20513), .A2(n20528), .B1(n20568), .B2(n20481), .ZN(
        n20468) );
  NAND3_X1 U23434 ( .A1(n20486), .A2(n20496), .A3(n20458), .ZN(n20460) );
  NAND2_X1 U23435 ( .A1(n20460), .A2(n20459), .ZN(n20463) );
  OR2_X1 U23436 ( .A1(n12324), .A2(n20461), .ZN(n20566) );
  OR2_X1 U23437 ( .A1(n20566), .A2(n20517), .ZN(n20465) );
  AOI22_X1 U23438 ( .A1(n20463), .A2(n20465), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20464), .ZN(n20462) );
  OAI211_X1 U23439 ( .C1(n20481), .C2(n20704), .A(n20526), .B(n20462), .ZN(
        n20483) );
  INV_X1 U23440 ( .A(n20463), .ZN(n20466) );
  OAI22_X1 U23441 ( .A1(n20466), .A2(n20465), .B1(n20464), .B2(n20519), .ZN(
        n20482) );
  AOI22_X1 U23442 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20483), .B1(
        n20569), .B2(n20482), .ZN(n20467) );
  OAI211_X1 U23443 ( .C1(n20531), .C2(n20486), .A(n20468), .B(n20467), .ZN(
        P1_U3129) );
  AOI22_X1 U23444 ( .A1(n20513), .A2(n20532), .B1(n20580), .B2(n20481), .ZN(
        n20470) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20483), .B1(
        n20581), .B2(n20482), .ZN(n20469) );
  OAI211_X1 U23446 ( .C1(n20535), .C2(n20486), .A(n20470), .B(n20469), .ZN(
        P1_U3130) );
  AOI22_X1 U23447 ( .A1(n20513), .A2(n20536), .B1(n20586), .B2(n20481), .ZN(
        n20472) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20483), .B1(
        n20587), .B2(n20482), .ZN(n20471) );
  OAI211_X1 U23449 ( .C1(n20539), .C2(n20486), .A(n20472), .B(n20471), .ZN(
        P1_U3131) );
  AOI22_X1 U23450 ( .A1(n20513), .A2(n20540), .B1(n20592), .B2(n20481), .ZN(
        n20474) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20483), .B1(
        n20593), .B2(n20482), .ZN(n20473) );
  OAI211_X1 U23452 ( .C1(n20543), .C2(n20486), .A(n20474), .B(n20473), .ZN(
        P1_U3132) );
  AOI22_X1 U23453 ( .A1(n20513), .A2(n20544), .B1(n20598), .B2(n20481), .ZN(
        n20476) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20483), .B1(
        n20599), .B2(n20482), .ZN(n20475) );
  OAI211_X1 U23455 ( .C1(n20547), .C2(n20486), .A(n20476), .B(n20475), .ZN(
        P1_U3133) );
  AOI22_X1 U23456 ( .A1(n20513), .A2(n20548), .B1(n20604), .B2(n20481), .ZN(
        n20478) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20483), .B1(
        n20605), .B2(n20482), .ZN(n20477) );
  OAI211_X1 U23458 ( .C1(n20551), .C2(n20486), .A(n20478), .B(n20477), .ZN(
        P1_U3134) );
  AOI22_X1 U23459 ( .A1(n20513), .A2(n20552), .B1(n20610), .B2(n20481), .ZN(
        n20480) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20483), .B1(
        n20611), .B2(n20482), .ZN(n20479) );
  OAI211_X1 U23461 ( .C1(n20555), .C2(n20486), .A(n20480), .B(n20479), .ZN(
        P1_U3135) );
  AOI22_X1 U23462 ( .A1(n20513), .A2(n20558), .B1(n20617), .B2(n20481), .ZN(
        n20485) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20483), .B1(
        n20619), .B2(n20482), .ZN(n20484) );
  OAI211_X1 U23464 ( .C1(n20563), .C2(n20486), .A(n20485), .B(n20484), .ZN(
        P1_U3136) );
  INV_X1 U23465 ( .A(n20572), .ZN(n20488) );
  INV_X1 U23466 ( .A(n20566), .ZN(n20518) );
  NOR2_X1 U23467 ( .A1(n20489), .A2(n20491), .ZN(n20511) );
  AOI21_X1 U23468 ( .B1(n20518), .B2(n20490), .A(n20511), .ZN(n20492) );
  OAI22_X1 U23469 ( .A1(n20492), .A2(n20565), .B1(n20491), .B2(n10613), .ZN(
        n20512) );
  AOI22_X1 U23470 ( .A1(n20569), .A2(n20512), .B1(n20568), .B2(n20511), .ZN(
        n20498) );
  INV_X1 U23471 ( .A(n20491), .ZN(n20495) );
  NAND2_X1 U23472 ( .A1(n20493), .A2(n20492), .ZN(n20494) );
  OAI221_X1 U23473 ( .B1(n20496), .B2(n20495), .C1(n20565), .C2(n20494), .A(
        n20573), .ZN(n20514) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20514), .B1(
        n20513), .B2(n20576), .ZN(n20497) );
  OAI211_X1 U23475 ( .C1(n20579), .C2(n20562), .A(n20498), .B(n20497), .ZN(
        P1_U3137) );
  AOI22_X1 U23476 ( .A1(n20581), .A2(n20512), .B1(n20580), .B2(n20511), .ZN(
        n20500) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20514), .B1(
        n20513), .B2(n20582), .ZN(n20499) );
  OAI211_X1 U23478 ( .C1(n20585), .C2(n20562), .A(n20500), .B(n20499), .ZN(
        P1_U3138) );
  AOI22_X1 U23479 ( .A1(n20587), .A2(n20512), .B1(n20586), .B2(n20511), .ZN(
        n20502) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20514), .B1(
        n20513), .B2(n20588), .ZN(n20501) );
  OAI211_X1 U23481 ( .C1(n20591), .C2(n20562), .A(n20502), .B(n20501), .ZN(
        P1_U3139) );
  AOI22_X1 U23482 ( .A1(n20593), .A2(n20512), .B1(n20592), .B2(n20511), .ZN(
        n20504) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20514), .B1(
        n20513), .B2(n20594), .ZN(n20503) );
  OAI211_X1 U23484 ( .C1(n20597), .C2(n20562), .A(n20504), .B(n20503), .ZN(
        P1_U3140) );
  AOI22_X1 U23485 ( .A1(n20599), .A2(n20512), .B1(n20598), .B2(n20511), .ZN(
        n20506) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20514), .B1(
        n20513), .B2(n20600), .ZN(n20505) );
  OAI211_X1 U23487 ( .C1(n20603), .C2(n20562), .A(n20506), .B(n20505), .ZN(
        P1_U3141) );
  AOI22_X1 U23488 ( .A1(n20605), .A2(n20512), .B1(n20604), .B2(n20511), .ZN(
        n20508) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20514), .B1(
        n20513), .B2(n20606), .ZN(n20507) );
  OAI211_X1 U23490 ( .C1(n20609), .C2(n20562), .A(n20508), .B(n20507), .ZN(
        P1_U3142) );
  AOI22_X1 U23491 ( .A1(n20611), .A2(n20512), .B1(n20610), .B2(n20511), .ZN(
        n20510) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20514), .B1(
        n20513), .B2(n20612), .ZN(n20509) );
  OAI211_X1 U23493 ( .C1(n20615), .C2(n20562), .A(n20510), .B(n20509), .ZN(
        P1_U3143) );
  AOI22_X1 U23494 ( .A1(n20619), .A2(n20512), .B1(n20617), .B2(n20511), .ZN(
        n20516) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20514), .B1(
        n20513), .B2(n20620), .ZN(n20515) );
  OAI211_X1 U23496 ( .C1(n20626), .C2(n20562), .A(n20516), .B(n20515), .ZN(
        P1_U3144) );
  NAND2_X1 U23497 ( .A1(n20518), .A2(n20517), .ZN(n20523) );
  OAI22_X1 U23498 ( .A1(n20523), .A2(n20565), .B1(n20520), .B2(n20519), .ZN(
        n20557) );
  NOR2_X1 U23499 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20570), .ZN(
        n20556) );
  AOI22_X1 U23500 ( .A1(n20569), .A2(n20557), .B1(n20568), .B2(n20556), .ZN(
        n20530) );
  INV_X1 U23501 ( .A(n20562), .ZN(n20522) );
  OAI21_X1 U23502 ( .B1(n20522), .B2(n20621), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20524) );
  AOI21_X1 U23503 ( .B1(n20524), .B2(n20523), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20527) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20559), .B1(
        n20621), .B2(n20528), .ZN(n20529) );
  OAI211_X1 U23505 ( .C1(n20531), .C2(n20562), .A(n20530), .B(n20529), .ZN(
        P1_U3145) );
  AOI22_X1 U23506 ( .A1(n20581), .A2(n20557), .B1(n20580), .B2(n20556), .ZN(
        n20534) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20559), .B1(
        n20621), .B2(n20532), .ZN(n20533) );
  OAI211_X1 U23508 ( .C1(n20535), .C2(n20562), .A(n20534), .B(n20533), .ZN(
        P1_U3146) );
  AOI22_X1 U23509 ( .A1(n20587), .A2(n20557), .B1(n20586), .B2(n20556), .ZN(
        n20538) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20559), .B1(
        n20621), .B2(n20536), .ZN(n20537) );
  OAI211_X1 U23511 ( .C1(n20539), .C2(n20562), .A(n20538), .B(n20537), .ZN(
        P1_U3147) );
  AOI22_X1 U23512 ( .A1(n20593), .A2(n20557), .B1(n20592), .B2(n20556), .ZN(
        n20542) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20559), .B1(
        n20621), .B2(n20540), .ZN(n20541) );
  OAI211_X1 U23514 ( .C1(n20543), .C2(n20562), .A(n20542), .B(n20541), .ZN(
        P1_U3148) );
  AOI22_X1 U23515 ( .A1(n20599), .A2(n20557), .B1(n20598), .B2(n20556), .ZN(
        n20546) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20559), .B1(
        n20621), .B2(n20544), .ZN(n20545) );
  OAI211_X1 U23517 ( .C1(n20547), .C2(n20562), .A(n20546), .B(n20545), .ZN(
        P1_U3149) );
  AOI22_X1 U23518 ( .A1(n20605), .A2(n20557), .B1(n20604), .B2(n20556), .ZN(
        n20550) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20559), .B1(
        n20621), .B2(n20548), .ZN(n20549) );
  OAI211_X1 U23520 ( .C1(n20551), .C2(n20562), .A(n20550), .B(n20549), .ZN(
        P1_U3150) );
  AOI22_X1 U23521 ( .A1(n20611), .A2(n20557), .B1(n20610), .B2(n20556), .ZN(
        n20554) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20559), .B1(
        n20621), .B2(n20552), .ZN(n20553) );
  OAI211_X1 U23523 ( .C1(n20555), .C2(n20562), .A(n20554), .B(n20553), .ZN(
        P1_U3151) );
  AOI22_X1 U23524 ( .A1(n20619), .A2(n20557), .B1(n20617), .B2(n20556), .ZN(
        n20561) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20559), .B1(
        n20621), .B2(n20558), .ZN(n20560) );
  OAI211_X1 U23526 ( .C1(n20563), .C2(n20562), .A(n20561), .B(n20560), .ZN(
        P1_U3152) );
  INV_X1 U23527 ( .A(n20616), .ZN(n20564) );
  OAI222_X1 U23528 ( .A1(n20567), .A2(n20566), .B1(n10613), .B2(n20570), .C1(
        n20565), .C2(n20564), .ZN(n20618) );
  AOI22_X1 U23529 ( .A1(n20569), .A2(n20618), .B1(n20568), .B2(n20616), .ZN(
        n20578) );
  INV_X1 U23530 ( .A(n20570), .ZN(n20575) );
  NOR2_X1 U23531 ( .A1(n20572), .A2(n20571), .ZN(n20574) );
  OAI21_X1 U23532 ( .B1(n20575), .B2(n20574), .A(n20573), .ZN(n20622) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20576), .ZN(n20577) );
  OAI211_X1 U23534 ( .C1(n20579), .C2(n20625), .A(n20578), .B(n20577), .ZN(
        P1_U3153) );
  AOI22_X1 U23535 ( .A1(n20581), .A2(n20618), .B1(n20580), .B2(n20616), .ZN(
        n20584) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20582), .ZN(n20583) );
  OAI211_X1 U23537 ( .C1(n20585), .C2(n20625), .A(n20584), .B(n20583), .ZN(
        P1_U3154) );
  AOI22_X1 U23538 ( .A1(n20587), .A2(n20618), .B1(n20586), .B2(n20616), .ZN(
        n20590) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20588), .ZN(n20589) );
  OAI211_X1 U23540 ( .C1(n20591), .C2(n20625), .A(n20590), .B(n20589), .ZN(
        P1_U3155) );
  AOI22_X1 U23541 ( .A1(n20593), .A2(n20618), .B1(n20592), .B2(n20616), .ZN(
        n20596) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20594), .ZN(n20595) );
  OAI211_X1 U23543 ( .C1(n20597), .C2(n20625), .A(n20596), .B(n20595), .ZN(
        P1_U3156) );
  AOI22_X1 U23544 ( .A1(n20599), .A2(n20618), .B1(n20598), .B2(n20616), .ZN(
        n20602) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20600), .ZN(n20601) );
  OAI211_X1 U23546 ( .C1(n20603), .C2(n20625), .A(n20602), .B(n20601), .ZN(
        P1_U3157) );
  AOI22_X1 U23547 ( .A1(n20605), .A2(n20618), .B1(n20604), .B2(n20616), .ZN(
        n20608) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20606), .ZN(n20607) );
  OAI211_X1 U23549 ( .C1(n20609), .C2(n20625), .A(n20608), .B(n20607), .ZN(
        P1_U3158) );
  AOI22_X1 U23550 ( .A1(n20611), .A2(n20618), .B1(n20610), .B2(n20616), .ZN(
        n20614) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20612), .ZN(n20613) );
  OAI211_X1 U23552 ( .C1(n20615), .C2(n20625), .A(n20614), .B(n20613), .ZN(
        P1_U3159) );
  AOI22_X1 U23553 ( .A1(n20619), .A2(n20618), .B1(n20617), .B2(n20616), .ZN(
        n20624) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20622), .B1(
        n20621), .B2(n20620), .ZN(n20623) );
  OAI211_X1 U23555 ( .C1(n20626), .C2(n20625), .A(n20624), .B(n20623), .ZN(
        P1_U3160) );
  NOR2_X1 U23556 ( .A1(n10081), .A2(n20627), .ZN(n20629) );
  OAI21_X1 U23557 ( .B1(n20629), .B2(n10613), .A(n20628), .ZN(P1_U3163) );
  AND2_X1 U23558 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20699), .ZN(
        P1_U3164) );
  AND2_X1 U23559 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20699), .ZN(
        P1_U3165) );
  AND2_X1 U23560 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20699), .ZN(
        P1_U3166) );
  AND2_X1 U23561 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20699), .ZN(
        P1_U3167) );
  AND2_X1 U23562 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20699), .ZN(
        P1_U3168) );
  AND2_X1 U23563 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20699), .ZN(
        P1_U3169) );
  AND2_X1 U23564 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20699), .ZN(
        P1_U3170) );
  AND2_X1 U23565 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20699), .ZN(
        P1_U3171) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20699), .ZN(
        P1_U3172) );
  AND2_X1 U23567 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20699), .ZN(
        P1_U3173) );
  AND2_X1 U23568 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20699), .ZN(
        P1_U3174) );
  AND2_X1 U23569 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20699), .ZN(
        P1_U3175) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20699), .ZN(
        P1_U3176) );
  AND2_X1 U23571 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20699), .ZN(
        P1_U3177) );
  AND2_X1 U23572 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20699), .ZN(
        P1_U3178) );
  AND2_X1 U23573 ( .A1(n20699), .A2(P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(
        P1_U3179) );
  AND2_X1 U23574 ( .A1(n20699), .A2(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(
        P1_U3180) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20699), .ZN(
        P1_U3181) );
  INV_X1 U23576 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20975) );
  NOR2_X1 U23577 ( .A1(n20703), .A2(n20975), .ZN(P1_U3182) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20699), .ZN(
        P1_U3183) );
  AND2_X1 U23579 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20699), .ZN(
        P1_U3184) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20699), .ZN(
        P1_U3185) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20699), .ZN(P1_U3186) );
  AND2_X1 U23582 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20699), .ZN(P1_U3187) );
  AND2_X1 U23583 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20699), .ZN(P1_U3188) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20699), .ZN(P1_U3189) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20699), .ZN(P1_U3190) );
  AND2_X1 U23586 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20699), .ZN(P1_U3191) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20699), .ZN(P1_U3192) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20699), .ZN(P1_U3193) );
  AOI21_X1 U23589 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20635), .A(n20630), 
        .ZN(n20641) );
  NOR2_X1 U23590 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20631) );
  OAI22_X1 U23591 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20986), .B1(n20631), 
        .B2(n20742), .ZN(n20632) );
  NOR2_X1 U23592 ( .A1(n20636), .A2(n20632), .ZN(n20633) );
  OAI22_X1 U23593 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20641), .B1(n20667), 
        .B2(n20633), .ZN(P1_U3194) );
  AOI21_X1 U23594 ( .B1(n20635), .B2(n20986), .A(n20634), .ZN(n20643) );
  OAI211_X1 U23595 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20636), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20642) );
  INV_X1 U23596 ( .A(n20637), .ZN(n20638) );
  AOI221_X1 U23597 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20986), .C1(n20639), 
        .C2(n20986), .A(n20638), .ZN(n20640) );
  OAI22_X1 U23598 ( .A1(n20643), .A2(n20642), .B1(n20641), .B2(n20640), .ZN(
        P1_U3196) );
  INV_X1 U23599 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20645) );
  AND2_X1 U23600 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20739), .ZN(n20691) );
  NOR2_X1 U23601 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20736), .ZN(n20687) );
  AOI22_X1 U23602 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20736), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20687), .ZN(n20644) );
  OAI21_X1 U23603 ( .B1(n20645), .B2(n20689), .A(n20644), .ZN(P1_U3197) );
  INV_X1 U23604 ( .A(n20687), .ZN(n20693) );
  AOI22_X1 U23605 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20736), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20691), .ZN(n20646) );
  OAI21_X1 U23606 ( .B1(n20649), .B2(n20693), .A(n20646), .ZN(P1_U3198) );
  OAI222_X1 U23607 ( .A1(n20689), .A2(n20649), .B1(n20648), .B2(n20739), .C1(
        n20647), .C2(n20693), .ZN(P1_U3199) );
  AOI222_X1 U23608 ( .A1(n20687), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20691), .ZN(n20650) );
  INV_X1 U23609 ( .A(n20650), .ZN(P1_U3200) );
  AOI222_X1 U23610 ( .A1(n20691), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20736), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20687), .ZN(n20651) );
  INV_X1 U23611 ( .A(n20651), .ZN(P1_U3201) );
  INV_X1 U23612 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20652) );
  OAI222_X1 U23613 ( .A1(n20689), .A2(n13022), .B1(n20652), .B2(n20667), .C1(
        n20654), .C2(n20693), .ZN(P1_U3202) );
  INV_X1 U23614 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20653) );
  OAI222_X1 U23615 ( .A1(n20689), .A2(n20654), .B1(n20653), .B2(n20667), .C1(
        n21024), .C2(n20693), .ZN(P1_U3203) );
  INV_X1 U23616 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20655) );
  OAI222_X1 U23617 ( .A1(n20693), .A2(n13104), .B1(n20655), .B2(n20667), .C1(
        n21024), .C2(n20689), .ZN(P1_U3204) );
  INV_X1 U23618 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20656) );
  OAI222_X1 U23619 ( .A1(n20689), .A2(n13104), .B1(n20656), .B2(n20667), .C1(
        n14388), .C2(n20693), .ZN(P1_U3205) );
  INV_X1 U23620 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20657) );
  OAI222_X1 U23621 ( .A1(n20689), .A2(n14388), .B1(n20657), .B2(n20667), .C1(
        n20659), .C2(n20693), .ZN(P1_U3206) );
  AOI22_X1 U23622 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20736), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20687), .ZN(n20658) );
  OAI21_X1 U23623 ( .B1(n20659), .B2(n20689), .A(n20658), .ZN(P1_U3207) );
  AOI22_X1 U23624 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20736), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20691), .ZN(n20660) );
  OAI21_X1 U23625 ( .B1(n20662), .B2(n20693), .A(n20660), .ZN(P1_U3208) );
  AOI22_X1 U23626 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20736), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20687), .ZN(n20661) );
  OAI21_X1 U23627 ( .B1(n20662), .B2(n20689), .A(n20661), .ZN(P1_U3209) );
  AOI22_X1 U23628 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20736), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20691), .ZN(n20663) );
  OAI21_X1 U23629 ( .B1(n20665), .B2(n20693), .A(n20663), .ZN(P1_U3210) );
  INV_X1 U23630 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20664) );
  OAI222_X1 U23631 ( .A1(n20689), .A2(n20665), .B1(n20664), .B2(n20667), .C1(
        n14355), .C2(n20693), .ZN(P1_U3211) );
  INV_X1 U23632 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20666) );
  OAI222_X1 U23633 ( .A1(n20689), .A2(n14355), .B1(n20666), .B2(n20667), .C1(
        n20669), .C2(n20693), .ZN(P1_U3212) );
  INV_X1 U23634 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20668) );
  OAI222_X1 U23635 ( .A1(n20689), .A2(n20669), .B1(n20668), .B2(n20667), .C1(
        n20671), .C2(n20693), .ZN(P1_U3213) );
  INV_X1 U23636 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20670) );
  OAI222_X1 U23637 ( .A1(n20689), .A2(n20671), .B1(n20670), .B2(n20739), .C1(
        n20672), .C2(n20693), .ZN(P1_U3214) );
  INV_X1 U23638 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20850) );
  OAI222_X1 U23639 ( .A1(n20693), .A2(n20674), .B1(n20850), .B2(n20739), .C1(
        n20672), .C2(n20689), .ZN(P1_U3215) );
  INV_X1 U23640 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20673) );
  OAI222_X1 U23641 ( .A1(n20689), .A2(n20674), .B1(n20673), .B2(n20739), .C1(
        n20676), .C2(n20693), .ZN(P1_U3216) );
  INV_X1 U23642 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20675) );
  OAI222_X1 U23643 ( .A1(n20689), .A2(n20676), .B1(n20675), .B2(n20739), .C1(
        n20677), .C2(n20693), .ZN(P1_U3217) );
  INV_X1 U23644 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20891) );
  INV_X1 U23645 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20679) );
  OAI222_X1 U23646 ( .A1(n20689), .A2(n20677), .B1(n20891), .B2(n20739), .C1(
        n20679), .C2(n20693), .ZN(P1_U3218) );
  INV_X1 U23647 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20678) );
  OAI222_X1 U23648 ( .A1(n20689), .A2(n20679), .B1(n20678), .B2(n20739), .C1(
        n20681), .C2(n20693), .ZN(P1_U3219) );
  INV_X1 U23649 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20680) );
  OAI222_X1 U23650 ( .A1(n20689), .A2(n20681), .B1(n20680), .B2(n20739), .C1(
        n20683), .C2(n20693), .ZN(P1_U3220) );
  INV_X1 U23651 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20682) );
  OAI222_X1 U23652 ( .A1(n20689), .A2(n20683), .B1(n20682), .B2(n20739), .C1(
        n20856), .C2(n20693), .ZN(P1_U3221) );
  INV_X1 U23653 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20684) );
  OAI222_X1 U23654 ( .A1(n20689), .A2(n20856), .B1(n20684), .B2(n20739), .C1(
        n20985), .C2(n20693), .ZN(P1_U3222) );
  INV_X1 U23655 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21040) );
  INV_X1 U23656 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n20686) );
  OAI222_X1 U23657 ( .A1(n20689), .A2(n20985), .B1(n21040), .B2(n20739), .C1(
        n20686), .C2(n20693), .ZN(P1_U3223) );
  INV_X1 U23658 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20685) );
  OAI222_X1 U23659 ( .A1(n20689), .A2(n20686), .B1(n20685), .B2(n20739), .C1(
        n20690), .C2(n20693), .ZN(P1_U3224) );
  AOI22_X1 U23660 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20687), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20736), .ZN(n20688) );
  OAI21_X1 U23661 ( .B1(n20690), .B2(n20689), .A(n20688), .ZN(P1_U3225) );
  AOI22_X1 U23662 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20691), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20736), .ZN(n20692) );
  OAI21_X1 U23663 ( .B1(n20694), .B2(n20693), .A(n20692), .ZN(P1_U3226) );
  MUX2_X1 U23664 ( .A(P1_BE_N_REG_3__SCAN_IN), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .S(n20739), .Z(P1_U3458) );
  MUX2_X1 U23665 ( .A(P1_BE_N_REG_2__SCAN_IN), .B(P1_BYTEENABLE_REG_2__SCAN_IN), .S(n20739), .Z(P1_U3459) );
  INV_X1 U23666 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20695) );
  AOI22_X1 U23667 ( .A1(n20739), .A2(n20696), .B1(n20695), .B2(n20736), .ZN(
        P1_U3460) );
  INV_X1 U23668 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20719) );
  INV_X1 U23669 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20697) );
  AOI22_X1 U23670 ( .A1(n20739), .A2(n20719), .B1(n20697), .B2(n20736), .ZN(
        P1_U3461) );
  INV_X1 U23671 ( .A(n20701), .ZN(n20698) );
  AOI21_X1 U23672 ( .B1(n20700), .B2(n20699), .A(n20698), .ZN(P1_U3464) );
  OAI21_X1 U23673 ( .B1(n20703), .B2(n20702), .A(n20701), .ZN(P1_U3465) );
  AOI21_X1 U23674 ( .B1(n20705), .B2(n20704), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n20707) );
  OAI22_X1 U23675 ( .A1(n20708), .A2(n20707), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20706), .ZN(n20710) );
  AOI22_X1 U23676 ( .A1(n20711), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20710), .B2(n20709), .ZN(n20712) );
  OAI21_X1 U23677 ( .B1(n20714), .B2(n20713), .A(n20712), .ZN(P1_U3474) );
  NAND2_X1 U23678 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20718) );
  INV_X1 U23679 ( .A(n20722), .ZN(n20715) );
  AOI211_X1 U23680 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(n20715), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20716) );
  AOI21_X1 U23681 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n20720), .A(n20716), 
        .ZN(n20717) );
  OAI21_X1 U23682 ( .B1(n20718), .B2(n20720), .A(n20717), .ZN(P1_U3481) );
  AOI22_X1 U23683 ( .A1(n20722), .A2(n20721), .B1(n20720), .B2(n20719), .ZN(
        P1_U3482) );
  INV_X1 U23684 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20723) );
  AOI22_X1 U23685 ( .A1(n20739), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20723), 
        .B2(n20736), .ZN(P1_U3483) );
  AOI211_X1 U23686 ( .C1(n20727), .C2(n20726), .A(n20725), .B(n20724), .ZN(
        n20735) );
  OAI211_X1 U23687 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20729), .A(n20728), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20732) );
  INV_X1 U23688 ( .A(n20730), .ZN(n20731) );
  AOI21_X1 U23689 ( .B1(n20732), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20731), 
        .ZN(n20734) );
  NAND2_X1 U23690 ( .A1(n20735), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20733) );
  OAI21_X1 U23691 ( .B1(n20735), .B2(n20734), .A(n20733), .ZN(P1_U3485) );
  AOI22_X1 U23692 ( .A1(n20739), .A2(n20738), .B1(n20737), .B2(n20736), .ZN(
        P1_U3486) );
  INV_X1 U23693 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20746) );
  AOI211_X1 U23694 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20742), .A(
        n20741), .B(n20740), .ZN(n20743) );
  AOI221_X1 U23695 ( .B1(n20746), .B2(n20745), .C1(n20744), .C2(n20745), .A(
        n20743), .ZN(n21136) );
  AOI22_X1 U23696 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(keyinput139), .B1(
        P1_INSTQUEUE_REG_14__0__SCAN_IN), .B2(keyinput243), .ZN(n20747) );
  OAI221_X1 U23697 ( .B1(P1_ADDRESS_REG_3__SCAN_IN), .B2(keyinput139), .C1(
        P1_INSTQUEUE_REG_14__0__SCAN_IN), .C2(keyinput243), .A(n20747), .ZN(
        n20754) );
  AOI22_X1 U23698 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(keyinput216), .B1(
        P1_INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput131), .ZN(n20748) );
  OAI221_X1 U23699 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(keyinput216), .C1(
        P1_INSTQUEUE_REG_7__5__SCAN_IN), .C2(keyinput131), .A(n20748), .ZN(
        n20753) );
  AOI22_X1 U23700 ( .A1(BUF2_REG_18__SCAN_IN), .A2(keyinput253), .B1(
        P2_STATE2_REG_0__SCAN_IN), .B2(keyinput215), .ZN(n20749) );
  OAI221_X1 U23701 ( .B1(BUF2_REG_18__SCAN_IN), .B2(keyinput253), .C1(
        P2_STATE2_REG_0__SCAN_IN), .C2(keyinput215), .A(n20749), .ZN(n20752)
         );
  AOI22_X1 U23702 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput170), .B1(
        P3_EAX_REG_3__SCAN_IN), .B2(keyinput238), .ZN(n20750) );
  OAI221_X1 U23703 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput170), .C1(
        P3_EAX_REG_3__SCAN_IN), .C2(keyinput238), .A(n20750), .ZN(n20751) );
  NOR4_X1 U23704 ( .A1(n20754), .A2(n20753), .A3(n20752), .A4(n20751), .ZN(
        n20782) );
  AOI22_X1 U23705 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput169), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput165), .ZN(n20755) );
  OAI221_X1 U23706 ( .B1(P2_DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput169), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput165), .A(n20755), .ZN(n20762) );
  AOI22_X1 U23707 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(keyinput181), .B1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput155), .ZN(n20756) );
  OAI221_X1 U23708 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(keyinput181), .C1(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(keyinput155), .A(n20756), 
        .ZN(n20761) );
  AOI22_X1 U23709 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput205), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput234), .ZN(n20757) );
  OAI221_X1 U23710 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput205), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput234), .A(n20757), .ZN(n20760)
         );
  AOI22_X1 U23711 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(keyinput133), 
        .B1(P2_EAX_REG_28__SCAN_IN), .B2(keyinput223), .ZN(n20758) );
  OAI221_X1 U23712 ( .B1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(keyinput133), 
        .C1(P2_EAX_REG_28__SCAN_IN), .C2(keyinput223), .A(n20758), .ZN(n20759)
         );
  NOR4_X1 U23713 ( .A1(n20762), .A2(n20761), .A3(n20760), .A4(n20759), .ZN(
        n20781) );
  AOI22_X1 U23714 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(keyinput247), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(keyinput128), .ZN(n20763) );
  OAI221_X1 U23715 ( .B1(P1_DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput247), .C1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(keyinput128), .A(n20763), 
        .ZN(n20770) );
  AOI22_X1 U23716 ( .A1(P1_EBX_REG_28__SCAN_IN), .A2(keyinput226), .B1(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .B2(keyinput197), .ZN(n20764) );
  OAI221_X1 U23717 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(keyinput226), .C1(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .C2(keyinput197), .A(n20764), .ZN(
        n20769) );
  AOI22_X1 U23718 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(keyinput210), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(keyinput246), .ZN(n20765) );
  OAI221_X1 U23719 ( .B1(P3_DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput210), .C1(
        P3_UWORD_REG_7__SCAN_IN), .C2(keyinput246), .A(n20765), .ZN(n20768) );
  AOI22_X1 U23720 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(keyinput239), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(keyinput245), .ZN(n20766) );
  OAI221_X1 U23721 ( .B1(P3_W_R_N_REG_SCAN_IN), .B2(keyinput239), .C1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .C2(keyinput245), .A(n20766), .ZN(
        n20767) );
  NOR4_X1 U23722 ( .A1(n20770), .A2(n20769), .A3(n20768), .A4(n20767), .ZN(
        n20780) );
  AOI22_X1 U23723 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput136), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput217), .ZN(n20771) );
  OAI221_X1 U23724 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput136), .C1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput217), .A(n20771), .ZN(
        n20778) );
  AOI22_X1 U23725 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(keyinput164), 
        .B1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B2(keyinput183), .ZN(n20772) );
  OAI221_X1 U23726 ( .B1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput164), 
        .C1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .C2(keyinput183), .A(n20772), 
        .ZN(n20777) );
  AOI22_X1 U23727 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(keyinput224), .B1(
        P3_STATE2_REG_0__SCAN_IN), .B2(keyinput129), .ZN(n20773) );
  OAI221_X1 U23728 ( .B1(P1_DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput224), .C1(
        P3_STATE2_REG_0__SCAN_IN), .C2(keyinput129), .A(n20773), .ZN(n20776)
         );
  AOI22_X1 U23729 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput132), .B1(
        P2_INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput206), .ZN(n20774) );
  OAI221_X1 U23730 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput132), .C1(
        P2_INSTQUEUE_REG_10__5__SCAN_IN), .C2(keyinput206), .A(n20774), .ZN(
        n20775) );
  NOR4_X1 U23731 ( .A1(n20778), .A2(n20777), .A3(n20776), .A4(n20775), .ZN(
        n20779) );
  NAND4_X1 U23732 ( .A1(n20782), .A2(n20781), .A3(n20780), .A4(n20779), .ZN(
        n20936) );
  AOI22_X1 U23733 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(keyinput218), 
        .B1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B2(keyinput207), .ZN(n20783) );
  OAI221_X1 U23734 ( .B1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B2(keyinput218), 
        .C1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .C2(keyinput207), .A(n20783), 
        .ZN(n20790) );
  AOI22_X1 U23735 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(keyinput244), .B1(
        NA), .B2(keyinput213), .ZN(n20784) );
  OAI221_X1 U23736 ( .B1(P3_DATAWIDTH_REG_27__SCAN_IN), .B2(keyinput244), .C1(
        NA), .C2(keyinput213), .A(n20784), .ZN(n20789) );
  AOI22_X1 U23737 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(keyinput178), .B1(
        P2_INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput222), .ZN(n20785) );
  OAI221_X1 U23738 ( .B1(P1_DATAWIDTH_REG_13__SCAN_IN), .B2(keyinput178), .C1(
        P2_INSTQUEUE_REG_12__0__SCAN_IN), .C2(keyinput222), .A(n20785), .ZN(
        n20788) );
  AOI22_X1 U23739 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(keyinput142), .B1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput147), .ZN(n20786) );
  OAI221_X1 U23740 ( .B1(P1_ADDRESS_REG_25__SCAN_IN), .B2(keyinput142), .C1(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(keyinput147), .A(n20786), 
        .ZN(n20787) );
  NOR4_X1 U23741 ( .A1(n20790), .A2(n20789), .A3(n20788), .A4(n20787), .ZN(
        n20822) );
  AOI22_X1 U23742 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput241), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(keyinput251), .ZN(n20791) );
  OAI221_X1 U23743 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput241), .C1(
        P1_UWORD_REG_4__SCAN_IN), .C2(keyinput251), .A(n20791), .ZN(n20798) );
  AOI22_X1 U23744 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(keyinput163), 
        .B1(P2_EAX_REG_15__SCAN_IN), .B2(keyinput182), .ZN(n20792) );
  OAI221_X1 U23745 ( .B1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput163), 
        .C1(P2_EAX_REG_15__SCAN_IN), .C2(keyinput182), .A(n20792), .ZN(n20797)
         );
  AOI22_X1 U23746 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(keyinput185), .B1(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput229), .ZN(n20793) );
  OAI221_X1 U23747 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(keyinput185), .C1(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(keyinput229), .A(n20793), .ZN(
        n20796) );
  AOI22_X1 U23748 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(keyinput248), 
        .B1(P2_REIP_REG_30__SCAN_IN), .B2(keyinput249), .ZN(n20794) );
  OAI221_X1 U23749 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(keyinput248), 
        .C1(P2_REIP_REG_30__SCAN_IN), .C2(keyinput249), .A(n20794), .ZN(n20795) );
  NOR4_X1 U23750 ( .A1(n20798), .A2(n20797), .A3(n20796), .A4(n20795), .ZN(
        n20821) );
  AOI22_X1 U23751 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(keyinput166), 
        .B1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(keyinput153), .ZN(n20799) );
  OAI221_X1 U23752 ( .B1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(keyinput166), 
        .C1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .C2(keyinput153), .A(n20799), 
        .ZN(n20806) );
  AOI22_X1 U23753 ( .A1(P3_ADDRESS_REG_26__SCAN_IN), .A2(keyinput154), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(keyinput137), .ZN(n20800) );
  OAI221_X1 U23754 ( .B1(P3_ADDRESS_REG_26__SCAN_IN), .B2(keyinput154), .C1(
        P1_REIP_REG_8__SCAN_IN), .C2(keyinput137), .A(n20800), .ZN(n20805) );
  AOI22_X1 U23755 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(keyinput171), 
        .B1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput203), .ZN(n20801)
         );
  OAI221_X1 U23756 ( .B1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(keyinput171), 
        .C1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput203), .A(n20801), 
        .ZN(n20804) );
  AOI22_X1 U23757 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(keyinput200), .B1(
        P1_INSTQUEUE_REG_3__1__SCAN_IN), .B2(keyinput221), .ZN(n20802) );
  OAI221_X1 U23758 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(keyinput200), .C1(
        P1_INSTQUEUE_REG_3__1__SCAN_IN), .C2(keyinput221), .A(n20802), .ZN(
        n20803) );
  NOR4_X1 U23759 ( .A1(n20806), .A2(n20805), .A3(n20804), .A4(n20803), .ZN(
        n20820) );
  AOI22_X1 U23760 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(keyinput161), 
        .B1(n20808), .B2(keyinput174), .ZN(n20807) );
  OAI221_X1 U23761 ( .B1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B2(keyinput161), 
        .C1(n20808), .C2(keyinput174), .A(n20807), .ZN(n20818) );
  AOI22_X1 U23762 ( .A1(n20954), .A2(keyinput162), .B1(n10025), .B2(
        keyinput173), .ZN(n20809) );
  OAI221_X1 U23763 ( .B1(n20954), .B2(keyinput162), .C1(n10025), .C2(
        keyinput173), .A(n20809), .ZN(n20817) );
  AOI22_X1 U23764 ( .A1(n20811), .A2(keyinput141), .B1(n21047), .B2(
        keyinput152), .ZN(n20810) );
  OAI221_X1 U23765 ( .B1(n20811), .B2(keyinput141), .C1(n21047), .C2(
        keyinput152), .A(n20810), .ZN(n20816) );
  AOI22_X1 U23766 ( .A1(n20814), .A2(keyinput160), .B1(keyinput158), .B2(
        n20813), .ZN(n20812) );
  OAI221_X1 U23767 ( .B1(n20814), .B2(keyinput160), .C1(n20813), .C2(
        keyinput158), .A(n20812), .ZN(n20815) );
  NOR4_X1 U23768 ( .A1(n20818), .A2(n20817), .A3(n20816), .A4(n20815), .ZN(
        n20819) );
  NAND4_X1 U23769 ( .A1(n20822), .A2(n20821), .A3(n20820), .A4(n20819), .ZN(
        n20935) );
  INV_X1 U23770 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n20953) );
  INV_X1 U23771 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20824) );
  AOI22_X1 U23772 ( .A1(n20953), .A2(keyinput193), .B1(n20824), .B2(
        keyinput194), .ZN(n20823) );
  OAI221_X1 U23773 ( .B1(n20953), .B2(keyinput193), .C1(n20824), .C2(
        keyinput194), .A(n20823), .ZN(n20834) );
  INV_X1 U23774 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n20826) );
  AOI22_X1 U23775 ( .A1(n20973), .A2(keyinput184), .B1(n20826), .B2(
        keyinput233), .ZN(n20825) );
  OAI221_X1 U23776 ( .B1(n20973), .B2(keyinput184), .C1(n20826), .C2(
        keyinput233), .A(n20825), .ZN(n20833) );
  AOI22_X1 U23777 ( .A1(n20948), .A2(keyinput212), .B1(n20828), .B2(
        keyinput176), .ZN(n20827) );
  OAI221_X1 U23778 ( .B1(n20948), .B2(keyinput212), .C1(n20828), .C2(
        keyinput176), .A(n20827), .ZN(n20832) );
  INV_X1 U23779 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20830) );
  AOI22_X1 U23780 ( .A1(n20830), .A2(keyinput172), .B1(n10032), .B2(
        keyinput235), .ZN(n20829) );
  OAI221_X1 U23781 ( .B1(n20830), .B2(keyinput172), .C1(n10032), .C2(
        keyinput235), .A(n20829), .ZN(n20831) );
  NOR4_X1 U23782 ( .A1(n20834), .A2(n20833), .A3(n20832), .A4(n20831), .ZN(
        n20877) );
  AOI22_X1 U23783 ( .A1(n20836), .A2(keyinput144), .B1(n21038), .B2(
        keyinput146), .ZN(n20835) );
  OAI221_X1 U23784 ( .B1(n20836), .B2(keyinput144), .C1(n21038), .C2(
        keyinput146), .A(n20835), .ZN(n20839) );
  XOR2_X1 U23785 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B(keyinput240), .Z(
        n20838) );
  XNOR2_X1 U23786 ( .A(n21040), .B(keyinput220), .ZN(n20837) );
  OR3_X1 U23787 ( .A1(n20839), .A2(n20838), .A3(n20837), .ZN(n20848) );
  AOI22_X1 U23788 ( .A1(n20842), .A2(keyinput148), .B1(n20841), .B2(
        keyinput156), .ZN(n20840) );
  OAI221_X1 U23789 ( .B1(n20842), .B2(keyinput148), .C1(n20841), .C2(
        keyinput156), .A(n20840), .ZN(n20847) );
  AOI22_X1 U23790 ( .A1(n20845), .A2(keyinput195), .B1(keyinput157), .B2(
        n20844), .ZN(n20843) );
  OAI221_X1 U23791 ( .B1(n20845), .B2(keyinput195), .C1(n20844), .C2(
        keyinput157), .A(n20843), .ZN(n20846) );
  NOR3_X1 U23792 ( .A1(n20848), .A2(n20847), .A3(n20846), .ZN(n20876) );
  INV_X1 U23793 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n20851) );
  AOI22_X1 U23794 ( .A1(n20851), .A2(keyinput237), .B1(n20850), .B2(
        keyinput211), .ZN(n20849) );
  OAI221_X1 U23795 ( .B1(n20851), .B2(keyinput237), .C1(n20850), .C2(
        keyinput211), .A(n20849), .ZN(n20863) );
  INV_X1 U23796 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20854) );
  AOI22_X1 U23797 ( .A1(n20854), .A2(keyinput214), .B1(n20853), .B2(
        keyinput151), .ZN(n20852) );
  OAI221_X1 U23798 ( .B1(n20854), .B2(keyinput214), .C1(n20853), .C2(
        keyinput151), .A(n20852), .ZN(n20862) );
  AOI22_X1 U23799 ( .A1(n20945), .A2(keyinput255), .B1(keyinput236), .B2(
        n20856), .ZN(n20855) );
  OAI221_X1 U23800 ( .B1(n20945), .B2(keyinput255), .C1(n20856), .C2(
        keyinput236), .A(n20855), .ZN(n20861) );
  INV_X1 U23801 ( .A(P3_LWORD_REG_11__SCAN_IN), .ZN(n20859) );
  AOI22_X1 U23802 ( .A1(n20859), .A2(keyinput189), .B1(keyinput228), .B2(
        n20858), .ZN(n20857) );
  OAI221_X1 U23803 ( .B1(n20859), .B2(keyinput189), .C1(n20858), .C2(
        keyinput228), .A(n20857), .ZN(n20860) );
  NOR4_X1 U23804 ( .A1(n20863), .A2(n20862), .A3(n20861), .A4(n20860), .ZN(
        n20875) );
  AOI22_X1 U23805 ( .A1(n13878), .A2(keyinput202), .B1(keyinput252), .B2(
        n21037), .ZN(n20864) );
  OAI221_X1 U23806 ( .B1(n13878), .B2(keyinput202), .C1(n21037), .C2(
        keyinput252), .A(n20864), .ZN(n20873) );
  INV_X1 U23807 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n21032) );
  AOI22_X1 U23808 ( .A1(n21032), .A2(keyinput204), .B1(n20866), .B2(
        keyinput201), .ZN(n20865) );
  OAI221_X1 U23809 ( .B1(n21032), .B2(keyinput204), .C1(n20866), .C2(
        keyinput201), .A(n20865), .ZN(n20872) );
  AOI22_X1 U23810 ( .A1(n14764), .A2(keyinput130), .B1(n10070), .B2(
        keyinput149), .ZN(n20867) );
  OAI221_X1 U23811 ( .B1(n14764), .B2(keyinput130), .C1(n10070), .C2(
        keyinput149), .A(n20867), .ZN(n20871) );
  AOI22_X1 U23812 ( .A1(n20982), .A2(keyinput186), .B1(keyinput140), .B2(
        n20869), .ZN(n20868) );
  OAI221_X1 U23813 ( .B1(n20982), .B2(keyinput186), .C1(n20869), .C2(
        keyinput140), .A(n20868), .ZN(n20870) );
  NOR4_X1 U23814 ( .A1(n20873), .A2(n20872), .A3(n20871), .A4(n20870), .ZN(
        n20874) );
  NAND4_X1 U23815 ( .A1(n20877), .A2(n20876), .A3(n20875), .A4(n20874), .ZN(
        n20934) );
  INV_X1 U23816 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20967) );
  AOI22_X1 U23817 ( .A1(n21014), .A2(keyinput180), .B1(n20967), .B2(
        keyinput199), .ZN(n20878) );
  OAI221_X1 U23818 ( .B1(n21014), .B2(keyinput180), .C1(n20967), .C2(
        keyinput199), .A(n20878), .ZN(n20888) );
  INV_X1 U23819 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n20972) );
  AOI22_X1 U23820 ( .A1(n20970), .A2(keyinput159), .B1(keyinput190), .B2(
        n20972), .ZN(n20879) );
  OAI221_X1 U23821 ( .B1(n20970), .B2(keyinput159), .C1(n20972), .C2(
        keyinput190), .A(n20879), .ZN(n20887) );
  AOI22_X1 U23822 ( .A1(n20882), .A2(keyinput167), .B1(keyinput198), .B2(
        n20881), .ZN(n20880) );
  OAI221_X1 U23823 ( .B1(n20882), .B2(keyinput167), .C1(n20881), .C2(
        keyinput198), .A(n20880), .ZN(n20886) );
  INV_X1 U23824 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n20947) );
  AOI22_X1 U23825 ( .A1(n20947), .A2(keyinput225), .B1(n20884), .B2(
        keyinput177), .ZN(n20883) );
  OAI221_X1 U23826 ( .B1(n20947), .B2(keyinput225), .C1(n20884), .C2(
        keyinput177), .A(n20883), .ZN(n20885) );
  NOR4_X1 U23827 ( .A1(n20888), .A2(n20887), .A3(n20886), .A4(n20885), .ZN(
        n20932) );
  INV_X1 U23828 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U23829 ( .A1(n20891), .A2(keyinput196), .B1(keyinput145), .B2(
        n20890), .ZN(n20889) );
  OAI221_X1 U23830 ( .B1(n20891), .B2(keyinput196), .C1(n20890), .C2(
        keyinput145), .A(n20889), .ZN(n20901) );
  INV_X1 U23831 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23832 ( .A1(n20894), .A2(keyinput168), .B1(keyinput179), .B2(
        n20893), .ZN(n20892) );
  OAI221_X1 U23833 ( .B1(n20894), .B2(keyinput168), .C1(n20893), .C2(
        keyinput179), .A(n20892), .ZN(n20900) );
  INV_X1 U23834 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21012) );
  AOI22_X1 U23835 ( .A1(n21012), .A2(keyinput242), .B1(keyinput134), .B2(
        n21043), .ZN(n20895) );
  OAI221_X1 U23836 ( .B1(n21012), .B2(keyinput242), .C1(n21043), .C2(
        keyinput134), .A(n20895), .ZN(n20899) );
  XOR2_X1 U23837 ( .A(n13881), .B(keyinput135), .Z(n20897) );
  XNOR2_X1 U23838 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B(keyinput209), .ZN(
        n20896) );
  NAND2_X1 U23839 ( .A1(n20897), .A2(n20896), .ZN(n20898) );
  NOR4_X1 U23840 ( .A1(n20901), .A2(n20900), .A3(n20899), .A4(n20898), .ZN(
        n20931) );
  INV_X1 U23841 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n20903) );
  AOI22_X1 U23842 ( .A1(n20904), .A2(keyinput191), .B1(keyinput188), .B2(
        n20903), .ZN(n20902) );
  OAI221_X1 U23843 ( .B1(n20904), .B2(keyinput191), .C1(n20903), .C2(
        keyinput188), .A(n20902), .ZN(n20915) );
  AOI22_X1 U23844 ( .A1(n20985), .A2(keyinput150), .B1(keyinput187), .B2(
        n20906), .ZN(n20905) );
  OAI221_X1 U23845 ( .B1(n20985), .B2(keyinput150), .C1(n20906), .C2(
        keyinput187), .A(n20905), .ZN(n20914) );
  INV_X1 U23846 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n20908) );
  AOI22_X1 U23847 ( .A1(n20968), .A2(keyinput143), .B1(n20908), .B2(
        keyinput175), .ZN(n20907) );
  OAI221_X1 U23848 ( .B1(n20968), .B2(keyinput143), .C1(n20908), .C2(
        keyinput175), .A(n20907), .ZN(n20913) );
  AOI22_X1 U23849 ( .A1(n20911), .A2(keyinput230), .B1(keyinput219), .B2(
        n20910), .ZN(n20909) );
  OAI221_X1 U23850 ( .B1(n20911), .B2(keyinput230), .C1(n20910), .C2(
        keyinput219), .A(n20909), .ZN(n20912) );
  NOR4_X1 U23851 ( .A1(n20915), .A2(n20914), .A3(n20913), .A4(n20912), .ZN(
        n20930) );
  AOI22_X1 U23852 ( .A1(n20918), .A2(keyinput232), .B1(keyinput227), .B2(
        n20917), .ZN(n20916) );
  OAI221_X1 U23853 ( .B1(n20918), .B2(keyinput232), .C1(n20917), .C2(
        keyinput227), .A(n20916), .ZN(n20928) );
  INV_X1 U23854 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20921) );
  INV_X1 U23855 ( .A(DATAI_17_), .ZN(n20920) );
  AOI22_X1 U23856 ( .A1(n20921), .A2(keyinput250), .B1(keyinput231), .B2(
        n20920), .ZN(n20919) );
  OAI221_X1 U23857 ( .B1(n20921), .B2(keyinput250), .C1(n20920), .C2(
        keyinput231), .A(n20919), .ZN(n20927) );
  AOI22_X1 U23858 ( .A1(n20959), .A2(keyinput208), .B1(n21044), .B2(
        keyinput138), .ZN(n20922) );
  OAI221_X1 U23859 ( .B1(n20959), .B2(keyinput208), .C1(n21044), .C2(
        keyinput138), .A(n20922), .ZN(n20926) );
  XOR2_X1 U23860 ( .A(n13309), .B(keyinput254), .Z(n20924) );
  XNOR2_X1 U23861 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput192), .ZN(
        n20923) );
  NAND2_X1 U23862 ( .A1(n20924), .A2(n20923), .ZN(n20925) );
  NOR4_X1 U23863 ( .A1(n20928), .A2(n20927), .A3(n20926), .A4(n20925), .ZN(
        n20929) );
  NAND4_X1 U23864 ( .A1(n20932), .A2(n20931), .A3(n20930), .A4(n20929), .ZN(
        n20933) );
  NOR4_X1 U23865 ( .A1(n20936), .A2(n20935), .A3(n20934), .A4(n20933), .ZN(
        n21134) );
  AOI22_X1 U23866 ( .A1(n20939), .A2(keyinput27), .B1(n20938), .B2(keyinput57), 
        .ZN(n20937) );
  OAI221_X1 U23867 ( .B1(n20939), .B2(keyinput27), .C1(n20938), .C2(keyinput57), .A(n20937), .ZN(n20943) );
  XOR2_X1 U23868 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput64), .Z(
        n20942) );
  XNOR2_X1 U23869 ( .A(n20940), .B(keyinput53), .ZN(n20941) );
  OR3_X1 U23870 ( .A1(n20943), .A2(n20942), .A3(n20941), .ZN(n20951) );
  AOI22_X1 U23871 ( .A1(n20945), .A2(keyinput127), .B1(keyinput7), .B2(n13881), 
        .ZN(n20944) );
  OAI221_X1 U23872 ( .B1(n20945), .B2(keyinput127), .C1(n13881), .C2(keyinput7), .A(n20944), .ZN(n20950) );
  AOI22_X1 U23873 ( .A1(n20948), .A2(keyinput84), .B1(n20947), .B2(keyinput97), 
        .ZN(n20946) );
  OAI221_X1 U23874 ( .B1(n20948), .B2(keyinput84), .C1(n20947), .C2(keyinput97), .A(n20946), .ZN(n20949) );
  NOR3_X1 U23875 ( .A1(n20951), .A2(n20950), .A3(n20949), .ZN(n21000) );
  AOI22_X1 U23876 ( .A1(n20954), .A2(keyinput34), .B1(keyinput65), .B2(n20953), 
        .ZN(n20952) );
  OAI221_X1 U23877 ( .B1(n20954), .B2(keyinput34), .C1(n20953), .C2(keyinput65), .A(n20952), .ZN(n20965) );
  AOI22_X1 U23878 ( .A1(n10581), .A2(keyinput5), .B1(keyinput42), .B2(n20956), 
        .ZN(n20955) );
  OAI221_X1 U23879 ( .B1(n10581), .B2(keyinput5), .C1(n20956), .C2(keyinput42), 
        .A(n20955), .ZN(n20964) );
  INV_X1 U23880 ( .A(P3_UWORD_REG_7__SCAN_IN), .ZN(n20958) );
  AOI22_X1 U23881 ( .A1(n20959), .A2(keyinput80), .B1(keyinput118), .B2(n20958), .ZN(n20957) );
  OAI221_X1 U23882 ( .B1(n20959), .B2(keyinput80), .C1(n20958), .C2(
        keyinput118), .A(n20957), .ZN(n20963) );
  XNOR2_X1 U23883 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B(keyinput79), .ZN(
        n20961) );
  XNOR2_X1 U23884 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput108), .ZN(n20960)
         );
  NAND2_X1 U23885 ( .A1(n20961), .A2(n20960), .ZN(n20962) );
  NOR4_X1 U23886 ( .A1(n20965), .A2(n20964), .A3(n20963), .A4(n20962), .ZN(
        n20999) );
  AOI22_X1 U23887 ( .A1(n20968), .A2(keyinput15), .B1(keyinput71), .B2(n20967), 
        .ZN(n20966) );
  OAI221_X1 U23888 ( .B1(n20968), .B2(keyinput15), .C1(n20967), .C2(keyinput71), .A(n20966), .ZN(n20980) );
  AOI22_X1 U23889 ( .A1(n13367), .A2(keyinput55), .B1(keyinput31), .B2(n20970), 
        .ZN(n20969) );
  OAI221_X1 U23890 ( .B1(n13367), .B2(keyinput55), .C1(n20970), .C2(keyinput31), .A(n20969), .ZN(n20979) );
  AOI22_X1 U23891 ( .A1(n20973), .A2(keyinput56), .B1(keyinput62), .B2(n20972), 
        .ZN(n20971) );
  OAI221_X1 U23892 ( .B1(n20973), .B2(keyinput56), .C1(n20972), .C2(keyinput62), .A(n20971), .ZN(n20978) );
  INV_X1 U23893 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n20976) );
  AOI22_X1 U23894 ( .A1(n20976), .A2(keyinput3), .B1(keyinput50), .B2(n20975), 
        .ZN(n20974) );
  OAI221_X1 U23895 ( .B1(n20976), .B2(keyinput3), .C1(n20975), .C2(keyinput50), 
        .A(n20974), .ZN(n20977) );
  NOR4_X1 U23896 ( .A1(n20980), .A2(n20979), .A3(n20978), .A4(n20977), .ZN(
        n20998) );
  AOI22_X1 U23897 ( .A1(n20983), .A2(keyinput26), .B1(n20982), .B2(keyinput58), 
        .ZN(n20981) );
  OAI221_X1 U23898 ( .B1(n20983), .B2(keyinput26), .C1(n20982), .C2(keyinput58), .A(n20981), .ZN(n20996) );
  AOI22_X1 U23899 ( .A1(n20986), .A2(keyinput85), .B1(n20985), .B2(keyinput22), 
        .ZN(n20984) );
  OAI221_X1 U23900 ( .B1(n20986), .B2(keyinput85), .C1(n20985), .C2(keyinput22), .A(n20984), .ZN(n20995) );
  AOI22_X1 U23901 ( .A1(n20989), .A2(keyinput123), .B1(keyinput111), .B2(
        n20988), .ZN(n20987) );
  OAI221_X1 U23902 ( .B1(n20989), .B2(keyinput123), .C1(n20988), .C2(
        keyinput111), .A(n20987), .ZN(n20994) );
  INV_X1 U23903 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n20992) );
  AOI22_X1 U23904 ( .A1(n20992), .A2(keyinput72), .B1(n20991), .B2(keyinput89), 
        .ZN(n20990) );
  OAI221_X1 U23905 ( .B1(n20992), .B2(keyinput72), .C1(n20991), .C2(keyinput89), .A(n20990), .ZN(n20993) );
  NOR4_X1 U23906 ( .A1(n20996), .A2(n20995), .A3(n20994), .A4(n20993), .ZN(
        n20997) );
  NAND4_X1 U23907 ( .A1(n21000), .A2(n20999), .A3(n20998), .A4(n20997), .ZN(
        n21133) );
  AOI22_X1 U23908 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(keyinput100), .B1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .B2(keyinput117), .ZN(n21001) );
  OAI221_X1 U23909 ( .B1(P2_DATAWIDTH_REG_31__SCAN_IN), .B2(keyinput100), .C1(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .C2(keyinput117), .A(n21001), .ZN(
        n21008) );
  AOI22_X1 U23910 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(keyinput39), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(keyinput25), .ZN(n21002) );
  OAI221_X1 U23911 ( .B1(P2_EAX_REG_9__SCAN_IN), .B2(keyinput39), .C1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .C2(keyinput25), .A(n21002), .ZN(
        n21007) );
  AOI22_X1 U23912 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(keyinput67), .B1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(keyinput38), .ZN(n21003) );
  OAI221_X1 U23913 ( .B1(P3_EAX_REG_19__SCAN_IN), .B2(keyinput67), .C1(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(keyinput38), .A(n21003), .ZN(
        n21006) );
  AOI22_X1 U23914 ( .A1(BUF1_REG_1__SCAN_IN), .A2(keyinput70), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(keyinput11), .ZN(n21004) );
  OAI221_X1 U23915 ( .B1(BUF1_REG_1__SCAN_IN), .B2(keyinput70), .C1(
        P1_ADDRESS_REG_3__SCAN_IN), .C2(keyinput11), .A(n21004), .ZN(n21005)
         );
  NOR4_X1 U23916 ( .A1(n21008), .A2(n21007), .A3(n21006), .A4(n21005), .ZN(
        n21131) );
  OAI22_X1 U23917 ( .A1(P2_ADDRESS_REG_5__SCAN_IN), .A2(keyinput104), .B1(
        BUF2_REG_18__SCAN_IN), .B2(keyinput125), .ZN(n21009) );
  AOI221_X1 U23918 ( .B1(P2_ADDRESS_REG_5__SCAN_IN), .B2(keyinput104), .C1(
        keyinput125), .C2(BUF2_REG_18__SCAN_IN), .A(n21009), .ZN(n21022) );
  OAI22_X1 U23919 ( .A1(n21012), .A2(keyinput114), .B1(n21011), .B2(
        keyinput120), .ZN(n21010) );
  AOI221_X1 U23920 ( .B1(n21012), .B2(keyinput114), .C1(keyinput120), .C2(
        n21011), .A(n21010), .ZN(n21021) );
  OAI22_X1 U23921 ( .A1(n21015), .A2(keyinput43), .B1(n21014), .B2(keyinput52), 
        .ZN(n21013) );
  AOI221_X1 U23922 ( .B1(n21015), .B2(keyinput43), .C1(keyinput52), .C2(n21014), .A(n21013), .ZN(n21020) );
  OAI22_X1 U23923 ( .A1(n21018), .A2(keyinput75), .B1(n21017), .B2(keyinput36), 
        .ZN(n21016) );
  AOI221_X1 U23924 ( .B1(n21018), .B2(keyinput75), .C1(keyinput36), .C2(n21017), .A(n21016), .ZN(n21019) );
  NAND4_X1 U23925 ( .A1(n21022), .A2(n21021), .A3(n21020), .A4(n21019), .ZN(
        n21055) );
  INV_X1 U23926 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n21025) );
  AOI22_X1 U23927 ( .A1(n21025), .A2(keyinput35), .B1(n21024), .B2(keyinput9), 
        .ZN(n21023) );
  OAI221_X1 U23928 ( .B1(n21025), .B2(keyinput35), .C1(n21024), .C2(keyinput9), 
        .A(n21023), .ZN(n21054) );
  OAI22_X1 U23929 ( .A1(n21028), .A2(keyinput121), .B1(n21027), .B2(keyinput37), .ZN(n21026) );
  AOI221_X1 U23930 ( .B1(n21028), .B2(keyinput121), .C1(keyinput37), .C2(
        n21027), .A(n21026), .ZN(n21035) );
  OAI22_X1 U23931 ( .A1(n10032), .A2(keyinput107), .B1(n21030), .B2(keyinput82), .ZN(n21029) );
  AOI221_X1 U23932 ( .B1(n10032), .B2(keyinput107), .C1(keyinput82), .C2(
        n21030), .A(n21029), .ZN(n21034) );
  OAI22_X1 U23933 ( .A1(n11599), .A2(keyinput0), .B1(n21032), .B2(keyinput76), 
        .ZN(n21031) );
  AOI221_X1 U23934 ( .B1(n11599), .B2(keyinput0), .C1(keyinput76), .C2(n21032), 
        .A(n21031), .ZN(n21033) );
  NAND3_X1 U23935 ( .A1(n21035), .A2(n21034), .A3(n21033), .ZN(n21053) );
  OAI22_X1 U23936 ( .A1(n21038), .A2(keyinput18), .B1(n21037), .B2(keyinput124), .ZN(n21036) );
  AOI221_X1 U23937 ( .B1(n21038), .B2(keyinput18), .C1(keyinput124), .C2(
        n21037), .A(n21036), .ZN(n21051) );
  INV_X1 U23938 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n21041) );
  OAI22_X1 U23939 ( .A1(n21041), .A2(keyinput33), .B1(n21040), .B2(keyinput92), 
        .ZN(n21039) );
  AOI221_X1 U23940 ( .B1(n21041), .B2(keyinput33), .C1(keyinput92), .C2(n21040), .A(n21039), .ZN(n21050) );
  OAI22_X1 U23941 ( .A1(n21044), .A2(keyinput10), .B1(n21043), .B2(keyinput6), 
        .ZN(n21042) );
  AOI221_X1 U23942 ( .B1(n21044), .B2(keyinput10), .C1(keyinput6), .C2(n21043), 
        .A(n21042), .ZN(n21049) );
  OAI22_X1 U23943 ( .A1(n21047), .A2(keyinput24), .B1(n21046), .B2(keyinput41), 
        .ZN(n21045) );
  AOI221_X1 U23944 ( .B1(n21047), .B2(keyinput24), .C1(keyinput41), .C2(n21046), .A(n21045), .ZN(n21048) );
  NAND4_X1 U23945 ( .A1(n21051), .A2(n21050), .A3(n21049), .A4(n21048), .ZN(
        n21052) );
  NOR4_X1 U23946 ( .A1(n21055), .A2(n21054), .A3(n21053), .A4(n21052), .ZN(
        n21130) );
  OAI22_X1 U23947 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(keyinput19), 
        .B1(keyinput98), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n21056) );
  AOI221_X1 U23948 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput19), 
        .C1(P1_EBX_REG_28__SCAN_IN), .C2(keyinput98), .A(n21056), .ZN(n21063)
         );
  OAI22_X1 U23949 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(keyinput109), 
        .B1(P3_REIP_REG_25__SCAN_IN), .B2(keyinput20), .ZN(n21057) );
  AOI221_X1 U23950 ( .B1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B2(keyinput109), 
        .C1(keyinput20), .C2(P3_REIP_REG_25__SCAN_IN), .A(n21057), .ZN(n21062)
         );
  OAI22_X1 U23951 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(keyinput45), 
        .B1(P3_LWORD_REG_11__SCAN_IN), .B2(keyinput61), .ZN(n21058) );
  AOI221_X1 U23952 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput45), 
        .C1(keyinput61), .C2(P3_LWORD_REG_11__SCAN_IN), .A(n21058), .ZN(n21061) );
  OAI22_X1 U23953 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(keyinput44), 
        .B1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B2(keyinput47), .ZN(n21059) );
  AOI221_X1 U23954 ( .B1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(keyinput44), 
        .C1(keyinput47), .C2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A(n21059), 
        .ZN(n21060) );
  NAND4_X1 U23955 ( .A1(n21063), .A2(n21062), .A3(n21061), .A4(n21060), .ZN(
        n21091) );
  OAI22_X1 U23956 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(keyinput74), 
        .B1(keyinput91), .B2(P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21064) );
  AOI221_X1 U23957 ( .B1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(keyinput74), 
        .C1(P2_DATAWIDTH_REG_19__SCAN_IN), .C2(keyinput91), .A(n21064), .ZN(
        n21071) );
  OAI22_X1 U23958 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(keyinput95), .B1(
        P2_EAX_REG_15__SCAN_IN), .B2(keyinput54), .ZN(n21065) );
  AOI221_X1 U23959 ( .B1(P2_EAX_REG_28__SCAN_IN), .B2(keyinput95), .C1(
        keyinput54), .C2(P2_EAX_REG_15__SCAN_IN), .A(n21065), .ZN(n21070) );
  OAI22_X1 U23960 ( .A1(BUF2_REG_25__SCAN_IN), .A2(keyinput2), .B1(keyinput110), .B2(P3_EAX_REG_3__SCAN_IN), .ZN(n21066) );
  AOI221_X1 U23961 ( .B1(BUF2_REG_25__SCAN_IN), .B2(keyinput2), .C1(
        P3_EAX_REG_3__SCAN_IN), .C2(keyinput110), .A(n21066), .ZN(n21069) );
  OAI22_X1 U23962 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(keyinput83), .B1(
        keyinput59), .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n21067) );
  AOI221_X1 U23963 ( .B1(P1_ADDRESS_REG_18__SCAN_IN), .B2(keyinput83), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput59), .A(n21067), .ZN(n21068) );
  NAND4_X1 U23964 ( .A1(n21071), .A2(n21070), .A3(n21069), .A4(n21068), .ZN(
        n21090) );
  OAI22_X1 U23965 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(keyinput1), .B1(
        keyinput86), .B2(P1_READREQUEST_REG_SCAN_IN), .ZN(n21072) );
  AOI221_X1 U23966 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(keyinput1), .C1(
        P1_READREQUEST_REG_SCAN_IN), .C2(keyinput86), .A(n21072), .ZN(n21079)
         );
  OAI22_X1 U23967 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(keyinput99), 
        .B1(keyinput116), .B2(P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n21073) );
  AOI221_X1 U23968 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput99), 
        .C1(P3_DATAWIDTH_REG_27__SCAN_IN), .C2(keyinput116), .A(n21073), .ZN(
        n21078) );
  OAI22_X1 U23969 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(keyinput87), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(keyinput4), .ZN(n21074) );
  AOI221_X1 U23970 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(keyinput87), .C1(
        keyinput4), .C2(P1_M_IO_N_REG_SCAN_IN), .A(n21074), .ZN(n21077) );
  OAI22_X1 U23971 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(keyinput14), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(keyinput60), .ZN(n21075) );
  AOI221_X1 U23972 ( .B1(P1_ADDRESS_REG_25__SCAN_IN), .B2(keyinput14), .C1(
        keyinput60), .C2(P1_UWORD_REG_6__SCAN_IN), .A(n21075), .ZN(n21076) );
  NAND4_X1 U23973 ( .A1(n21079), .A2(n21078), .A3(n21077), .A4(n21076), .ZN(
        n21089) );
  OAI22_X1 U23974 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(keyinput126), 
        .B1(keyinput49), .B2(P1_EAX_REG_22__SCAN_IN), .ZN(n21080) );
  AOI221_X1 U23975 ( .B1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput126), 
        .C1(P1_EAX_REG_22__SCAN_IN), .C2(keyinput49), .A(n21080), .ZN(n21087)
         );
  OAI22_X1 U23976 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(keyinput40), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(keyinput77), .ZN(n21081) );
  AOI221_X1 U23977 ( .B1(P2_REIP_REG_11__SCAN_IN), .B2(keyinput40), .C1(
        keyinput77), .C2(P1_DATAO_REG_30__SCAN_IN), .A(n21081), .ZN(n21086) );
  OAI22_X1 U23978 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(keyinput66), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(keyinput13), .ZN(n21082) );
  AOI221_X1 U23979 ( .B1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(keyinput66), 
        .C1(keyinput13), .C2(P1_DATAO_REG_3__SCAN_IN), .A(n21082), .ZN(n21085)
         );
  OAI22_X1 U23980 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(keyinput73), 
        .B1(P3_REIP_REG_22__SCAN_IN), .B2(keyinput16), .ZN(n21083) );
  AOI221_X1 U23981 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput73), 
        .C1(keyinput16), .C2(P3_REIP_REG_22__SCAN_IN), .A(n21083), .ZN(n21084)
         );
  NAND4_X1 U23982 ( .A1(n21087), .A2(n21086), .A3(n21085), .A4(n21084), .ZN(
        n21088) );
  NOR4_X1 U23983 ( .A1(n21091), .A2(n21090), .A3(n21089), .A4(n21088), .ZN(
        n21129) );
  OAI22_X1 U23984 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(keyinput105), .B1(
        keyinput96), .B2(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21092) );
  AOI221_X1 U23985 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(keyinput105), .C1(
        P1_DATAWIDTH_REG_15__SCAN_IN), .C2(keyinput96), .A(n21092), .ZN(n21099) );
  OAI22_X1 U23986 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(keyinput88), .B1(
        keyinput119), .B2(P1_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21093) );
  AOI221_X1 U23987 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(keyinput88), .C1(
        P1_DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput119), .A(n21093), .ZN(
        n21098) );
  OAI22_X1 U23988 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(keyinput46), .B1(
        keyinput23), .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n21094) );
  AOI221_X1 U23989 ( .B1(P3_REIP_REG_2__SCAN_IN), .B2(keyinput46), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput23), .A(n21094), .ZN(n21097) );
  OAI22_X1 U23990 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(keyinput48), .B1(
        P3_INSTQUEUE_REG_4__3__SCAN_IN), .B2(keyinput90), .ZN(n21095) );
  AOI221_X1 U23991 ( .B1(P1_EAX_REG_20__SCAN_IN), .B2(keyinput48), .C1(
        keyinput90), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(n21095), .ZN(
        n21096) );
  NAND4_X1 U23992 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        n21127) );
  OAI22_X1 U23993 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(keyinput122), 
        .B1(BUF2_REG_7__SCAN_IN), .B2(keyinput28), .ZN(n21100) );
  AOI221_X1 U23994 ( .B1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B2(keyinput122), 
        .C1(keyinput28), .C2(BUF2_REG_7__SCAN_IN), .A(n21100), .ZN(n21107) );
  OAI22_X1 U23995 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(keyinput93), .B1(
        keyinput68), .B2(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21101) );
  AOI221_X1 U23996 ( .B1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B2(keyinput93), 
        .C1(P1_ADDRESS_REG_21__SCAN_IN), .C2(keyinput68), .A(n21101), .ZN(
        n21106) );
  OAI22_X1 U23997 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput101), 
        .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput12), .ZN(n21102) );
  AOI221_X1 U23998 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput101), 
        .C1(keyinput12), .C2(P2_DATAO_REG_12__SCAN_IN), .A(n21102), .ZN(n21105) );
  OAI22_X1 U23999 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(keyinput63), .B1(
        keyinput29), .B2(P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21103) );
  AOI221_X1 U24000 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(keyinput63), .C1(
        P3_DATAWIDTH_REG_15__SCAN_IN), .C2(keyinput29), .A(n21103), .ZN(n21104) );
  NAND4_X1 U24001 ( .A1(n21107), .A2(n21106), .A3(n21105), .A4(n21104), .ZN(
        n21126) );
  OAI22_X1 U24002 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(keyinput115), 
        .B1(keyinput51), .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n21108) );
  AOI221_X1 U24003 ( .B1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B2(keyinput115), 
        .C1(P3_DATAO_REG_14__SCAN_IN), .C2(keyinput51), .A(n21108), .ZN(n21115) );
  OAI22_X1 U24004 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(keyinput21), .B1(
        P1_INSTQUEUE_REG_10__7__SCAN_IN), .B2(keyinput112), .ZN(n21109) );
  AOI221_X1 U24005 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(keyinput21), .C1(
        keyinput112), .C2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(n21109), .ZN(
        n21114) );
  OAI22_X1 U24006 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(keyinput113), .B1(
        P2_W_R_N_REG_SCAN_IN), .B2(keyinput30), .ZN(n21110) );
  AOI221_X1 U24007 ( .B1(P1_DATAO_REG_21__SCAN_IN), .B2(keyinput113), .C1(
        keyinput30), .C2(P2_W_R_N_REG_SCAN_IN), .A(n21110), .ZN(n21113) );
  OAI22_X1 U24008 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(keyinput94), 
        .B1(keyinput32), .B2(P1_EBX_REG_2__SCAN_IN), .ZN(n21111) );
  AOI221_X1 U24009 ( .B1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput94), 
        .C1(P1_EBX_REG_2__SCAN_IN), .C2(keyinput32), .A(n21111), .ZN(n21112)
         );
  NAND4_X1 U24010 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21125) );
  OAI22_X1 U24011 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(keyinput17), .B1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput8), .ZN(n21116) );
  AOI221_X1 U24012 ( .B1(P2_UWORD_REG_5__SCAN_IN), .B2(keyinput17), .C1(
        keyinput8), .C2(P1_BYTEENABLE_REG_1__SCAN_IN), .A(n21116), .ZN(n21123)
         );
  OAI22_X1 U24013 ( .A1(DATAI_17_), .A2(keyinput103), .B1(
        P2_DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput102), .ZN(n21117) );
  AOI221_X1 U24014 ( .B1(DATAI_17_), .B2(keyinput103), .C1(keyinput102), .C2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A(n21117), .ZN(n21122) );
  OAI22_X1 U24015 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(keyinput81), .B1(
        keyinput78), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n21118) );
  AOI221_X1 U24016 ( .B1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput81), 
        .C1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .C2(keyinput78), .A(n21118), 
        .ZN(n21121) );
  OAI22_X1 U24017 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(keyinput69), .B1(
        keyinput106), .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n21119) );
  AOI221_X1 U24018 ( .B1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B2(keyinput69), 
        .C1(P2_DATAO_REG_27__SCAN_IN), .C2(keyinput106), .A(n21119), .ZN(
        n21120) );
  NAND4_X1 U24019 ( .A1(n21123), .A2(n21122), .A3(n21121), .A4(n21120), .ZN(
        n21124) );
  NOR4_X1 U24020 ( .A1(n21127), .A2(n21126), .A3(n21125), .A4(n21124), .ZN(
        n21128) );
  NAND4_X1 U24021 ( .A1(n21131), .A2(n21130), .A3(n21129), .A4(n21128), .ZN(
        n21132) );
  NOR3_X1 U24022 ( .A1(n21134), .A2(n21133), .A3(n21132), .ZN(n21135) );
  XNOR2_X1 U24023 ( .A(n21136), .B(n21135), .ZN(P2_U3209) );
  AND2_X1 U12719 ( .A1(n10256), .A2(n12376), .ZN(n10350) );
  INV_X1 U11748 ( .A(n10431), .ZN(n20070) );
  INV_X2 U11366 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11599) );
  CLKBUF_X2 U13140 ( .A(n10433), .Z(n20079) );
  BUF_X1 U11354 ( .A(n13271), .Z(n14018) );
  CLKBUF_X1 U11248 ( .A(n10403), .Z(n11084) );
  INV_X1 U16483 ( .A(n13363), .ZN(n19144) );
  OR2_X1 U16443 ( .A1(n13244), .A2(n13246), .ZN(n13305) );
  AND2_X1 U16852 ( .A1(n14614), .A2(n14615), .ZN(n14617) );
  OR2_X1 U12703 ( .A1(n13244), .A2(n13256), .ZN(n15435) );
  BUF_X2 U11230 ( .A(n11566), .Z(n9798) );
  BUF_X2 U11251 ( .A(n10997), .Z(n11079) );
  CLKBUF_X1 U11268 ( .A(n11085), .Z(n9810) );
  NAND2_X1 U11282 ( .A1(n13754), .A2(n9902), .ZN(n13850) );
  AOI21_X1 U11361 ( .B1(n12462), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n12448), .ZN(n12677) );
  CLKBUF_X1 U11437 ( .A(n11492), .Z(n9789) );
  CLKBUF_X2 U11525 ( .A(n11454), .Z(n14070) );
  CLKBUF_X1 U12345 ( .A(n14121), .Z(n14122) );
  NAND2_X1 U12382 ( .A1(n14992), .A2(n13550), .ZN(n14993) );
  CLKBUF_X1 U12737 ( .A(n17334), .Z(n17343) );
  CLKBUF_X1 U13793 ( .A(n16378), .Z(n16384) );
  NOR2_X2 U15509 ( .A1(n15429), .A2(n15430), .ZN(n19174) );
  NAND3_X2 U16813 ( .A1(n19771), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19624), 
        .ZN(n15430) );
endmodule

